module aes_cipher_top (
	clk, 
	rst, 
	ld, 
	done, 
	key_127_, 
	key_126_, 
	key_125_, 
	key_124_, 
	key_123_, 
	key_122_, 
	key_121_, 
	key_120_, 
	key_119_, 
	key_118_, 
	key_117_, 
	key_116_, 
	key_115_, 
	key_114_, 
	key_113_, 
	key_112_, 
	key_111_, 
	key_110_, 
	key_109_, 
	key_108_, 
	key_107_, 
	key_106_, 
	key_105_, 
	key_104_, 
	key_103_, 
	key_102_, 
	key_101_, 
	key_100_, 
	key_99_, 
	key_98_, 
	key_97_, 
	key_96_, 
	key_95_, 
	key_94_, 
	key_93_, 
	key_92_, 
	key_91_, 
	key_90_, 
	key_89_, 
	key_88_, 
	key_87_, 
	key_86_, 
	key_85_, 
	key_84_, 
	key_83_, 
	key_82_, 
	key_81_, 
	key_80_, 
	key_79_, 
	key_78_, 
	key_77_, 
	key_76_, 
	key_75_, 
	key_74_, 
	key_73_, 
	key_72_, 
	key_71_, 
	key_70_, 
	key_69_, 
	key_68_, 
	key_67_, 
	key_66_, 
	key_65_, 
	key_64_, 
	key_63_, 
	key_62_, 
	key_61_, 
	key_60_, 
	key_59_, 
	key_58_, 
	key_57_, 
	key_56_, 
	key_55_, 
	key_54_, 
	key_53_, 
	key_52_, 
	key_51_, 
	key_50_, 
	key_49_, 
	key_48_, 
	key_47_, 
	key_46_, 
	key_45_, 
	key_44_, 
	key_43_, 
	key_42_, 
	key_41_, 
	key_40_, 
	key_39_, 
	key_38_, 
	key_37_, 
	key_36_, 
	key_35_, 
	key_34_, 
	key_33_, 
	key_32_, 
	key_31_, 
	key_30_, 
	key_29_, 
	key_28_, 
	key_27_, 
	key_26_, 
	key_25_, 
	key_24_, 
	key_23_, 
	key_22_, 
	key_21_, 
	key_20_, 
	key_19_, 
	key_18_, 
	key_17_, 
	key_16_, 
	key_15_, 
	key_14_, 
	key_13_, 
	key_12_, 
	key_11_, 
	key_10_, 
	key_9_, 
	key_8_, 
	key_7_, 
	key_6_, 
	key_5_, 
	key_4_, 
	key_3_, 
	key_2_, 
	key_1_, 
	key_0_, 
	text_in_127_, 
	text_in_126_, 
	text_in_125_, 
	text_in_124_, 
	text_in_123_, 
	text_in_122_, 
	text_in_121_, 
	text_in_120_, 
	text_in_119_, 
	text_in_118_, 
	text_in_117_, 
	text_in_116_, 
	text_in_115_, 
	text_in_114_, 
	text_in_113_, 
	text_in_112_, 
	text_in_111_, 
	text_in_110_, 
	text_in_109_, 
	text_in_108_, 
	text_in_107_, 
	text_in_106_, 
	text_in_105_, 
	text_in_104_, 
	text_in_103_, 
	text_in_102_, 
	text_in_101_, 
	text_in_100_, 
	text_in_99_, 
	text_in_98_, 
	text_in_97_, 
	text_in_96_, 
	text_in_95_, 
	text_in_94_, 
	text_in_93_, 
	text_in_92_, 
	text_in_91_, 
	text_in_90_, 
	text_in_89_, 
	text_in_88_, 
	text_in_87_, 
	text_in_86_, 
	text_in_85_, 
	text_in_84_, 
	text_in_83_, 
	text_in_82_, 
	text_in_81_, 
	text_in_80_, 
	text_in_79_, 
	text_in_78_, 
	text_in_77_, 
	text_in_76_, 
	text_in_75_, 
	text_in_74_, 
	text_in_73_, 
	text_in_72_, 
	text_in_71_, 
	text_in_70_, 
	text_in_69_, 
	text_in_68_, 
	text_in_67_, 
	text_in_66_, 
	text_in_65_, 
	text_in_64_, 
	text_in_63_, 
	text_in_62_, 
	text_in_61_, 
	text_in_60_, 
	text_in_59_, 
	text_in_58_, 
	text_in_57_, 
	text_in_56_, 
	text_in_55_, 
	text_in_54_, 
	text_in_53_, 
	text_in_52_, 
	text_in_51_, 
	text_in_50_, 
	text_in_49_, 
	text_in_48_, 
	text_in_47_, 
	text_in_46_, 
	text_in_45_, 
	text_in_44_, 
	text_in_43_, 
	text_in_42_, 
	text_in_41_, 
	text_in_40_, 
	text_in_39_, 
	text_in_38_, 
	text_in_37_, 
	text_in_36_, 
	text_in_35_, 
	text_in_34_, 
	text_in_33_, 
	text_in_32_, 
	text_in_31_, 
	text_in_30_, 
	text_in_29_, 
	text_in_28_, 
	text_in_27_, 
	text_in_26_, 
	text_in_25_, 
	text_in_24_, 
	text_in_23_, 
	text_in_22_, 
	text_in_21_, 
	text_in_20_, 
	text_in_19_, 
	text_in_18_, 
	text_in_17_, 
	text_in_16_, 
	text_in_15_, 
	text_in_14_, 
	text_in_13_, 
	text_in_12_, 
	text_in_11_, 
	text_in_10_, 
	text_in_9_, 
	text_in_8_, 
	text_in_7_, 
	text_in_6_, 
	text_in_5_, 
	text_in_4_, 
	text_in_3_, 
	text_in_2_, 
	text_in_1_, 
	text_in_0_, 
	text_out_127_, 
	text_out_126_, 
	text_out_125_, 
	text_out_124_, 
	text_out_123_, 
	text_out_122_, 
	text_out_121_, 
	text_out_120_, 
	text_out_119_, 
	text_out_118_, 
	text_out_117_, 
	text_out_116_, 
	text_out_115_, 
	text_out_114_, 
	text_out_113_, 
	text_out_112_, 
	text_out_111_, 
	text_out_110_, 
	text_out_109_, 
	text_out_108_, 
	text_out_107_, 
	text_out_106_, 
	text_out_105_, 
	text_out_104_, 
	text_out_103_, 
	text_out_102_, 
	text_out_101_, 
	text_out_100_, 
	text_out_99_, 
	text_out_98_, 
	text_out_97_, 
	text_out_96_, 
	text_out_95_, 
	text_out_94_, 
	text_out_93_, 
	text_out_92_, 
	text_out_91_, 
	text_out_90_, 
	text_out_89_, 
	text_out_88_, 
	text_out_87_, 
	text_out_86_, 
	text_out_85_, 
	text_out_84_, 
	text_out_83_, 
	text_out_82_, 
	text_out_81_, 
	text_out_80_, 
	text_out_79_, 
	text_out_78_, 
	text_out_77_, 
	text_out_76_, 
	text_out_75_, 
	text_out_74_, 
	text_out_73_, 
	text_out_72_, 
	text_out_71_, 
	text_out_70_, 
	text_out_69_, 
	text_out_68_, 
	text_out_67_, 
	text_out_66_, 
	text_out_65_, 
	text_out_64_, 
	text_out_63_, 
	text_out_62_, 
	text_out_61_, 
	text_out_60_, 
	text_out_59_, 
	text_out_58_, 
	text_out_57_, 
	text_out_56_, 
	text_out_55_, 
	text_out_54_, 
	text_out_53_, 
	text_out_52_, 
	text_out_51_, 
	text_out_50_, 
	text_out_49_, 
	text_out_48_, 
	text_out_47_, 
	text_out_46_, 
	text_out_45_, 
	text_out_44_, 
	text_out_43_, 
	text_out_42_, 
	text_out_41_, 
	text_out_40_, 
	text_out_39_, 
	text_out_38_, 
	text_out_37_, 
	text_out_36_, 
	text_out_35_, 
	text_out_34_, 
	text_out_33_, 
	text_out_32_, 
	text_out_31_, 
	text_out_30_, 
	text_out_29_, 
	text_out_28_, 
	text_out_27_, 
	text_out_26_, 
	text_out_25_, 
	text_out_24_, 
	text_out_23_, 
	text_out_22_, 
	text_out_21_, 
	text_out_20_, 
	text_out_19_, 
	text_out_18_, 
	text_out_17_, 
	text_out_16_, 
	text_out_15_, 
	text_out_14_, 
	text_out_13_, 
	text_out_12_, 
	text_out_11_, 
	text_out_10_, 
	text_out_9_, 
	text_out_8_, 
	text_out_7_, 
	text_out_6_, 
	text_out_5_, 
	text_out_4_, 
	text_out_3_, 
	text_out_2_, 
	text_out_1_, 
	text_out_0_, 
	SE, 
	SI, 
	SO);
   input clk;
   input rst;
   input ld;
   output done;
   input key_127_;
   input key_126_;
   input key_125_;
   input key_124_;
   input key_123_;
   input key_122_;
   input key_121_;
   input key_120_;
   input key_119_;
   input key_118_;
   input key_117_;
   input key_116_;
   input key_115_;
   input key_114_;
   input key_113_;
   input key_112_;
   input key_111_;
   input key_110_;
   input key_109_;
   input key_108_;
   input key_107_;
   input key_106_;
   input key_105_;
   input key_104_;
   input key_103_;
   input key_102_;
   input key_101_;
   input key_100_;
   input key_99_;
   input key_98_;
   input key_97_;
   input key_96_;
   input key_95_;
   input key_94_;
   input key_93_;
   input key_92_;
   input key_91_;
   input key_90_;
   input key_89_;
   input key_88_;
   input key_87_;
   input key_86_;
   input key_85_;
   input key_84_;
   input key_83_;
   input key_82_;
   input key_81_;
   input key_80_;
   input key_79_;
   input key_78_;
   input key_77_;
   input key_76_;
   input key_75_;
   input key_74_;
   input key_73_;
   input key_72_;
   input key_71_;
   input key_70_;
   input key_69_;
   input key_68_;
   input key_67_;
   input key_66_;
   input key_65_;
   input key_64_;
   input key_63_;
   input key_62_;
   input key_61_;
   input key_60_;
   input key_59_;
   input key_58_;
   input key_57_;
   input key_56_;
   input key_55_;
   input key_54_;
   input key_53_;
   input key_52_;
   input key_51_;
   input key_50_;
   input key_49_;
   input key_48_;
   input key_47_;
   input key_46_;
   input key_45_;
   input key_44_;
   input key_43_;
   input key_42_;
   input key_41_;
   input key_40_;
   input key_39_;
   input key_38_;
   input key_37_;
   input key_36_;
   input key_35_;
   input key_34_;
   input key_33_;
   input key_32_;
   input key_31_;
   input key_30_;
   input key_29_;
   input key_28_;
   input key_27_;
   input key_26_;
   input key_25_;
   input key_24_;
   input key_23_;
   input key_22_;
   input key_21_;
   input key_20_;
   input key_19_;
   input key_18_;
   input key_17_;
   input key_16_;
   input key_15_;
   input key_14_;
   input key_13_;
   input key_12_;
   input key_11_;
   input key_10_;
   input key_9_;
   input key_8_;
   input key_7_;
   input key_6_;
   input key_5_;
   input key_4_;
   input key_3_;
   input key_2_;
   input key_1_;
   input key_0_;
   input text_in_127_;
   input text_in_126_;
   input text_in_125_;
   input text_in_124_;
   input text_in_123_;
   input text_in_122_;
   input text_in_121_;
   input text_in_120_;
   input text_in_119_;
   input text_in_118_;
   input text_in_117_;
   input text_in_116_;
   input text_in_115_;
   input text_in_114_;
   input text_in_113_;
   input text_in_112_;
   input text_in_111_;
   input text_in_110_;
   input text_in_109_;
   input text_in_108_;
   input text_in_107_;
   input text_in_106_;
   input text_in_105_;
   input text_in_104_;
   input text_in_103_;
   input text_in_102_;
   input text_in_101_;
   input text_in_100_;
   input text_in_99_;
   input text_in_98_;
   input text_in_97_;
   input text_in_96_;
   input text_in_95_;
   input text_in_94_;
   input text_in_93_;
   input text_in_92_;
   input text_in_91_;
   input text_in_90_;
   input text_in_89_;
   input text_in_88_;
   input text_in_87_;
   input text_in_86_;
   input text_in_85_;
   input text_in_84_;
   input text_in_83_;
   input text_in_82_;
   input text_in_81_;
   input text_in_80_;
   input text_in_79_;
   input text_in_78_;
   input text_in_77_;
   input text_in_76_;
   input text_in_75_;
   input text_in_74_;
   input text_in_73_;
   input text_in_72_;
   input text_in_71_;
   input text_in_70_;
   input text_in_69_;
   input text_in_68_;
   input text_in_67_;
   input text_in_66_;
   input text_in_65_;
   input text_in_64_;
   input text_in_63_;
   input text_in_62_;
   input text_in_61_;
   input text_in_60_;
   input text_in_59_;
   input text_in_58_;
   input text_in_57_;
   input text_in_56_;
   input text_in_55_;
   input text_in_54_;
   input text_in_53_;
   input text_in_52_;
   input text_in_51_;
   input text_in_50_;
   input text_in_49_;
   input text_in_48_;
   input text_in_47_;
   input text_in_46_;
   input text_in_45_;
   input text_in_44_;
   input text_in_43_;
   input text_in_42_;
   input text_in_41_;
   input text_in_40_;
   input text_in_39_;
   input text_in_38_;
   input text_in_37_;
   input text_in_36_;
   input text_in_35_;
   input text_in_34_;
   input text_in_33_;
   input text_in_32_;
   input text_in_31_;
   input text_in_30_;
   input text_in_29_;
   input text_in_28_;
   input text_in_27_;
   input text_in_26_;
   input text_in_25_;
   input text_in_24_;
   input text_in_23_;
   input text_in_22_;
   input text_in_21_;
   input text_in_20_;
   input text_in_19_;
   input text_in_18_;
   input text_in_17_;
   input text_in_16_;
   input text_in_15_;
   input text_in_14_;
   input text_in_13_;
   input text_in_12_;
   input text_in_11_;
   input text_in_10_;
   input text_in_9_;
   input text_in_8_;
   input text_in_7_;
   input text_in_6_;
   input text_in_5_;
   input text_in_4_;
   input text_in_3_;
   input text_in_2_;
   input text_in_1_;
   input text_in_0_;
   output text_out_127_;
   output text_out_126_;
   output text_out_125_;
   output text_out_124_;
   output text_out_123_;
   output text_out_122_;
   output text_out_121_;
   output text_out_120_;
   output text_out_119_;
   output text_out_118_;
   output text_out_117_;
   output text_out_116_;
   output text_out_115_;
   output text_out_114_;
   output text_out_113_;
   output text_out_112_;
   output text_out_111_;
   output text_out_110_;
   output text_out_109_;
   output text_out_108_;
   output text_out_107_;
   output text_out_106_;
   output text_out_105_;
   output text_out_104_;
   output text_out_103_;
   output text_out_102_;
   output text_out_101_;
   output text_out_100_;
   output text_out_99_;
   output text_out_98_;
   output text_out_97_;
   output text_out_96_;
   output text_out_95_;
   output text_out_94_;
   output text_out_93_;
   output text_out_92_;
   output text_out_91_;
   output text_out_90_;
   output text_out_89_;
   output text_out_88_;
   output text_out_87_;
   output text_out_86_;
   output text_out_85_;
   output text_out_84_;
   output text_out_83_;
   output text_out_82_;
   output text_out_81_;
   output text_out_80_;
   output text_out_79_;
   output text_out_78_;
   output text_out_77_;
   output text_out_76_;
   output text_out_75_;
   output text_out_74_;
   output text_out_73_;
   output text_out_72_;
   output text_out_71_;
   output text_out_70_;
   output text_out_69_;
   output text_out_68_;
   output text_out_67_;
   output text_out_66_;
   output text_out_65_;
   output text_out_64_;
   output text_out_63_;
   output text_out_62_;
   output text_out_61_;
   output text_out_60_;
   output text_out_59_;
   output text_out_58_;
   output text_out_57_;
   output text_out_56_;
   output text_out_55_;
   output text_out_54_;
   output text_out_53_;
   output text_out_52_;
   output text_out_51_;
   output text_out_50_;
   output text_out_49_;
   output text_out_48_;
   output text_out_47_;
   output text_out_46_;
   output text_out_45_;
   output text_out_44_;
   output text_out_43_;
   output text_out_42_;
   output text_out_41_;
   output text_out_40_;
   output text_out_39_;
   output text_out_38_;
   output text_out_37_;
   output text_out_36_;
   output text_out_35_;
   output text_out_34_;
   output text_out_33_;
   output text_out_32_;
   output text_out_31_;
   output text_out_30_;
   output text_out_29_;
   output text_out_28_;
   output text_out_27_;
   output text_out_26_;
   output text_out_25_;
   output text_out_24_;
   output text_out_23_;
   output text_out_22_;
   output text_out_21_;
   output text_out_20_;
   output text_out_19_;
   output text_out_18_;
   output text_out_17_;
   output text_out_16_;
   output text_out_15_;
   output text_out_14_;
   output text_out_13_;
   output text_out_12_;
   output text_out_11_;
   output text_out_10_;
   output text_out_9_;
   output text_out_8_;
   output text_out_7_;
   output text_out_6_;
   output text_out_5_;
   output text_out_4_;
   output text_out_3_;
   output text_out_2_;
   output text_out_1_;
   output text_out_0_;
   input SE;
   input SI;
   output SO;

   // Internal wires
   wire FE_PSN8338_n19791;
   wire FE_PSN8337_n16909;
   wire FE_PSN8336_n23340;
   wire FE_PSN8335_n17606;
   wire FE_PSN8334_n15539;
   wire FE_PSN8333_n18478;
   wire FE_PSN8332_n23879;
   wire FE_PSN8331_n24113;
   wire FE_PSN8330_n17761;
   wire FE_PSN8329_n21638;
   wire FE_PSN8328_n20260;
   wire FE_PSN8327_n24562;
   wire FE_PSN8326_n21455;
   wire FE_PSN8325_FE_OFN28811_n19170;
   wire FE_PSN8324_n15987;
   wire FE_PSN8323_n22543;
   wire FE_PSN8322_n25105;
   wire FE_PSN8321_n26520;
   wire FE_PSN8320_n18176;
   wire FE_PSN8319_n21725;
   wire FE_PSN8318_n21455;
   wire FE_PSN8317_n20850;
   wire FE_PSN8316_n23781;
   wire FE_PSN8315_FE_OFN16135_sa22_4;
   wire FE_PSN8314_n25722;
   wire FE_PSN8313_FE_OCPN29469_n17747;
   wire FE_PSN8312_n21442;
   wire FE_PSN8311_n25105;
   wire FE_PSN8310_n17473;
   wire FE_PSN8309_n21372;
   wire FE_PSN8308_n22624;
   wire FE_PSN8307_FE_OFN27207_w3_30;
   wire FE_PSN8306_FE_OFN28689_sa03_5;
   wire FE_PSN8305_n21217;
   wire FE_PSN8304_n24565;
   wire FE_PSN8303_n19222;
   wire FE_PSN8302_n24562;
   wire FE_PSN8301_n23197;
   wire FE_PSN8300_n26482;
   wire FE_PSN8299_FE_OFN4_w3_22;
   wire FE_PSN8298_FE_OFN27151_n;
   wire FE_PSN8297_FE_OFN8_w3_14;
   wire FE_PSN8296_FE_OFN26588_n24062;
   wire FE_PSN8295_FE_OFN28669_sa31_5;
   wire FE_PSN8294_n22310;
   wire FE_PSN8293_n25317;
   wire FE_PSN8292_FE_OFN26041_w3_17;
   wire FE_PSN8291_n26404;
   wire FE_PSN8290_n21439;
   wire FE_PSN8289_FE_OFN28514_sa00_1;
   wire FE_PSN8288_n17275;
   wire FE_PSN8287_FE_OCPN27494_n26479;
   wire FE_PSN8286_FE_OCPN29260_sa00_5;
   wire FE_PSN8285_FE_OCPN29463_n;
   wire FE_PSN8284_n21438;
   wire FE_PSN8283_n22629;
   wire FE_PSN8282_n21154;
   wire FE_PSN8281_n25118;
   wire FE_PSN8280_n15660;
   wire FE_PSN8279_FE_OCPN27292_n25389;
   wire FE_PSN8278_n25605;
   wire FE_PSN8277_n16099;
   wire FE_PSN8276_FE_OFN28712_n;
   wire FE_PSN8275_FE_OCPN27818_n17267;
   wire FE_PSN8274_n21164;
   wire FE_PSN8273_n24087;
   wire FE_PSN8272_n20428;
   wire FE_PSN8271_n15924;
   wire FE_PSN8270_n26027;
   wire FE_OCPN8269_FE_OFN16136_sa02_5;
   wire FE_OCPN8268_n26632;
   wire FE_OCPN8267_n16069;
   wire FE_OCPN8266_sa21_2;
   wire FE_OCPN8265_n24362;
   wire FE_OCPN8264_n13890;
   wire FE_OCPN8263_n25039;
   wire FE_OCPN8262_n21726;
   wire FE_OCPN8261_n26513;
   wire FE_OCPN8260_n26335;
   wire FE_OCPN8259_FE_OFN28686_FE_OCPN27812;
   wire FE_OCPN8258_n26572;
   wire FE_OCPN8257_n18178;
   wire FE_OCPN8256_n16873;
   wire FE_OCPN8255_n21002;
   wire FE_OCPN8254_w3_3;
   wire FE_OCPN8253_n17149;
   wire FE_OCPN8252_FE_OFN28661_w3_7;
   wire FE_OCPN8251_FE_OFN28672_sa01_2;
   wire FE_OCPN8250_n22692;
   wire FE_OCPN8249_n26944;
   wire FE_OCPN8248_n16145;
   wire FE_OCPN8247_n21317;
   wire FE_OCPN8246_n27143;
   wire FE_OCPN8245_n25295;
   wire FE_OCPN8244_n25778;
   wire FE_OCPN8243_n24899;
   wire FE_OCPN8242_n20527;
   wire FE_OCPN8241_n22041;
   wire FE_OCPN8240_n17618;
   wire FE_OCPN8239_n24844;
   wire FE_OCPN8238_n26472;
   wire FE_OCPN8237_n21561;
   wire FE_OCPN8236_n22438;
   wire FE_OCPN8235_n24589;
   wire FE_OCPN8234_n25199;
   wire FE_OCPN8233_n21647;
   wire FE_OCPN8232_FE_OFN27206_w3_30;
   wire FE_OCPN8231_n20522;
   wire FE_OCPN8230_n20993;
   wire FE_OCPN8229_n25750;
   wire FE_OCPN8228_n24165;
   wire FE_OCPN8227_n25950;
   wire FE_OCPN8226_n23113;
   wire FE_OCPN8225_n26172;
   wire FE_OCPN8224_n22773;
   wire FE_OCPN8223_n16063;
   wire FE_OCPN8222_n27006;
   wire FE_OCPN8221_n26825;
   wire FE_OCPN8220_n26198;
   wire FE_OCPN8219_n22197;
   wire FE_OCPN8218_n25507;
   wire FE_OCPN8217_n26319;
   wire FE_OCPN8216_n13916;
   wire FE_OCPN8215_n25287;
   wire FE_OCPN8214_n27185;
   wire FE_OCPN8213_FE_OFN29234_n16996;
   wire FE_OCPN8212_n26261;
   wire FE_OCPN8211_n24166;
   wire FE_OCPN8210_n25287;
   wire FE_OCPN8209_n26051;
   wire FE_OCPN8208_n27094;
   wire FE_OCPN8207_n18497;
   wire FE_OCPN8206_n25544;
   wire FE_OCPN29590_n449;
   wire FE_OCPN29589_n426;
   wire FE_OCPN29588_n457;
   wire FE_OCPN29587_n26857;
   wire FE_OCPN29586_n26857;
   wire FE_RN_287_0;
   wire FE_RN_286_0;
   wire FE_RN_285_0;
   wire FE_RN_284_0;
   wire FE_RN_283_0;
   wire FE_OCPN29585_n22281;
   wire FE_RN_282_0;
   wire FE_OCPN29584_n;
   wire FE_OCPN29583_n15422;
   wire FE_RN_281_0;
   wire FE_RN_280_0;
   wire FE_RN_279_0;
   wire FE_RN_278_0;
   wire FE_OCPN29581_n16097;
   wire FE_OCPN29580_n;
   wire FE_OCPN29579_n18837;
   wire FE_OCPN29578_FE_OFN27214_w3_17;
   wire FE_OCPN29577_n24298;
   wire FE_OCPN29576_n26930;
   wire FE_OCPN29574_n484;
   wire FE_OCPN29573_n15184;
   wire FE_OCPN29572_n24468;
   wire FE_OCPN29571_n26355;
   wire FE_OCPN29570_n15423;
   wire FE_OCPN29569_n18947;
   wire FE_RN_277_0;
   wire FE_RN_276_0;
   wire FE_OCPN29568_n18257;
   wire FE_OCPN29567_n23806;
   wire FE_OCPN29565_n432;
   wire FE_OCPN29564_n16012;
   wire FE_OCPN29563_n18602;
   wire FE_RN_275_0;
   wire FE_RN_274_0;
   wire FE_RN_273_0;
   wire FE_RN_272_0;
   wire FE_RN_271_0;
   wire FE_OCPN29562_n25138;
   wire FE_OCPN29561_n23532;
   wire FE_OCPN29559_n17900;
   wire FE_OCPN29557_n18161;
   wire FE_OCPN29556_n383;
   wire FE_OCPN29555_n20593;
   wire FE_OCPN29554_n22507;
   wire FE_OCPN29553_n19602;
   wire FE_OCPN29552_n393;
   wire FE_OCPN29551_n;
   wire FE_RN_270_0;
   wire FE_OCPN29550_n16114;
   wire FE_OCPN29548_n25717;
   wire FE_OCPN29547_n15183;
   wire FE_RN_268_0;
   wire FE_OCPN29546_n;
   wire FE_OCPN29545_n22529;
   wire FE_OCPN29544_n20527;
   wire FE_OCPN29543_FE_OFN28862_n;
   wire FE_OCPN29542_n21151;
   wire FE_OCPN29541_n25870;
   wire FE_RN_267_0;
   wire FE_OCPN29540_FE_OFN25927_n26527;
   wire FE_OCPN29539_n24927;
   wire FE_OCPN29538_n24927;
   wire FE_OCPN29537_FE_OFN28699_w3_6;
   wire FE_OCPN29536_FE_OFN8_w3_14;
   wire FE_OCPN29535_FE_OFN8_w3_14;
   wire FE_OCPN29534_FE_OFN8_w3_14;
   wire FE_OCPN29533_n26971;
   wire FE_OCPN29532_n25697;
   wire FE_OCPN29531_FE_OFN25926_n26922;
   wire FE_OCPN29529_n23125;
   wire FE_OCPN29528_n24138;
   wire FE_OCPN29527_n24138;
   wire FE_OCPN29526_sa31_4;
   wire FE_OCPN29525_n18947;
   wire FE_OCPN29524_n25029;
   wire FE_OCPN29523_n25544;
   wire FE_OCPN29521_n24755;
   wire FE_OCPN29520_n24755;
   wire FE_OCPN29519_n;
   wire FE_OCPN29517_n;
   wire FE_OCPN29515_n27136;
   wire FE_OCPN29514_n27136;
   wire FE_OCPN29513_n17447;
   wire FE_OCPN29512_n16750;
   wire FE_OCPN29511_n22226;
   wire FE_OCPN29510_n16996;
   wire FE_OCPN29509_FE_OFN16184_w3_9;
   wire FE_OCPN29508_FE_OFN16184_w3_9;
   wire FE_OCPN29506_FE_OFN16184_w3_9;
   wire FE_OCPN29505_n22457;
   wire FE_OCPN29504_sa11_4;
   wire FE_OCPN29503_n24627;
   wire FE_OCPN29502_w3_23;
   wire FE_OCPN29501_FE_OFN28662_w3_7;
   wire FE_OCPN29500_FE_OFN28662_w3_7;
   wire FE_OCPN29499_FE_OFN16131_sa12_1;
   wire FE_OCPN29498_n16581;
   wire FE_OCPN29497_sa21_1;
   wire FE_OCPN29496_n24789;
   wire FE_OCPN29494_sa12_4;
   wire FE_OCPN29493_sa12_4;
   wire FE_OCPN29492_sa12_4;
   wire FE_OCPN29491_sa12_4;
   wire FE_OCPN29490_n17001;
   wire FE_OCPN29489_sa23_3;
   wire FE_OCPN29488_FE_OFN25883_n22945;
   wire FE_OCPN29487_FE_OFN28694_sa33_4;
   wire FE_OCPN29486_sa12_3;
   wire FE_OCPN29485_sa12_3;
   wire FE_OCPN29484_sa12_3;
   wire FE_OCPN29483_FE_OFN26014_sa31_3;
   wire FE_OCPN29482_FE_OFN26014_sa31_3;
   wire FE_OCPN29481_n26537;
   wire FE_OCPN29480_n20913;
   wire FE_OCPN29478_n23306;
   wire FE_OCPN29477_sa12_5;
   wire FE_OCPN29476_sa12_5;
   wire FE_OCPN29475_n25054;
   wire FE_OCPN29474_n19119;
   wire FE_OCPN29473_n26579;
   wire FE_OCPN29471_n24175;
   wire FE_OCPN29470_n24175;
   wire FE_OCPN29469_n17747;
   wire FE_OCPN29468_n15919;
   wire FE_OCPN29467_n25102;
   wire FE_OCPN29464_n;
   wire FE_OCPN29463_n;
   wire FE_OCPN29461_n22197;
   wire FE_OCPN29460_n26227;
   wire FE_OCPN29459_n;
   wire FE_OCPN29458_n26442;
   wire FE_OCPN29457_n25722;
   wire FE_OCPN29455_n18671;
   wire FE_OCPN29454_n18671;
   wire FE_OCPN29453_sa12_4;
   wire FE_OCPN29452_n16240;
   wire FE_OCPN29451_n;
   wire FE_OCPN29450_sa21_0;
   wire FE_OCPN29449_n17521;
   wire FE_OCPN29448_n27189;
   wire FE_OCPN29447_n27189;
   wire FE_OCPN29446_n17115;
   wire FE_OCPN29445_n27203;
   wire FE_OCPN29444_n25507;
   wire FE_OCPN29443_n25507;
   wire FE_OCPN29442_n458;
   wire FE_OCPN29441_sa23_4;
   wire FE_OCPN29440_sa23_4;
   wire FE_OCPN29439_n17447;
   wire FE_OCPN29438_sa33_2;
   wire FE_OCPN29437_n25864;
   wire FE_OCPN29436_n22080;
   wire FE_OCPN29435_n17445;
   wire FE_OCPN29434_n408;
   wire FE_OCPN29433_n25040;
   wire FE_OCPN29432_sa30_3;
   wire FE_OCPN29431_sa30_3;
   wire FE_OCPN29430_FE_OFN31_sa20_0;
   wire FE_OCPN29429_FE_OFN16141_sa01_3;
   wire FE_OCPN29428_FE_OFN27131_w3_29;
   wire FE_OCPN29427_w3_15;
   wire FE_OCPN29426_FE_OFN16444_sa13_1;
   wire FE_OCPN29425_n24172;
   wire FE_OCPN29424_FE_OFN26039_sa10_2;
   wire FE_OCPN29423_n26970;
   wire FE_OCPN29422_n23397;
   wire FE_OCPN29421_FE_OFN16128_sa32_2;
   wire FE_OCPN29420_FE_OFN16128_sa32_2;
   wire FE_OCPN29419_FE_OFN16128_sa32_2;
   wire FE_OCPN29418_n;
   wire FE_OCPN29417_n455;
   wire FE_OCPN29416_n22516;
   wire FE_OCPN29415_n17237;
   wire FE_OCPN29414_n;
   wire FE_OCPN29413_sa30_5;
   wire FE_OCPN29412_sa30_5;
   wire FE_OCPN29411_n;
   wire FE_OCPN29409_n22461;
   wire FE_OCPN29408_n22461;
   wire FE_RN_266_0;
   wire FE_OCPN29407_FE_OFN142_sa10_0;
   wire FE_RN_265_0;
   wire FE_RN_264_0;
   wire FE_RN_263_0;
   wire FE_OCPN29406_n18710;
   wire FE_OCPN29405_FE_OFN27148_sa32_3;
   wire FE_OCPN29404_FE_OFN27148_sa32_3;
   wire FE_OCPN29400_sa30_3;
   wire FE_OCPN29399_sa30_3;
   wire FE_OCPN29398_sa30_3;
   wire FE_OCPN29397_n26502;
   wire FE_OCPN29396_n19149;
   wire FE_OCPN29394_n479;
   wire FE_OCPN29393_n483;
   wire FE_OCPN29391_FE_OFN29162_sa33_2;
   wire FE_OCPN29390_n26528;
   wire FE_OCPN29389_n26528;
   wire FE_OCPN29388_n22461;
   wire FE_RN_262_0;
   wire FE_RN_261_0;
   wire FE_RN_260_0;
   wire FE_OCPN29387_n25273;
   wire FE_OCPN29386_n16073;
   wire FE_OCPN29385_n;
   wire FE_OCPN29383_n26674;
   wire FE_OCPN29382_n26674;
   wire FE_OCPN29381_n26796;
   wire FE_OCPN29380_sa20_1;
   wire FE_OCPN29379_sa20_1;
   wire FE_OCPN29378_n23266;
   wire FE_OCPN29376_n24099;
   wire FE_OCPN29374_FE_OFN29191_sa23_2;
   wire FE_OCPN29373_FE_OFN29191_sa23_2;
   wire FE_OCPN29371_n16191;
   wire FE_OCPN29370_FE_OFN28744;
   wire FE_OCPN29369_n16982;
   wire FE_OCPN29368_FE_OFN16247_sa30_1;
   wire FE_RN_259_0;
   wire FE_OCPN29365_n24639;
   wire FE_OCPN29364_n448;
   wire FE_OCPN29363_n14011;
   wire FE_OCPN29361_n25696;
   wire FE_OCPN29359_n26586;
   wire FE_OCPN29358_n17159;
   wire FE_OCPN29356_n27110;
   wire FE_OCPN29355_n492;
   wire FE_OCPN29353_n26586;
   wire FE_OCPN29352_n25173;
   wire FE_OCPN29351_FE_OFN26116_sa13_1;
   wire FE_OCPN29350_w3_25;
   wire CTS_40;
   wire CTS_39;
   wire CTS_38;
   wire CTS_37;
   wire CTS_36;
   wire CTS_35;
   wire CTS_34;
   wire CTS_33;
   wire CTS_32;
   wire CTS_31;
   wire FE_OCPN7662_n26633;
   wire FE_OCPN29349_FE_OCPN27405_sa03_4;
   wire FE_OCPN7660_FE_OFN28720_sa20_1;
   wire FE_OCPN7658_n27056;
   wire FE_OCPN7657_n26213;
   wire FE_OCPN7656_n24301;
   wire FE_OCPN7653_n24270;
   wire FE_OCPN7650_n27110;
   wire FE_OCPN7649_n23259;
   wire FE_OCPN7647_FE_OFN141_sa03_1;
   wire FE_OCPN7645_n20962;
   wire FE_OCPN7644_n21523;
   wire FE_OCPN7643_n17646;
   wire FE_OCPN7642_n26319;
   wire FE_OCPN7641_n25778;
   wire FE_OCPN7640_n18765;
   wire FE_OCPN7638_n26183;
   wire FE_OCPN7637_n25422;
   wire FE_OCPN7636_n25940;
   wire FE_OCPN7633_n26815;
   wire FE_OCPN7631_n24750;
   wire FE_OCPN7629_FE_OFN105_n27178;
   wire FE_OCPN7626_n18582;
   wire FE_OCPN7625_n26501;
   wire FE_OCPN7623_FE_OFN4_w3_22;
   wire FE_OCPN7622_n24526;
   wire FE_OCPN7621_n26898;
   wire FE_OCPN7620_n25761;
   wire FE_OCPN7619_FE_OFN28689_sa03_5;
   wire FE_OCPN7618_n21027;
   wire FE_OCPN7617_n26009;
   wire FE_OCPN7616_FE_OFN16184_w3_9;
   wire FE_OCPN7613_n24166;
   wire FE_OCPN7612_n25229;
   wire FE_OCPN7610_n25861;
   wire FE_OCPN7609_n26145;
   wire FE_OCPN7607_n23539;
   wire FE_OCPN7605_n26234;
   wire FE_OCPN7599_n26721;
   wire FE_OCPN7598_n25174;
   wire FE_OCPN7597_n21981;
   wire FE_OCPN7596_n24647;
   wire FE_OCPN7595_n17426;
   wire FE_OCPN7589_n26420;
   wire FE_OCPN7586_n17693;
   wire FE_OCPN7585_FE_OFN25926_n26922;
   wire FE_OCPN7584_n23447;
   wire FE_OCPN7583_n26983;
   wire FE_OCPN29348_n17592;
   wire FE_RN_258_0;
   wire FE_OCPN29346_n12998;
   wire FE_OCPN29342_n25357;
   wire FE_OCPN29341_FE_OFN29148_n;
   wire FE_OCPN29340_n17079;
   wire FE_OCPN7556_n26504;
   wire FE_OCPN29335_n;
   wire FE_OCPN29334_n17330;
   wire FE_OCPN29333_n17330;
   wire FE_RN_257_0;
   wire FE_OCPN29331_n20933;
   wire FE_OCPN29330_n26459;
   wire FE_OCPN29329_n15517;
   wire FE_RN_256_0;
   wire FE_RN_255_0;
   wire FE_RN_254_0;
   wire FE_RN_253_0;
   wire FE_OCPN29327_n21017;
   wire FE_OCPN29324_n23216;
   wire FE_OCPN29323_n19721;
   wire FE_RN_252_0;
   wire FE_RN_251_0;
   wire FE_RN_250_0;
   wire FE_RN_249_0;
   wire FE_RN_248_0;
   wire FE_RN_247_0;
   wire FE_RN_243_0;
   wire FE_RN_242_0;
   wire FE_OCPN29321_n17876;
   wire FE_OCPN29320_n22461;
   wire FE_OCPN29318_n25524;
   wire FE_OCPN29314_n;
   wire FE_OCPN29309_n26452;
   wire FE_OCPN29308_n;
   wire FE_OCPN29307_FE_OFN25989_sa21_4;
   wire FE_OCPN29305_n23302;
   wire FE_OCPN29304_n17526;
   wire FE_OCPN29302_sa00_4;
   wire FE_OCPN29299_FE_OFN29232_n16875;
   wire FE_OCPN29298_n25028;
   wire FE_OCPN29295_n18739;
   wire FE_OCPN29294_n23925;
   wire FE_OCPN29293_FE_OFN28678_sa21_3;
   wire FE_OCPN29292_n18640;
   wire FE_OCPN29291_n17282;
   wire FE_OCPN29289_n22162;
   wire FE_OCPN29287_n27210;
   wire FE_OCPN29284_n19821;
   wire FE_OCPN29283_n23439;
   wire FE_OCPN29281_sa22_0;
   wire FE_OCPN29279_n25353;
   wire FE_OCPN29277_n26713;
   wire FE_OCPN29274_n26478;
   wire FE_OCPN29269_sa22_1;
   wire FE_OCPN29267_n25935;
   wire FE_OCPN29265_FE_OFN28698_sa21_1;
   wire FE_OCPN29263_n24537;
   wire FE_OCPN29262_n24750;
   wire FE_OCPN29260_sa00_5;
   wire FE_OCPN29258_n27171;
   wire FE_RN_241_0;
   wire FE_RN_240_0;
   wire FE_RN_239_0;
   wire FE_RN_238_0;
   wire FE_OCPN29257_n474;
   wire FE_OCPN29256_n418;
   wire FE_RN_237_0;
   wire FE_RN_236_0;
   wire FE_RN_235_0;
   wire FE_RN_234_0;
   wire FE_OFN29255_n;
   wire FE_OFN29254_n;
   wire FE_OFN29251_n18536;
   wire FE_OFN29250_FE_OCPN27371_sa20_2;
   wire FE_OFN29249_n;
   wire FE_OFN29246_n;
   wire FE_OFN29243_n17065;
   wire FE_OFN29242_n26856;
   wire FE_OFN29241_n22811;
   wire FE_OFN29238_n22811;
   wire FE_OFN29237_n22811;
   wire FE_OFN29235_n;
   wire FE_OFN29234_n16996;
   wire FE_OFN29228_n25218;
   wire FE_OFN29227_n24510;
   wire FE_OFN29226_n16793;
   wire FE_OFN29225_sa12_0;
   wire FE_OFN29224_FE_OCPN28074_n27049;
   wire FE_OFN29223_sa20_0;
   wire FE_OFN29215_n24262;
   wire FE_OFN29211_n23587;
   wire FE_OFN29210_FE_OCPN27261_sa02_0;
   wire FE_OFN29209_FE_OCPN27978_w3_3;
   wire FE_OFN29208_n16436;
   wire FE_OFN29207_n;
   wire FE_OFN29204_sa10_2;
   wire FE_OFN29200_n18521;
   wire FE_OFN29199_FE_OCPN27726_n;
   wire FE_OFN29195_n22850;
   wire FE_OFN29192_n13870;
   wire FE_OFN29191_sa23_2;
   wire FE_OFN29189_sa23_0;
   wire FE_OFN29187_FE_OCPN27571_n20235;
   wire FE_OFN29184_n17744;
   wire FE_OFN29182_n21708;
   wire FE_OFN29181_n24479;
   wire FE_OFN29180_n26222;
   wire FE_OFN29179_n;
   wire FE_OFN29178_sa20_4;
   wire FE_OFN29177_sa20_4;
   wire FE_OFN29175_n21755;
   wire FE_OFN29173_n;
   wire FE_OFN29172_sa00_4;
   wire FE_OFN29171_n17510;
   wire FE_OFN29170_n17510;
   wire FE_OFN29169_n17510;
   wire FE_OFN29164_sa33_2;
   wire FE_OFN29163_sa33_2;
   wire FE_OFN29162_sa33_2;
   wire FE_OFN29161_n;
   wire FE_OFN29160_n25363;
   wire FE_OFN29159_n21892;
   wire FE_OFN29158_n18860;
   wire FE_OFN29154_n19753;
   wire FE_OFN29153_n19753;
   wire FE_OFN29152_sa22_0;
   wire FE_OFN29151_n22988;
   wire FE_OFN29150_sa20_5;
   wire FE_OFN29148_n;
   wire FE_OFN29147_sa31_1;
   wire FE_OFN29145_sa31_1;
   wire FE_OFN29144_n17747;
   wire FE_OFN29143_n25444;
   wire FE_OFN29142_n27049;
   wire FE_OFN29141_n26574;
   wire FE_OFN29140_n18527;
   wire FE_OFN29139_n18527;
   wire FE_OFN29137_FE_OCPN27228_sa11_2;
   wire FE_OFN29136_n;
   wire FE_OFN29135_n21551;
   wire FE_OFN29134_sa33_0;
   wire FE_OFN29131_FE_OCPN27371_sa20_2;
   wire FE_OFN29125_n;
   wire FE_OFN29124_n;
   wire FE_OFN29123_n;
   wire FE_OFN29122_n;
   wire FE_OFN29121_n26026;
   wire FE_OFN29117_n;
   wire FE_OFN29112_FE_OCPN27870_n18527;
   wire FE_OFN29109_n;
   wire FE_OFN29102_FE_OCPN27261_sa02_0;
   wire FE_OFN29101_n16418;
   wire FE_OFN29096_n25188;
   wire FE_OFN29094_n21607;
   wire FE_OFN29091_n;
   wire FE_OFN29087_n;
   wire FE_OFN29081_n18526;
   wire FE_OFN29080_n22310;
   wire FE_OFN29079_FE_OCPN27518_n17251;
   wire FE_OFN29076_n18540;
   wire FE_OFN29075_n22745;
   wire FE_OFN29074_n17170;
   wire FE_OFN29067_n;
   wire FE_OFN29066_FE_OCPN27328_sa21_2;
   wire FE_OFN29063_n25433;
   wire FE_OFN29062_n18651;
   wire FE_OFN29061_n22505;
   wire FE_OFN29054_n17453;
   wire FE_OFN29052_w3_5;
   wire FE_OFN29051_n25465;
   wire FE_OFN29049_n17756;
   wire FE_OFN29048_n17756;
   wire FE_OFN29047_n21980;
   wire FE_OFN29044_n19967;
   wire FE_OFN29043_n;
   wire FE_OFN29042_n;
   wire FE_OFN29041_n21415;
   wire FE_OFN29040_n17404;
   wire FE_OFN29039_n26763;
   wire FE_OFN29037_n;
   wire FE_OFN29036_n20806;
   wire FE_OFN29035_n17116;
   wire FE_OFN29034_FE_OCPN27414_n23359;
   wire FE_OFN29033_FE_OCPN27414_n23359;
   wire FE_OFN29032_FE_OCPN27728_n21981;
   wire FE_OFN29031_n23968;
   wire FE_OFN29029_n26579;
   wire FE_OFN29027_n19135;
   wire FE_OFN29026_n20911;
   wire FE_OFN29024_n;
   wire FE_OFN29023_n16750;
   wire FE_OFN29021_sa20_3;
   wire FE_OFN29020_n25146;
   wire FE_OFN29018_n15921;
   wire FE_OFN29017_n15921;
   wire FE_OFN29016_n16512;
   wire FE_OFN29015_n25040;
   wire FE_OFN29011_n27113;
   wire FE_OFN29010_n27113;
   wire FE_OFN29005_n23558;
   wire FE_OFN29003_n23491;
   wire FE_OFN29001_n23491;
   wire FE_OFN29000_n18698;
   wire FE_OFN28999_n16923;
   wire FE_OFN28998_n16923;
   wire FE_OFN28997_sa03_4;
   wire FE_OFN28996_n17464;
   wire FE_OFN28995_n16850;
   wire FE_OFN28994_FE_OCPN5176_n25870;
   wire FE_OFN28991_n19938;
   wire FE_OFN28990_n26276;
   wire FE_OFN28988_n18597;
   wire FE_OFN28987_n18597;
   wire FE_OFN28986_n18597;
   wire FE_OFN28985_sa21_5;
   wire FE_OFN28984_n20851;
   wire FE_OFN28981_n16767;
   wire FE_OFN28980_n18169;
   wire FE_OFN28979_n;
   wire FE_OFN28977_n;
   wire FE_OFN28976_n;
   wire FE_OFN28973_n25273;
   wire FE_OFN28972_n27021;
   wire FE_OFN28971_n23947;
   wire FE_OFN28970_n19890;
   wire FE_OFN28969_n19890;
   wire FE_OFN28968_n26780;
   wire FE_OFN28966_n23329;
   wire FE_OFN28965_n24869;
   wire FE_OFN28964_n16273;
   wire FE_OFN28963_n24480;
   wire FE_OFN28962_n17744;
   wire FE_OFN28961_n17744;
   wire FE_OFN28960_n25379;
   wire FE_OFN28958_n17261;
   wire FE_OFN28956_n18011;
   wire FE_OFN28955_n18011;
   wire FE_OFN28954_n18011;
   wire FE_OFN28953_n18011;
   wire FE_OFN28952_n18011;
   wire FE_OFN28951_n18011;
   wire FE_OFN28950_n18011;
   wire FE_OFN28949_n18011;
   wire FE_OFN28948_n18011;
   wire FE_OFN28947_sa12_5;
   wire FE_OFN28946_n23135;
   wire FE_OFN28942_n21456;
   wire FE_OFN28941_sa02_2;
   wire FE_OFN28939_n21129;
   wire FE_OFN28936_n18104;
   wire FE_OFN28935_n18104;
   wire FE_OFN28934_n24552;
   wire FE_OFN28933_n16321;
   wire FE_OFN28931_n17897;
   wire FE_OFN28930_n22836;
   wire FE_OFN28929_n15182;
   wire FE_OFN28928_n22374;
   wire FE_OFN28927_n22374;
   wire FE_OFN28925_sa30_0;
   wire FE_OFN28924_n25912;
   wire FE_OFN28923_n21873;
   wire FE_OFN28922_n24249;
   wire FE_OFN28921_n20660;
   wire FE_OFN28920_n24254;
   wire FE_OFN28919_n24155;
   wire FE_OFN28918_n16949;
   wire FE_OFN28916_sa10_4;
   wire FE_OFN28915_FE_OCPN27241_sa11_1;
   wire FE_OFN28914_n20007;
   wire FE_OFN28913_n18247;
   wire FE_OFN28912_n16534;
   wire FE_OFN28911_n16534;
   wire FE_OFN28910_n16534;
   wire FE_OFN28909_w3_23;
   wire FE_OFN28908_w3_23;
   wire FE_OFN28907_n26049;
   wire FE_OFN28904_n25733;
   wire FE_OFN28903_sa21_0;
   wire FE_OFN28902_n25414;
   wire FE_OFN28901_sa30_4;
   wire FE_OFN28898_n13805;
   wire FE_OFN28897_n20132;
   wire FE_OFN28896_sa30_2;
   wire FE_OFN28895_sa30_2;
   wire FE_OFN28894_n;
   wire FE_OFN28893_n;
   wire FE_OFN28892_n;
   wire FE_OFN28891_n;
   wire FE_OFN28890_n;
   wire FE_OFN28889_n15845;
   wire FE_OFN28886_FE_OCPN27675_n17986;
   wire FE_OFN28884_n;
   wire FE_OFN28883_n;
   wire FE_OFN28882_FE_OCPN27356_sa12_0;
   wire FE_OFN28877_FE_OCPN27730_n17464;
   wire FE_OFN28874_FE_OCPN27551_sa11_4;
   wire FE_OFN28869_FE_OCPN27715_n23875;
   wire FE_OFN28868_FE_OCPN27715_n23875;
   wire FE_OFN28862_n;
   wire FE_OFN28859_FE_OCPN27664_w3_25;
   wire FE_OFN28858_FE_OCPN27664_w3_25;
   wire FE_OFN28856_n15450;
   wire FE_OFN28853_FE_OCPN28408;
   wire FE_OFN28850_FE_OCPN27840;
   wire FE_OFN28848_n14912;
   wire FE_OFN28846_n26367;
   wire FE_OFN28844_FE_OCPN27570_n17791;
   wire FE_OFN28841_n22980;
   wire FE_OFN28840_n;
   wire FE_OFN28836_FE_OCPN27631_n16774;
   wire FE_OFN28835_n;
   wire FE_OFN28834_FE_OCPN28371_n17900;
   wire FE_OFN28832_n19789;
   wire FE_OFN28831_n15838;
   wire FE_OFN28829_n;
   wire FE_OFN28827_n15683;
   wire FE_OFN28823_n17860;
   wire FE_OFN28820_n;
   wire FE_OFN28818_n17602;
   wire FE_OFN28817_n;
   wire FE_OFN28815_n18523;
   wire FE_OFN28813_n15414;
   wire FE_OFN28812_FE_OCPN27261_sa02_0;
   wire FE_OFN28811_n19170;
   wire FE_OFN28809_n;
   wire FE_OFN28808_n26291;
   wire FE_OFN28807_n24944;
   wire FE_OFN28806_n24944;
   wire FE_OFN28801_n16978;
   wire FE_OFN28800_n22526;
   wire FE_OFN28798_FE_OCPN27947_n18177;
   wire FE_OFN28796_n17301;
   wire FE_OFN28792_n15787;
   wire FE_OFN28791_n;
   wire FE_OFN28790_n;
   wire FE_OFN28787_n19000;
   wire FE_OFN28783_n26099;
   wire FE_OFN28779_n24257;
   wire FE_OFN28778_FE_OCPN28352_n16748;
   wire FE_OFN28776_n18532;
   wire FE_OFN28775_n16992;
   wire FE_OFN28771_n;
   wire FE_OFN28769_n15478;
   wire FE_OFN28767_n26103;
   wire FE_OFN28764_n17928;
   wire FE_OFN28758_n15422;
   wire FE_OFN28753_sa31_2;
   wire FE_OFN28752_n;
   wire FE_OFN28751_n;
   wire FE_OFN28749_n;
   wire FE_OFN28747_n;
   wire FE_OFN28744_FE_OCPN27908;
   wire FE_OFN28741_n;
   wire FE_OFN28739_n17898;
   wire FE_OFN28738_n16989;
   wire FE_OFN28736_FE_OCPN28216_sa01_5;
   wire FE_OFN28734_n;
   wire FE_OFN28732_n;
   wire FE_OFN28730_FE_OCPN28416_sa02_3;
   wire FE_OFN28729_n20617;
   wire FE_OFN28727_sa33_1;
   wire FE_OFN28725_n16982;
   wire FE_OFN28723_n22750;
   wire FE_OFN28722_sa10_3;
   wire FE_OFN28721_n;
   wire FE_OFN28720_sa20_1;
   wire FE_OFN28719_n20025;
   wire FE_OFN28718_sa01_1;
   wire FE_OFN28717_n15158;
   wire FE_OFN28715_w3_15;
   wire FE_OFN28713_n;
   wire FE_OFN28712_n;
   wire FE_OFN28711_n;
   wire FE_OFN28710_n20841;
   wire FE_OFN28707_n;
   wire FE_OFN28706_n;
   wire FE_OFN28704_FE_OCPN27740_sa02_4;
   wire FE_OFN28703_FE_OCPN27740_sa02_4;
   wire FE_OFN28701_w3_16;
   wire FE_OFN28699_w3_6;
   wire FE_OFN28698_sa21_1;
   wire FE_OFN28696_sa32_4;
   wire FE_OFN28695_n;
   wire FE_OFN28694_sa33_4;
   wire FE_OFN28691_n13725;
   wire FE_OFN28690_n25979;
   wire FE_OFN28689_sa03_5;
   wire FE_OFN28688_sa22_2;
   wire FE_OFN28686_FE_OCPN27812;
   wire FE_OFN28683_w3_21;
   wire FE_OFN28682_n15888;
   wire FE_OFN28680_n;
   wire FE_OFN28679_sa33_5;
   wire FE_OFN28678_sa21_3;
   wire FE_OFN28677_n17998;
   wire FE_OFN28676_sa12_5;
   wire FE_OFN28674_n;
   wire FE_OFN28673_n;
   wire FE_OFN28672_sa01_2;
   wire FE_OFN28671_FE_OCPN28076;
   wire FE_OFN28669_sa31_5;
   wire FE_OFN28665_FE_OCPN27566;
   wire FE_OFN28663_n;
   wire FE_OFN28662_w3_7;
   wire FE_OFN28661_w3_7;
   wire FE_OFN28660_w3_7;
   wire FE_OFN28659_n15934;
   wire FE_OFN28658_n15934;
   wire FE_OFN28656_FE_OFN25986_n21012;
   wire FE_OFN28655_FE_OFN25986_n21012;
   wire FE_OFN28654_n22751;
   wire FE_OFN28652_n21642;
   wire FE_OFN28651_FE_OFN26140_n23585;
   wire FE_OFN28650_n23802;
   wire FE_OFN28649_n23802;
   wire FE_OFN28648_n23549;
   wire FE_OFN28647_n21764;
   wire FE_OFN28643_sa33_0;
   wire FE_OFN28637_n25102;
   wire FE_OFN28635_n21034;
   wire FE_OFN28633_n17716;
   wire FE_OFN28630_n23385;
   wire FE_OFN28628_n15667;
   wire FE_OFN28627_n21377;
   wire FE_OFN28626_n22094;
   wire FE_OFN28625_n26101;
   wire FE_OFN28624_n13874;
   wire FE_OFN28623_n13874;
   wire FE_OFN28622_n25870;
   wire FE_OFN28619_n20437;
   wire FE_OFN28618_n25322;
   wire FE_OFN28616_n26191;
   wire FE_OFN28615_n26191;
   wire FE_OFN28614_n21715;
   wire FE_OFN28610_n22125;
   wire FE_OFN28609_n19730;
   wire FE_OFN28608_n21027;
   wire FE_OFN28607_n23884;
   wire FE_OFN28605_n23949;
   wire FE_OFN28604_n14534;
   wire FE_OFN28603_n14534;
   wire FE_OFN28602_n14534;
   wire FE_OFN28600_n14289;
   wire FE_OFN28598_n20933;
   wire FE_OFN28596_n23948;
   wire FE_OFN28595_n20189;
   wire FE_OFN28594_n26454;
   wire FE_OFN28593_n18627;
   wire FE_OFN28592_n16427;
   wire FE_OFN28590_n24391;
   wire FE_OFN28589_n21048;
   wire FE_OFN28588_n21048;
   wire FE_OFN28586_n24736;
   wire FE_OFN28584_n17001;
   wire FE_OFN28583_n17001;
   wire FE_OFN28582_n25657;
   wire FE_OFN28581_n23491;
   wire FE_OFN28580_n23491;
   wire FE_OFN28579_n23491;
   wire FE_OFN28578_FE_OFN16316_n24840;
   wire FE_OFN28576_n27003;
   wire FE_OFN28574_n16016;
   wire FE_OFN28573_n26748;
   wire FE_OFN28572_n21723;
   wire FE_OFN28571_w3_28;
   wire FE_OFN28570_n19172;
   wire FE_OFN28569_n18755;
   wire FE_OFN28567_n19514;
   wire FE_OFN28566_n21491;
   wire FE_OFN28565_n26845;
   wire FE_OFN28564_n18308;
   wire FE_OFN28563_n20480;
   wire FE_OFN28562_n19342;
   wire FE_OFN28561_n25419;
   wire FE_OFN28560_n22749;
   wire FE_OFN28559_n18278;
   wire FE_OFN28558_n23073;
   wire FE_OFN28557_n25031;
   wire FE_OFN28556_n24516;
   wire FE_OFN28554_n21876;
   wire FE_OFN28553_n25599;
   wire FE_OFN28552_n20105;
   wire FE_OFN28551_FE_OFN26114_n;
   wire FE_OFN28549_n21934;
   wire FE_OFN28548_n27092;
   wire FE_OFN28546_n26091;
   wire FE_OFN28544_n13805;
   wire FE_OFN28543_FE_OFN109_n15994;
   wire FE_OFN28542_n15433;
   wire FE_OFN28541_n16476;
   wire FE_OFN28540_n21599;
   wire FE_OFN28539_n22336;
   wire FE_OFN28538_n16166;
   wire FE_OFN28537_sa20_2;
   wire FE_OFN28536_sa20_2;
   wire FE_OFN28535_n19738;
   wire FE_OFN28534_n21462;
   wire FE_OFN28533_n24995;
   wire FE_OFN28531_FE_OFN56_n14826;
   wire FE_OFN28530_n14593;
   wire FE_OFN28529_n16774;
   wire FE_OFN28528_n25241;
   wire FE_OFN28525_n25751;
   wire FE_OFN28523_sa03_1;
   wire FE_OFN28522_n17261;
   wire FE_OFN28521_n26007;
   wire FE_OFN28520_n22753;
   wire FE_OFN28516_FE_OFN27192_sa31_2;
   wire FE_OFN28515_n22062;
   wire FE_OFN28514_sa00_1;
   wire FE_OFN28513_n20470;
   wire FE_OFN28512_n27020;
   wire FE_OFN28511_n25088;
   wire FE_OFN28510_n21215;
   wire FE_OFN28508_sa11_0;
   wire FE_OFN28507_sa11_0;
   wire FE_OFN28506_n26996;
   wire FE_OFN28505_n23296;
   wire FE_OFN28504_n25956;
   wire FE_OFN28503_n26596;
   wire FE_OFN28502_n25865;
   wire FE_OFN28501_FE_OFN26020_n14010;
   wire FE_OFN28500_FE_OCPN5078_n25823;
   wire FE_OFN28499_sa00_6;
   wire FE_OFN28496_n15201;
   wire FE_OFN28495_n24584;
   wire FE_OFN28492_sa31_0;
   wire FE_OFN28491_sa13_3;
   wire FE_OFN28490_ld_r;
   wire FE_OFN28489_ld_r;
   wire FE_OFN28487_ld_r;
   wire FE_OFN28486_ld_r;
   wire FE_OFN28485_ld_r;
   wire FE_OFN28484_ld_r;
   wire FE_OFN28483_ld_r;
   wire FE_OFN28482_ld_r;
   wire FE_OFN28481_n15298;
   wire FE_OFN28480_sa30_7;
   wire FE_OFN28479_sa13_2;
   wire FE_OFN28478_sa13_2;
   wire FE_OFN28477_n23853;
   wire FE_OFN28476_sa12_0;
   wire FE_OFN28475_n23573;
   wire FE_OFN28474_FE_OCPN5038_n26735;
   wire FE_OFN28473_n26911;
   wire FE_OFN28472_ld;
   wire FE_OFN28471_ld;
   wire FE_OFN28470_ld;
   wire FE_OFN28469_ld;
   wire FE_OFN28468_ld;
   wire FE_OFN28467_ld;
   wire FE_OFN28466_ld;
   wire FE_OFN28465_ld;
   wire FE_OFN28464_ld;
   wire FE_OFN28463_ld;
   wire FE_OFN28462_ld;
   wire FE_OFN28461_ld;
   wire FE_OFN28460_ld;
   wire FE_OFN28459_ld;
   wire FE_OFN28458_ld;
   wire FE_OFN28457_ld;
   wire FE_OFN28456_n13348;
   wire FE_OFN28455_n13348;
   wire FE_OFN28454_n13348;
   wire FE_OFN28453_n13348;
   wire FE_OFN28452_w3_29;
   wire FE_OFN28451_n26990;
   wire FE_RN_233_0;
   wire FE_RN_232_0;
   wire FE_RN_231_0;
   wire FE_RN_230_0;
   wire FE_OCPN5199_n21457;
   wire FE_OCPN5198_n25566;
   wire FE_OCPN5195_FE_OFN25874_sa03_2;
   wire FE_OCPN5191_n20272;
   wire FE_OCPN5188_n22414;
   wire FE_OCPN5182_n21090;
   wire FE_OCPN5178_n25039;
   wire FE_OCPN5172_n26281;
   wire FE_OCPN5167_n22336;
   wire FE_OCPN5166_n27203;
   wire FE_OCPN5158_n24742;
   wire FE_OCPN5156_n23958;
   wire FE_OCPN5153_n23127;
   wire FE_OCPN5147_n18548;
   wire FE_OCPN5146_n26207;
   wire FE_OCPN5143_n19361;
   wire FE_OCPN5140_n21049;
   wire FE_OCPN5139_n24167;
   wire FE_OCPN5137_n23600;
   wire FE_OCPN5133_n26620;
   wire FE_OCPN5132_n23890;
   wire FE_OCPN5131_n25916;
   wire FE_OCPN5129_sa32_3;
   wire FE_OCPN5126_sa21_2;
   wire FE_OCPN5119_n25762;
   wire FE_OCPN5116_n25443;
   wire FE_OCPN5115_n25574;
   wire FE_OCPN5112_n25135;
   wire FE_OCPN5110_n23721;
   wire FE_OCPN5109_n26551;
   wire FE_OCPN5107_n24418;
   wire FE_OCPN5106_n25999;
   wire FE_OCPN5105_n25099;
   wire FE_OCPN5099_n24677;
   wire FE_OCPN5088_n27079;
   wire FE_OCPN5086_n26050;
   wire FE_OCPN5083_sa21_2;
   wire FE_OCPN5082_n22663;
   wire FE_OCPN5080_n25758;
   wire FE_OCPN5079_n20287;
   wire FE_OCPN5077_n25855;
   wire FE_OCPN5076_n24192;
   wire FE_OCPN5073_n24996;
   wire FE_OCPN5072_n23451;
   wire FE_OCPN5068_n25984;
   wire FE_OCPN5062_n20505;
   wire FE_OCPN5056_n26535;
   wire FE_OCPN5053_n25832;
   wire FE_OCPN5051_n25883;
   wire FE_OCPN5045_n26098;
   wire FE_OCPN5043_n26230;
   wire FE_OCPN5041_n26726;
   wire FE_OCPN5038_n26735;
   wire FE_OCPN5022_n26716;
   wire FE_OCPN5021_n17446;
   wire FE_OCPN5020_n27079;
   wire FE_OCPN5015_n23031;
   wire FE_RN_229_0;
   wire FE_RN_228_0;
   wire FE_RN_227_0;
   wire FE_RN_226_0;
   wire FE_RN_224_0;
   wire FE_OCPN28447_n23392;
   wire FE_RN_223_0;
   wire FE_OCPN28444_n428;
   wire FE_OCPN28442_n27056;
   wire FE_OCPN28438_n27080;
   wire FE_OCPN28437_n23932;
   wire FE_RN_222_0;
   wire FE_OCPN28434_n17546;
   wire FE_OCPN28432_n23829;
   wire FE_OCPN28431_n21734;
   wire FE_OCPN28427_n25064;
   wire FE_OCPN28425_n18597;
   wire FE_OCPN28423_n18836;
   wire FE_RN_220_0;
   wire FE_OCPN28418_n19586;
   wire FE_OCPN28417_n21396;
   wire FE_OCPN28408_FE_OFN16433_w3_11;
   wire FE_OCPN28407_FE_OFN16433_w3_11;
   wire FE_OCPN28404_n13874;
   wire FE_RN_219_0;
   wire FE_OCPN28402_w3_13;
   wire FE_OCPN28398_n15808;
   wire FE_OCPN4698_n25497;
   wire FE_OCPN4686_n19142;
   wire FE_OCPN4685_n15658;
   wire FE_OCPN4680_n21317;
   wire FE_OCPN28397_n23082;
   wire FE_OCPN28394_FE_OFN27043_n;
   wire FE_OCPN28392_n22380;
   wire FE_OCPN28389_n21479;
   wire FE_OCPN28386_n17899;
   wire FE_OCPN28383_n24808;
   wire FE_OCPN28381_n26660;
   wire FE_OCPN28380_n22433;
   wire FE_OCPN28378_n22632;
   wire FE_RN_218_0;
   wire FE_OCPN28366_n25329;
   wire FE_OCPN28365_n21549;
   wire FE_OCPN28363_n22979;
   wire FE_OCPN28358_n21899;
   wire FE_OCPN28357_n22882;
   wire FE_OCPN28355_n26909;
   wire FE_OCPN28354_n16677;
   wire FE_OCPN28353_n18534;
   wire FE_RN_217_0;
   wire FE_OCPN28346_n24051;
   wire FE_OCPN28334_n16497;
   wire FE_OCPN28328_n25953;
   wire FE_OCPN28327_n15899;
   wire FE_RN_216_0;
   wire FE_OCPN28323_FE_OFN16427_sa10_3;
   wire FE_OCPN28322_n18141;
   wire FE_OCPN28321_n21341;
   wire FE_OCPN28320_n25954;
   wire FE_OCPN28316_n26980;
   wire FE_OCPN28314_n20842;
   wire FE_OCPN28312_n20842;
   wire FE_OCPN28311_n26789;
   wire FE_OCPN28310_n22585;
   wire FE_OCPN28309_n22779;
   wire FE_OCPN28307_n26491;
   wire FE_OCPN28305_n26451;
   wire FE_OCPN28303_n20961;
   wire FE_RN_215_0;
   wire FE_RN_214_0;
   wire FE_RN_213_0;
   wire FE_RN_212_0;
   wire FE_RN_211_0;
   wire FE_RN_210_0;
   wire FE_RN_209_0;
   wire FE_RN_208_0;
   wire FE_RN_207_0;
   wire FE_RN_206_0;
   wire FE_RN_205_0;
   wire FE_RN_204_0;
   wire FE_OCPN28301_n22448;
   wire FE_RN_203_0;
   wire FE_RN_202_0;
   wire FE_RN_201_0;
   wire FE_RN_200_0;
   wire FE_RN_198_0;
   wire FE_RN_197_0;
   wire FE_RN_196_0;
   wire FE_RN_195_0;
   wire FE_RN_194_0;
   wire FE_RN_193_0;
   wire FE_RN_192_0;
   wire FE_RN_191_0;
   wire FE_RN_190_0;
   wire FE_RN_188_0;
   wire FE_RN_187_0;
   wire FE_RN_186_0;
   wire FE_RN_185_0;
   wire FE_RN_184_0;
   wire FE_RN_183_0;
   wire FE_RN_182_0;
   wire FE_RN_181_0;
   wire FE_RN_180_0;
   wire FE_RN_179_0;
   wire FE_OCPN28299_n;
   wire FE_OCPN28298_n;
   wire FE_OCPN28297_n23417;
   wire FE_RN_178_0;
   wire FE_RN_177_0;
   wire FE_RN_175_0;
   wire FE_RN_174_0;
   wire FE_RN_173_0;
   wire FE_RN_171_0;
   wire FE_RN_170_0;
   wire FE_RN_169_0;
   wire FE_RN_168_0;
   wire FE_RN_166_0;
   wire FE_RN_165_0;
   wire FE_RN_164_0;
   wire FE_RN_163_0;
   wire FE_RN_162_0;
   wire FE_RN_161_0;
   wire FE_RN_160_0;
   wire FE_RN_159_0;
   wire FE_OCPN28296_n15386;
   wire FE_RN_158_0;
   wire FE_RN_157_0;
   wire FE_RN_156_0;
   wire FE_RN_155_0;
   wire FE_RN_154_0;
   wire FE_RN_153_0;
   wire FE_RN_152_0;
   wire FE_RN_151_0;
   wire FE_RN_150_0;
   wire FE_RN_149_0;
   wire FE_RN_148_0;
   wire FE_RN_147_0;
   wire FE_RN_146_0;
   wire FE_RN_145_0;
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_142_0;
   wire FE_OCPN28289_n20235;
   wire FE_OCPN28279_n;
   wire FE_OCPN28278_n15512;
   wire FE_RN_141_0;
   wire FE_RN_140_0;
   wire FE_RN_139_0;
   wire FE_RN_138_0;
   wire FE_RN_137_0;
   wire FE_RN_136_0;
   wire FE_RN_135_0;
   wire FE_RN_134_0;
   wire FE_RN_133_0;
   wire FE_RN_132_0;
   wire FE_RN_131_0;
   wire FE_RN_130_0;
   wire FE_RN_129_0;
   wire FE_RN_128_0;
   wire FE_RN_127_0;
   wire FE_RN_126_0;
   wire FE_RN_125_0;
   wire FE_OCPN28270_n17237;
   wire FE_RN_124_0;
   wire FE_OCPN28268_n19911;
   wire FE_OCPN28266_n20920;
   wire FE_RN_123_0;
   wire FE_RN_122_0;
   wire FE_OCPN28257_n23689;
   wire FE_RN_121_0;
   wire FE_OCPN28250_n19573;
   wire FE_OCPN28248_n17971;
   wire FE_OCPN28246_n;
   wire FE_OCPN28245_n;
   wire FE_OCPN28241_n22142;
   wire FE_RN_120_0;
   wire FE_RN_119_0;
   wire FE_OCPN28235_n26631;
   wire FE_OCPN28232_n17949;
   wire FE_RN_118_0;
   wire FE_OCPN28230_n23644;
   wire FE_OCPN28229_n17529;
   wire FE_OCPN28223_FE_OFN27219_n18522;
   wire FE_RN_117_0;
   wire FE_OCPN28217_sa01_5;
   wire FE_OCPN28214_n21500;
   wire FE_OCPN28212_n16980;
   wire FE_OCPN28204_n20526;
   wire FE_OCPN28202_n16991;
   wire FE_RN_116_0;
   wire FE_RN_115_0;
   wire FE_RN_114_0;
   wire FE_RN_113_0;
   wire FE_RN_112_0;
   wire FE_RN_111_0;
   wire FE_RN_110_0;
   wire FE_RN_109_0;
   wire FE_RN_108_0;
   wire FE_OCPN28198_n22776;
   wire FE_OCPN28196_n22547;
   wire FE_OCPN28189_n20491;
   wire FE_OCPN28187_n16806;
   wire FE_OCPN28186_n16123;
   wire FE_OCPN28184_n18020;
   wire FE_OCPN28179_n16535;
   wire FE_OCPN28175_n21818;
   wire FE_OCPN28173_n27153;
   wire FE_OCPN28172_n20449;
   wire FE_RN_107_0;
   wire FE_OCPN28169_n25121;
   wire FE_OCPN28167_n21472;
   wire FE_OCPN28163_FE_OFN99_sa20_5;
   wire FE_OCPN28158_n;
   wire FE_OCPN28157_n16534;
   wire FE_OCPN28156_n26304;
   wire FE_OCPN28150_n27152;
   wire FE_OCPN28149_n17121;
   wire FE_OCPN28145_n16535;
   wire FE_OCPN28141_n;
   wire FE_OCPN28140_FE_OFN133_n24306;
   wire FE_OCPN28138_n26654;
   wire FE_OCPN28137_n17170;
   wire FE_OCPN28135_sa12_3;
   wire FE_RN_106_0;
   wire FE_RN_105_0;
   wire FE_RN_104_0;
   wire FE_RN_103_0;
   wire FE_RN_102_0;
   wire FE_RN_101_0;
   wire FE_RN_100_0;
   wire FE_RN_99_0;
   wire FE_RN_98_0;
   wire FE_RN_97_0;
   wire FE_RN_96_0;
   wire FE_RN_95_0;
   wire FE_RN_94_0;
   wire FE_RN_93_0;
   wire FE_RN_92_0;
   wire FE_RN_91_0;
   wire FE_RN_90_0;
   wire FE_RN_89_0;
   wire FE_RN_88_0;
   wire FE_RN_87_0;
   wire FE_RN_86_0;
   wire FE_RN_85_0;
   wire FE_RN_84_0;
   wire FE_RN_83_0;
   wire FE_RN_82_0;
   wire FE_RN_81_0;
   wire FE_RN_80_0;
   wire FE_RN_79_0;
   wire FE_RN_78_0;
   wire FE_RN_77_0;
   wire FE_OCPN28131_n26796;
   wire FE_OCPN28127_n16872;
   wire FE_OCPN28123_n27047;
   wire FE_OCPN28122_n27157;
   wire FE_RN_76_0;
   wire FE_OCPN28121_n16975;
   wire FE_OCPN28120_n16975;
   wire FE_OCPN28119_n26955;
   wire FE_RN_74_0;
   wire FE_RN_73_0;
   wire FE_RN_71_0;
   wire FE_RN_69_0;
   wire FE_RN_68_0;
   wire FE_RN_67_0;
   wire FE_RN_66_0;
   wire FE_OCPN28115_n25293;
   wire FE_RN_65_0;
   wire FE_RN_64_0;
   wire FE_RN_63_0;
   wire FE_OCPN28112_n26664;
   wire FE_OCPN28111_n19091;
   wire FE_OCPN28110_n;
   wire FE_OCPN28107_n23504;
   wire FE_OCPN28106_FE_OFN25876_n25462;
   wire FE_OCPN28100_n25470;
   wire FE_OCPN28098_n20907;
   wire FE_OCPN28096_w3_31;
   wire FE_OCPN28093_FE_OFN26534_w3_19;
   wire FE_OCPN28089_n23913;
   wire FE_OCPN28086_n22034;
   wire FE_OCPN28083_n26574;
   wire FE_OCPN28082_n21860;
   wire FE_OCPN28078_n24296;
   wire FE_OCPN28077_n;
   wire FE_OCPN28076_FE_OFN9_w3_6;
   wire FE_OCPN28075_n16048;
   wire FE_OCPN28073_n27049;
   wire FE_OCPN28072_w3_3;
   wire FE_OCPN28071_n25092;
   wire FE_RN_62_0;
   wire FE_RN_61_0;
   wire FE_RN_60_0;
   wire FE_OCPN28065_n15774;
   wire FE_RN_58_0;
   wire FE_OCPN28061_n20076;
   wire FE_OCPN28057_n17603;
   wire FE_OCPN28054_n26501;
   wire FE_OCPN28053_sa10_1;
   wire FE_OCPN28052_sa10_1;
   wire FE_OCPN28049_sa30_0;
   wire FE_OCPN28040_n19766;
   wire FE_OCPN28038_n23252;
   wire FE_OCPN28037_n22855;
   wire FE_OCPN28027_n22125;
   wire FE_OCPN28024_n26427;
   wire FE_OCPN28023_n25770;
   wire FE_OCPN28021_n21445;
   wire FE_OCPN28017_n18548;
   wire FE_OCPN28016_n21124;
   wire FE_OCPN28008_n16290;
   wire FE_OCPN28006_n17454;
   wire FE_RN_54_0;
   wire FE_OCPN28001_n21310;
   wire FE_OCPN28000_n22450;
   wire FE_OCPN27998_n18019;
   wire FE_OCPN27991_n26336;
   wire FE_OCPN27990_FE_OFN16132_sa03_5;
   wire FE_OCPN27988_n26454;
   wire FE_OCPN27987_FE_OFN4_w3_22;
   wire FE_OCPN27986_n18970;
   wire FE_OCPN27985_n24831;
   wire FE_RN_53_0;
   wire FE_OCPN27979_FE_OFN16147_sa22_1;
   wire FE_OCPN27978_w3_3;
   wire FE_OCPN27975_n18871;
   wire FE_OCPN27972_n20988;
   wire FE_OCPN27971_n21627;
   wire FE_OCPN27968_n21154;
   wire FE_OCPN27966_n18473;
   wire FE_OCPN27956_n;
   wire FE_OCPN27955_n22945;
   wire FE_OCPN27954_n22945;
   wire FE_OCPN27953_n22945;
   wire FE_OCPN27951_n19098;
   wire FE_OCPN27948_FE_OFN26173_n21511;
   wire FE_OCPN27947_n18177;
   wire FE_RN_52_0;
   wire FE_OCPN27941_n;
   wire FE_OCPN27940_n26842;
   wire FE_OCPN27937_n18841;
   wire FE_OCPN27935_n26773;
   wire FE_OCPN27933_n23328;
   wire FE_OCPN27929_FE_OFN4_w3_22;
   wire FE_OCPN27928_FE_OFN4_w3_22;
   wire FE_OCPN27922_n26712;
   wire FE_OCPN27919_n20155;
   wire FE_OCPN27918_n21042;
   wire FE_OCPN27916_n;
   wire FE_OCPN27908_FE_OFN16156_sa00_2;
   wire FE_OCPN27906_n23131;
   wire FE_OCPN27903_n19223;
   wire FE_OCPN27902_n20514;
   wire FE_OCPN27900_n23949;
   wire FE_OCPN27896_n18583;
   wire FE_OCPN27891_n18561;
   wire FE_OCPN27888_sa12_2;
   wire FE_OCPN27887_n17331;
   wire FE_OCPN27884_n26717;
   wire FE_OCPN27882_n18829;
   wire FE_OCPN27881_FE_OFN27126_sa23_3;
   wire FE_OCPN27877_n21980;
   wire FE_OCPN27871_n17317;
   wire FE_OCPN27870_n18527;
   wire FE_OCPN27866_n;
   wire FE_OCPN27859_n25868;
   wire FE_OCPN27848_n23255;
   wire FE_OCPN27843_n18750;
   wire FE_OCPN27840_FE_OFN27078_sa23_5;
   wire FE_OCPN27838_n17747;
   wire FE_OCPN27836_n16976;
   wire FE_OCPN27829_n25102;
   wire FE_OCPN27825_n25169;
   wire FE_OCPN27819_n17245;
   wire FE_OCPN27818_n17267;
   wire FE_OCPN27817_n21921;
   wire FE_OCPN27815_n25769;
   wire FE_OCPN27812_FE_OFN16463_sa32_0;
   wire FE_OCPN27810_n;
   wire FE_OCPN27809_n26938;
   wire FE_OCPN27807_n23375;
   wire FE_OCPN27806_n25497;
   wire FE_OCPN27804_sa12_1;
   wire FE_OCPN27803_sa23_4;
   wire FE_OCPN27800_n;
   wire FE_RN_51_0;
   wire FE_RN_50_0;
   wire FE_RN_49_0;
   wire FE_RN_48_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_OCPN27796_n26659;
   wire FE_OCPN27792_n18333;
   wire FE_OCPN27787_n26728;
   wire FE_OCPN27786_n16490;
   wire FE_OCPN27782_n16873;
   wire FE_OCPN27780_n20083;
   wire FE_OCPN27778_n25621;
   wire FE_OCPN27774_n25351;
   wire FE_OCPN27773_n22070;
   wire FE_OCPN27772_n24234;
   wire FE_OCPN27771_n19275;
   wire FE_OCPN27770_n26049;
   wire FE_OCPN27765_FE_OFN16265_n26527;
   wire FE_OCPN27764_n22152;
   wire FE_OCPN27761_n16977;
   wire FE_OCPN27757_n21819;
   wire FE_OCPN27753_n26685;
   wire FE_OCPN27750_n22293;
   wire FE_OCPN27744_n26362;
   wire FE_OCPN27743_n22009;
   wire FE_OCPN27741_n;
   wire FE_OCPN27740_sa02_4;
   wire FE_OCPN27735_n16750;
   wire FE_OCPN27733_n17996;
   wire FE_OCPN27730_n17464;
   wire FE_OCPN27729_n24362;
   wire FE_OCPN27727_n22964;
   wire FE_OCPN27726_n;
   wire FE_OCPN27723_n;
   wire FE_OCPN27722_n23336;
   wire FE_OCPN27721_n23336;
   wire FE_OCPN27720_n23306;
   wire FE_OCPN27719_n23306;
   wire FE_OCPN27715_n23875;
   wire FE_OCPN27712_sa01_4;
   wire FE_OCPN27710_n19011;
   wire FE_OCPN27703_n19847;
   wire FE_OCPN27697_n16309;
   wire FE_OCPN27690_n16757;
   wire FE_OCPN27689_n20172;
   wire FE_OCPN27685_n26968;
   wire FE_OCPN27684_n17139;
   wire FE_OCPN27682_n25414;
   wire FE_OCPN27679_n18631;
   wire FE_OCPN27678_n26227;
   wire FE_OCPN27675_n17986;
   wire FE_OCPN27673_n18163;
   wire FE_OCPN27666_n17418;
   wire FE_OCPN27665_w3_25;
   wire FE_OCPN27664_w3_25;
   wire FE_OCPN27659_w3_25;
   wire FE_OCPN27656_w3_25;
   wire FE_OCPN27655_w3_25;
   wire FE_OCPN27652_n20176;
   wire FE_RN_44_0;
   wire FE_OCPN27649_n17236;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_RN_38_0;
   wire FE_OCPN27642_n16758;
   wire FE_OCPN27641_n27121;
   wire FE_OCPN27637_n26428;
   wire FE_OCPN27636_sa10_4;
   wire FE_OCPN27635_sa10_4;
   wire FE_OCPN27634_n20169;
   wire FE_OCPN27633_sa20_5;
   wire FE_OCPN27632_n16774;
   wire FE_OCPN27631_n16774;
   wire FE_OCPN27629_n25589;
   wire FE_OCPN27628_n23455;
   wire FE_OCPN27627_sa23_1;
   wire FE_OCPN27625_sa11_5;
   wire FE_OCPN27624_n26971;
   wire FE_OCPN27617_n18016;
   wire FE_OCPN27616_n16760;
   wire FE_OCPN27611_n23426;
   wire FE_OCPN27606_n23869;
   wire FE_OCPN27605_n23357;
   wire FE_OCPN27604_n16421;
   wire FE_OCPN27601_n17475;
   wire FE_OCPN27599_n18875;
   wire FE_OCPN27593_n16908;
   wire FE_OCPN27592_n17501;
   wire FE_OCPN27591_n23742;
   wire FE_RN_37_0;
   wire FE_OCPN27589_n25987;
   wire FE_OCPN27588_n19824;
   wire FE_OCPN27585_sa02_1;
   wire FE_OCPN27584_n22497;
   wire FE_OCPN27583_n26193;
   wire FE_OCPN27580_n;
   wire FE_OCPN27579_FE_OFN16138_sa02_5;
   wire FE_OCPN27577_sa23_4;
   wire FE_OCPN27574_n20196;
   wire FE_OCPN27573_n20196;
   wire FE_OCPN27572_sa02_1;
   wire FE_OCPN27570_n17791;
   wire FE_OCPN27568_sa33_3;
   wire FE_OCPN27566_FE_OFN16138_sa02_5;
   wire FE_OCPN27562_n17447;
   wire FE_RN_35_0;
   wire FE_OCPN27560_n25755;
   wire FE_OCPN27558_sa20_4;
   wire FE_OCPN27557_sa20_4;
   wire FE_OCPN27556_n17843;
   wire FE_OCPN27555_n16422;
   wire FE_OCPN27554_n20007;
   wire FE_OCPN27553_n19975;
   wire FE_RN_27_0;
   wire FE_RN_26_0;
   wire FE_OCPN27546_sa33_4;
   wire FE_OCPN27544_sa33_4;
   wire FE_OCPN27542_sa20_3;
   wire FE_OCPN27541_n26748;
   wire FE_OCPN27539_n16875;
   wire FE_OCPN27538_n25383;
   wire FE_OCPN27535_n;
   wire FE_OCPN27534_n;
   wire FE_OCPN27532_n21643;
   wire FE_OCPN27531_n21643;
   wire FE_OCPN27530_n362;
   wire FE_RN_24_0;
   wire FE_RN_23_0;
   wire FE_OCPN27525_n26434;
   wire FE_OCPN27522_n25921;
   wire FE_OCPN27521_n18163;
   wire FE_OCPN27519_n25407;
   wire FE_OCPN27518_n17251;
   wire FE_OCPN27516_n26292;
   wire FE_OCPN27514_n25981;
   wire FE_OCPN27512_sa11_2;
   wire FE_OCPN27508_n20339;
   wire FE_OCPN27507_n25695;
   wire FE_OCPN27505_n24684;
   wire FE_OCPN27503_n20195;
   wire FE_OCPN27500_n19834;
   wire FE_OCPN27499_FE_OFN16151_sa32_5;
   wire FE_OCPN27498_sa23_2;
   wire FE_OCPN27497_n25431;
   wire FE_OCPN27496_n21820;
   wire FE_OCPN27494_n26479;
   wire FE_OCPN27491_n26351;
   wire FE_OCPN27490_n18798;
   wire FE_RN_21_0;
   wire FE_OCPN27483_FE_OFN16132_sa03_5;
   wire FE_OCPN27482_sa23_5;
   wire FE_OCPN27478_n25011;
   wire FE_OCPN27476_n26852;
   wire FE_OCPN27467_n25483;
   wire FE_OCPN27462_n26215;
   wire FE_OCPN27460_n16913;
   wire FE_OCPN27458_n24891;
   wire FE_OCPN27456_n27189;
   wire FE_OCPN27454_n16789;
   wire FE_OCPN27451_n26236;
   wire FE_OCPN27447_n26638;
   wire FE_OCPN27446_n24847;
   wire FE_OCPN27445_n26837;
   wire FE_OCPN27444_n20064;
   wire FE_OCPN27442_n27202;
   wire FE_OCPN27441_n25688;
   wire FE_OCPN27439_n27030;
   wire FE_OCPN27435_n26790;
   wire FE_OCPN27433_n21571;
   wire FE_OCPN27430_n26334;
   wire FE_OCPN27429_sa12_3;
   wire FE_OCPN27428_n26027;
   wire FE_OCPN27424_n22560;
   wire FE_OCPN27423_sa01_0;
   wire FE_OCPN27421_n25768;
   wire FE_OCPN27420_n18794;
   wire FE_OCPN27419_n26602;
   wire FE_OCPN27414_n23359;
   wire FE_OCPN27412_n24491;
   wire FE_OCPN27405_sa03_4;
   wire FE_OCPN27403_sa01_5;
   wire FE_OCPN27402_n24523;
   wire FE_OCPN27399_n22598;
   wire FE_OCPN27394_n26223;
   wire FE_OCPN27393_sa03_0;
   wire FE_OCPN27391_n27079;
   wire FE_OCPN27388_FE_OFN25990_sa21_4;
   wire FE_OCPN27384_n22888;
   wire FE_OCPN27379_n26809;
   wire FE_OCPN27377_n26853;
   wire FE_OCPN27375_n26860;
   wire FE_OCPN27374_n26394;
   wire FE_OCPN27373_n26172;
   wire FE_OCPN27371_sa20_2;
   wire FE_OCPN27368_sa12_3;
   wire FE_OCPN27367_sa21_0;
   wire FE_OCPN27366_n26326;
   wire FE_OCPN27365_sa11_4;
   wire FE_OCPN27363_n26649;
   wire FE_OCPN27362_n25679;
   wire FE_OCPN27361_n24719;
   wire FE_OCPN27359_n26726;
   wire FE_OCPN27358_n26586;
   wire FE_OCPN27357_n26369;
   wire FE_OCPN27354_n26982;
   wire FE_OCPN27338_n19149;
   wire FE_OCPN27337_n19149;
   wire FE_OCPN27333_n25250;
   wire FE_OCPN27330_n;
   wire FE_OCPN27328_sa21_2;
   wire FE_OCPN27327_sa21_2;
   wire FE_OCPN27322_n25755;
   wire FE_OCPN27321_n26380;
   wire FE_OCPN27320_n410;
   wire FE_OCPN27316_n25849;
   wire FE_OCPN27314_n26113;
   wire FE_OCPN27313_n21845;
   wire FE_OCPN27310_n26389;
   wire FE_OCPN27306_n334;
   wire FE_OCPN27302_n26910;
   wire FE_OCPN27295_n26851;
   wire FE_OCPN27292_n25389;
   wire FE_OCPN27289_sa21_5;
   wire FE_OCPN27288_n25091;
   wire FE_OCPN27285_n18011;
   wire FE_OCPN27284_n26633;
   wire FE_OCPN27283_n26867;
   wire FE_OCPN27282_n25437;
   wire FE_OCPN27276_sa02_0;
   wire FE_OCPN27274_n26394;
   wire FE_OCPN27273_sa02_3;
   wire FE_OCPN27271_n26961;
   wire FE_OCPN27267_n18794;
   wire FE_OCPN27261_sa02_0;
   wire FE_OCPN27253_n17923;
   wire FE_OCPN27252_n22753;
   wire FE_OCPN27246_n22663;
   wire FE_OCPN27242_sa11_1;
   wire FE_OCPN27241_sa11_1;
   wire FE_OCPN27235_n27143;
   wire FE_OCPN27234_n26837;
   wire FE_RN_19_0;
   wire FE_RN_18_0;
   wire FE_RN_17_0;
   wire FE_RN_16_0;
   wire FE_RN_15_0;
   wire FE_OCPN27230_sa32_3;
   wire FE_OCPN27229_sa11_2;
   wire FE_OCPN27228_sa11_2;
   wire FE_OCPN27227_sa00_5;
   wire FE_RN_12_0;
   wire FE_RN_11_0;
   wire FE_RN_10_0;
   wire FE_OCPN27226_n25357;
   wire FE_OCPN27224_sa00_5;
   wire FE_RN_9_0;
   wire FE_RN_8_0;
   wire FE_RN_7_0;
   wire FE_RN_6_0;
   wire FE_RN_4_0;
   wire FE_RN_3_0;
   wire FE_RN_2_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire FE_OFN27222_n14593;
   wire FE_OFN27218_n14745;
   wire FE_OFN27216_n14091;
   wire FE_OFN27214_w3_17;
   wire FE_OFN27212_w3_30;
   wire FE_OFN27211_w3_30;
   wire FE_OFN27210_w3_30;
   wire FE_OFN27209_w3_30;
   wire FE_OFN27208_w3_30;
   wire FE_OFN27207_w3_30;
   wire FE_OFN27206_w3_30;
   wire FE_OFN27202_n;
   wire FE_OFN27200_n;
   wire FE_OFN27196_n;
   wire FE_OFN27189_n;
   wire FE_OFN27186_sa13_4;
   wire FE_OFN27179_n20327;
   wire FE_OFN27176_n;
   wire FE_OFN27173_n;
   wire FE_OFN27172_n17441;
   wire FE_OFN27169_n26683;
   wire FE_OFN27168_n16334;
   wire FE_OFN27165_n;
   wire FE_OFN27163_n20304;
   wire FE_OFN27157_n23928;
   wire FE_OFN27156_n;
   wire FE_OFN27155_sa21_4;
   wire FE_OFN27152_n17315;
   wire FE_OFN27151_n;
   wire FE_OFN27150_n22175;
   wire FE_OFN27148_sa32_3;
   wire FE_OFN27147_n25284;
   wire FE_OFN27145_n23216;
   wire FE_OFN27142_n25934;
   wire FE_OFN27140_n20007;
   wire FE_OFN27138_n24012;
   wire FE_OFN27136_n15992;
   wire FE_OFN27135_n15992;
   wire FE_OFN27133_n21725;
   wire FE_OFN27131_w3_29;
   wire FE_OFN27130_w3_28;
   wire FE_OFN27129_w3_28;
   wire FE_OFN27128_sa23_3;
   wire FE_OFN27127_sa23_3;
   wire FE_OFN27126_sa23_3;
   wire FE_OFN27125_n21057;
   wire FE_OFN27124_w3_1;
   wire FE_OFN27123_n26275;
   wire FE_OFN27116_n16293;
   wire FE_OFN27115_n;
   wire FE_OFN27111_n;
   wire FE_OFN27100_n25675;
   wire FE_OFN27096_n;
   wire FE_OFN27094_n24956;
   wire FE_OFN27090_n23558;
   wire FE_OFN27089_n23558;
   wire FE_OFN27088_n23754;
   wire FE_OFN27085_n;
   wire FE_OFN27083_n;
   wire FE_OFN27082_n25377;
   wire FE_OFN27078_sa23_5;
   wire FE_OFN27075_n23409;
   wire FE_OFN27074_n13868;
   wire FE_OFN27072_n18671;
   wire FE_OFN27070_n;
   wire FE_OFN27069_n24478;
   wire FE_OFN27066_n13869;
   wire FE_OFN27065_n17059;
   wire FE_OFN27064_n22438;
   wire FE_OFN27062_n16438;
   wire FE_OFN27061_n15239;
   wire FE_OFN27058_n22094;
   wire FE_OFN27057_n13662;
   wire FE_OFN27056_n22995;
   wire FE_OFN27052_n21551;
   wire FE_OFN27048_n23045;
   wire FE_OFN27046_n22024;
   wire FE_OFN27045_n;
   wire FE_OFN27044_n15236;
   wire FE_OFN27043_n;
   wire FE_OFN26651_n19573;
   wire FE_OFN26650_n27164;
   wire FE_OFN26649_n22206;
   wire FE_OFN26648_n22197;
   wire FE_OFN26646_n16159;
   wire FE_OFN26645_n;
   wire FE_OFN26644_n19599;
   wire FE_OFN26642_w3_14;
   wire FE_OFN26641_w3_14;
   wire FE_OFN26640_w3_14;
   wire FE_OFN26639_w3_14;
   wire FE_OFN26638_w3_14;
   wire FE_OFN26637_w3_14;
   wire FE_OFN26636_w3_14;
   wire FE_OFN26635_w3_14;
   wire FE_OFN26634_w3_14;
   wire FE_OFN26633_w3_14;
   wire FE_OFN26630_n16190;
   wire FE_OFN26629_sa31_4;
   wire FE_OFN26628_n;
   wire FE_OFN26624_n15376;
   wire FE_OFN26614_n;
   wire FE_OFN26600_sa13_0;
   wire FE_OFN26597_n;
   wire FE_OFN26595_sa31_4;
   wire FE_OFN26591_w3_3;
   wire FE_OFN26589_sa12_1;
   wire FE_OFN26588_n24062;
   wire FE_OFN26587_n23011;
   wire FE_OFN26585_n23011;
   wire FE_OFN26584_n20059;
   wire FE_OFN26581_n21317;
   wire FE_OFN26578_n23913;
   wire FE_OFN26577_n;
   wire FE_OFN26575_n20369;
   wire FE_OFN26572_n19405;
   wire FE_OFN26570_n20866;
   wire FE_OFN26569_n20866;
   wire FE_OFN26567_n;
   wire FE_OFN26566_n24208;
   wire FE_OFN26564_n;
   wire FE_OFN26559_n26754;
   wire FE_OFN26558_n26911;
   wire FE_OFN26557_n19302;
   wire FE_OFN26556_n23236;
   wire FE_OFN26554_n19170;
   wire FE_OFN26553_n24644;
   wire FE_OFN26552_n14545;
   wire FE_OFN26550_n16331;
   wire FE_OFN26549_n16248;
   wire FE_OFN26548_n18206;
   wire FE_OFN26546_n24537;
   wire FE_OFN26545_n16447;
   wire FE_OFN26542_n26155;
   wire FE_OFN26541_n16100;
   wire FE_OFN26539_w3_19;
   wire FE_OFN26538_w3_19;
   wire FE_OFN26535_w3_19;
   wire FE_OFN26534_w3_19;
   wire FE_OFN26533_n21922;
   wire FE_OFN26532_n13766;
   wire FE_OFN26531_n;
   wire FE_OFN26528_n23302;
   wire FE_OFN26172_n19609;
   wire FE_OFN26170_n19361;
   wire FE_OFN26166_n24855;
   wire FE_OFN26164_w3_13;
   wire FE_OFN26163_w3_13;
   wire FE_OFN26162_w3_13;
   wire FE_OFN26161_sa10_4;
   wire FE_OFN26160_sa10_4;
   wire FE_OFN26159_n22080;
   wire FE_OFN26158_n22224;
   wire FE_OFN26154_n16132;
   wire FE_OFN26150_n21253;
   wire FE_OFN26149_n26245;
   wire FE_OFN26148_n26245;
   wire FE_OFN26147_n27041;
   wire FE_OFN26146_n18774;
   wire FE_OFN26141_n23307;
   wire FE_OFN26140_n23585;
   wire FE_OFN26139_n16125;
   wire FE_OFN26137_n16125;
   wire FE_OFN26136_sa22_3;
   wire FE_OFN26133_sa22_3;
   wire FE_OFN26132_sa01_3;
   wire FE_OFN26131_n15376;
   wire FE_OFN26129_w3_15;
   wire FE_OFN26127_n22925;
   wire FE_OFN26125_n22742;
   wire FE_OFN26121_n16107;
   wire FE_OFN26120_n;
   wire FE_OFN26114_n;
   wire FE_OFN26112_n13288;
   wire FE_OFN26111_n13288;
   wire FE_OFN26110_n15848;
   wire FE_OFN26107_sa31_5;
   wire FE_OFN26104_n13659;
   wire FE_OFN26096_n16294;
   wire FE_OFN26095_n16293;
   wire FE_OFN26091_n24663;
   wire FE_OFN26084_n15106;
   wire FE_OFN26078_sa33_2;
   wire FE_OFN26077_n;
   wire FE_OFN26076_w3_30;
   wire FE_OFN26073_n;
   wire FE_OFN26072_n26720;
   wire FE_OFN26062_n16435;
   wire FE_OFN26061_n;
   wire FE_OFN26060_sa31_4;
   wire FE_OFN26059_n;
   wire FE_OFN26058_w3_1;
   wire FE_OFN26057_w3_1;
   wire FE_OFN26055_n;
   wire FE_OFN26054_sa01_3;
   wire FE_OFN26053_n25415;
   wire FE_OFN26051_w3_27;
   wire FE_OFN26049_w3_27;
   wire FE_OFN26048_w3_27;
   wire FE_OFN26045_n25377;
   wire FE_OFN26041_w3_17;
   wire FE_OFN26039_sa10_2;
   wire FE_OFN26038_n24887;
   wire FE_OFN26037_n22144;
   wire FE_OFN26035_n;
   wire FE_OFN26033_n20197;
   wire FE_OFN26032_n20230;
   wire FE_OFN26031_n22499;
   wire FE_OFN26030_n25368;
   wire FE_OFN26024_n26115;
   wire FE_OFN26023_n20807;
   wire FE_OFN26021_n16253;
   wire FE_OFN26020_n14010;
   wire FE_OFN26019_n26319;
   wire FE_OFN26015_sa31_3;
   wire FE_OFN26014_sa31_3;
   wire FE_OFN26012_n27208;
   wire FE_OFN26009_n18213;
   wire FE_OFN26007_n16010;
   wire FE_OFN26005_n17451;
   wire FE_OFN26003_n15992;
   wire FE_OFN26001_n24836;
   wire FE_OFN25999_n25875;
   wire FE_OFN25998_n17781;
   wire FE_OFN25997_n;
   wire FE_OFN25996_n26006;
   wire FE_OFN25993_n16767;
   wire FE_OFN25989_sa21_4;
   wire FE_OFN25987_n23322;
   wire FE_OFN25986_n21012;
   wire FE_OFN25985_n15997;
   wire FE_OFN25981_n13868;
   wire FE_OFN25980_n19087;
   wire FE_OFN25979_n;
   wire FE_OFN25977_n18922;
   wire FE_OFN25975_n16217;
   wire FE_OFN25973_n26087;
   wire FE_OFN25972_n20056;
   wire FE_OFN25971_n14472;
   wire FE_OFN25970_n;
   wire FE_OFN25968_n22668;
   wire FE_OFN25966_n13646;
   wire FE_OFN25963_n27123;
   wire FE_OFN25961_w3_8;
   wire FE_OFN25960_n;
   wire FE_OFN25959_n23011;
   wire FE_OFN25958_sa30_3;
   wire FE_OFN25956_n16575;
   wire FE_OFN25955_n25122;
   wire FE_OFN25954_n18719;
   wire FE_OFN25952_n22312;
   wire FE_OFN25950_sa01_2;
   wire FE_OFN25949_n21475;
   wire FE_OFN25946_sa32_6;
   wire FE_OFN25941_n22857;
   wire FE_OFN25940_n24621;
   wire FE_OFN25939_n26275;
   wire FE_OFN25938_sa33_3;
   wire FE_OFN25937_n23943;
   wire FE_OFN25934_n;
   wire FE_OFN25929_n16073;
   wire FE_OFN25928_n15779;
   wire FE_OFN25927_n26527;
   wire FE_OFN25926_n26922;
   wire FE_OFN25920_n15995;
   wire FE_OFN25918_n15813;
   wire FE_OFN25917_n21591;
   wire FE_OFN25915_n15514;
   wire FE_OFN25912_n15848;
   wire FE_OFN25911_n26491;
   wire FE_OFN25909_w3_20;
   wire FE_OFN25908_sa12_2;
   wire FE_OFN25907_sa12_2;
   wire FE_OFN25906_sa12_2;
   wire FE_OFN25904_n16143;
   wire FE_OFN25901_n22133;
   wire FE_OFN25900_w3_4;
   wire FE_OFN25899_w3_4;
   wire FE_OFN25897_w3_4;
   wire FE_OFN25896_w3_4;
   wire FE_OFN25895_n13662;
   wire FE_OFN25893_n15214;
   wire FE_OFN25892_n16264;
   wire FE_OFN25891_n15770;
   wire FE_OFN25890_n23497;
   wire FE_OFN25889_n20913;
   wire FE_OFN25887_w3_3;
   wire FE_OFN25886_w3_3;
   wire FE_OFN25883_n22945;
   wire FE_OFN25882_n16262;
   wire FE_OFN25881_w3_24;
   wire FE_OFN25880_w3_24;
   wire FE_OFN25879_sa11_0;
   wire FE_OFN25878_n17329;
   wire FE_OFN25875_n15227;
   wire FE_OFN21730_sa03_3;
   wire FE_OFN16463_sa32_0;
   wire FE_OFN16459_n;
   wire FE_OFN16451_n;
   wire FE_OFN16450_n23315;
   wire FE_OFN16448_n;
   wire FE_OFN16447_n16749;
   wire FE_OFN16445_sa13_1;
   wire FE_OFN16444_sa13_1;
   wire FE_OFN16441_w3_21;
   wire FE_OFN16437_n;
   wire FE_OFN16436_w3_11;
   wire FE_OFN16432_w3_16;
   wire FE_OFN16431_w3_16;
   wire FE_OFN16430_sa33_3;
   wire FE_OFN16426_w3_20;
   wire FE_OFN16423_n24831;
   wire FE_OFN16421_n23974;
   wire FE_OFN16417_n;
   wire FE_OFN16415_sa31_2;
   wire FE_OFN16413_n26687;
   wire FE_OFN16412_w3_26;
   wire FE_OFN16411_n15884;
   wire FE_OFN16407_n23322;
   wire FE_OFN16405_n16117;
   wire FE_OFN16403_n16117;
   wire FE_OFN16402_n19704;
   wire FE_OFN16400_n17404;
   wire FE_OFN16398_n24241;
   wire FE_OFN16396_n25869;
   wire FE_OFN16395_n26801;
   wire FE_OFN16392_n24102;
   wire FE_OFN16391_n22490;
   wire FE_OFN16389_n19359;
   wire FE_OFN16385_n18525;
   wire FE_OFN16380_n20584;
   wire FE_OFN16378_n23030;
   wire FE_OFN16377_n23998;
   wire FE_OFN16375_n25750;
   wire FE_OFN16370_n16261;
   wire FE_OFN16369_n16717;
   wire FE_OFN16368_n18545;
   wire FE_OFN16367_n21973;
   wire FE_OFN16361_n16263;
   wire FE_OFN16360_n16051;
   wire FE_OFN16356_n22874;
   wire FE_OFN16353_n25672;
   wire FE_OFN16352_n14289;
   wire FE_OFN16351_n26084;
   wire FE_OFN16349_n19960;
   wire FE_OFN16348_n15949;
   wire FE_OFN16341_n27008;
   wire FE_OFN16340_n26317;
   wire FE_OFN16334_n25823;
   wire FE_OFN16333_sa30_4;
   wire FE_OFN16331_n27151;
   wire FE_OFN16329_n27151;
   wire FE_OFN16328_n23821;
   wire FE_OFN16326_n19058;
   wire FE_OFN16324_n25832;
   wire FE_OFN16322_n25946;
   wire FE_OFN16319_n20527;
   wire FE_OFN16316_n24840;
   wire FE_OFN16315_sa31_5;
   wire FE_OFN16313_w3_0;
   wire FE_OFN16311_n26252;
   wire FE_OFN16307_n27010;
   wire FE_OFN16306_n27041;
   wire FE_OFN16305_n15984;
   wire FE_OFN16304_n22808;
   wire FE_OFN16301_n25905;
   wire FE_OFN16300_n14826;
   wire FE_OFN16298_sa13_2;
   wire FE_OFN16297_n24803;
   wire FE_OFN16295_n23837;
   wire FE_OFN16294_n19461;
   wire FE_OFN16292_n25175;
   wire FE_OFN16291_n23142;
   wire FE_OFN16287_n16230;
   wire FE_OFN16283_n26788;
   wire FE_OFN16281_n26011;
   wire FE_OFN16278_w3_5;
   wire FE_OFN16276_w3_5;
   wire FE_OFN16275_n26536;
   wire FE_OFN16274_n14664;
   wire FE_OFN16273_n14664;
   wire FE_OFN16272_n24767;
   wire FE_OFN16271_n26814;
   wire FE_OFN16269_n15808;
   wire FE_OFN16268_sa13_3;
   wire FE_OFN16267_sa21_4;
   wire FE_OFN16265_n26527;
   wire FE_OFN16263_n25976;
   wire FE_OFN16262_n16052;
   wire FE_OFN16260_n24927;
   wire FE_OFN16255_n26684;
   wire FE_OFN16254_n14008;
   wire FE_OFN16253_n16189;
   wire FE_OFN16252_n27003;
   wire FE_OFN16251_n16162;
   wire FE_OFN16250_n26165;
   wire FE_OFN16249_n25956;
   wire FE_OFN16248_n20235;
   wire FE_OFN16247_sa30_1;
   wire FE_OFN16246_n16113;
   wire FE_OFN16241_n23552;
   wire FE_OFN16240_n14011;
   wire FE_OFN16239_n14005;
   wire FE_OFN16236_n13655;
   wire FE_OFN16235_n15055;
   wire FE_OFN16234_sa02_2;
   wire FE_OFN16232_n17691;
   wire FE_OFN16231_n17691;
   wire FE_OFN16229_sa20_4;
   wire FE_OFN16227_n26602;
   wire FE_OFN16225_n15195;
   wire FE_OFN16221_n21234;
   wire FE_OFN16220_n25219;
   wire FE_OFN16218_n18418;
   wire FE_OFN16216_n19573;
   wire FE_OFN16215_ld_r;
   wire FE_OFN16214_ld_r;
   wire FE_OFN16213_ld_r;
   wire FE_OFN16211_n13876;
   wire FE_OFN16210_n13876;
   wire FE_OFN16208_n23101;
   wire FE_OFN16206_n15240;
   wire FE_OFN16203_n22313;
   wire FE_OFN16202_n19806;
   wire FE_OFN16201_n15197;
   wire FE_OFN16200_sa30_2;
   wire FE_OFN16197_sa31_6;
   wire FE_OFN16195_n13771;
   wire FE_OFN16193_n15200;
   wire FE_OFN16192_n17524;
   wire FE_OFN16189_n25672;
   wire FE_OFN16184_w3_9;
   wire FE_OFN16182_w3_9;
   wire FE_OFN16181_sa13_5;
   wire FE_OFN16180_n26542;
   wire FE_OFN16179_w3_19;
   wire FE_OFN16178_w3_19;
   wire FE_OFN16177_n27207;
   wire FE_OFN16176_n27207;
   wire FE_OFN16170_n26637;
   wire FE_OFN16169_n26567;
   wire FE_OFN16164_n25081;
   wire FE_OFN16163_n26584;
   wire FE_OFN16162_n25869;
   wire FE_OFN16159_w3_24;
   wire FE_OFN16158_n26959;
   wire FE_OFN16153_n16747;
   wire FE_OFN16150_sa10_4;
   wire FE_OFN16148_n25466;
   wire FE_OFN16145_n15214;
   wire FE_OFN16141_sa01_3;
   wire FE_OFN16136_sa02_5;
   wire FE_OFN16135_sa22_4;
   wire FE_OFN16131_sa12_1;
   wire FE_OFN16130_n19119;
   wire FE_OFN16128_sa32_2;
   wire FE_OFN175_sa12_6;
   wire FE_OFN174_sa33_6;
   wire FE_OFN173_sa33_6;
   wire FE_OFN171_n26739;
   wire FE_OFN169_n23992;
   wire FE_OFN168_n24268;
   wire FE_OFN167_sa21_7;
   wire FE_OFN166_sa12_7;
   wire FE_OFN165_sa12_7;
   wire FE_OFN164_n24529;
   wire FE_OFN163_sa00_7;
   wire FE_OFN162_sa23_7;
   wire FE_OFN161_n26440;
   wire FE_OFN160_n26440;
   wire FE_OFN156_sa03_6;
   wire FE_OFN155_n26788;
   wire FE_OFN154_n26788;
   wire FE_OFN152_n20170;
   wire FE_OFN150_sa11_7;
   wire FE_OFN148_sa00_1;
   wire FE_OFN142_sa10_0;
   wire FE_OFN141_sa03_1;
   wire FE_OFN140_w3_2;
   wire FE_OFN138_sa11_0;
   wire FE_OFN136_sa32_7;
   wire FE_OFN135_n26172;
   wire FE_OFN134_sa31_6;
   wire FE_OFN133_n24306;
   wire FE_OFN132_n18247;
   wire FE_OFN131_sa10_6;
   wire FE_OFN130_sa10_5;
   wire FE_OFN128_sa13_7;
   wire FE_OFN127_sa13_7;
   wire FE_OFN125_sa01_1;
   wire FE_OFN122_n22751;
   wire FE_OFN118_sa03_7;
   wire FE_OFN117_n24628;
   wire FE_OFN116_n27187;
   wire FE_OFN115_n27187;
   wire FE_OFN114_n22512;
   wire FE_OFN112_n15994;
   wire FE_OFN109_n15994;
   wire FE_OFN108_n26971;
   wire FE_OFN107_n22745;
   wire FE_OFN106_n24511;
   wire FE_OFN105_n27178;
   wire FE_OFN104_n27179;
   wire FE_OFN102_w3_12;
   wire FE_OFN101_w3_12;
   wire FE_OFN100_sa31_1;
   wire FE_OFN97_n20994;
   wire FE_OFN95_n19498;
   wire FE_OFN94_sa11_5;
   wire FE_OFN90_sa33_7;
   wire FE_OFN87_n21551;
   wire FE_OFN86_n26674;
   wire FE_OFN85_n23588;
   wire FE_OFN79_n16857;
   wire FE_OFN78_n22457;
   wire FE_OFN75_n15253;
   wire FE_OFN73_sa12_5;
   wire FE_OFN72_n15506;
   wire FE_OFN70_w2_20;
   wire FE_OFN69_sa32_4;
   wire FE_OFN68_sa02_6;
   wire FE_OFN66_w1_25;
   wire FE_OFN65_n21412;
   wire FE_OFN64_w0_31;
   wire FE_OFN62_sa21_3;
   wire FE_OFN60_n27007;
   wire FE_OFN59_sa10_7;
   wire FE_OFN58_w1_4;
   wire FE_OFN57_n19754;
   wire FE_OFN56_n14826;
   wire FE_OFN55_sa22_5;
   wire FE_OFN54_sa22_2;
   wire FE_OFN53_w0_8;
   wire FE_OFN51_w3_18;
   wire FE_OFN50_w3_18;
   wire FE_OFN49_w0_23;
   wire FE_OFN48_w0_2;
   wire FE_OFN47_w1_2;
   wire FE_OFN46_w0_12;
   wire FE_OFN45_sa23_6;
   wire FE_OFN44_w0_9;
   wire FE_OFN43_w0_10;
   wire FE_OFN42_sa00_0;
   wire FE_OFN41_n20971;
   wire FE_OFN40_w0_19;
   wire FE_OFN39_w0_21;
   wire FE_OFN38_w0_17;
   wire FE_OFN37_w3_23;
   wire FE_OFN34_w3_22;
   wire FE_OFN31_sa20_0;
   wire FE_OFN30_n25256;
   wire FE_OFN28_w3_23;
   wire FE_OFN27_n16125;
   wire FE_OFN26_n16125;
   wire FE_OFN25_n16125;
   wire FE_OFN24_n16125;
   wire FE_OFN23_n16125;
   wire FE_OFN22_n16125;
   wire FE_OFN21_n16125;
   wire FE_OFN20_n16125;
   wire FE_OFN19_n16125;
   wire FE_OFN18_n16125;
   wire FE_OFN17_FE_DBTN0_ld_r;
   wire FE_OFN16_FE_DBTN0_ld_r;
   wire FE_OFN15_FE_DBTN0_ld_r;
   wire FE_OFN14_FE_DBTN0_ld_r;
   wire FE_OFN13_FE_DBTN0_ld_r;
   wire FE_OFN12_FE_DBTN0_ld_r;
   wire FE_OFN8_w3_14;
   wire FE_OFN7_w3_22;
   wire FE_OFN6_w3_22;
   wire FE_OFN5_w3_22;
   wire FE_OFN4_w3_22;
   wire FE_OFN3_ld_r;
   wire FE_OFN2_ld_r;
   wire FE_OFN1_ld_r;
   wire FE_OFN0_ld;
   wire FE_DBTN0_ld_r;
   wire dcnt_3_;
   wire dcnt_2_;
   wire dcnt_1_;
   wire dcnt_0_;
   wire text_in_r_127_;
   wire text_in_r_126_;
   wire text_in_r_125_;
   wire text_in_r_124_;
   wire text_in_r_123_;
   wire text_in_r_122_;
   wire text_in_r_121_;
   wire text_in_r_120_;
   wire text_in_r_119_;
   wire text_in_r_118_;
   wire text_in_r_117_;
   wire text_in_r_116_;
   wire text_in_r_115_;
   wire text_in_r_114_;
   wire text_in_r_113_;
   wire text_in_r_112_;
   wire text_in_r_111_;
   wire text_in_r_110_;
   wire text_in_r_109_;
   wire text_in_r_108_;
   wire text_in_r_107_;
   wire text_in_r_106_;
   wire text_in_r_105_;
   wire text_in_r_104_;
   wire text_in_r_103_;
   wire text_in_r_102_;
   wire text_in_r_101_;
   wire text_in_r_100_;
   wire text_in_r_99_;
   wire text_in_r_98_;
   wire text_in_r_97_;
   wire text_in_r_96_;
   wire text_in_r_95_;
   wire text_in_r_94_;
   wire text_in_r_93_;
   wire text_in_r_92_;
   wire text_in_r_91_;
   wire text_in_r_90_;
   wire text_in_r_89_;
   wire text_in_r_88_;
   wire text_in_r_87_;
   wire text_in_r_86_;
   wire text_in_r_85_;
   wire text_in_r_84_;
   wire text_in_r_83_;
   wire text_in_r_82_;
   wire text_in_r_81_;
   wire text_in_r_80_;
   wire text_in_r_79_;
   wire text_in_r_78_;
   wire text_in_r_77_;
   wire text_in_r_76_;
   wire text_in_r_75_;
   wire text_in_r_74_;
   wire text_in_r_73_;
   wire text_in_r_72_;
   wire text_in_r_71_;
   wire text_in_r_70_;
   wire text_in_r_69_;
   wire text_in_r_68_;
   wire text_in_r_67_;
   wire text_in_r_66_;
   wire text_in_r_65_;
   wire text_in_r_64_;
   wire text_in_r_63_;
   wire text_in_r_62_;
   wire text_in_r_61_;
   wire text_in_r_60_;
   wire text_in_r_59_;
   wire text_in_r_58_;
   wire text_in_r_57_;
   wire text_in_r_56_;
   wire text_in_r_55_;
   wire text_in_r_54_;
   wire text_in_r_53_;
   wire text_in_r_52_;
   wire text_in_r_51_;
   wire text_in_r_50_;
   wire text_in_r_49_;
   wire text_in_r_48_;
   wire text_in_r_47_;
   wire text_in_r_46_;
   wire text_in_r_45_;
   wire text_in_r_44_;
   wire text_in_r_43_;
   wire text_in_r_42_;
   wire text_in_r_41_;
   wire text_in_r_40_;
   wire text_in_r_39_;
   wire text_in_r_38_;
   wire text_in_r_37_;
   wire text_in_r_36_;
   wire text_in_r_35_;
   wire text_in_r_34_;
   wire text_in_r_33_;
   wire text_in_r_32_;
   wire text_in_r_31_;
   wire text_in_r_30_;
   wire text_in_r_29_;
   wire text_in_r_28_;
   wire text_in_r_27_;
   wire text_in_r_26_;
   wire text_in_r_25_;
   wire text_in_r_24_;
   wire text_in_r_23_;
   wire text_in_r_22_;
   wire text_in_r_21_;
   wire text_in_r_20_;
   wire text_in_r_19_;
   wire text_in_r_18_;
   wire text_in_r_17_;
   wire text_in_r_16_;
   wire text_in_r_15_;
   wire text_in_r_14_;
   wire text_in_r_13_;
   wire text_in_r_12_;
   wire text_in_r_11_;
   wire text_in_r_10_;
   wire text_in_r_9_;
   wire text_in_r_8_;
   wire text_in_r_7_;
   wire text_in_r_6_;
   wire text_in_r_5_;
   wire text_in_r_4_;
   wire text_in_r_3_;
   wire text_in_r_2_;
   wire text_in_r_1_;
   wire text_in_r_0_;
   wire ld_r;
   wire w3_31_;
   wire w3_30_;
   wire w3_29_;
   wire w3_28_;
   wire w3_27_;
   wire w3_26_;
   wire w3_25_;
   wire w3_24_;
   wire w3_23_;
   wire w3_22_;
   wire w3_21_;
   wire w3_20_;
   wire w3_19_;
   wire w3_18_;
   wire w3_17_;
   wire w3_16_;
   wire w3_15_;
   wire w3_14_;
   wire w3_13_;
   wire w3_12_;
   wire w3_11_;
   wire w3_10_;
   wire w3_9_;
   wire w3_8_;
   wire w3_7_;
   wire w3_6_;
   wire w3_5_;
   wire w3_4_;
   wire w3_3_;
   wire w3_2_;
   wire w3_1_;
   wire w3_0_;
   wire sa33_7_;
   wire sa33_6_;
   wire sa33_5_;
   wire sa33_4_;
   wire sa33_3_;
   wire sa33_2_;
   wire sa33_1_;
   wire sa33_0_;
   wire sa23_7_;
   wire sa23_6_;
   wire sa23_5_;
   wire sa23_4_;
   wire sa23_3_;
   wire sa23_2_;
   wire sa23_1_;
   wire sa23_0_;
   wire sa13_7_;
   wire sa13_6_;
   wire sa13_5_;
   wire sa13_4_;
   wire sa13_3_;
   wire sa13_2_;
   wire sa13_1_;
   wire sa13_0_;
   wire sa03_7_;
   wire sa03_6_;
   wire sa03_5_;
   wire sa03_4_;
   wire sa03_3_;
   wire sa03_2_;
   wire sa03_1_;
   wire sa03_0_;
   wire w2_31_;
   wire w2_30_;
   wire w2_29_;
   wire w2_28_;
   wire w2_27_;
   wire w2_26_;
   wire w2_25_;
   wire w2_24_;
   wire w2_23_;
   wire w2_22_;
   wire w2_21_;
   wire w2_20_;
   wire w2_19_;
   wire w2_18_;
   wire w2_17_;
   wire w2_16_;
   wire w2_15_;
   wire w2_14_;
   wire w2_13_;
   wire w2_12_;
   wire w2_11_;
   wire w2_10_;
   wire w2_9_;
   wire w2_8_;
   wire w2_7_;
   wire w2_6_;
   wire w2_5_;
   wire w2_4_;
   wire w2_3_;
   wire w2_2_;
   wire w2_1_;
   wire w2_0_;
   wire sa32_7_;
   wire sa32_6_;
   wire sa32_5_;
   wire sa32_4_;
   wire sa32_3_;
   wire sa32_2_;
   wire sa32_1_;
   wire sa32_0_;
   wire sa22_7_;
   wire sa22_6_;
   wire sa22_5_;
   wire sa22_4_;
   wire sa22_3_;
   wire sa22_2_;
   wire sa22_1_;
   wire sa22_0_;
   wire sa12_7_;
   wire sa12_6_;
   wire sa12_5_;
   wire sa12_4_;
   wire sa12_3_;
   wire sa12_2_;
   wire sa12_1_;
   wire sa12_0_;
   wire sa02_7_;
   wire sa02_6_;
   wire sa02_5_;
   wire sa02_4_;
   wire sa02_3_;
   wire sa02_2_;
   wire sa02_1_;
   wire sa02_0_;
   wire w1_31_;
   wire w1_30_;
   wire w1_29_;
   wire w1_28_;
   wire w1_27_;
   wire w1_26_;
   wire w1_25_;
   wire w1_24_;
   wire w1_23_;
   wire w1_22_;
   wire w1_21_;
   wire w1_20_;
   wire w1_19_;
   wire w1_18_;
   wire w1_17_;
   wire w1_16_;
   wire w1_15_;
   wire w1_14_;
   wire w1_13_;
   wire w1_12_;
   wire w1_11_;
   wire w1_10_;
   wire w1_9_;
   wire w1_8_;
   wire w1_7_;
   wire w1_6_;
   wire w1_5_;
   wire w1_4_;
   wire w1_3_;
   wire w1_2_;
   wire w1_1_;
   wire w1_0_;
   wire sa31_7_;
   wire sa31_6_;
   wire sa31_5_;
   wire sa31_4_;
   wire sa31_3_;
   wire sa31_2_;
   wire sa31_1_;
   wire sa31_0_;
   wire sa21_7_;
   wire sa21_6_;
   wire sa21_5_;
   wire sa21_4_;
   wire sa21_3_;
   wire sa21_2_;
   wire sa21_1_;
   wire sa21_0_;
   wire sa11_7_;
   wire sa11_6_;
   wire sa11_5_;
   wire sa11_4_;
   wire sa11_3_;
   wire sa11_2_;
   wire sa11_1_;
   wire sa11_0_;
   wire sa01_7_;
   wire sa01_6_;
   wire sa01_5_;
   wire sa01_4_;
   wire sa01_3_;
   wire sa01_2_;
   wire sa01_1_;
   wire sa01_0_;
   wire w0_31_;
   wire w0_30_;
   wire w0_29_;
   wire w0_28_;
   wire w0_27_;
   wire w0_26_;
   wire w0_25_;
   wire w0_24_;
   wire w0_23_;
   wire w0_22_;
   wire w0_21_;
   wire w0_20_;
   wire w0_19_;
   wire w0_18_;
   wire w0_17_;
   wire w0_16_;
   wire w0_15_;
   wire w0_14_;
   wire w0_13_;
   wire w0_12_;
   wire w0_11_;
   wire w0_10_;
   wire w0_9_;
   wire w0_8_;
   wire w0_7_;
   wire w0_6_;
   wire w0_5_;
   wire w0_4_;
   wire w0_3_;
   wire w0_2_;
   wire w0_1_;
   wire w0_0_;
   wire sa30_7_;
   wire sa30_6_;
   wire sa30_5_;
   wire sa30_4_;
   wire sa30_3_;
   wire sa30_2_;
   wire sa30_1_;
   wire sa30_0_;
   wire sa20_7_;
   wire sa20_6_;
   wire sa20_5_;
   wire sa20_4_;
   wire sa20_3_;
   wire sa20_2_;
   wire sa20_1_;
   wire sa20_0_;
   wire sa10_7_;
   wire sa10_6_;
   wire sa10_5_;
   wire sa10_4_;
   wire sa10_3_;
   wire sa10_2_;
   wire sa10_1_;
   wire sa10_0_;
   wire sa00_7_;
   wire sa00_6_;
   wire sa00_5_;
   wire sa00_4_;
   wire sa00_3_;
   wire sa00_2_;
   wire sa00_1_;
   wire sa00_0_;
   wire u0_rcon_24_;
   wire u0_rcon_25_;
   wire u0_rcon_26_;
   wire u0_rcon_27_;
   wire u0_rcon_28_;
   wire u0_rcon_29_;
   wire u0_rcon_30_;
   wire u0_rcon_31_;
   wire u0_r0_rcnt_0_;
   wire u0_r0_rcnt_1_;
   wire u0_r0_rcnt_2_;
   wire u0_r0_rcnt_3_;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n669;
   wire n671;
   wire n673;
   wire n675;
   wire n677;
   wire n679;
   wire n681;
   wire n683;
   wire n685;
   wire n687;
   wire n689;
   wire n691;
   wire n693;
   wire n695;
   wire n697;
   wire n699;
   wire n701;
   wire n703;
   wire n705;
   wire n707;
   wire n709;
   wire n711;
   wire n713;
   wire n715;
   wire n717;
   wire n719;
   wire n721;
   wire n723;
   wire n725;
   wire n727;
   wire n729;
   wire n731;
   wire n733;
   wire n735;
   wire n737;
   wire n739;
   wire n741;
   wire n743;
   wire n745;
   wire n747;
   wire n749;
   wire n751;
   wire n753;
   wire n755;
   wire n757;
   wire n759;
   wire n761;
   wire n763;
   wire n765;
   wire n767;
   wire n769;
   wire n771;
   wire n773;
   wire n775;
   wire n777;
   wire n779;
   wire n781;
   wire n783;
   wire n785;
   wire n787;
   wire n789;
   wire n791;
   wire n793;
   wire n795;
   wire n797;
   wire n799;
   wire n801;
   wire n803;
   wire n805;
   wire n807;
   wire n809;
   wire n811;
   wire n813;
   wire n815;
   wire n817;
   wire n819;
   wire n821;
   wire n823;
   wire n825;
   wire n827;
   wire n829;
   wire n831;
   wire n833;
   wire n835;
   wire n837;
   wire n839;
   wire n841;
   wire n843;
   wire n845;
   wire n847;
   wire n849;
   wire n851;
   wire n853;
   wire n855;
   wire n857;
   wire n859;
   wire n861;
   wire n863;
   wire n865;
   wire n867;
   wire n869;
   wire n871;
   wire n873;
   wire n875;
   wire n877;
   wire n879;
   wire n881;
   wire n883;
   wire n885;
   wire n887;
   wire n889;
   wire n891;
   wire n893;
   wire n895;
   wire n897;
   wire n899;
   wire n901;
   wire n903;
   wire n905;
   wire n907;
   wire n909;
   wire n911;
   wire n913;
   wire n915;
   wire n917;
   wire n919;
   wire n921;
   wire n923;
   wire n924;
   wire n926;
   wire n928;
   wire n930;
   wire n12994;
   wire n12998;
   wire n12999;
   wire n13000;
   wire n13001;
   wire n13002;
   wire n13003;
   wire n13004;
   wire n13005;
   wire n13006;
   wire n13007;
   wire n13008;
   wire n13009;
   wire n13010;
   wire n13011;
   wire n13012;
   wire n13013;
   wire n13014;
   wire n13015;
   wire n13016;
   wire n13017;
   wire n13018;
   wire n13019;
   wire n13020;
   wire n13021;
   wire n13022;
   wire n13023;
   wire n13024;
   wire n13025;
   wire n13026;
   wire n13027;
   wire n13028;
   wire n13029;
   wire n13030;
   wire n13031;
   wire n13032;
   wire n13033;
   wire n13034;
   wire n13035;
   wire n13036;
   wire n13037;
   wire n13038;
   wire n13039;
   wire n13040;
   wire n13041;
   wire n13042;
   wire n13043;
   wire n13044;
   wire n13045;
   wire n13046;
   wire n13047;
   wire n13048;
   wire n13049;
   wire n13050;
   wire n13051;
   wire n13052;
   wire n13053;
   wire n13054;
   wire n13055;
   wire n13056;
   wire n13057;
   wire n13058;
   wire n13059;
   wire n13060;
   wire n13061;
   wire n13062;
   wire n13063;
   wire n13064;
   wire n13065;
   wire n13066;
   wire n13067;
   wire n13068;
   wire n13069;
   wire n13070;
   wire n13071;
   wire n13072;
   wire n13073;
   wire n13074;
   wire n13075;
   wire n13076;
   wire n13077;
   wire n13078;
   wire n13079;
   wire n13080;
   wire n13081;
   wire n13082;
   wire n13083;
   wire n13084;
   wire n13085;
   wire n13086;
   wire n13087;
   wire n13088;
   wire n13089;
   wire n13090;
   wire n13091;
   wire n13092;
   wire n13093;
   wire n13094;
   wire n13095;
   wire n13096;
   wire n13097;
   wire n13098;
   wire n13099;
   wire n13100;
   wire n13101;
   wire n13102;
   wire n13103;
   wire n13104;
   wire n13105;
   wire n13106;
   wire n13107;
   wire n13108;
   wire n13109;
   wire n13110;
   wire n13111;
   wire n13112;
   wire n13113;
   wire n13114;
   wire n13115;
   wire n13116;
   wire n13117;
   wire n13118;
   wire n13119;
   wire n13120;
   wire n13121;
   wire n13122;
   wire n13123;
   wire n13124;
   wire n13125;
   wire n13126;
   wire n13127;
   wire n13128;
   wire n13129;
   wire n13130;
   wire n13131;
   wire n13132;
   wire n13133;
   wire n13134;
   wire n13135;
   wire n13136;
   wire n13137;
   wire n13138;
   wire n13139;
   wire n13140;
   wire n13141;
   wire n13142;
   wire n13143;
   wire n13144;
   wire n13145;
   wire n13146;
   wire n13147;
   wire n13148;
   wire n13149;
   wire n13150;
   wire n13151;
   wire n13152;
   wire n13153;
   wire n13154;
   wire n13155;
   wire n13156;
   wire n13157;
   wire n13158;
   wire n13159;
   wire n13160;
   wire n13161;
   wire n13162;
   wire n13163;
   wire n13164;
   wire n13165;
   wire n13166;
   wire n13167;
   wire n13168;
   wire n13169;
   wire n13170;
   wire n13171;
   wire n13172;
   wire n13173;
   wire n13174;
   wire n13175;
   wire n13176;
   wire n13177;
   wire n13178;
   wire n13179;
   wire n13180;
   wire n13181;
   wire n13182;
   wire n13183;
   wire n13184;
   wire n13185;
   wire n13186;
   wire n13187;
   wire n13188;
   wire n13189;
   wire n13190;
   wire n13191;
   wire n13192;
   wire n13193;
   wire n13194;
   wire n13195;
   wire n13196;
   wire n13197;
   wire n13198;
   wire n13199;
   wire n13200;
   wire n13201;
   wire n13202;
   wire n13203;
   wire n13204;
   wire n13205;
   wire n13206;
   wire n13207;
   wire n13208;
   wire n13209;
   wire n13210;
   wire n13211;
   wire n13212;
   wire n13213;
   wire n13214;
   wire n13215;
   wire n13216;
   wire n13217;
   wire n13218;
   wire n13219;
   wire n13220;
   wire n13221;
   wire n13222;
   wire n13223;
   wire n13224;
   wire n13225;
   wire n13226;
   wire n13227;
   wire n13228;
   wire n13229;
   wire n13230;
   wire n13231;
   wire n13232;
   wire n13233;
   wire n13234;
   wire n13235;
   wire n13236;
   wire n13237;
   wire n13238;
   wire n13239;
   wire n13240;
   wire n13241;
   wire n13242;
   wire n13243;
   wire n13244;
   wire n13245;
   wire n13246;
   wire n13247;
   wire n13248;
   wire n13249;
   wire n13250;
   wire n13251;
   wire n13252;
   wire n13253;
   wire n13254;
   wire n13255;
   wire n13256;
   wire n13257;
   wire n13258;
   wire n13259;
   wire n13260;
   wire n13261;
   wire n13262;
   wire n13263;
   wire n13264;
   wire n13265;
   wire n13266;
   wire n13267;
   wire n13268;
   wire n13269;
   wire n13270;
   wire n13271;
   wire n13272;
   wire n13273;
   wire n13274;
   wire n13275;
   wire n13276;
   wire n13277;
   wire n13278;
   wire n13279;
   wire n13280;
   wire n13281;
   wire n13282;
   wire n13283;
   wire n13284;
   wire n13285;
   wire n13286;
   wire n13287;
   wire n13288;
   wire n13289;
   wire n13290;
   wire n13291;
   wire n13292;
   wire n13293;
   wire n13294;
   wire n13295;
   wire n13296;
   wire n13297;
   wire n13298;
   wire n13299;
   wire n13300;
   wire n13301;
   wire n13302;
   wire n13303;
   wire n13304;
   wire n13305;
   wire n13306;
   wire n13307;
   wire n13308;
   wire n13309;
   wire n13310;
   wire n13311;
   wire n13312;
   wire n13313;
   wire n13314;
   wire n13315;
   wire n13316;
   wire n13317;
   wire n13318;
   wire n13319;
   wire n13320;
   wire n13321;
   wire n13322;
   wire n13323;
   wire n13324;
   wire n13325;
   wire n13326;
   wire n13327;
   wire n13328;
   wire n13329;
   wire n13330;
   wire n13331;
   wire n13332;
   wire n13333;
   wire n13334;
   wire n13335;
   wire n13336;
   wire n13337;
   wire n13338;
   wire n13339;
   wire n13340;
   wire n13341;
   wire n13342;
   wire n13343;
   wire n13344;
   wire n13345;
   wire n13346;
   wire n13347;
   wire n13348;
   wire n13349;
   wire n13350;
   wire n13351;
   wire n13352;
   wire n13353;
   wire n13354;
   wire n13355;
   wire n13356;
   wire n13357;
   wire n13358;
   wire n13359;
   wire n13360;
   wire n13361;
   wire n13362;
   wire n13363;
   wire n13364;
   wire n13365;
   wire n13366;
   wire n13367;
   wire n13368;
   wire n13369;
   wire n13370;
   wire n13371;
   wire n13372;
   wire n13373;
   wire n13374;
   wire n13375;
   wire n13376;
   wire n13377;
   wire n13378;
   wire n13379;
   wire n13380;
   wire n13381;
   wire n13382;
   wire n13383;
   wire n13384;
   wire n13385;
   wire n13386;
   wire n13387;
   wire n13388;
   wire n13389;
   wire n13390;
   wire n13391;
   wire n13392;
   wire n13393;
   wire n13394;
   wire n13395;
   wire n13396;
   wire n13397;
   wire n13398;
   wire n13399;
   wire n13400;
   wire n13401;
   wire n13402;
   wire n13403;
   wire n13404;
   wire n13405;
   wire n13406;
   wire n13407;
   wire n13408;
   wire n13409;
   wire n13410;
   wire n13411;
   wire n13412;
   wire n13413;
   wire n13414;
   wire n13415;
   wire n13416;
   wire n13417;
   wire n13418;
   wire n13419;
   wire n13420;
   wire n13421;
   wire n13422;
   wire n13423;
   wire n13424;
   wire n13425;
   wire n13426;
   wire n13427;
   wire n13428;
   wire n13429;
   wire n13430;
   wire n13431;
   wire n13432;
   wire n13433;
   wire n13434;
   wire n13435;
   wire n13436;
   wire n13437;
   wire n13438;
   wire n13439;
   wire n13440;
   wire n13441;
   wire n13442;
   wire n13443;
   wire n13444;
   wire n13445;
   wire n13446;
   wire n13447;
   wire n13448;
   wire n13449;
   wire n13450;
   wire n13451;
   wire n13452;
   wire n13453;
   wire n13454;
   wire n13455;
   wire n13456;
   wire n13457;
   wire n13458;
   wire n13459;
   wire n13460;
   wire n13461;
   wire n13462;
   wire n13463;
   wire n13464;
   wire n13465;
   wire n13466;
   wire n13467;
   wire n13468;
   wire n13469;
   wire n13470;
   wire n13471;
   wire n13472;
   wire n13473;
   wire n13474;
   wire n13475;
   wire n13476;
   wire n13477;
   wire n13478;
   wire n13479;
   wire n13480;
   wire n13481;
   wire n13482;
   wire n13483;
   wire n13484;
   wire n13485;
   wire n13486;
   wire n13487;
   wire n13488;
   wire n13489;
   wire n13490;
   wire n13491;
   wire n13492;
   wire n13493;
   wire n13494;
   wire n13495;
   wire n13496;
   wire n13497;
   wire n13498;
   wire n13499;
   wire n13500;
   wire n13501;
   wire n13502;
   wire n13503;
   wire n13504;
   wire n13505;
   wire n13506;
   wire n13507;
   wire n13508;
   wire n13509;
   wire n13510;
   wire n13511;
   wire n13514;
   wire n13515;
   wire n13516;
   wire n13517;
   wire n13518;
   wire n13519;
   wire n13520;
   wire n13521;
   wire n13522;
   wire n13523;
   wire n13524;
   wire n13525;
   wire n13526;
   wire n13527;
   wire n13528;
   wire n13529;
   wire n13530;
   wire n13531;
   wire n13532;
   wire n13533;
   wire n13534;
   wire n13535;
   wire n13536;
   wire n13537;
   wire n13538;
   wire n13539;
   wire n13540;
   wire n13541;
   wire n13542;
   wire n13543;
   wire n13544;
   wire n13545;
   wire n13546;
   wire n13547;
   wire n13548;
   wire n13549;
   wire n13550;
   wire n13551;
   wire n13552;
   wire n13553;
   wire n13554;
   wire n13555;
   wire n13556;
   wire n13557;
   wire n13558;
   wire n13559;
   wire n13560;
   wire n13561;
   wire n13562;
   wire n13563;
   wire n13564;
   wire n13565;
   wire n13566;
   wire n13567;
   wire n13568;
   wire n13569;
   wire n13570;
   wire n13571;
   wire n13572;
   wire n13573;
   wire n13574;
   wire n13575;
   wire n13576;
   wire n13577;
   wire n13578;
   wire n13579;
   wire n13580;
   wire n13581;
   wire n13582;
   wire n13583;
   wire n13584;
   wire n13585;
   wire n13586;
   wire n13587;
   wire n13588;
   wire n13589;
   wire n13590;
   wire n13591;
   wire n13592;
   wire n13593;
   wire n13594;
   wire n13595;
   wire n13596;
   wire n13597;
   wire n13599;
   wire n13600;
   wire n13601;
   wire n13602;
   wire n13603;
   wire n13604;
   wire n13605;
   wire n13606;
   wire n13607;
   wire n13608;
   wire n13609;
   wire n13610;
   wire n13611;
   wire n13612;
   wire n13613;
   wire n13614;
   wire n13615;
   wire n13616;
   wire n13617;
   wire n13618;
   wire n13619;
   wire n13620;
   wire n13621;
   wire n13622;
   wire n13623;
   wire n13624;
   wire n13625;
   wire n13626;
   wire n13627;
   wire n13628;
   wire n13629;
   wire n13630;
   wire n13631;
   wire n13632;
   wire n13633;
   wire n13634;
   wire n13635;
   wire n13636;
   wire n13637;
   wire n13638;
   wire n13639;
   wire n13640;
   wire n13641;
   wire n13642;
   wire n13643;
   wire n13644;
   wire n13645;
   wire n13646;
   wire n13647;
   wire n13648;
   wire n13649;
   wire n13650;
   wire n13651;
   wire n13652;
   wire n13653;
   wire n13654;
   wire n13655;
   wire n13656;
   wire n13657;
   wire n13658;
   wire n13659;
   wire n13660;
   wire n13661;
   wire n13662;
   wire n13663;
   wire n13664;
   wire n13665;
   wire n13666;
   wire n13667;
   wire n13668;
   wire n13669;
   wire n13670;
   wire n13671;
   wire n13672;
   wire n13673;
   wire n13674;
   wire n13675;
   wire n13676;
   wire n13677;
   wire n13678;
   wire n13679;
   wire n13680;
   wire n13681;
   wire n13682;
   wire n13683;
   wire n13684;
   wire n13685;
   wire n13686;
   wire n13687;
   wire n13688;
   wire n13689;
   wire n13690;
   wire n13691;
   wire n13692;
   wire n13693;
   wire n13694;
   wire n13695;
   wire n13696;
   wire n13697;
   wire n13698;
   wire n13699;
   wire n13700;
   wire n13701;
   wire n13702;
   wire n13703;
   wire n13704;
   wire n13705;
   wire n13706;
   wire n13707;
   wire n13708;
   wire n13709;
   wire n13710;
   wire n13711;
   wire n13712;
   wire n13713;
   wire n13714;
   wire n13715;
   wire n13716;
   wire n13717;
   wire n13718;
   wire n13719;
   wire n13720;
   wire n13721;
   wire n13722;
   wire n13723;
   wire n13724;
   wire n13725;
   wire n13726;
   wire n13727;
   wire n13728;
   wire n13729;
   wire n13730;
   wire n13731;
   wire n13732;
   wire n13733;
   wire n13734;
   wire n13735;
   wire n13736;
   wire n13737;
   wire n13738;
   wire n13739;
   wire n13740;
   wire n13741;
   wire n13742;
   wire n13743;
   wire n13744;
   wire n13745;
   wire n13746;
   wire n13747;
   wire n13748;
   wire n13749;
   wire n13750;
   wire n13751;
   wire n13752;
   wire n13753;
   wire n13754;
   wire n13755;
   wire n13756;
   wire n13757;
   wire n13758;
   wire n13759;
   wire n13760;
   wire n13761;
   wire n13762;
   wire n13763;
   wire n13764;
   wire n13765;
   wire n13766;
   wire n13767;
   wire n13768;
   wire n13769;
   wire n13770;
   wire n13771;
   wire n13772;
   wire n13773;
   wire n13774;
   wire n13775;
   wire n13776;
   wire n13777;
   wire n13778;
   wire n13779;
   wire n13780;
   wire n13781;
   wire n13782;
   wire n13783;
   wire n13784;
   wire n13785;
   wire n13786;
   wire n13787;
   wire n13788;
   wire n13789;
   wire n13790;
   wire n13791;
   wire n13792;
   wire n13793;
   wire n13794;
   wire n13795;
   wire n13796;
   wire n13797;
   wire n13798;
   wire n13799;
   wire n13800;
   wire n13801;
   wire n13802;
   wire n13803;
   wire n13804;
   wire n13805;
   wire n13806;
   wire n13807;
   wire n13808;
   wire n13809;
   wire n13810;
   wire n13811;
   wire n13812;
   wire n13813;
   wire n13814;
   wire n13815;
   wire n13816;
   wire n13817;
   wire n13818;
   wire n13819;
   wire n13820;
   wire n13821;
   wire n13822;
   wire n13823;
   wire n13824;
   wire n13825;
   wire n13826;
   wire n13827;
   wire n13828;
   wire n13829;
   wire n13830;
   wire n13831;
   wire n13832;
   wire n13833;
   wire n13834;
   wire n13835;
   wire n13836;
   wire n13837;
   wire n13838;
   wire n13839;
   wire n13840;
   wire n13841;
   wire n13842;
   wire n13843;
   wire n13844;
   wire n13845;
   wire n13846;
   wire n13847;
   wire n13848;
   wire n13849;
   wire n13850;
   wire n13851;
   wire n13852;
   wire n13853;
   wire n13854;
   wire n13855;
   wire n13856;
   wire n13857;
   wire n13858;
   wire n13859;
   wire n13860;
   wire n13861;
   wire n13862;
   wire n13863;
   wire n13864;
   wire n13865;
   wire n13866;
   wire n13867;
   wire n13868;
   wire n13869;
   wire n13870;
   wire n13871;
   wire n13872;
   wire n13873;
   wire n13874;
   wire n13875;
   wire n13876;
   wire n13877;
   wire n13878;
   wire n13879;
   wire n13880;
   wire n13881;
   wire n13882;
   wire n13883;
   wire n13884;
   wire n13885;
   wire n13886;
   wire n13887;
   wire n13888;
   wire n13889;
   wire n13890;
   wire n13891;
   wire n13892;
   wire n13893;
   wire n13894;
   wire n13895;
   wire n13896;
   wire n13897;
   wire n13898;
   wire n13899;
   wire n13900;
   wire n13901;
   wire n13902;
   wire n13903;
   wire n13904;
   wire n13905;
   wire n13906;
   wire n13907;
   wire n13908;
   wire n13909;
   wire n13910;
   wire n13911;
   wire n13912;
   wire n13913;
   wire n13914;
   wire n13915;
   wire n13916;
   wire n13917;
   wire n13918;
   wire n13919;
   wire n13920;
   wire n13921;
   wire n13922;
   wire n13923;
   wire n13924;
   wire n13925;
   wire n13926;
   wire n13927;
   wire n13928;
   wire n13929;
   wire n13930;
   wire n13931;
   wire n13932;
   wire n13933;
   wire n13934;
   wire n13935;
   wire n13936;
   wire n13937;
   wire n13938;
   wire n13939;
   wire n13940;
   wire n13941;
   wire n13942;
   wire n13943;
   wire n13944;
   wire n13945;
   wire n13946;
   wire n13947;
   wire n13948;
   wire n13949;
   wire n13950;
   wire n13951;
   wire n13952;
   wire n13953;
   wire n13954;
   wire n13955;
   wire n13956;
   wire n13957;
   wire n13958;
   wire n13959;
   wire n13960;
   wire n13961;
   wire n13962;
   wire n13963;
   wire n13964;
   wire n13965;
   wire n13966;
   wire n13967;
   wire n13968;
   wire n13969;
   wire n13970;
   wire n13971;
   wire n13972;
   wire n13973;
   wire n13974;
   wire n13975;
   wire n13976;
   wire n13977;
   wire n13978;
   wire n13979;
   wire n13980;
   wire n13981;
   wire n13982;
   wire n13983;
   wire n13984;
   wire n13985;
   wire n13986;
   wire n13987;
   wire n13988;
   wire n13989;
   wire n13990;
   wire n13991;
   wire n13992;
   wire n13993;
   wire n13994;
   wire n13995;
   wire n13996;
   wire n13997;
   wire n13998;
   wire n13999;
   wire n14000;
   wire n14001;
   wire n14002;
   wire n14003;
   wire n14004;
   wire n14005;
   wire n14006;
   wire n14007;
   wire n14008;
   wire n14009;
   wire n14011;
   wire n14012;
   wire n14013;
   wire n14014;
   wire n14015;
   wire n14016;
   wire n14017;
   wire n14018;
   wire n14019;
   wire n14020;
   wire n14021;
   wire n14022;
   wire n14023;
   wire n14024;
   wire n14025;
   wire n14026;
   wire n14027;
   wire n14028;
   wire n14029;
   wire n14030;
   wire n14031;
   wire n14032;
   wire n14033;
   wire n14034;
   wire n14035;
   wire n14036;
   wire n14037;
   wire n14038;
   wire n14039;
   wire n14040;
   wire n14041;
   wire n14042;
   wire n14043;
   wire n14044;
   wire n14045;
   wire n14046;
   wire n14047;
   wire n14048;
   wire n14049;
   wire n14050;
   wire n14051;
   wire n14052;
   wire n14053;
   wire n14054;
   wire n14055;
   wire n14056;
   wire n14057;
   wire n14058;
   wire n14059;
   wire n14060;
   wire n14061;
   wire n14062;
   wire n14063;
   wire n14064;
   wire n14065;
   wire n14066;
   wire n14067;
   wire n14068;
   wire n14069;
   wire n14070;
   wire n14071;
   wire n14072;
   wire n14073;
   wire n14074;
   wire n14075;
   wire n14076;
   wire n14077;
   wire n14078;
   wire n14079;
   wire n14080;
   wire n14081;
   wire n14082;
   wire n14083;
   wire n14084;
   wire n14085;
   wire n14086;
   wire n14087;
   wire n14088;
   wire n14089;
   wire n14090;
   wire n14091;
   wire n14092;
   wire n14093;
   wire n14094;
   wire n14095;
   wire n14096;
   wire n14097;
   wire n14098;
   wire n14099;
   wire n14100;
   wire n14101;
   wire n14102;
   wire n14103;
   wire n14104;
   wire n14105;
   wire n14106;
   wire n14107;
   wire n14108;
   wire n14109;
   wire n14110;
   wire n14111;
   wire n14112;
   wire n14113;
   wire n14114;
   wire n14115;
   wire n14116;
   wire n14117;
   wire n14118;
   wire n14119;
   wire n14120;
   wire n14121;
   wire n14122;
   wire n14123;
   wire n14124;
   wire n14125;
   wire n14126;
   wire n14127;
   wire n14128;
   wire n14129;
   wire n14130;
   wire n14131;
   wire n14132;
   wire n14133;
   wire n14134;
   wire n14135;
   wire n14136;
   wire n14137;
   wire n14138;
   wire n14140;
   wire n14141;
   wire n14142;
   wire n14143;
   wire n14144;
   wire n14145;
   wire n14146;
   wire n14147;
   wire n14148;
   wire n14149;
   wire n14150;
   wire n14151;
   wire n14152;
   wire n14153;
   wire n14154;
   wire n14155;
   wire n14156;
   wire n14157;
   wire n14158;
   wire n14159;
   wire n14160;
   wire n14161;
   wire n14162;
   wire n14163;
   wire n14164;
   wire n14165;
   wire n14166;
   wire n14167;
   wire n14168;
   wire n14169;
   wire n14170;
   wire n14171;
   wire n14172;
   wire n14173;
   wire n14174;
   wire n14175;
   wire n14176;
   wire n14177;
   wire n14178;
   wire n14179;
   wire n14180;
   wire n14181;
   wire n14182;
   wire n14183;
   wire n14184;
   wire n14185;
   wire n14186;
   wire n14187;
   wire n14188;
   wire n14189;
   wire n14190;
   wire n14191;
   wire n14192;
   wire n14193;
   wire n14194;
   wire n14195;
   wire n14196;
   wire n14197;
   wire n14198;
   wire n14199;
   wire n14200;
   wire n14201;
   wire n14202;
   wire n14203;
   wire n14204;
   wire n14205;
   wire n14206;
   wire n14207;
   wire n14208;
   wire n14209;
   wire n14210;
   wire n14211;
   wire n14212;
   wire n14213;
   wire n14214;
   wire n14215;
   wire n14216;
   wire n14217;
   wire n14218;
   wire n14219;
   wire n14220;
   wire n14221;
   wire n14222;
   wire n14223;
   wire n14224;
   wire n14225;
   wire n14226;
   wire n14227;
   wire n14228;
   wire n14229;
   wire n14230;
   wire n14231;
   wire n14232;
   wire n14233;
   wire n14234;
   wire n14235;
   wire n14236;
   wire n14237;
   wire n14238;
   wire n14239;
   wire n14240;
   wire n14241;
   wire n14242;
   wire n14243;
   wire n14244;
   wire n14245;
   wire n14246;
   wire n14247;
   wire n14248;
   wire n14249;
   wire n14250;
   wire n14251;
   wire n14252;
   wire n14253;
   wire n14254;
   wire n14255;
   wire n14256;
   wire n14257;
   wire n14258;
   wire n14259;
   wire n14260;
   wire n14261;
   wire n14262;
   wire n14263;
   wire n14264;
   wire n14265;
   wire n14266;
   wire n14267;
   wire n14268;
   wire n14269;
   wire n14270;
   wire n14271;
   wire n14272;
   wire n14273;
   wire n14274;
   wire n14275;
   wire n14276;
   wire n14277;
   wire n14278;
   wire n14279;
   wire n14280;
   wire n14281;
   wire n14282;
   wire n14283;
   wire n14284;
   wire n14285;
   wire n14286;
   wire n14287;
   wire n14288;
   wire n14289;
   wire n14290;
   wire n14291;
   wire n14292;
   wire n14293;
   wire n14294;
   wire n14295;
   wire n14296;
   wire n14297;
   wire n14298;
   wire n14299;
   wire n14300;
   wire n14301;
   wire n14302;
   wire n14303;
   wire n14304;
   wire n14305;
   wire n14306;
   wire n14307;
   wire n14308;
   wire n14309;
   wire n14310;
   wire n14311;
   wire n14312;
   wire n14313;
   wire n14314;
   wire n14315;
   wire n14316;
   wire n14317;
   wire n14318;
   wire n14319;
   wire n14320;
   wire n14321;
   wire n14322;
   wire n14323;
   wire n14324;
   wire n14325;
   wire n14326;
   wire n14327;
   wire n14328;
   wire n14329;
   wire n14330;
   wire n14331;
   wire n14332;
   wire n14333;
   wire n14334;
   wire n14335;
   wire n14336;
   wire n14337;
   wire n14338;
   wire n14339;
   wire n14340;
   wire n14341;
   wire n14342;
   wire n14343;
   wire n14344;
   wire n14345;
   wire n14346;
   wire n14348;
   wire n14349;
   wire n14350;
   wire n14351;
   wire n14352;
   wire n14353;
   wire n14354;
   wire n14355;
   wire n14356;
   wire n14357;
   wire n14358;
   wire n14359;
   wire n14360;
   wire n14361;
   wire n14362;
   wire n14363;
   wire n14364;
   wire n14365;
   wire n14366;
   wire n14367;
   wire n14368;
   wire n14369;
   wire n14370;
   wire n14371;
   wire n14372;
   wire n14373;
   wire n14374;
   wire n14375;
   wire n14376;
   wire n14377;
   wire n14378;
   wire n14379;
   wire n14380;
   wire n14381;
   wire n14382;
   wire n14383;
   wire n14384;
   wire n14385;
   wire n14386;
   wire n14387;
   wire n14388;
   wire n14389;
   wire n14390;
   wire n14391;
   wire n14392;
   wire n14393;
   wire n14394;
   wire n14395;
   wire n14396;
   wire n14397;
   wire n14398;
   wire n14399;
   wire n14400;
   wire n14401;
   wire n14402;
   wire n14403;
   wire n14404;
   wire n14405;
   wire n14406;
   wire n14407;
   wire n14408;
   wire n14409;
   wire n14410;
   wire n14411;
   wire n14412;
   wire n14413;
   wire n14414;
   wire n14415;
   wire n14416;
   wire n14417;
   wire n14418;
   wire n14419;
   wire n14420;
   wire n14421;
   wire n14422;
   wire n14423;
   wire n14424;
   wire n14425;
   wire n14426;
   wire n14427;
   wire n14428;
   wire n14429;
   wire n14430;
   wire n14431;
   wire n14432;
   wire n14433;
   wire n14434;
   wire n14435;
   wire n14436;
   wire n14437;
   wire n14438;
   wire n14439;
   wire n14440;
   wire n14441;
   wire n14442;
   wire n14443;
   wire n14444;
   wire n14445;
   wire n14446;
   wire n14447;
   wire n14448;
   wire n14449;
   wire n14450;
   wire n14451;
   wire n14452;
   wire n14453;
   wire n14454;
   wire n14455;
   wire n14456;
   wire n14457;
   wire n14458;
   wire n14459;
   wire n14460;
   wire n14461;
   wire n14462;
   wire n14463;
   wire n14464;
   wire n14465;
   wire n14466;
   wire n14467;
   wire n14468;
   wire n14469;
   wire n14470;
   wire n14471;
   wire n14472;
   wire n14473;
   wire n14474;
   wire n14475;
   wire n14476;
   wire n14477;
   wire n14478;
   wire n14479;
   wire n14480;
   wire n14481;
   wire n14482;
   wire n14483;
   wire n14484;
   wire n14485;
   wire n14486;
   wire n14487;
   wire n14488;
   wire n14489;
   wire n14490;
   wire n14491;
   wire n14492;
   wire n14493;
   wire n14494;
   wire n14495;
   wire n14496;
   wire n14497;
   wire n14498;
   wire n14499;
   wire n14500;
   wire n14501;
   wire n14502;
   wire n14503;
   wire n14504;
   wire n14505;
   wire n14506;
   wire n14507;
   wire n14508;
   wire n14509;
   wire n14510;
   wire n14511;
   wire n14512;
   wire n14513;
   wire n14514;
   wire n14515;
   wire n14516;
   wire n14517;
   wire n14518;
   wire n14520;
   wire n14522;
   wire n14523;
   wire n14524;
   wire n14525;
   wire n14526;
   wire n14527;
   wire n14528;
   wire n14529;
   wire n14530;
   wire n14531;
   wire n14532;
   wire n14533;
   wire n14534;
   wire n14535;
   wire n14536;
   wire n14537;
   wire n14538;
   wire n14539;
   wire n14540;
   wire n14541;
   wire n14542;
   wire n14543;
   wire n14544;
   wire n14545;
   wire n14546;
   wire n14547;
   wire n14548;
   wire n14549;
   wire n14550;
   wire n14551;
   wire n14552;
   wire n14553;
   wire n14554;
   wire n14555;
   wire n14556;
   wire n14557;
   wire n14558;
   wire n14559;
   wire n14560;
   wire n14561;
   wire n14562;
   wire n14563;
   wire n14564;
   wire n14565;
   wire n14566;
   wire n14567;
   wire n14568;
   wire n14569;
   wire n14570;
   wire n14571;
   wire n14572;
   wire n14573;
   wire n14574;
   wire n14575;
   wire n14576;
   wire n14577;
   wire n14578;
   wire n14579;
   wire n14580;
   wire n14581;
   wire n14582;
   wire n14583;
   wire n14584;
   wire n14585;
   wire n14586;
   wire n14587;
   wire n14588;
   wire n14589;
   wire n14590;
   wire n14591;
   wire n14592;
   wire n14593;
   wire n14595;
   wire n14596;
   wire n14597;
   wire n14598;
   wire n14599;
   wire n14600;
   wire n14601;
   wire n14602;
   wire n14603;
   wire n14604;
   wire n14605;
   wire n14606;
   wire n14607;
   wire n14608;
   wire n14609;
   wire n14610;
   wire n14611;
   wire n14612;
   wire n14613;
   wire n14614;
   wire n14615;
   wire n14616;
   wire n14617;
   wire n14618;
   wire n14619;
   wire n14620;
   wire n14621;
   wire n14622;
   wire n14623;
   wire n14624;
   wire n14625;
   wire n14626;
   wire n14627;
   wire n14628;
   wire n14629;
   wire n14630;
   wire n14631;
   wire n14632;
   wire n14633;
   wire n14634;
   wire n14635;
   wire n14636;
   wire n14637;
   wire n14638;
   wire n14639;
   wire n14640;
   wire n14641;
   wire n14642;
   wire n14643;
   wire n14644;
   wire n14645;
   wire n14646;
   wire n14647;
   wire n14648;
   wire n14649;
   wire n14650;
   wire n14651;
   wire n14652;
   wire n14653;
   wire n14654;
   wire n14655;
   wire n14656;
   wire n14657;
   wire n14658;
   wire n14659;
   wire n14660;
   wire n14661;
   wire n14662;
   wire n14663;
   wire n14664;
   wire n14665;
   wire n14666;
   wire n14667;
   wire n14668;
   wire n14669;
   wire n14670;
   wire n14671;
   wire n14672;
   wire n14673;
   wire n14674;
   wire n14675;
   wire n14676;
   wire n14677;
   wire n14678;
   wire n14679;
   wire n14680;
   wire n14681;
   wire n14682;
   wire n14683;
   wire n14684;
   wire n14685;
   wire n14686;
   wire n14687;
   wire n14688;
   wire n14689;
   wire n14690;
   wire n14691;
   wire n14692;
   wire n14693;
   wire n14694;
   wire n14695;
   wire n14696;
   wire n14697;
   wire n14698;
   wire n14699;
   wire n14700;
   wire n14701;
   wire n14702;
   wire n14703;
   wire n14704;
   wire n14705;
   wire n14706;
   wire n14707;
   wire n14708;
   wire n14709;
   wire n14710;
   wire n14711;
   wire n14712;
   wire n14713;
   wire n14714;
   wire n14715;
   wire n14716;
   wire n14717;
   wire n14718;
   wire n14719;
   wire n14720;
   wire n14721;
   wire n14722;
   wire n14723;
   wire n14724;
   wire n14725;
   wire n14726;
   wire n14727;
   wire n14728;
   wire n14729;
   wire n14730;
   wire n14731;
   wire n14732;
   wire n14733;
   wire n14734;
   wire n14735;
   wire n14736;
   wire n14737;
   wire n14738;
   wire n14739;
   wire n14740;
   wire n14741;
   wire n14742;
   wire n14743;
   wire n14744;
   wire n14745;
   wire n14746;
   wire n14747;
   wire n14748;
   wire n14749;
   wire n14750;
   wire n14751;
   wire n14752;
   wire n14753;
   wire n14754;
   wire n14755;
   wire n14756;
   wire n14757;
   wire n14758;
   wire n14759;
   wire n14760;
   wire n14761;
   wire n14762;
   wire n14763;
   wire n14764;
   wire n14765;
   wire n14766;
   wire n14767;
   wire n14768;
   wire n14769;
   wire n14770;
   wire n14771;
   wire n14772;
   wire n14773;
   wire n14774;
   wire n14775;
   wire n14776;
   wire n14777;
   wire n14778;
   wire n14779;
   wire n14780;
   wire n14781;
   wire n14782;
   wire n14783;
   wire n14784;
   wire n14785;
   wire n14786;
   wire n14787;
   wire n14788;
   wire n14789;
   wire n14790;
   wire n14791;
   wire n14792;
   wire n14793;
   wire n14794;
   wire n14795;
   wire n14796;
   wire n14797;
   wire n14798;
   wire n14799;
   wire n14800;
   wire n14801;
   wire n14802;
   wire n14803;
   wire n14804;
   wire n14805;
   wire n14806;
   wire n14807;
   wire n14808;
   wire n14809;
   wire n14810;
   wire n14811;
   wire n14812;
   wire n14813;
   wire n14814;
   wire n14815;
   wire n14816;
   wire n14817;
   wire n14818;
   wire n14819;
   wire n14820;
   wire n14821;
   wire n14822;
   wire n14823;
   wire n14824;
   wire n14826;
   wire n14827;
   wire n14829;
   wire n14830;
   wire n14831;
   wire n14832;
   wire n14833;
   wire n14834;
   wire n14835;
   wire n14836;
   wire n14837;
   wire n14838;
   wire n14839;
   wire n14840;
   wire n14841;
   wire n14842;
   wire n14843;
   wire n14844;
   wire n14845;
   wire n14846;
   wire n14847;
   wire n14848;
   wire n14849;
   wire n14850;
   wire n14851;
   wire n14852;
   wire n14853;
   wire n14854;
   wire n14855;
   wire n14856;
   wire n14857;
   wire n14858;
   wire n14859;
   wire n14860;
   wire n14861;
   wire n14862;
   wire n14863;
   wire n14864;
   wire n14865;
   wire n14866;
   wire n14867;
   wire n14868;
   wire n14869;
   wire n14870;
   wire n14871;
   wire n14872;
   wire n14873;
   wire n14874;
   wire n14875;
   wire n14876;
   wire n14877;
   wire n14878;
   wire n14879;
   wire n14880;
   wire n14881;
   wire n14882;
   wire n14883;
   wire n14884;
   wire n14885;
   wire n14886;
   wire n14887;
   wire n14888;
   wire n14889;
   wire n14890;
   wire n14891;
   wire n14892;
   wire n14893;
   wire n14894;
   wire n14895;
   wire n14896;
   wire n14897;
   wire n14898;
   wire n14899;
   wire n14900;
   wire n14901;
   wire n14902;
   wire n14903;
   wire n14904;
   wire n14905;
   wire n14906;
   wire n14907;
   wire n14908;
   wire n14909;
   wire n14910;
   wire n14911;
   wire n14912;
   wire n14913;
   wire n14914;
   wire n14915;
   wire n14916;
   wire n14917;
   wire n14918;
   wire n14919;
   wire n14920;
   wire n14921;
   wire n14922;
   wire n14923;
   wire n14924;
   wire n14925;
   wire n14926;
   wire n14927;
   wire n14928;
   wire n14929;
   wire n14930;
   wire n14931;
   wire n14932;
   wire n14933;
   wire n14934;
   wire n14935;
   wire n14936;
   wire n14937;
   wire n14938;
   wire n14939;
   wire n14940;
   wire n14941;
   wire n14942;
   wire n14943;
   wire n14944;
   wire n14945;
   wire n14946;
   wire n14947;
   wire n14948;
   wire n14949;
   wire n14950;
   wire n14951;
   wire n14952;
   wire n14953;
   wire n14954;
   wire n14955;
   wire n14956;
   wire n14957;
   wire n14958;
   wire n14959;
   wire n14960;
   wire n14961;
   wire n14962;
   wire n14963;
   wire n14964;
   wire n14965;
   wire n14966;
   wire n14967;
   wire n14968;
   wire n14969;
   wire n14970;
   wire n14971;
   wire n14972;
   wire n14973;
   wire n14974;
   wire n14975;
   wire n14976;
   wire n14977;
   wire n14978;
   wire n14979;
   wire n14980;
   wire n14981;
   wire n14982;
   wire n14983;
   wire n14984;
   wire n14985;
   wire n14986;
   wire n14987;
   wire n14988;
   wire n14989;
   wire n14990;
   wire n14991;
   wire n14992;
   wire n14993;
   wire n14994;
   wire n14995;
   wire n14996;
   wire n14997;
   wire n14998;
   wire n14999;
   wire n15000;
   wire n15001;
   wire n15002;
   wire n15003;
   wire n15004;
   wire n15005;
   wire n15006;
   wire n15007;
   wire n15008;
   wire n15009;
   wire n15010;
   wire n15011;
   wire n15012;
   wire n15013;
   wire n15014;
   wire n15015;
   wire n15016;
   wire n15017;
   wire n15018;
   wire n15019;
   wire n15020;
   wire n15021;
   wire n15022;
   wire n15023;
   wire n15024;
   wire n15025;
   wire n15026;
   wire n15027;
   wire n15028;
   wire n15029;
   wire n15030;
   wire n15031;
   wire n15032;
   wire n15033;
   wire n15034;
   wire n15035;
   wire n15036;
   wire n15037;
   wire n15038;
   wire n15039;
   wire n15040;
   wire n15041;
   wire n15042;
   wire n15043;
   wire n15044;
   wire n15045;
   wire n15046;
   wire n15047;
   wire n15048;
   wire n15049;
   wire n15050;
   wire n15051;
   wire n15052;
   wire n15053;
   wire n15054;
   wire n15056;
   wire n15057;
   wire n15058;
   wire n15059;
   wire n15060;
   wire n15061;
   wire n15062;
   wire n15063;
   wire n15064;
   wire n15065;
   wire n15066;
   wire n15067;
   wire n15068;
   wire n15069;
   wire n15070;
   wire n15071;
   wire n15072;
   wire n15073;
   wire n15074;
   wire n15075;
   wire n15076;
   wire n15077;
   wire n15078;
   wire n15079;
   wire n15080;
   wire n15081;
   wire n15082;
   wire n15083;
   wire n15084;
   wire n15085;
   wire n15086;
   wire n15087;
   wire n15088;
   wire n15089;
   wire n15090;
   wire n15091;
   wire n15092;
   wire n15093;
   wire n15094;
   wire n15095;
   wire n15096;
   wire n15097;
   wire n15098;
   wire n15099;
   wire n15100;
   wire n15101;
   wire n15102;
   wire n15103;
   wire n15104;
   wire n15105;
   wire n15107;
   wire n15108;
   wire n15109;
   wire n15110;
   wire n15111;
   wire n15112;
   wire n15113;
   wire n15114;
   wire n15115;
   wire n15116;
   wire n15117;
   wire n15118;
   wire n15119;
   wire n15120;
   wire n15121;
   wire n15122;
   wire n15123;
   wire n15124;
   wire n15125;
   wire n15126;
   wire n15127;
   wire n15128;
   wire n15129;
   wire n15130;
   wire n15131;
   wire n15132;
   wire n15133;
   wire n15134;
   wire n15135;
   wire n15136;
   wire n15137;
   wire n15138;
   wire n15139;
   wire n15140;
   wire n15141;
   wire n15142;
   wire n15143;
   wire n15145;
   wire n15146;
   wire n15148;
   wire n15149;
   wire n15150;
   wire n15151;
   wire n15152;
   wire n15153;
   wire n15154;
   wire n15155;
   wire n15156;
   wire n15157;
   wire n15158;
   wire n15159;
   wire n15160;
   wire n15161;
   wire n15162;
   wire n15163;
   wire n15164;
   wire n15165;
   wire n15166;
   wire n15167;
   wire n15168;
   wire n15169;
   wire n15170;
   wire n15171;
   wire n15172;
   wire n15173;
   wire n15174;
   wire n15175;
   wire n15176;
   wire n15177;
   wire n15178;
   wire n15179;
   wire n15180;
   wire n15181;
   wire n15182;
   wire n15183;
   wire n15184;
   wire n15185;
   wire n15186;
   wire n15187;
   wire n15188;
   wire n15189;
   wire n15190;
   wire n15191;
   wire n15192;
   wire n15193;
   wire n15194;
   wire n15195;
   wire n15196;
   wire n15197;
   wire n15198;
   wire n15199;
   wire n15200;
   wire n15201;
   wire n15202;
   wire n15203;
   wire n15205;
   wire n15206;
   wire n15207;
   wire n15208;
   wire n15209;
   wire n15210;
   wire n15211;
   wire n15212;
   wire n15213;
   wire n15215;
   wire n15216;
   wire n15217;
   wire n15218;
   wire n15219;
   wire n15220;
   wire n15221;
   wire n15222;
   wire n15223;
   wire n15224;
   wire n15225;
   wire n15226;
   wire n15228;
   wire n15229;
   wire n15230;
   wire n15231;
   wire n15232;
   wire n15233;
   wire n15234;
   wire n15235;
   wire n15236;
   wire n15237;
   wire n15238;
   wire n15239;
   wire n15240;
   wire n15241;
   wire n15242;
   wire n15243;
   wire n15244;
   wire n15245;
   wire n15246;
   wire n15247;
   wire n15248;
   wire n15249;
   wire n15250;
   wire n15251;
   wire n15252;
   wire n15253;
   wire n15254;
   wire n15255;
   wire n15256;
   wire n15257;
   wire n15258;
   wire n15259;
   wire n15260;
   wire n15261;
   wire n15262;
   wire n15263;
   wire n15264;
   wire n15265;
   wire n15266;
   wire n15267;
   wire n15268;
   wire n15269;
   wire n15270;
   wire n15271;
   wire n15272;
   wire n15273;
   wire n15274;
   wire n15275;
   wire n15276;
   wire n15277;
   wire n15278;
   wire n15279;
   wire n15280;
   wire n15281;
   wire n15282;
   wire n15283;
   wire n15284;
   wire n15285;
   wire n15286;
   wire n15287;
   wire n15288;
   wire n15289;
   wire n15290;
   wire n15291;
   wire n15292;
   wire n15293;
   wire n15294;
   wire n15295;
   wire n15296;
   wire n15297;
   wire n15298;
   wire n15299;
   wire n15300;
   wire n15301;
   wire n15302;
   wire n15303;
   wire n15304;
   wire n15305;
   wire n15306;
   wire n15307;
   wire n15308;
   wire n15309;
   wire n15310;
   wire n15311;
   wire n15312;
   wire n15313;
   wire n15314;
   wire n15315;
   wire n15316;
   wire n15317;
   wire n15318;
   wire n15319;
   wire n15320;
   wire n15321;
   wire n15322;
   wire n15323;
   wire n15324;
   wire n15325;
   wire n15326;
   wire n15327;
   wire n15329;
   wire n15330;
   wire n15331;
   wire n15332;
   wire n15333;
   wire n15334;
   wire n15335;
   wire n15336;
   wire n15337;
   wire n15338;
   wire n15339;
   wire n15340;
   wire n15341;
   wire n15342;
   wire n15343;
   wire n15344;
   wire n15345;
   wire n15346;
   wire n15347;
   wire n15348;
   wire n15349;
   wire n15350;
   wire n15351;
   wire n15352;
   wire n15353;
   wire n15354;
   wire n15355;
   wire n15356;
   wire n15357;
   wire n15358;
   wire n15359;
   wire n15360;
   wire n15361;
   wire n15362;
   wire n15363;
   wire n15364;
   wire n15365;
   wire n15366;
   wire n15367;
   wire n15368;
   wire n15369;
   wire n15370;
   wire n15371;
   wire n15372;
   wire n15373;
   wire n15374;
   wire n15375;
   wire n15376;
   wire n15377;
   wire n15378;
   wire n15379;
   wire n15380;
   wire n15381;
   wire n15382;
   wire n15383;
   wire n15384;
   wire n15385;
   wire n15386;
   wire n15387;
   wire n15388;
   wire n15389;
   wire n15390;
   wire n15391;
   wire n15392;
   wire n15393;
   wire n15394;
   wire n15395;
   wire n15396;
   wire n15397;
   wire n15398;
   wire n15399;
   wire n15400;
   wire n15401;
   wire n15402;
   wire n15403;
   wire n15404;
   wire n15405;
   wire n15406;
   wire n15407;
   wire n15408;
   wire n15409;
   wire n15410;
   wire n15411;
   wire n15412;
   wire n15413;
   wire n15414;
   wire n15415;
   wire n15416;
   wire n15417;
   wire n15418;
   wire n15419;
   wire n15420;
   wire n15421;
   wire n15422;
   wire n15423;
   wire n15424;
   wire n15425;
   wire n15426;
   wire n15427;
   wire n15428;
   wire n15429;
   wire n15430;
   wire n15431;
   wire n15432;
   wire n15433;
   wire n15434;
   wire n15435;
   wire n15436;
   wire n15437;
   wire n15438;
   wire n15439;
   wire n15440;
   wire n15441;
   wire n15442;
   wire n15443;
   wire n15444;
   wire n15445;
   wire n15446;
   wire n15447;
   wire n15448;
   wire n15449;
   wire n15450;
   wire n15451;
   wire n15452;
   wire n15453;
   wire n15454;
   wire n15455;
   wire n15456;
   wire n15457;
   wire n15458;
   wire n15459;
   wire n15460;
   wire n15461;
   wire n15462;
   wire n15463;
   wire n15464;
   wire n15465;
   wire n15466;
   wire n15467;
   wire n15468;
   wire n15469;
   wire n15470;
   wire n15471;
   wire n15472;
   wire n15473;
   wire n15474;
   wire n15475;
   wire n15476;
   wire n15477;
   wire n15478;
   wire n15479;
   wire n15480;
   wire n15481;
   wire n15482;
   wire n15483;
   wire n15484;
   wire n15485;
   wire n15486;
   wire n15487;
   wire n15488;
   wire n15489;
   wire n15490;
   wire n15491;
   wire n15492;
   wire n15493;
   wire n15494;
   wire n15495;
   wire n15496;
   wire n15497;
   wire n15498;
   wire n15499;
   wire n15500;
   wire n15501;
   wire n15502;
   wire n15503;
   wire n15504;
   wire n15505;
   wire n15506;
   wire n15507;
   wire n15508;
   wire n15509;
   wire n15510;
   wire n15511;
   wire n15512;
   wire n15513;
   wire n15514;
   wire n15515;
   wire n15516;
   wire n15517;
   wire n15518;
   wire n15519;
   wire n15520;
   wire n15521;
   wire n15522;
   wire n15523;
   wire n15524;
   wire n15525;
   wire n15526;
   wire n15527;
   wire n15528;
   wire n15529;
   wire n15530;
   wire n15531;
   wire n15532;
   wire n15533;
   wire n15534;
   wire n15536;
   wire n15537;
   wire n15538;
   wire n15539;
   wire n15540;
   wire n15541;
   wire n15542;
   wire n15543;
   wire n15544;
   wire n15545;
   wire n15546;
   wire n15547;
   wire n15548;
   wire n15549;
   wire n15550;
   wire n15551;
   wire n15552;
   wire n15553;
   wire n15554;
   wire n15555;
   wire n15556;
   wire n15557;
   wire n15558;
   wire n15559;
   wire n15560;
   wire n15561;
   wire n15562;
   wire n15563;
   wire n15564;
   wire n15565;
   wire n15566;
   wire n15567;
   wire n15568;
   wire n15569;
   wire n15570;
   wire n15571;
   wire n15572;
   wire n15573;
   wire n15574;
   wire n15575;
   wire n15576;
   wire n15577;
   wire n15578;
   wire n15579;
   wire n15580;
   wire n15581;
   wire n15582;
   wire n15583;
   wire n15584;
   wire n15585;
   wire n15586;
   wire n15587;
   wire n15588;
   wire n15589;
   wire n15590;
   wire n15591;
   wire n15592;
   wire n15593;
   wire n15594;
   wire n15595;
   wire n15596;
   wire n15597;
   wire n15598;
   wire n15599;
   wire n15600;
   wire n15601;
   wire n15602;
   wire n15603;
   wire n15604;
   wire n15605;
   wire n15606;
   wire n15607;
   wire n15608;
   wire n15609;
   wire n15610;
   wire n15611;
   wire n15612;
   wire n15613;
   wire n15614;
   wire n15615;
   wire n15616;
   wire n15617;
   wire n15619;
   wire n15620;
   wire n15621;
   wire n15622;
   wire n15623;
   wire n15624;
   wire n15625;
   wire n15626;
   wire n15627;
   wire n15628;
   wire n15629;
   wire n15630;
   wire n15631;
   wire n15632;
   wire n15633;
   wire n15634;
   wire n15635;
   wire n15636;
   wire n15637;
   wire n15638;
   wire n15639;
   wire n15640;
   wire n15641;
   wire n15642;
   wire n15643;
   wire n15644;
   wire n15645;
   wire n15646;
   wire n15647;
   wire n15648;
   wire n15649;
   wire n15650;
   wire n15651;
   wire n15652;
   wire n15653;
   wire n15654;
   wire n15655;
   wire n15656;
   wire n15657;
   wire n15658;
   wire n15659;
   wire n15660;
   wire n15661;
   wire n15662;
   wire n15663;
   wire n15664;
   wire n15665;
   wire n15666;
   wire n15667;
   wire n15668;
   wire n15669;
   wire n15670;
   wire n15671;
   wire n15672;
   wire n15673;
   wire n15674;
   wire n15675;
   wire n15676;
   wire n15677;
   wire n15678;
   wire n15679;
   wire n15680;
   wire n15681;
   wire n15682;
   wire n15683;
   wire n15684;
   wire n15685;
   wire n15686;
   wire n15687;
   wire n15688;
   wire n15689;
   wire n15690;
   wire n15691;
   wire n15692;
   wire n15693;
   wire n15694;
   wire n15695;
   wire n15696;
   wire n15697;
   wire n15698;
   wire n15699;
   wire n15700;
   wire n15701;
   wire n15702;
   wire n15703;
   wire n15704;
   wire n15705;
   wire n15706;
   wire n15707;
   wire n15708;
   wire n15709;
   wire n15710;
   wire n15711;
   wire n15712;
   wire n15713;
   wire n15714;
   wire n15715;
   wire n15717;
   wire n15718;
   wire n15719;
   wire n15720;
   wire n15721;
   wire n15722;
   wire n15723;
   wire n15724;
   wire n15726;
   wire n15727;
   wire n15728;
   wire n15729;
   wire n15730;
   wire n15731;
   wire n15732;
   wire n15733;
   wire n15734;
   wire n15735;
   wire n15736;
   wire n15737;
   wire n15738;
   wire n15739;
   wire n15741;
   wire n15742;
   wire n15743;
   wire n15744;
   wire n15745;
   wire n15746;
   wire n15747;
   wire n15748;
   wire n15749;
   wire n15750;
   wire n15751;
   wire n15752;
   wire n15753;
   wire n15754;
   wire n15755;
   wire n15756;
   wire n15757;
   wire n15758;
   wire n15759;
   wire n15760;
   wire n15761;
   wire n15762;
   wire n15763;
   wire n15764;
   wire n15765;
   wire n15766;
   wire n15767;
   wire n15768;
   wire n15769;
   wire n15770;
   wire n15771;
   wire n15772;
   wire n15773;
   wire n15774;
   wire n15775;
   wire n15776;
   wire n15777;
   wire n15778;
   wire n15779;
   wire n15780;
   wire n15781;
   wire n15782;
   wire n15783;
   wire n15784;
   wire n15785;
   wire n15786;
   wire n15787;
   wire n15788;
   wire n15789;
   wire n15790;
   wire n15791;
   wire n15792;
   wire n15793;
   wire n15794;
   wire n15795;
   wire n15796;
   wire n15797;
   wire n15798;
   wire n15799;
   wire n15800;
   wire n15801;
   wire n15802;
   wire n15803;
   wire n15804;
   wire n15805;
   wire n15806;
   wire n15807;
   wire n15808;
   wire n15809;
   wire n15810;
   wire n15811;
   wire n15812;
   wire n15813;
   wire n15814;
   wire n15815;
   wire n15816;
   wire n15817;
   wire n15818;
   wire n15819;
   wire n15820;
   wire n15821;
   wire n15822;
   wire n15823;
   wire n15824;
   wire n15825;
   wire n15827;
   wire n15828;
   wire n15829;
   wire n15830;
   wire n15831;
   wire n15832;
   wire n15833;
   wire n15834;
   wire n15835;
   wire n15837;
   wire n15838;
   wire n15839;
   wire n15840;
   wire n15841;
   wire n15842;
   wire n15843;
   wire n15844;
   wire n15845;
   wire n15846;
   wire n15847;
   wire n15848;
   wire n15849;
   wire n15850;
   wire n15851;
   wire n15852;
   wire n15853;
   wire n15854;
   wire n15855;
   wire n15856;
   wire n15857;
   wire n15858;
   wire n15859;
   wire n15860;
   wire n15861;
   wire n15862;
   wire n15863;
   wire n15864;
   wire n15865;
   wire n15866;
   wire n15867;
   wire n15868;
   wire n15869;
   wire n15870;
   wire n15871;
   wire n15872;
   wire n15873;
   wire n15874;
   wire n15875;
   wire n15876;
   wire n15877;
   wire n15878;
   wire n15879;
   wire n15880;
   wire n15881;
   wire n15882;
   wire n15883;
   wire n15884;
   wire n15885;
   wire n15886;
   wire n15887;
   wire n15888;
   wire n15889;
   wire n15890;
   wire n15891;
   wire n15892;
   wire n15893;
   wire n15894;
   wire n15895;
   wire n15896;
   wire n15897;
   wire n15898;
   wire n15899;
   wire n15900;
   wire n15901;
   wire n15902;
   wire n15903;
   wire n15904;
   wire n15905;
   wire n15906;
   wire n15907;
   wire n15908;
   wire n15909;
   wire n15910;
   wire n15911;
   wire n15912;
   wire n15913;
   wire n15914;
   wire n15915;
   wire n15916;
   wire n15917;
   wire n15918;
   wire n15919;
   wire n15920;
   wire n15921;
   wire n15922;
   wire n15923;
   wire n15924;
   wire n15925;
   wire n15926;
   wire n15927;
   wire n15928;
   wire n15929;
   wire n15930;
   wire n15931;
   wire n15932;
   wire n15933;
   wire n15934;
   wire n15935;
   wire n15936;
   wire n15937;
   wire n15938;
   wire n15939;
   wire n15940;
   wire n15941;
   wire n15942;
   wire n15943;
   wire n15944;
   wire n15945;
   wire n15946;
   wire n15947;
   wire n15948;
   wire n15949;
   wire n15950;
   wire n15951;
   wire n15952;
   wire n15953;
   wire n15954;
   wire n15955;
   wire n15956;
   wire n15957;
   wire n15958;
   wire n15959;
   wire n15960;
   wire n15961;
   wire n15962;
   wire n15963;
   wire n15964;
   wire n15965;
   wire n15966;
   wire n15967;
   wire n15968;
   wire n15969;
   wire n15970;
   wire n15971;
   wire n15972;
   wire n15973;
   wire n15974;
   wire n15975;
   wire n15976;
   wire n15977;
   wire n15978;
   wire n15979;
   wire n15980;
   wire n15981;
   wire n15982;
   wire n15983;
   wire n15984;
   wire n15985;
   wire n15986;
   wire n15987;
   wire n15988;
   wire n15989;
   wire n15990;
   wire n15991;
   wire n15992;
   wire n15993;
   wire n15994;
   wire n15995;
   wire n15996;
   wire n15997;
   wire n15998;
   wire n15999;
   wire n16000;
   wire n16001;
   wire n16002;
   wire n16003;
   wire n16004;
   wire n16005;
   wire n16006;
   wire n16007;
   wire n16008;
   wire n16009;
   wire n16010;
   wire n16012;
   wire n16013;
   wire n16014;
   wire n16015;
   wire n16016;
   wire n16017;
   wire n16018;
   wire n16019;
   wire n16020;
   wire n16021;
   wire n16022;
   wire n16023;
   wire n16024;
   wire n16025;
   wire n16026;
   wire n16027;
   wire n16028;
   wire n16029;
   wire n16030;
   wire n16031;
   wire n16032;
   wire n16033;
   wire n16034;
   wire n16035;
   wire n16036;
   wire n16037;
   wire n16038;
   wire n16039;
   wire n16040;
   wire n16041;
   wire n16042;
   wire n16043;
   wire n16044;
   wire n16045;
   wire n16046;
   wire n16047;
   wire n16048;
   wire n16049;
   wire n16050;
   wire n16052;
   wire n16053;
   wire n16054;
   wire n16055;
   wire n16056;
   wire n16057;
   wire n16058;
   wire n16059;
   wire n16060;
   wire n16061;
   wire n16062;
   wire n16063;
   wire n16064;
   wire n16065;
   wire n16066;
   wire n16067;
   wire n16068;
   wire n16069;
   wire n16070;
   wire n16071;
   wire n16073;
   wire n16074;
   wire n16075;
   wire n16076;
   wire n16077;
   wire n16078;
   wire n16079;
   wire n16080;
   wire n16081;
   wire n16082;
   wire n16083;
   wire n16084;
   wire n16085;
   wire n16086;
   wire n16087;
   wire n16088;
   wire n16089;
   wire n16090;
   wire n16091;
   wire n16092;
   wire n16093;
   wire n16094;
   wire n16095;
   wire n16096;
   wire n16097;
   wire n16098;
   wire n16099;
   wire n16100;
   wire n16101;
   wire n16102;
   wire n16103;
   wire n16104;
   wire n16105;
   wire n16106;
   wire n16108;
   wire n16109;
   wire n16110;
   wire n16111;
   wire n16112;
   wire n16113;
   wire n16114;
   wire n16115;
   wire n16117;
   wire n16118;
   wire n16119;
   wire n16120;
   wire n16121;
   wire n16122;
   wire n16123;
   wire n16124;
   wire n16125;
   wire n16126;
   wire n16127;
   wire n16128;
   wire n16129;
   wire n16130;
   wire n16131;
   wire n16133;
   wire n16134;
   wire n16135;
   wire n16136;
   wire n16137;
   wire n16138;
   wire n16139;
   wire n16140;
   wire n16141;
   wire n16142;
   wire n16143;
   wire n16144;
   wire n16145;
   wire n16146;
   wire n16147;
   wire n16148;
   wire n16149;
   wire n16150;
   wire n16151;
   wire n16152;
   wire n16153;
   wire n16154;
   wire n16155;
   wire n16156;
   wire n16157;
   wire n16158;
   wire n16159;
   wire n16160;
   wire n16161;
   wire n16162;
   wire n16163;
   wire n16164;
   wire n16165;
   wire n16166;
   wire n16167;
   wire n16168;
   wire n16170;
   wire n16171;
   wire n16172;
   wire n16174;
   wire n16175;
   wire n16176;
   wire n16177;
   wire n16178;
   wire n16179;
   wire n16180;
   wire n16181;
   wire n16182;
   wire n16183;
   wire n16184;
   wire n16185;
   wire n16186;
   wire n16187;
   wire n16188;
   wire n16189;
   wire n16191;
   wire n16192;
   wire n16193;
   wire n16194;
   wire n16195;
   wire n16196;
   wire n16197;
   wire n16198;
   wire n16199;
   wire n16200;
   wire n16201;
   wire n16202;
   wire n16203;
   wire n16204;
   wire n16205;
   wire n16206;
   wire n16207;
   wire n16208;
   wire n16209;
   wire n16210;
   wire n16211;
   wire n16212;
   wire n16213;
   wire n16214;
   wire n16215;
   wire n16216;
   wire n16218;
   wire n16219;
   wire n16220;
   wire n16221;
   wire n16222;
   wire n16223;
   wire n16224;
   wire n16225;
   wire n16226;
   wire n16227;
   wire n16228;
   wire n16229;
   wire n16230;
   wire n16231;
   wire n16232;
   wire n16233;
   wire n16234;
   wire n16235;
   wire n16236;
   wire n16237;
   wire n16238;
   wire n16239;
   wire n16240;
   wire n16242;
   wire n16243;
   wire n16244;
   wire n16245;
   wire n16246;
   wire n16247;
   wire n16248;
   wire n16249;
   wire n16250;
   wire n16251;
   wire n16252;
   wire n16253;
   wire n16254;
   wire n16255;
   wire n16257;
   wire n16258;
   wire n16259;
   wire n16260;
   wire n16261;
   wire n16262;
   wire n16263;
   wire n16265;
   wire n16266;
   wire n16267;
   wire n16268;
   wire n16269;
   wire n16270;
   wire n16271;
   wire n16272;
   wire n16273;
   wire n16274;
   wire n16275;
   wire n16276;
   wire n16278;
   wire n16279;
   wire n16280;
   wire n16281;
   wire n16282;
   wire n16283;
   wire n16284;
   wire n16285;
   wire n16286;
   wire n16287;
   wire n16288;
   wire n16289;
   wire n16290;
   wire n16291;
   wire n16295;
   wire n16296;
   wire n16297;
   wire n16298;
   wire n16299;
   wire n16300;
   wire n16301;
   wire n16302;
   wire n16303;
   wire n16304;
   wire n16305;
   wire n16306;
   wire n16307;
   wire n16308;
   wire n16309;
   wire n16310;
   wire n16311;
   wire n16312;
   wire n16313;
   wire n16314;
   wire n16315;
   wire n16316;
   wire n16317;
   wire n16318;
   wire n16319;
   wire n16320;
   wire n16321;
   wire n16322;
   wire n16323;
   wire n16324;
   wire n16326;
   wire n16327;
   wire n16328;
   wire n16329;
   wire n16330;
   wire n16331;
   wire n16332;
   wire n16333;
   wire n16334;
   wire n16335;
   wire n16336;
   wire n16337;
   wire n16338;
   wire n16339;
   wire n16340;
   wire n16341;
   wire n16342;
   wire n16343;
   wire n16344;
   wire n16345;
   wire n16346;
   wire n16347;
   wire n16348;
   wire n16349;
   wire n16350;
   wire n16351;
   wire n16352;
   wire n16353;
   wire n16354;
   wire n16355;
   wire n16356;
   wire n16357;
   wire n16358;
   wire n16359;
   wire n16360;
   wire n16361;
   wire n16362;
   wire n16363;
   wire n16364;
   wire n16365;
   wire n16366;
   wire n16367;
   wire n16368;
   wire n16369;
   wire n16370;
   wire n16371;
   wire n16372;
   wire n16373;
   wire n16374;
   wire n16375;
   wire n16376;
   wire n16377;
   wire n16378;
   wire n16379;
   wire n16380;
   wire n16381;
   wire n16382;
   wire n16385;
   wire n16386;
   wire n16387;
   wire n16388;
   wire n16389;
   wire n16390;
   wire n16391;
   wire n16392;
   wire n16393;
   wire n16394;
   wire n16395;
   wire n16396;
   wire n16397;
   wire n16398;
   wire n16399;
   wire n16400;
   wire n16401;
   wire n16402;
   wire n16403;
   wire n16404;
   wire n16405;
   wire n16406;
   wire n16407;
   wire n16408;
   wire n16409;
   wire n16410;
   wire n16411;
   wire n16412;
   wire n16413;
   wire n16414;
   wire n16415;
   wire n16416;
   wire n16417;
   wire n16418;
   wire n16419;
   wire n16421;
   wire n16422;
   wire n16423;
   wire n16424;
   wire n16425;
   wire n16426;
   wire n16427;
   wire n16429;
   wire n16430;
   wire n16432;
   wire n16433;
   wire n16434;
   wire n16436;
   wire n16437;
   wire n16438;
   wire n16439;
   wire n16440;
   wire n16441;
   wire n16442;
   wire n16443;
   wire n16444;
   wire n16445;
   wire n16446;
   wire n16447;
   wire n16448;
   wire n16449;
   wire n16450;
   wire n16451;
   wire n16452;
   wire n16453;
   wire n16454;
   wire n16455;
   wire n16456;
   wire n16457;
   wire n16458;
   wire n16459;
   wire n16460;
   wire n16461;
   wire n16462;
   wire n16463;
   wire n16464;
   wire n16465;
   wire n16466;
   wire n16467;
   wire n16468;
   wire n16469;
   wire n16470;
   wire n16471;
   wire n16472;
   wire n16473;
   wire n16474;
   wire n16475;
   wire n16476;
   wire n16477;
   wire n16478;
   wire n16479;
   wire n16480;
   wire n16481;
   wire n16482;
   wire n16483;
   wire n16484;
   wire n16485;
   wire n16486;
   wire n16487;
   wire n16488;
   wire n16489;
   wire n16490;
   wire n16491;
   wire n16492;
   wire n16493;
   wire n16494;
   wire n16495;
   wire n16496;
   wire n16497;
   wire n16498;
   wire n16499;
   wire n16500;
   wire n16501;
   wire n16502;
   wire n16503;
   wire n16504;
   wire n16505;
   wire n16506;
   wire n16507;
   wire n16508;
   wire n16509;
   wire n16510;
   wire n16511;
   wire n16512;
   wire n16513;
   wire n16514;
   wire n16515;
   wire n16516;
   wire n16517;
   wire n16518;
   wire n16519;
   wire n16520;
   wire n16521;
   wire n16522;
   wire n16523;
   wire n16524;
   wire n16525;
   wire n16526;
   wire n16527;
   wire n16528;
   wire n16529;
   wire n16530;
   wire n16531;
   wire n16533;
   wire n16534;
   wire n16536;
   wire n16537;
   wire n16538;
   wire n16539;
   wire n16540;
   wire n16541;
   wire n16542;
   wire n16543;
   wire n16544;
   wire n16545;
   wire n16546;
   wire n16547;
   wire n16548;
   wire n16549;
   wire n16550;
   wire n16551;
   wire n16552;
   wire n16553;
   wire n16554;
   wire n16555;
   wire n16556;
   wire n16557;
   wire n16558;
   wire n16559;
   wire n16560;
   wire n16561;
   wire n16562;
   wire n16563;
   wire n16564;
   wire n16565;
   wire n16566;
   wire n16567;
   wire n16568;
   wire n16569;
   wire n16570;
   wire n16571;
   wire n16572;
   wire n16573;
   wire n16574;
   wire n16575;
   wire n16576;
   wire n16577;
   wire n16578;
   wire n16579;
   wire n16580;
   wire n16581;
   wire n16582;
   wire n16583;
   wire n16584;
   wire n16585;
   wire n16586;
   wire n16587;
   wire n16588;
   wire n16589;
   wire n16590;
   wire n16591;
   wire n16592;
   wire n16593;
   wire n16594;
   wire n16596;
   wire n16597;
   wire n16598;
   wire n16599;
   wire n16600;
   wire n16601;
   wire n16602;
   wire n16603;
   wire n16604;
   wire n16605;
   wire n16606;
   wire n16607;
   wire n16608;
   wire n16609;
   wire n16610;
   wire n16611;
   wire n16612;
   wire n16613;
   wire n16614;
   wire n16615;
   wire n16616;
   wire n16617;
   wire n16618;
   wire n16619;
   wire n16620;
   wire n16621;
   wire n16622;
   wire n16623;
   wire n16624;
   wire n16625;
   wire n16626;
   wire n16627;
   wire n16628;
   wire n16629;
   wire n16630;
   wire n16631;
   wire n16632;
   wire n16633;
   wire n16634;
   wire n16635;
   wire n16636;
   wire n16637;
   wire n16638;
   wire n16639;
   wire n16640;
   wire n16641;
   wire n16642;
   wire n16643;
   wire n16644;
   wire n16645;
   wire n16646;
   wire n16647;
   wire n16648;
   wire n16649;
   wire n16650;
   wire n16651;
   wire n16652;
   wire n16653;
   wire n16654;
   wire n16655;
   wire n16656;
   wire n16658;
   wire n16659;
   wire n16660;
   wire n16661;
   wire n16662;
   wire n16663;
   wire n16664;
   wire n16665;
   wire n16666;
   wire n16667;
   wire n16668;
   wire n16669;
   wire n16670;
   wire n16671;
   wire n16672;
   wire n16673;
   wire n16674;
   wire n16675;
   wire n16676;
   wire n16677;
   wire n16678;
   wire n16679;
   wire n16680;
   wire n16681;
   wire n16682;
   wire n16683;
   wire n16684;
   wire n16685;
   wire n16686;
   wire n16687;
   wire n16688;
   wire n16689;
   wire n16690;
   wire n16691;
   wire n16692;
   wire n16693;
   wire n16694;
   wire n16695;
   wire n16696;
   wire n16697;
   wire n16698;
   wire n16699;
   wire n16700;
   wire n16701;
   wire n16702;
   wire n16703;
   wire n16704;
   wire n16705;
   wire n16706;
   wire n16707;
   wire n16708;
   wire n16709;
   wire n16710;
   wire n16711;
   wire n16712;
   wire n16713;
   wire n16714;
   wire n16715;
   wire n16716;
   wire n16717;
   wire n16718;
   wire n16719;
   wire n16720;
   wire n16721;
   wire n16722;
   wire n16723;
   wire n16724;
   wire n16725;
   wire n16726;
   wire n16727;
   wire n16728;
   wire n16729;
   wire n16730;
   wire n16731;
   wire n16732;
   wire n16733;
   wire n16734;
   wire n16735;
   wire n16736;
   wire n16737;
   wire n16738;
   wire n16739;
   wire n16740;
   wire n16741;
   wire n16742;
   wire n16743;
   wire n16744;
   wire n16745;
   wire n16746;
   wire n16747;
   wire n16748;
   wire n16749;
   wire n16750;
   wire n16751;
   wire n16752;
   wire n16753;
   wire n16754;
   wire n16755;
   wire n16756;
   wire n16757;
   wire n16758;
   wire n16759;
   wire n16760;
   wire n16761;
   wire n16762;
   wire n16763;
   wire n16764;
   wire n16765;
   wire n16766;
   wire n16767;
   wire n16768;
   wire n16769;
   wire n16770;
   wire n16771;
   wire n16772;
   wire n16773;
   wire n16774;
   wire n16775;
   wire n16776;
   wire n16777;
   wire n16779;
   wire n16780;
   wire n16781;
   wire n16782;
   wire n16783;
   wire n16784;
   wire n16785;
   wire n16786;
   wire n16787;
   wire n16788;
   wire n16789;
   wire n16790;
   wire n16791;
   wire n16793;
   wire n16794;
   wire n16795;
   wire n16796;
   wire n16797;
   wire n16798;
   wire n16799;
   wire n16800;
   wire n16801;
   wire n16802;
   wire n16803;
   wire n16804;
   wire n16805;
   wire n16806;
   wire n16807;
   wire n16808;
   wire n16809;
   wire n16810;
   wire n16811;
   wire n16812;
   wire n16814;
   wire n16815;
   wire n16816;
   wire n16817;
   wire n16818;
   wire n16819;
   wire n16820;
   wire n16821;
   wire n16822;
   wire n16823;
   wire n16824;
   wire n16825;
   wire n16826;
   wire n16827;
   wire n16828;
   wire n16829;
   wire n16830;
   wire n16831;
   wire n16832;
   wire n16833;
   wire n16834;
   wire n16835;
   wire n16836;
   wire n16837;
   wire n16838;
   wire n16839;
   wire n16840;
   wire n16841;
   wire n16842;
   wire n16843;
   wire n16844;
   wire n16845;
   wire n16846;
   wire n16847;
   wire n16848;
   wire n16849;
   wire n16850;
   wire n16851;
   wire n16852;
   wire n16853;
   wire n16854;
   wire n16855;
   wire n16856;
   wire n16857;
   wire n16858;
   wire n16859;
   wire n16860;
   wire n16861;
   wire n16862;
   wire n16863;
   wire n16864;
   wire n16865;
   wire n16867;
   wire n16868;
   wire n16869;
   wire n16870;
   wire n16871;
   wire n16872;
   wire n16873;
   wire n16874;
   wire n16875;
   wire n16877;
   wire n16878;
   wire n16879;
   wire n16880;
   wire n16881;
   wire n16882;
   wire n16883;
   wire n16884;
   wire n16885;
   wire n16886;
   wire n16887;
   wire n16888;
   wire n16889;
   wire n16890;
   wire n16891;
   wire n16893;
   wire n16894;
   wire n16895;
   wire n16896;
   wire n16897;
   wire n16898;
   wire n16899;
   wire n16900;
   wire n16901;
   wire n16902;
   wire n16903;
   wire n16904;
   wire n16905;
   wire n16906;
   wire n16907;
   wire n16908;
   wire n16909;
   wire n16910;
   wire n16911;
   wire n16912;
   wire n16913;
   wire n16914;
   wire n16915;
   wire n16916;
   wire n16917;
   wire n16918;
   wire n16919;
   wire n16920;
   wire n16921;
   wire n16922;
   wire n16923;
   wire n16924;
   wire n16925;
   wire n16926;
   wire n16927;
   wire n16928;
   wire n16929;
   wire n16930;
   wire n16931;
   wire n16932;
   wire n16933;
   wire n16934;
   wire n16935;
   wire n16936;
   wire n16937;
   wire n16938;
   wire n16939;
   wire n16940;
   wire n16941;
   wire n16942;
   wire n16943;
   wire n16944;
   wire n16945;
   wire n16946;
   wire n16947;
   wire n16948;
   wire n16949;
   wire n16950;
   wire n16951;
   wire n16952;
   wire n16953;
   wire n16954;
   wire n16955;
   wire n16956;
   wire n16957;
   wire n16958;
   wire n16959;
   wire n16960;
   wire n16961;
   wire n16962;
   wire n16963;
   wire n16964;
   wire n16965;
   wire n16966;
   wire n16967;
   wire n16968;
   wire n16969;
   wire n16970;
   wire n16971;
   wire n16972;
   wire n16973;
   wire n16974;
   wire n16975;
   wire n16976;
   wire n16977;
   wire n16978;
   wire n16980;
   wire n16981;
   wire n16982;
   wire n16983;
   wire n16984;
   wire n16985;
   wire n16986;
   wire n16987;
   wire n16988;
   wire n16989;
   wire n16990;
   wire n16991;
   wire n16992;
   wire n16993;
   wire n16994;
   wire n16995;
   wire n16996;
   wire n16997;
   wire n16998;
   wire n16999;
   wire n17000;
   wire n17001;
   wire n17002;
   wire n17003;
   wire n17004;
   wire n17005;
   wire n17006;
   wire n17007;
   wire n17008;
   wire n17009;
   wire n17010;
   wire n17011;
   wire n17012;
   wire n17013;
   wire n17014;
   wire n17015;
   wire n17016;
   wire n17017;
   wire n17018;
   wire n17019;
   wire n17020;
   wire n17021;
   wire n17022;
   wire n17023;
   wire n17024;
   wire n17025;
   wire n17026;
   wire n17027;
   wire n17028;
   wire n17029;
   wire n17030;
   wire n17031;
   wire n17033;
   wire n17034;
   wire n17035;
   wire n17036;
   wire n17037;
   wire n17038;
   wire n17039;
   wire n17040;
   wire n17041;
   wire n17042;
   wire n17043;
   wire n17044;
   wire n17045;
   wire n17046;
   wire n17047;
   wire n17048;
   wire n17049;
   wire n17050;
   wire n17051;
   wire n17052;
   wire n17053;
   wire n17054;
   wire n17055;
   wire n17056;
   wire n17057;
   wire n17058;
   wire n17059;
   wire n17060;
   wire n17061;
   wire n17062;
   wire n17063;
   wire n17064;
   wire n17065;
   wire n17066;
   wire n17067;
   wire n17068;
   wire n17069;
   wire n17070;
   wire n17071;
   wire n17072;
   wire n17073;
   wire n17074;
   wire n17075;
   wire n17076;
   wire n17077;
   wire n17078;
   wire n17079;
   wire n17080;
   wire n17081;
   wire n17082;
   wire n17083;
   wire n17084;
   wire n17085;
   wire n17086;
   wire n17087;
   wire n17088;
   wire n17089;
   wire n17090;
   wire n17091;
   wire n17092;
   wire n17093;
   wire n17094;
   wire n17095;
   wire n17096;
   wire n17097;
   wire n17098;
   wire n17099;
   wire n17100;
   wire n17101;
   wire n17102;
   wire n17103;
   wire n17104;
   wire n17105;
   wire n17106;
   wire n17107;
   wire n17108;
   wire n17109;
   wire n17110;
   wire n17111;
   wire n17112;
   wire n17113;
   wire n17114;
   wire n17115;
   wire n17116;
   wire n17117;
   wire n17118;
   wire n17119;
   wire n17120;
   wire n17121;
   wire n17122;
   wire n17123;
   wire n17124;
   wire n17125;
   wire n17126;
   wire n17127;
   wire n17128;
   wire n17129;
   wire n17130;
   wire n17131;
   wire n17132;
   wire n17133;
   wire n17134;
   wire n17135;
   wire n17136;
   wire n17137;
   wire n17138;
   wire n17139;
   wire n17140;
   wire n17141;
   wire n17142;
   wire n17143;
   wire n17144;
   wire n17145;
   wire n17146;
   wire n17147;
   wire n17148;
   wire n17149;
   wire n17150;
   wire n17151;
   wire n17152;
   wire n17153;
   wire n17154;
   wire n17155;
   wire n17156;
   wire n17157;
   wire n17158;
   wire n17159;
   wire n17160;
   wire n17161;
   wire n17162;
   wire n17163;
   wire n17164;
   wire n17165;
   wire n17166;
   wire n17167;
   wire n17168;
   wire n17169;
   wire n17170;
   wire n17171;
   wire n17172;
   wire n17173;
   wire n17174;
   wire n17175;
   wire n17176;
   wire n17179;
   wire n17180;
   wire n17181;
   wire n17182;
   wire n17183;
   wire n17184;
   wire n17185;
   wire n17186;
   wire n17187;
   wire n17188;
   wire n17189;
   wire n17190;
   wire n17191;
   wire n17192;
   wire n17193;
   wire n17194;
   wire n17195;
   wire n17196;
   wire n17197;
   wire n17198;
   wire n17199;
   wire n17200;
   wire n17201;
   wire n17202;
   wire n17203;
   wire n17204;
   wire n17205;
   wire n17206;
   wire n17207;
   wire n17208;
   wire n17209;
   wire n17210;
   wire n17211;
   wire n17212;
   wire n17213;
   wire n17214;
   wire n17215;
   wire n17216;
   wire n17217;
   wire n17218;
   wire n17219;
   wire n17220;
   wire n17221;
   wire n17222;
   wire n17223;
   wire n17224;
   wire n17225;
   wire n17226;
   wire n17227;
   wire n17228;
   wire n17229;
   wire n17230;
   wire n17231;
   wire n17232;
   wire n17233;
   wire n17234;
   wire n17236;
   wire n17237;
   wire n17239;
   wire n17240;
   wire n17241;
   wire n17242;
   wire n17243;
   wire n17244;
   wire n17245;
   wire n17246;
   wire n17247;
   wire n17248;
   wire n17249;
   wire n17250;
   wire n17251;
   wire n17252;
   wire n17253;
   wire n17254;
   wire n17255;
   wire n17256;
   wire n17257;
   wire n17258;
   wire n17259;
   wire n17260;
   wire n17261;
   wire n17262;
   wire n17263;
   wire n17264;
   wire n17265;
   wire n17266;
   wire n17268;
   wire n17269;
   wire n17270;
   wire n17271;
   wire n17272;
   wire n17273;
   wire n17274;
   wire n17275;
   wire n17276;
   wire n17277;
   wire n17278;
   wire n17279;
   wire n17280;
   wire n17281;
   wire n17282;
   wire n17283;
   wire n17284;
   wire n17285;
   wire n17286;
   wire n17287;
   wire n17288;
   wire n17289;
   wire n17290;
   wire n17291;
   wire n17292;
   wire n17293;
   wire n17294;
   wire n17295;
   wire n17296;
   wire n17297;
   wire n17298;
   wire n17299;
   wire n17300;
   wire n17301;
   wire n17302;
   wire n17303;
   wire n17304;
   wire n17305;
   wire n17306;
   wire n17307;
   wire n17308;
   wire n17309;
   wire n17310;
   wire n17312;
   wire n17313;
   wire n17314;
   wire n17317;
   wire n17318;
   wire n17320;
   wire n17321;
   wire n17322;
   wire n17323;
   wire n17324;
   wire n17325;
   wire n17326;
   wire n17327;
   wire n17328;
   wire n17329;
   wire n17330;
   wire n17331;
   wire n17332;
   wire n17333;
   wire n17334;
   wire n17335;
   wire n17336;
   wire n17337;
   wire n17338;
   wire n17339;
   wire n17340;
   wire n17341;
   wire n17342;
   wire n17343;
   wire n17344;
   wire n17345;
   wire n17346;
   wire n17347;
   wire n17348;
   wire n17349;
   wire n17350;
   wire n17351;
   wire n17352;
   wire n17353;
   wire n17354;
   wire n17355;
   wire n17356;
   wire n17357;
   wire n17358;
   wire n17359;
   wire n17360;
   wire n17361;
   wire n17362;
   wire n17363;
   wire n17364;
   wire n17365;
   wire n17366;
   wire n17367;
   wire n17368;
   wire n17369;
   wire n17370;
   wire n17371;
   wire n17372;
   wire n17373;
   wire n17374;
   wire n17375;
   wire n17376;
   wire n17377;
   wire n17378;
   wire n17379;
   wire n17380;
   wire n17381;
   wire n17382;
   wire n17383;
   wire n17384;
   wire n17385;
   wire n17386;
   wire n17387;
   wire n17388;
   wire n17389;
   wire n17390;
   wire n17391;
   wire n17392;
   wire n17393;
   wire n17394;
   wire n17395;
   wire n17396;
   wire n17397;
   wire n17398;
   wire n17399;
   wire n17401;
   wire n17402;
   wire n17403;
   wire n17404;
   wire n17405;
   wire n17406;
   wire n17407;
   wire n17408;
   wire n17409;
   wire n17410;
   wire n17411;
   wire n17412;
   wire n17413;
   wire n17414;
   wire n17415;
   wire n17416;
   wire n17417;
   wire n17418;
   wire n17419;
   wire n17420;
   wire n17421;
   wire n17422;
   wire n17423;
   wire n17424;
   wire n17425;
   wire n17426;
   wire n17428;
   wire n17429;
   wire n17430;
   wire n17431;
   wire n17432;
   wire n17433;
   wire n17434;
   wire n17435;
   wire n17436;
   wire n17437;
   wire n17438;
   wire n17439;
   wire n17440;
   wire n17441;
   wire n17442;
   wire n17443;
   wire n17444;
   wire n17445;
   wire n17446;
   wire n17447;
   wire n17449;
   wire n17450;
   wire n17451;
   wire n17452;
   wire n17453;
   wire n17454;
   wire n17455;
   wire n17456;
   wire n17457;
   wire n17458;
   wire n17459;
   wire n17460;
   wire n17461;
   wire n17462;
   wire n17463;
   wire n17464;
   wire n17465;
   wire n17466;
   wire n17467;
   wire n17468;
   wire n17469;
   wire n17470;
   wire n17471;
   wire n17472;
   wire n17473;
   wire n17474;
   wire n17475;
   wire n17476;
   wire n17477;
   wire n17479;
   wire n17480;
   wire n17481;
   wire n17482;
   wire n17483;
   wire n17484;
   wire n17485;
   wire n17486;
   wire n17487;
   wire n17488;
   wire n17489;
   wire n17490;
   wire n17491;
   wire n17492;
   wire n17493;
   wire n17494;
   wire n17495;
   wire n17496;
   wire n17497;
   wire n17498;
   wire n17499;
   wire n17500;
   wire n17501;
   wire n17502;
   wire n17503;
   wire n17504;
   wire n17505;
   wire n17506;
   wire n17507;
   wire n17508;
   wire n17509;
   wire n17510;
   wire n17511;
   wire n17512;
   wire n17513;
   wire n17514;
   wire n17515;
   wire n17516;
   wire n17517;
   wire n17518;
   wire n17519;
   wire n17520;
   wire n17521;
   wire n17522;
   wire n17525;
   wire n17526;
   wire n17527;
   wire n17528;
   wire n17529;
   wire n17530;
   wire n17531;
   wire n17532;
   wire n17533;
   wire n17534;
   wire n17535;
   wire n17536;
   wire n17537;
   wire n17538;
   wire n17539;
   wire n17540;
   wire n17542;
   wire n17543;
   wire n17544;
   wire n17545;
   wire n17546;
   wire n17547;
   wire n17548;
   wire n17549;
   wire n17550;
   wire n17551;
   wire n17552;
   wire n17553;
   wire n17554;
   wire n17555;
   wire n17556;
   wire n17557;
   wire n17558;
   wire n17559;
   wire n17560;
   wire n17561;
   wire n17562;
   wire n17563;
   wire n17564;
   wire n17565;
   wire n17566;
   wire n17567;
   wire n17568;
   wire n17569;
   wire n17570;
   wire n17571;
   wire n17572;
   wire n17573;
   wire n17574;
   wire n17575;
   wire n17576;
   wire n17577;
   wire n17578;
   wire n17579;
   wire n17580;
   wire n17581;
   wire n17582;
   wire n17583;
   wire n17584;
   wire n17585;
   wire n17586;
   wire n17587;
   wire n17588;
   wire n17589;
   wire n17590;
   wire n17591;
   wire n17592;
   wire n17593;
   wire n17594;
   wire n17595;
   wire n17596;
   wire n17597;
   wire n17598;
   wire n17599;
   wire n17600;
   wire n17601;
   wire n17602;
   wire n17603;
   wire n17604;
   wire n17605;
   wire n17606;
   wire n17607;
   wire n17608;
   wire n17609;
   wire n17610;
   wire n17611;
   wire n17612;
   wire n17613;
   wire n17614;
   wire n17615;
   wire n17616;
   wire n17617;
   wire n17618;
   wire n17619;
   wire n17620;
   wire n17621;
   wire n17622;
   wire n17623;
   wire n17624;
   wire n17625;
   wire n17626;
   wire n17627;
   wire n17628;
   wire n17629;
   wire n17630;
   wire n17631;
   wire n17632;
   wire n17633;
   wire n17634;
   wire n17635;
   wire n17636;
   wire n17637;
   wire n17638;
   wire n17639;
   wire n17640;
   wire n17641;
   wire n17642;
   wire n17643;
   wire n17644;
   wire n17645;
   wire n17646;
   wire n17647;
   wire n17648;
   wire n17649;
   wire n17650;
   wire n17651;
   wire n17652;
   wire n17653;
   wire n17654;
   wire n17655;
   wire n17656;
   wire n17657;
   wire n17658;
   wire n17659;
   wire n17660;
   wire n17661;
   wire n17662;
   wire n17663;
   wire n17664;
   wire n17665;
   wire n17666;
   wire n17667;
   wire n17668;
   wire n17669;
   wire n17670;
   wire n17671;
   wire n17672;
   wire n17673;
   wire n17674;
   wire n17675;
   wire n17678;
   wire n17679;
   wire n17680;
   wire n17681;
   wire n17682;
   wire n17683;
   wire n17684;
   wire n17685;
   wire n17686;
   wire n17687;
   wire n17688;
   wire n17689;
   wire n17690;
   wire n17691;
   wire n17692;
   wire n17693;
   wire n17694;
   wire n17695;
   wire n17696;
   wire n17697;
   wire n17698;
   wire n17699;
   wire n17700;
   wire n17701;
   wire n17702;
   wire n17703;
   wire n17704;
   wire n17705;
   wire n17706;
   wire n17707;
   wire n17708;
   wire n17709;
   wire n17710;
   wire n17711;
   wire n17712;
   wire n17713;
   wire n17714;
   wire n17715;
   wire n17716;
   wire n17717;
   wire n17718;
   wire n17719;
   wire n17720;
   wire n17721;
   wire n17722;
   wire n17723;
   wire n17724;
   wire n17725;
   wire n17726;
   wire n17727;
   wire n17728;
   wire n17729;
   wire n17730;
   wire n17731;
   wire n17732;
   wire n17733;
   wire n17734;
   wire n17735;
   wire n17736;
   wire n17737;
   wire n17738;
   wire n17740;
   wire n17741;
   wire n17742;
   wire n17743;
   wire n17744;
   wire n17745;
   wire n17747;
   wire n17748;
   wire n17749;
   wire n17750;
   wire n17751;
   wire n17752;
   wire n17753;
   wire n17754;
   wire n17755;
   wire n17756;
   wire n17757;
   wire n17758;
   wire n17759;
   wire n17760;
   wire n17761;
   wire n17762;
   wire n17763;
   wire n17764;
   wire n17765;
   wire n17766;
   wire n17767;
   wire n17768;
   wire n17769;
   wire n17770;
   wire n17771;
   wire n17772;
   wire n17773;
   wire n17774;
   wire n17775;
   wire n17776;
   wire n17777;
   wire n17778;
   wire n17780;
   wire n17782;
   wire n17783;
   wire n17784;
   wire n17785;
   wire n17786;
   wire n17787;
   wire n17788;
   wire n17789;
   wire n17790;
   wire n17791;
   wire n17792;
   wire n17793;
   wire n17794;
   wire n17795;
   wire n17796;
   wire n17797;
   wire n17798;
   wire n17799;
   wire n17801;
   wire n17802;
   wire n17803;
   wire n17804;
   wire n17805;
   wire n17806;
   wire n17807;
   wire n17808;
   wire n17809;
   wire n17810;
   wire n17811;
   wire n17812;
   wire n17813;
   wire n17814;
   wire n17815;
   wire n17816;
   wire n17817;
   wire n17818;
   wire n17819;
   wire n17820;
   wire n17821;
   wire n17822;
   wire n17823;
   wire n17824;
   wire n17825;
   wire n17826;
   wire n17827;
   wire n17828;
   wire n17829;
   wire n17830;
   wire n17831;
   wire n17832;
   wire n17833;
   wire n17834;
   wire n17835;
   wire n17836;
   wire n17837;
   wire n17838;
   wire n17840;
   wire n17841;
   wire n17842;
   wire n17843;
   wire n17844;
   wire n17845;
   wire n17846;
   wire n17847;
   wire n17848;
   wire n17849;
   wire n17850;
   wire n17851;
   wire n17852;
   wire n17853;
   wire n17854;
   wire n17855;
   wire n17856;
   wire n17857;
   wire n17858;
   wire n17859;
   wire n17860;
   wire n17861;
   wire n17862;
   wire n17863;
   wire n17864;
   wire n17865;
   wire n17866;
   wire n17867;
   wire n17868;
   wire n17869;
   wire n17870;
   wire n17871;
   wire n17872;
   wire n17873;
   wire n17874;
   wire n17875;
   wire n17876;
   wire n17877;
   wire n17878;
   wire n17879;
   wire n17880;
   wire n17881;
   wire n17882;
   wire n17883;
   wire n17884;
   wire n17885;
   wire n17886;
   wire n17887;
   wire n17888;
   wire n17889;
   wire n17890;
   wire n17891;
   wire n17892;
   wire n17893;
   wire n17894;
   wire n17895;
   wire n17896;
   wire n17898;
   wire n17899;
   wire n17900;
   wire n17901;
   wire n17902;
   wire n17903;
   wire n17904;
   wire n17906;
   wire n17907;
   wire n17908;
   wire n17909;
   wire n17910;
   wire n17912;
   wire n17913;
   wire n17914;
   wire n17915;
   wire n17916;
   wire n17917;
   wire n17918;
   wire n17919;
   wire n17920;
   wire n17921;
   wire n17922;
   wire n17923;
   wire n17925;
   wire n17926;
   wire n17927;
   wire n17928;
   wire n17929;
   wire n17930;
   wire n17931;
   wire n17932;
   wire n17933;
   wire n17934;
   wire n17935;
   wire n17936;
   wire n17937;
   wire n17938;
   wire n17939;
   wire n17940;
   wire n17941;
   wire n17942;
   wire n17943;
   wire n17944;
   wire n17945;
   wire n17946;
   wire n17947;
   wire n17948;
   wire n17949;
   wire n17950;
   wire n17951;
   wire n17952;
   wire n17953;
   wire n17954;
   wire n17955;
   wire n17956;
   wire n17957;
   wire n17958;
   wire n17959;
   wire n17960;
   wire n17961;
   wire n17962;
   wire n17963;
   wire n17964;
   wire n17965;
   wire n17966;
   wire n17967;
   wire n17968;
   wire n17969;
   wire n17970;
   wire n17971;
   wire n17972;
   wire n17973;
   wire n17974;
   wire n17975;
   wire n17976;
   wire n17977;
   wire n17978;
   wire n17979;
   wire n17980;
   wire n17981;
   wire n17982;
   wire n17983;
   wire n17984;
   wire n17986;
   wire n17989;
   wire n17990;
   wire n17991;
   wire n17992;
   wire n17993;
   wire n17994;
   wire n17995;
   wire n17996;
   wire n17997;
   wire n17998;
   wire n17999;
   wire n18000;
   wire n18001;
   wire n18002;
   wire n18003;
   wire n18004;
   wire n18005;
   wire n18006;
   wire n18007;
   wire n18008;
   wire n18009;
   wire n18010;
   wire n18011;
   wire n18012;
   wire n18013;
   wire n18014;
   wire n18015;
   wire n18016;
   wire n18017;
   wire n18018;
   wire n18019;
   wire n18020;
   wire n18021;
   wire n18022;
   wire n18023;
   wire n18024;
   wire n18025;
   wire n18026;
   wire n18027;
   wire n18028;
   wire n18029;
   wire n18031;
   wire n18032;
   wire n18033;
   wire n18034;
   wire n18035;
   wire n18036;
   wire n18037;
   wire n18038;
   wire n18039;
   wire n18040;
   wire n18041;
   wire n18042;
   wire n18043;
   wire n18044;
   wire n18045;
   wire n18046;
   wire n18047;
   wire n18048;
   wire n18049;
   wire n18050;
   wire n18051;
   wire n18052;
   wire n18053;
   wire n18054;
   wire n18055;
   wire n18056;
   wire n18057;
   wire n18058;
   wire n18059;
   wire n18060;
   wire n18061;
   wire n18062;
   wire n18063;
   wire n18064;
   wire n18065;
   wire n18066;
   wire n18067;
   wire n18068;
   wire n18069;
   wire n18070;
   wire n18071;
   wire n18072;
   wire n18073;
   wire n18074;
   wire n18075;
   wire n18076;
   wire n18077;
   wire n18078;
   wire n18079;
   wire n18080;
   wire n18081;
   wire n18082;
   wire n18083;
   wire n18084;
   wire n18085;
   wire n18086;
   wire n18087;
   wire n18088;
   wire n18089;
   wire n18090;
   wire n18091;
   wire n18092;
   wire n18093;
   wire n18094;
   wire n18095;
   wire n18096;
   wire n18097;
   wire n18098;
   wire n18099;
   wire n18100;
   wire n18101;
   wire n18102;
   wire n18103;
   wire n18104;
   wire n18105;
   wire n18106;
   wire n18107;
   wire n18108;
   wire n18109;
   wire n18110;
   wire n18111;
   wire n18112;
   wire n18113;
   wire n18114;
   wire n18115;
   wire n18116;
   wire n18117;
   wire n18118;
   wire n18119;
   wire n18120;
   wire n18121;
   wire n18122;
   wire n18123;
   wire n18124;
   wire n18125;
   wire n18126;
   wire n18127;
   wire n18128;
   wire n18129;
   wire n18130;
   wire n18131;
   wire n18132;
   wire n18133;
   wire n18134;
   wire n18135;
   wire n18136;
   wire n18137;
   wire n18138;
   wire n18139;
   wire n18140;
   wire n18141;
   wire n18142;
   wire n18143;
   wire n18144;
   wire n18145;
   wire n18146;
   wire n18147;
   wire n18148;
   wire n18149;
   wire n18150;
   wire n18151;
   wire n18152;
   wire n18153;
   wire n18154;
   wire n18155;
   wire n18156;
   wire n18157;
   wire n18158;
   wire n18159;
   wire n18160;
   wire n18161;
   wire n18162;
   wire n18164;
   wire n18165;
   wire n18166;
   wire n18167;
   wire n18168;
   wire n18169;
   wire n18170;
   wire n18171;
   wire n18172;
   wire n18173;
   wire n18174;
   wire n18175;
   wire n18176;
   wire n18177;
   wire n18178;
   wire n18179;
   wire n18180;
   wire n18181;
   wire n18182;
   wire n18183;
   wire n18184;
   wire n18185;
   wire n18186;
   wire n18187;
   wire n18188;
   wire n18189;
   wire n18190;
   wire n18191;
   wire n18192;
   wire n18193;
   wire n18194;
   wire n18195;
   wire n18196;
   wire n18197;
   wire n18198;
   wire n18199;
   wire n18200;
   wire n18201;
   wire n18202;
   wire n18203;
   wire n18204;
   wire n18205;
   wire n18206;
   wire n18207;
   wire n18208;
   wire n18209;
   wire n18210;
   wire n18211;
   wire n18212;
   wire n18213;
   wire n18214;
   wire n18215;
   wire n18216;
   wire n18217;
   wire n18218;
   wire n18219;
   wire n18221;
   wire n18222;
   wire n18223;
   wire n18224;
   wire n18225;
   wire n18226;
   wire n18227;
   wire n18228;
   wire n18229;
   wire n18230;
   wire n18231;
   wire n18232;
   wire n18233;
   wire n18234;
   wire n18235;
   wire n18236;
   wire n18237;
   wire n18238;
   wire n18239;
   wire n18240;
   wire n18241;
   wire n18242;
   wire n18244;
   wire n18245;
   wire n18246;
   wire n18247;
   wire n18248;
   wire n18249;
   wire n18250;
   wire n18251;
   wire n18252;
   wire n18253;
   wire n18254;
   wire n18255;
   wire n18256;
   wire n18257;
   wire n18258;
   wire n18259;
   wire n18260;
   wire n18261;
   wire n18262;
   wire n18263;
   wire n18264;
   wire n18265;
   wire n18267;
   wire n18268;
   wire n18269;
   wire n18270;
   wire n18271;
   wire n18272;
   wire n18273;
   wire n18274;
   wire n18275;
   wire n18276;
   wire n18277;
   wire n18278;
   wire n18279;
   wire n18280;
   wire n18281;
   wire n18282;
   wire n18283;
   wire n18284;
   wire n18286;
   wire n18287;
   wire n18288;
   wire n18289;
   wire n18290;
   wire n18291;
   wire n18292;
   wire n18293;
   wire n18294;
   wire n18295;
   wire n18296;
   wire n18297;
   wire n18298;
   wire n18299;
   wire n18300;
   wire n18301;
   wire n18302;
   wire n18303;
   wire n18304;
   wire n18305;
   wire n18306;
   wire n18307;
   wire n18308;
   wire n18309;
   wire n18311;
   wire n18312;
   wire n18313;
   wire n18314;
   wire n18315;
   wire n18316;
   wire n18317;
   wire n18318;
   wire n18319;
   wire n18320;
   wire n18321;
   wire n18322;
   wire n18323;
   wire n18324;
   wire n18325;
   wire n18326;
   wire n18327;
   wire n18328;
   wire n18329;
   wire n18330;
   wire n18331;
   wire n18332;
   wire n18333;
   wire n18334;
   wire n18335;
   wire n18336;
   wire n18337;
   wire n18338;
   wire n18339;
   wire n18340;
   wire n18341;
   wire n18342;
   wire n18343;
   wire n18344;
   wire n18345;
   wire n18346;
   wire n18347;
   wire n18348;
   wire n18349;
   wire n18351;
   wire n18352;
   wire n18353;
   wire n18354;
   wire n18355;
   wire n18356;
   wire n18357;
   wire n18359;
   wire n18360;
   wire n18361;
   wire n18362;
   wire n18363;
   wire n18364;
   wire n18365;
   wire n18366;
   wire n18367;
   wire n18368;
   wire n18369;
   wire n18370;
   wire n18371;
   wire n18372;
   wire n18373;
   wire n18374;
   wire n18375;
   wire n18376;
   wire n18377;
   wire n18378;
   wire n18379;
   wire n18380;
   wire n18381;
   wire n18382;
   wire n18383;
   wire n18384;
   wire n18385;
   wire n18386;
   wire n18387;
   wire n18388;
   wire n18389;
   wire n18390;
   wire n18391;
   wire n18392;
   wire n18393;
   wire n18394;
   wire n18395;
   wire n18396;
   wire n18397;
   wire n18398;
   wire n18399;
   wire n18400;
   wire n18401;
   wire n18402;
   wire n18403;
   wire n18404;
   wire n18405;
   wire n18406;
   wire n18407;
   wire n18408;
   wire n18409;
   wire n18410;
   wire n18411;
   wire n18412;
   wire n18413;
   wire n18414;
   wire n18415;
   wire n18416;
   wire n18417;
   wire n18418;
   wire n18419;
   wire n18420;
   wire n18421;
   wire n18422;
   wire n18423;
   wire n18424;
   wire n18425;
   wire n18426;
   wire n18427;
   wire n18428;
   wire n18429;
   wire n18430;
   wire n18431;
   wire n18433;
   wire n18434;
   wire n18435;
   wire n18436;
   wire n18437;
   wire n18438;
   wire n18439;
   wire n18441;
   wire n18442;
   wire n18443;
   wire n18444;
   wire n18445;
   wire n18446;
   wire n18447;
   wire n18448;
   wire n18450;
   wire n18451;
   wire n18452;
   wire n18453;
   wire n18454;
   wire n18455;
   wire n18456;
   wire n18457;
   wire n18458;
   wire n18459;
   wire n18460;
   wire n18461;
   wire n18462;
   wire n18463;
   wire n18465;
   wire n18466;
   wire n18467;
   wire n18468;
   wire n18469;
   wire n18470;
   wire n18471;
   wire n18472;
   wire n18473;
   wire n18474;
   wire n18475;
   wire n18476;
   wire n18477;
   wire n18478;
   wire n18479;
   wire n18480;
   wire n18481;
   wire n18482;
   wire n18483;
   wire n18484;
   wire n18485;
   wire n18486;
   wire n18487;
   wire n18488;
   wire n18489;
   wire n18490;
   wire n18491;
   wire n18492;
   wire n18493;
   wire n18494;
   wire n18495;
   wire n18496;
   wire n18497;
   wire n18498;
   wire n18499;
   wire n18500;
   wire n18501;
   wire n18502;
   wire n18503;
   wire n18504;
   wire n18505;
   wire n18506;
   wire n18507;
   wire n18508;
   wire n18509;
   wire n18510;
   wire n18511;
   wire n18512;
   wire n18513;
   wire n18514;
   wire n18515;
   wire n18516;
   wire n18517;
   wire n18518;
   wire n18519;
   wire n18520;
   wire n18521;
   wire n18522;
   wire n18523;
   wire n18524;
   wire n18526;
   wire n18527;
   wire n18528;
   wire n18529;
   wire n18530;
   wire n18531;
   wire n18532;
   wire n18533;
   wire n18534;
   wire n18535;
   wire n18536;
   wire n18537;
   wire n18538;
   wire n18539;
   wire n18540;
   wire n18541;
   wire n18542;
   wire n18543;
   wire n18544;
   wire n18546;
   wire n18547;
   wire n18548;
   wire n18549;
   wire n18550;
   wire n18551;
   wire n18552;
   wire n18553;
   wire n18554;
   wire n18555;
   wire n18556;
   wire n18557;
   wire n18558;
   wire n18559;
   wire n18560;
   wire n18561;
   wire n18562;
   wire n18563;
   wire n18564;
   wire n18565;
   wire n18566;
   wire n18567;
   wire n18568;
   wire n18569;
   wire n18570;
   wire n18571;
   wire n18572;
   wire n18573;
   wire n18574;
   wire n18575;
   wire n18576;
   wire n18577;
   wire n18578;
   wire n18579;
   wire n18580;
   wire n18581;
   wire n18582;
   wire n18583;
   wire n18584;
   wire n18585;
   wire n18586;
   wire n18587;
   wire n18588;
   wire n18589;
   wire n18590;
   wire n18591;
   wire n18592;
   wire n18593;
   wire n18594;
   wire n18595;
   wire n18596;
   wire n18597;
   wire n18598;
   wire n18599;
   wire n18600;
   wire n18601;
   wire n18602;
   wire n18603;
   wire n18604;
   wire n18605;
   wire n18606;
   wire n18607;
   wire n18608;
   wire n18609;
   wire n18610;
   wire n18611;
   wire n18612;
   wire n18613;
   wire n18614;
   wire n18615;
   wire n18616;
   wire n18617;
   wire n18618;
   wire n18619;
   wire n18620;
   wire n18621;
   wire n18622;
   wire n18623;
   wire n18624;
   wire n18625;
   wire n18626;
   wire n18627;
   wire n18628;
   wire n18629;
   wire n18630;
   wire n18631;
   wire n18632;
   wire n18633;
   wire n18634;
   wire n18635;
   wire n18636;
   wire n18637;
   wire n18638;
   wire n18639;
   wire n18640;
   wire n18641;
   wire n18642;
   wire n18643;
   wire n18644;
   wire n18645;
   wire n18646;
   wire n18647;
   wire n18648;
   wire n18649;
   wire n18650;
   wire n18651;
   wire n18652;
   wire n18653;
   wire n18654;
   wire n18655;
   wire n18656;
   wire n18657;
   wire n18658;
   wire n18660;
   wire n18661;
   wire n18662;
   wire n18663;
   wire n18664;
   wire n18665;
   wire n18666;
   wire n18667;
   wire n18668;
   wire n18669;
   wire n18670;
   wire n18671;
   wire n18672;
   wire n18673;
   wire n18674;
   wire n18675;
   wire n18676;
   wire n18677;
   wire n18678;
   wire n18679;
   wire n18680;
   wire n18681;
   wire n18682;
   wire n18683;
   wire n18684;
   wire n18685;
   wire n18686;
   wire n18687;
   wire n18688;
   wire n18689;
   wire n18690;
   wire n18691;
   wire n18692;
   wire n18693;
   wire n18694;
   wire n18695;
   wire n18696;
   wire n18697;
   wire n18698;
   wire n18699;
   wire n18700;
   wire n18701;
   wire n18702;
   wire n18703;
   wire n18704;
   wire n18705;
   wire n18706;
   wire n18707;
   wire n18708;
   wire n18709;
   wire n18710;
   wire n18711;
   wire n18712;
   wire n18713;
   wire n18714;
   wire n18715;
   wire n18716;
   wire n18717;
   wire n18718;
   wire n18719;
   wire n18720;
   wire n18721;
   wire n18722;
   wire n18723;
   wire n18724;
   wire n18725;
   wire n18726;
   wire n18727;
   wire n18728;
   wire n18729;
   wire n18730;
   wire n18731;
   wire n18732;
   wire n18733;
   wire n18734;
   wire n18735;
   wire n18736;
   wire n18737;
   wire n18738;
   wire n18739;
   wire n18740;
   wire n18741;
   wire n18742;
   wire n18743;
   wire n18744;
   wire n18745;
   wire n18746;
   wire n18747;
   wire n18748;
   wire n18749;
   wire n18750;
   wire n18751;
   wire n18752;
   wire n18753;
   wire n18754;
   wire n18755;
   wire n18756;
   wire n18757;
   wire n18758;
   wire n18759;
   wire n18760;
   wire n18761;
   wire n18762;
   wire n18763;
   wire n18764;
   wire n18765;
   wire n18766;
   wire n18767;
   wire n18768;
   wire n18769;
   wire n18770;
   wire n18771;
   wire n18772;
   wire n18773;
   wire n18774;
   wire n18775;
   wire n18776;
   wire n18777;
   wire n18778;
   wire n18779;
   wire n18780;
   wire n18781;
   wire n18782;
   wire n18783;
   wire n18784;
   wire n18785;
   wire n18786;
   wire n18787;
   wire n18788;
   wire n18789;
   wire n18790;
   wire n18791;
   wire n18792;
   wire n18793;
   wire n18794;
   wire n18795;
   wire n18796;
   wire n18797;
   wire n18798;
   wire n18799;
   wire n18800;
   wire n18801;
   wire n18802;
   wire n18803;
   wire n18804;
   wire n18805;
   wire n18806;
   wire n18807;
   wire n18808;
   wire n18809;
   wire n18810;
   wire n18811;
   wire n18812;
   wire n18813;
   wire n18814;
   wire n18815;
   wire n18816;
   wire n18817;
   wire n18818;
   wire n18819;
   wire n18820;
   wire n18821;
   wire n18822;
   wire n18823;
   wire n18824;
   wire n18825;
   wire n18826;
   wire n18827;
   wire n18828;
   wire n18829;
   wire n18830;
   wire n18831;
   wire n18832;
   wire n18833;
   wire n18834;
   wire n18835;
   wire n18836;
   wire n18837;
   wire n18838;
   wire n18839;
   wire n18840;
   wire n18841;
   wire n18842;
   wire n18843;
   wire n18844;
   wire n18845;
   wire n18846;
   wire n18847;
   wire n18848;
   wire n18849;
   wire n18850;
   wire n18851;
   wire n18852;
   wire n18853;
   wire n18854;
   wire n18855;
   wire n18856;
   wire n18857;
   wire n18858;
   wire n18859;
   wire n18860;
   wire n18861;
   wire n18862;
   wire n18863;
   wire n18864;
   wire n18865;
   wire n18866;
   wire n18867;
   wire n18868;
   wire n18869;
   wire n18870;
   wire n18871;
   wire n18872;
   wire n18873;
   wire n18874;
   wire n18875;
   wire n18876;
   wire n18877;
   wire n18878;
   wire n18879;
   wire n18880;
   wire n18881;
   wire n18882;
   wire n18883;
   wire n18884;
   wire n18885;
   wire n18886;
   wire n18887;
   wire n18888;
   wire n18889;
   wire n18890;
   wire n18891;
   wire n18892;
   wire n18893;
   wire n18894;
   wire n18895;
   wire n18896;
   wire n18897;
   wire n18898;
   wire n18899;
   wire n18900;
   wire n18901;
   wire n18902;
   wire n18903;
   wire n18904;
   wire n18905;
   wire n18906;
   wire n18907;
   wire n18908;
   wire n18909;
   wire n18910;
   wire n18911;
   wire n18912;
   wire n18913;
   wire n18914;
   wire n18915;
   wire n18916;
   wire n18917;
   wire n18918;
   wire n18919;
   wire n18920;
   wire n18921;
   wire n18922;
   wire n18923;
   wire n18924;
   wire n18925;
   wire n18926;
   wire n18927;
   wire n18928;
   wire n18929;
   wire n18930;
   wire n18931;
   wire n18932;
   wire n18933;
   wire n18934;
   wire n18936;
   wire n18937;
   wire n18938;
   wire n18939;
   wire n18940;
   wire n18941;
   wire n18942;
   wire n18943;
   wire n18944;
   wire n18945;
   wire n18946;
   wire n18947;
   wire n18948;
   wire n18949;
   wire n18950;
   wire n18951;
   wire n18952;
   wire n18953;
   wire n18954;
   wire n18955;
   wire n18956;
   wire n18957;
   wire n18958;
   wire n18959;
   wire n18960;
   wire n18961;
   wire n18962;
   wire n18963;
   wire n18964;
   wire n18965;
   wire n18966;
   wire n18967;
   wire n18968;
   wire n18970;
   wire n18971;
   wire n18972;
   wire n18973;
   wire n18974;
   wire n18975;
   wire n18976;
   wire n18977;
   wire n18978;
   wire n18979;
   wire n18980;
   wire n18981;
   wire n18983;
   wire n18984;
   wire n18985;
   wire n18986;
   wire n18987;
   wire n18988;
   wire n18989;
   wire n18990;
   wire n18991;
   wire n18992;
   wire n18993;
   wire n18994;
   wire n18995;
   wire n18996;
   wire n18997;
   wire n18998;
   wire n18999;
   wire n19000;
   wire n19001;
   wire n19002;
   wire n19003;
   wire n19004;
   wire n19006;
   wire n19007;
   wire n19009;
   wire n19010;
   wire n19011;
   wire n19012;
   wire n19013;
   wire n19014;
   wire n19015;
   wire n19016;
   wire n19017;
   wire n19018;
   wire n19019;
   wire n19020;
   wire n19021;
   wire n19022;
   wire n19023;
   wire n19024;
   wire n19025;
   wire n19026;
   wire n19027;
   wire n19028;
   wire n19029;
   wire n19030;
   wire n19031;
   wire n19032;
   wire n19033;
   wire n19034;
   wire n19035;
   wire n19036;
   wire n19037;
   wire n19038;
   wire n19039;
   wire n19040;
   wire n19041;
   wire n19042;
   wire n19043;
   wire n19044;
   wire n19045;
   wire n19046;
   wire n19047;
   wire n19048;
   wire n19049;
   wire n19050;
   wire n19051;
   wire n19052;
   wire n19053;
   wire n19054;
   wire n19055;
   wire n19056;
   wire n19057;
   wire n19058;
   wire n19059;
   wire n19060;
   wire n19061;
   wire n19063;
   wire n19066;
   wire n19067;
   wire n19068;
   wire n19069;
   wire n19070;
   wire n19071;
   wire n19072;
   wire n19073;
   wire n19074;
   wire n19075;
   wire n19076;
   wire n19077;
   wire n19078;
   wire n19079;
   wire n19080;
   wire n19081;
   wire n19082;
   wire n19083;
   wire n19084;
   wire n19085;
   wire n19086;
   wire n19087;
   wire n19088;
   wire n19089;
   wire n19090;
   wire n19091;
   wire n19092;
   wire n19093;
   wire n19094;
   wire n19095;
   wire n19096;
   wire n19097;
   wire n19098;
   wire n19099;
   wire n19100;
   wire n19101;
   wire n19102;
   wire n19103;
   wire n19104;
   wire n19105;
   wire n19106;
   wire n19107;
   wire n19108;
   wire n19109;
   wire n19110;
   wire n19111;
   wire n19112;
   wire n19113;
   wire n19114;
   wire n19115;
   wire n19116;
   wire n19117;
   wire n19118;
   wire n19119;
   wire n19120;
   wire n19121;
   wire n19122;
   wire n19123;
   wire n19124;
   wire n19125;
   wire n19126;
   wire n19127;
   wire n19128;
   wire n19129;
   wire n19130;
   wire n19131;
   wire n19132;
   wire n19133;
   wire n19137;
   wire n19138;
   wire n19139;
   wire n19140;
   wire n19141;
   wire n19142;
   wire n19143;
   wire n19144;
   wire n19145;
   wire n19146;
   wire n19147;
   wire n19148;
   wire n19149;
   wire n19150;
   wire n19151;
   wire n19152;
   wire n19153;
   wire n19154;
   wire n19155;
   wire n19156;
   wire n19157;
   wire n19158;
   wire n19159;
   wire n19160;
   wire n19161;
   wire n19162;
   wire n19163;
   wire n19164;
   wire n19165;
   wire n19166;
   wire n19167;
   wire n19168;
   wire n19169;
   wire n19170;
   wire n19171;
   wire n19172;
   wire n19173;
   wire n19174;
   wire n19175;
   wire n19176;
   wire n19177;
   wire n19178;
   wire n19179;
   wire n19180;
   wire n19181;
   wire n19182;
   wire n19183;
   wire n19184;
   wire n19185;
   wire n19186;
   wire n19187;
   wire n19188;
   wire n19189;
   wire n19190;
   wire n19191;
   wire n19192;
   wire n19193;
   wire n19194;
   wire n19195;
   wire n19196;
   wire n19197;
   wire n19198;
   wire n19199;
   wire n19200;
   wire n19201;
   wire n19202;
   wire n19203;
   wire n19204;
   wire n19205;
   wire n19206;
   wire n19207;
   wire n19208;
   wire n19209;
   wire n19210;
   wire n19211;
   wire n19212;
   wire n19213;
   wire n19214;
   wire n19215;
   wire n19216;
   wire n19217;
   wire n19218;
   wire n19219;
   wire n19220;
   wire n19221;
   wire n19222;
   wire n19223;
   wire n19224;
   wire n19225;
   wire n19226;
   wire n19227;
   wire n19228;
   wire n19229;
   wire n19230;
   wire n19231;
   wire n19232;
   wire n19233;
   wire n19234;
   wire n19235;
   wire n19236;
   wire n19237;
   wire n19238;
   wire n19239;
   wire n19240;
   wire n19241;
   wire n19242;
   wire n19243;
   wire n19244;
   wire n19245;
   wire n19246;
   wire n19247;
   wire n19248;
   wire n19249;
   wire n19250;
   wire n19251;
   wire n19252;
   wire n19253;
   wire n19254;
   wire n19255;
   wire n19256;
   wire n19257;
   wire n19258;
   wire n19259;
   wire n19260;
   wire n19261;
   wire n19263;
   wire n19264;
   wire n19265;
   wire n19266;
   wire n19267;
   wire n19268;
   wire n19269;
   wire n19270;
   wire n19271;
   wire n19272;
   wire n19273;
   wire n19274;
   wire n19275;
   wire n19276;
   wire n19277;
   wire n19278;
   wire n19279;
   wire n19280;
   wire n19281;
   wire n19282;
   wire n19283;
   wire n19284;
   wire n19285;
   wire n19286;
   wire n19287;
   wire n19288;
   wire n19289;
   wire n19290;
   wire n19291;
   wire n19292;
   wire n19293;
   wire n19294;
   wire n19295;
   wire n19296;
   wire n19297;
   wire n19298;
   wire n19299;
   wire n19300;
   wire n19301;
   wire n19302;
   wire n19303;
   wire n19304;
   wire n19305;
   wire n19306;
   wire n19307;
   wire n19308;
   wire n19309;
   wire n19310;
   wire n19311;
   wire n19312;
   wire n19313;
   wire n19314;
   wire n19315;
   wire n19316;
   wire n19317;
   wire n19318;
   wire n19319;
   wire n19320;
   wire n19321;
   wire n19322;
   wire n19323;
   wire n19324;
   wire n19325;
   wire n19326;
   wire n19327;
   wire n19328;
   wire n19329;
   wire n19330;
   wire n19331;
   wire n19332;
   wire n19333;
   wire n19334;
   wire n19335;
   wire n19336;
   wire n19337;
   wire n19338;
   wire n19339;
   wire n19340;
   wire n19341;
   wire n19342;
   wire n19343;
   wire n19344;
   wire n19345;
   wire n19346;
   wire n19347;
   wire n19348;
   wire n19349;
   wire n19350;
   wire n19351;
   wire n19352;
   wire n19353;
   wire n19354;
   wire n19355;
   wire n19356;
   wire n19357;
   wire n19358;
   wire n19359;
   wire n19360;
   wire n19361;
   wire n19362;
   wire n19363;
   wire n19364;
   wire n19365;
   wire n19366;
   wire n19367;
   wire n19368;
   wire n19369;
   wire n19370;
   wire n19371;
   wire n19372;
   wire n19373;
   wire n19374;
   wire n19375;
   wire n19376;
   wire n19377;
   wire n19378;
   wire n19379;
   wire n19380;
   wire n19381;
   wire n19382;
   wire n19383;
   wire n19384;
   wire n19385;
   wire n19386;
   wire n19387;
   wire n19388;
   wire n19389;
   wire n19390;
   wire n19391;
   wire n19392;
   wire n19393;
   wire n19394;
   wire n19395;
   wire n19396;
   wire n19397;
   wire n19398;
   wire n19399;
   wire n19400;
   wire n19401;
   wire n19402;
   wire n19403;
   wire n19404;
   wire n19405;
   wire n19406;
   wire n19407;
   wire n19408;
   wire n19409;
   wire n19410;
   wire n19411;
   wire n19412;
   wire n19413;
   wire n19414;
   wire n19415;
   wire n19417;
   wire n19418;
   wire n19419;
   wire n19420;
   wire n19421;
   wire n19422;
   wire n19423;
   wire n19424;
   wire n19425;
   wire n19427;
   wire n19428;
   wire n19429;
   wire n19430;
   wire n19431;
   wire n19432;
   wire n19433;
   wire n19434;
   wire n19435;
   wire n19436;
   wire n19437;
   wire n19438;
   wire n19439;
   wire n19440;
   wire n19441;
   wire n19442;
   wire n19443;
   wire n19444;
   wire n19445;
   wire n19446;
   wire n19447;
   wire n19448;
   wire n19449;
   wire n19450;
   wire n19451;
   wire n19452;
   wire n19453;
   wire n19454;
   wire n19455;
   wire n19456;
   wire n19457;
   wire n19458;
   wire n19459;
   wire n19460;
   wire n19461;
   wire n19462;
   wire n19463;
   wire n19464;
   wire n19465;
   wire n19466;
   wire n19467;
   wire n19468;
   wire n19469;
   wire n19470;
   wire n19471;
   wire n19472;
   wire n19473;
   wire n19474;
   wire n19475;
   wire n19476;
   wire n19477;
   wire n19478;
   wire n19479;
   wire n19480;
   wire n19481;
   wire n19482;
   wire n19483;
   wire n19484;
   wire n19485;
   wire n19486;
   wire n19487;
   wire n19488;
   wire n19489;
   wire n19490;
   wire n19491;
   wire n19492;
   wire n19493;
   wire n19494;
   wire n19495;
   wire n19496;
   wire n19497;
   wire n19498;
   wire n19499;
   wire n19500;
   wire n19501;
   wire n19502;
   wire n19503;
   wire n19504;
   wire n19505;
   wire n19506;
   wire n19507;
   wire n19508;
   wire n19509;
   wire n19510;
   wire n19511;
   wire n19512;
   wire n19513;
   wire n19514;
   wire n19515;
   wire n19516;
   wire n19517;
   wire n19518;
   wire n19519;
   wire n19520;
   wire n19521;
   wire n19523;
   wire n19524;
   wire n19525;
   wire n19526;
   wire n19527;
   wire n19528;
   wire n19530;
   wire n19531;
   wire n19532;
   wire n19533;
   wire n19534;
   wire n19535;
   wire n19536;
   wire n19537;
   wire n19538;
   wire n19539;
   wire n19540;
   wire n19541;
   wire n19542;
   wire n19543;
   wire n19544;
   wire n19545;
   wire n19546;
   wire n19547;
   wire n19548;
   wire n19549;
   wire n19550;
   wire n19551;
   wire n19552;
   wire n19553;
   wire n19554;
   wire n19555;
   wire n19556;
   wire n19557;
   wire n19558;
   wire n19559;
   wire n19560;
   wire n19561;
   wire n19562;
   wire n19563;
   wire n19564;
   wire n19565;
   wire n19566;
   wire n19567;
   wire n19568;
   wire n19569;
   wire n19570;
   wire n19571;
   wire n19572;
   wire n19573;
   wire n19574;
   wire n19575;
   wire n19576;
   wire n19577;
   wire n19578;
   wire n19579;
   wire n19580;
   wire n19581;
   wire n19582;
   wire n19583;
   wire n19584;
   wire n19585;
   wire n19586;
   wire n19587;
   wire n19588;
   wire n19589;
   wire n19590;
   wire n19591;
   wire n19592;
   wire n19593;
   wire n19594;
   wire n19595;
   wire n19596;
   wire n19597;
   wire n19598;
   wire n19600;
   wire n19601;
   wire n19602;
   wire n19603;
   wire n19604;
   wire n19605;
   wire n19606;
   wire n19607;
   wire n19608;
   wire n19609;
   wire n19610;
   wire n19611;
   wire n19612;
   wire n19613;
   wire n19614;
   wire n19615;
   wire n19616;
   wire n19617;
   wire n19618;
   wire n19619;
   wire n19620;
   wire n19621;
   wire n19622;
   wire n19623;
   wire n19624;
   wire n19625;
   wire n19627;
   wire n19628;
   wire n19629;
   wire n19630;
   wire n19632;
   wire n19633;
   wire n19634;
   wire n19635;
   wire n19636;
   wire n19637;
   wire n19638;
   wire n19639;
   wire n19640;
   wire n19641;
   wire n19642;
   wire n19643;
   wire n19644;
   wire n19645;
   wire n19646;
   wire n19647;
   wire n19648;
   wire n19649;
   wire n19650;
   wire n19651;
   wire n19652;
   wire n19653;
   wire n19654;
   wire n19655;
   wire n19656;
   wire n19657;
   wire n19658;
   wire n19659;
   wire n19660;
   wire n19661;
   wire n19662;
   wire n19663;
   wire n19664;
   wire n19665;
   wire n19666;
   wire n19667;
   wire n19668;
   wire n19669;
   wire n19670;
   wire n19671;
   wire n19672;
   wire n19673;
   wire n19674;
   wire n19675;
   wire n19676;
   wire n19677;
   wire n19678;
   wire n19679;
   wire n19680;
   wire n19681;
   wire n19682;
   wire n19683;
   wire n19684;
   wire n19685;
   wire n19686;
   wire n19687;
   wire n19688;
   wire n19689;
   wire n19690;
   wire n19691;
   wire n19692;
   wire n19693;
   wire n19694;
   wire n19695;
   wire n19696;
   wire n19697;
   wire n19698;
   wire n19699;
   wire n19700;
   wire n19701;
   wire n19702;
   wire n19703;
   wire n19704;
   wire n19706;
   wire n19707;
   wire n19708;
   wire n19709;
   wire n19710;
   wire n19711;
   wire n19712;
   wire n19713;
   wire n19714;
   wire n19715;
   wire n19716;
   wire n19717;
   wire n19718;
   wire n19719;
   wire n19720;
   wire n19721;
   wire n19722;
   wire n19723;
   wire n19724;
   wire n19725;
   wire n19726;
   wire n19727;
   wire n19728;
   wire n19729;
   wire n19730;
   wire n19731;
   wire n19732;
   wire n19733;
   wire n19734;
   wire n19735;
   wire n19736;
   wire n19737;
   wire n19738;
   wire n19739;
   wire n19740;
   wire n19741;
   wire n19742;
   wire n19743;
   wire n19744;
   wire n19745;
   wire n19746;
   wire n19747;
   wire n19748;
   wire n19749;
   wire n19750;
   wire n19751;
   wire n19752;
   wire n19753;
   wire n19754;
   wire n19755;
   wire n19756;
   wire n19758;
   wire n19759;
   wire n19760;
   wire n19761;
   wire n19762;
   wire n19763;
   wire n19764;
   wire n19765;
   wire n19766;
   wire n19767;
   wire n19768;
   wire n19769;
   wire n19770;
   wire n19771;
   wire n19772;
   wire n19773;
   wire n19774;
   wire n19775;
   wire n19776;
   wire n19777;
   wire n19778;
   wire n19779;
   wire n19781;
   wire n19782;
   wire n19783;
   wire n19784;
   wire n19785;
   wire n19786;
   wire n19787;
   wire n19788;
   wire n19789;
   wire n19790;
   wire n19791;
   wire n19792;
   wire n19793;
   wire n19794;
   wire n19795;
   wire n19796;
   wire n19797;
   wire n19798;
   wire n19799;
   wire n19800;
   wire n19801;
   wire n19802;
   wire n19803;
   wire n19804;
   wire n19805;
   wire n19807;
   wire n19808;
   wire n19809;
   wire n19810;
   wire n19811;
   wire n19812;
   wire n19813;
   wire n19814;
   wire n19815;
   wire n19816;
   wire n19817;
   wire n19818;
   wire n19819;
   wire n19820;
   wire n19821;
   wire n19822;
   wire n19823;
   wire n19824;
   wire n19825;
   wire n19826;
   wire n19827;
   wire n19828;
   wire n19829;
   wire n19830;
   wire n19831;
   wire n19832;
   wire n19833;
   wire n19834;
   wire n19835;
   wire n19836;
   wire n19837;
   wire n19838;
   wire n19839;
   wire n19840;
   wire n19841;
   wire n19842;
   wire n19843;
   wire n19844;
   wire n19845;
   wire n19846;
   wire n19847;
   wire n19848;
   wire n19849;
   wire n19850;
   wire n19851;
   wire n19852;
   wire n19853;
   wire n19854;
   wire n19855;
   wire n19856;
   wire n19857;
   wire n19858;
   wire n19859;
   wire n19860;
   wire n19861;
   wire n19862;
   wire n19863;
   wire n19864;
   wire n19865;
   wire n19866;
   wire n19867;
   wire n19868;
   wire n19869;
   wire n19870;
   wire n19871;
   wire n19872;
   wire n19873;
   wire n19874;
   wire n19875;
   wire n19876;
   wire n19877;
   wire n19878;
   wire n19879;
   wire n19880;
   wire n19881;
   wire n19882;
   wire n19883;
   wire n19884;
   wire n19885;
   wire n19886;
   wire n19887;
   wire n19888;
   wire n19889;
   wire n19890;
   wire n19892;
   wire n19893;
   wire n19894;
   wire n19895;
   wire n19896;
   wire n19897;
   wire n19898;
   wire n19899;
   wire n19900;
   wire n19901;
   wire n19902;
   wire n19903;
   wire n19904;
   wire n19905;
   wire n19906;
   wire n19907;
   wire n19908;
   wire n19909;
   wire n19910;
   wire n19911;
   wire n19913;
   wire n19914;
   wire n19915;
   wire n19916;
   wire n19917;
   wire n19918;
   wire n19919;
   wire n19920;
   wire n19921;
   wire n19922;
   wire n19923;
   wire n19924;
   wire n19925;
   wire n19926;
   wire n19927;
   wire n19928;
   wire n19929;
   wire n19930;
   wire n19932;
   wire n19933;
   wire n19934;
   wire n19935;
   wire n19936;
   wire n19937;
   wire n19938;
   wire n19940;
   wire n19941;
   wire n19942;
   wire n19943;
   wire n19944;
   wire n19945;
   wire n19946;
   wire n19947;
   wire n19948;
   wire n19949;
   wire n19950;
   wire n19951;
   wire n19953;
   wire n19954;
   wire n19955;
   wire n19956;
   wire n19957;
   wire n19958;
   wire n19959;
   wire n19961;
   wire n19962;
   wire n19963;
   wire n19964;
   wire n19965;
   wire n19966;
   wire n19967;
   wire n19968;
   wire n19969;
   wire n19970;
   wire n19971;
   wire n19972;
   wire n19973;
   wire n19974;
   wire n19975;
   wire n19976;
   wire n19977;
   wire n19978;
   wire n19979;
   wire n19981;
   wire n19982;
   wire n19983;
   wire n19984;
   wire n19985;
   wire n19986;
   wire n19987;
   wire n19988;
   wire n19989;
   wire n19990;
   wire n19991;
   wire n19992;
   wire n19993;
   wire n19994;
   wire n19995;
   wire n19996;
   wire n19997;
   wire n19998;
   wire n19999;
   wire n20000;
   wire n20001;
   wire n20002;
   wire n20003;
   wire n20004;
   wire n20005;
   wire n20006;
   wire n20007;
   wire n20008;
   wire n20009;
   wire n20010;
   wire n20011;
   wire n20012;
   wire n20013;
   wire n20014;
   wire n20015;
   wire n20016;
   wire n20017;
   wire n20018;
   wire n20019;
   wire n20020;
   wire n20021;
   wire n20022;
   wire n20023;
   wire n20024;
   wire n20026;
   wire n20027;
   wire n20028;
   wire n20030;
   wire n20031;
   wire n20032;
   wire n20033;
   wire n20034;
   wire n20035;
   wire n20036;
   wire n20037;
   wire n20038;
   wire n20039;
   wire n20040;
   wire n20041;
   wire n20042;
   wire n20043;
   wire n20044;
   wire n20045;
   wire n20046;
   wire n20047;
   wire n20048;
   wire n20049;
   wire n20050;
   wire n20051;
   wire n20052;
   wire n20053;
   wire n20054;
   wire n20055;
   wire n20056;
   wire n20057;
   wire n20058;
   wire n20059;
   wire n20060;
   wire n20061;
   wire n20062;
   wire n20063;
   wire n20064;
   wire n20065;
   wire n20066;
   wire n20067;
   wire n20068;
   wire n20069;
   wire n20070;
   wire n20071;
   wire n20072;
   wire n20073;
   wire n20074;
   wire n20075;
   wire n20076;
   wire n20077;
   wire n20078;
   wire n20079;
   wire n20080;
   wire n20081;
   wire n20082;
   wire n20083;
   wire n20084;
   wire n20085;
   wire n20086;
   wire n20087;
   wire n20088;
   wire n20089;
   wire n20090;
   wire n20091;
   wire n20092;
   wire n20093;
   wire n20094;
   wire n20095;
   wire n20096;
   wire n20097;
   wire n20098;
   wire n20099;
   wire n20100;
   wire n20101;
   wire n20102;
   wire n20103;
   wire n20104;
   wire n20105;
   wire n20106;
   wire n20107;
   wire n20108;
   wire n20109;
   wire n20110;
   wire n20111;
   wire n20112;
   wire n20113;
   wire n20114;
   wire n20115;
   wire n20116;
   wire n20117;
   wire n20118;
   wire n20119;
   wire n20120;
   wire n20121;
   wire n20122;
   wire n20123;
   wire n20124;
   wire n20125;
   wire n20126;
   wire n20127;
   wire n20128;
   wire n20129;
   wire n20130;
   wire n20131;
   wire n20132;
   wire n20133;
   wire n20134;
   wire n20135;
   wire n20136;
   wire n20137;
   wire n20138;
   wire n20139;
   wire n20140;
   wire n20141;
   wire n20142;
   wire n20143;
   wire n20144;
   wire n20145;
   wire n20146;
   wire n20147;
   wire n20148;
   wire n20149;
   wire n20150;
   wire n20151;
   wire n20152;
   wire n20153;
   wire n20154;
   wire n20155;
   wire n20156;
   wire n20157;
   wire n20158;
   wire n20159;
   wire n20160;
   wire n20161;
   wire n20162;
   wire n20163;
   wire n20164;
   wire n20165;
   wire n20166;
   wire n20167;
   wire n20168;
   wire n20169;
   wire n20170;
   wire n20171;
   wire n20172;
   wire n20173;
   wire n20174;
   wire n20175;
   wire n20176;
   wire n20177;
   wire n20178;
   wire n20179;
   wire n20180;
   wire n20181;
   wire n20182;
   wire n20183;
   wire n20184;
   wire n20185;
   wire n20186;
   wire n20187;
   wire n20188;
   wire n20189;
   wire n20190;
   wire n20191;
   wire n20192;
   wire n20193;
   wire n20194;
   wire n20195;
   wire n20196;
   wire n20197;
   wire n20198;
   wire n20199;
   wire n20200;
   wire n20201;
   wire n20202;
   wire n20203;
   wire n20204;
   wire n20205;
   wire n20206;
   wire n20208;
   wire n20209;
   wire n20210;
   wire n20211;
   wire n20212;
   wire n20213;
   wire n20214;
   wire n20216;
   wire n20217;
   wire n20218;
   wire n20219;
   wire n20220;
   wire n20221;
   wire n20222;
   wire n20223;
   wire n20224;
   wire n20225;
   wire n20226;
   wire n20227;
   wire n20228;
   wire n20229;
   wire n20230;
   wire n20231;
   wire n20232;
   wire n20233;
   wire n20234;
   wire n20235;
   wire n20236;
   wire n20237;
   wire n20238;
   wire n20239;
   wire n20240;
   wire n20241;
   wire n20242;
   wire n20243;
   wire n20244;
   wire n20245;
   wire n20246;
   wire n20247;
   wire n20248;
   wire n20249;
   wire n20250;
   wire n20251;
   wire n20252;
   wire n20253;
   wire n20254;
   wire n20255;
   wire n20256;
   wire n20257;
   wire n20258;
   wire n20259;
   wire n20260;
   wire n20261;
   wire n20262;
   wire n20263;
   wire n20264;
   wire n20265;
   wire n20266;
   wire n20267;
   wire n20268;
   wire n20269;
   wire n20270;
   wire n20271;
   wire n20272;
   wire n20273;
   wire n20274;
   wire n20275;
   wire n20276;
   wire n20277;
   wire n20278;
   wire n20279;
   wire n20280;
   wire n20281;
   wire n20282;
   wire n20283;
   wire n20284;
   wire n20285;
   wire n20286;
   wire n20287;
   wire n20288;
   wire n20289;
   wire n20290;
   wire n20291;
   wire n20292;
   wire n20293;
   wire n20294;
   wire n20295;
   wire n20296;
   wire n20297;
   wire n20298;
   wire n20299;
   wire n20300;
   wire n20301;
   wire n20302;
   wire n20303;
   wire n20304;
   wire n20305;
   wire n20306;
   wire n20307;
   wire n20308;
   wire n20309;
   wire n20310;
   wire n20311;
   wire n20312;
   wire n20313;
   wire n20314;
   wire n20315;
   wire n20316;
   wire n20317;
   wire n20318;
   wire n20319;
   wire n20320;
   wire n20321;
   wire n20322;
   wire n20323;
   wire n20324;
   wire n20325;
   wire n20326;
   wire n20327;
   wire n20328;
   wire n20329;
   wire n20330;
   wire n20331;
   wire n20332;
   wire n20333;
   wire n20334;
   wire n20335;
   wire n20336;
   wire n20337;
   wire n20338;
   wire n20339;
   wire n20340;
   wire n20341;
   wire n20342;
   wire n20343;
   wire n20344;
   wire n20345;
   wire n20346;
   wire n20347;
   wire n20348;
   wire n20349;
   wire n20350;
   wire n20351;
   wire n20352;
   wire n20353;
   wire n20354;
   wire n20355;
   wire n20356;
   wire n20357;
   wire n20358;
   wire n20359;
   wire n20360;
   wire n20361;
   wire n20362;
   wire n20363;
   wire n20364;
   wire n20365;
   wire n20366;
   wire n20367;
   wire n20368;
   wire n20369;
   wire n20370;
   wire n20371;
   wire n20373;
   wire n20374;
   wire n20375;
   wire n20376;
   wire n20377;
   wire n20378;
   wire n20379;
   wire n20380;
   wire n20381;
   wire n20382;
   wire n20383;
   wire n20384;
   wire n20385;
   wire n20386;
   wire n20387;
   wire n20388;
   wire n20389;
   wire n20390;
   wire n20391;
   wire n20392;
   wire n20393;
   wire n20394;
   wire n20395;
   wire n20396;
   wire n20397;
   wire n20398;
   wire n20399;
   wire n20400;
   wire n20401;
   wire n20402;
   wire n20403;
   wire n20404;
   wire n20405;
   wire n20406;
   wire n20407;
   wire n20408;
   wire n20409;
   wire n20410;
   wire n20411;
   wire n20412;
   wire n20413;
   wire n20414;
   wire n20415;
   wire n20416;
   wire n20417;
   wire n20418;
   wire n20419;
   wire n20420;
   wire n20421;
   wire n20422;
   wire n20423;
   wire n20424;
   wire n20425;
   wire n20426;
   wire n20427;
   wire n20428;
   wire n20429;
   wire n20430;
   wire n20431;
   wire n20432;
   wire n20433;
   wire n20434;
   wire n20435;
   wire n20436;
   wire n20437;
   wire n20438;
   wire n20439;
   wire n20440;
   wire n20441;
   wire n20442;
   wire n20443;
   wire n20444;
   wire n20445;
   wire n20446;
   wire n20447;
   wire n20448;
   wire n20449;
   wire n20450;
   wire n20451;
   wire n20452;
   wire n20453;
   wire n20454;
   wire n20455;
   wire n20456;
   wire n20457;
   wire n20458;
   wire n20459;
   wire n20460;
   wire n20461;
   wire n20462;
   wire n20463;
   wire n20464;
   wire n20465;
   wire n20466;
   wire n20467;
   wire n20468;
   wire n20469;
   wire n20470;
   wire n20471;
   wire n20472;
   wire n20473;
   wire n20474;
   wire n20475;
   wire n20476;
   wire n20477;
   wire n20478;
   wire n20479;
   wire n20480;
   wire n20481;
   wire n20482;
   wire n20483;
   wire n20484;
   wire n20485;
   wire n20486;
   wire n20487;
   wire n20488;
   wire n20489;
   wire n20490;
   wire n20491;
   wire n20492;
   wire n20493;
   wire n20494;
   wire n20495;
   wire n20496;
   wire n20497;
   wire n20498;
   wire n20499;
   wire n20500;
   wire n20501;
   wire n20502;
   wire n20503;
   wire n20504;
   wire n20505;
   wire n20506;
   wire n20507;
   wire n20509;
   wire n20510;
   wire n20512;
   wire n20513;
   wire n20514;
   wire n20515;
   wire n20516;
   wire n20517;
   wire n20518;
   wire n20519;
   wire n20520;
   wire n20521;
   wire n20522;
   wire n20523;
   wire n20524;
   wire n20525;
   wire n20526;
   wire n20527;
   wire n20528;
   wire n20529;
   wire n20530;
   wire n20531;
   wire n20532;
   wire n20533;
   wire n20534;
   wire n20535;
   wire n20536;
   wire n20537;
   wire n20538;
   wire n20539;
   wire n20540;
   wire n20541;
   wire n20542;
   wire n20543;
   wire n20544;
   wire n20545;
   wire n20546;
   wire n20547;
   wire n20548;
   wire n20549;
   wire n20550;
   wire n20551;
   wire n20552;
   wire n20553;
   wire n20554;
   wire n20555;
   wire n20556;
   wire n20557;
   wire n20558;
   wire n20559;
   wire n20560;
   wire n20561;
   wire n20562;
   wire n20563;
   wire n20564;
   wire n20565;
   wire n20566;
   wire n20567;
   wire n20568;
   wire n20569;
   wire n20570;
   wire n20571;
   wire n20572;
   wire n20573;
   wire n20574;
   wire n20575;
   wire n20576;
   wire n20577;
   wire n20578;
   wire n20579;
   wire n20580;
   wire n20581;
   wire n20582;
   wire n20583;
   wire n20584;
   wire n20585;
   wire n20588;
   wire n20589;
   wire n20590;
   wire n20591;
   wire n20592;
   wire n20593;
   wire n20594;
   wire n20595;
   wire n20596;
   wire n20597;
   wire n20598;
   wire n20599;
   wire n20600;
   wire n20601;
   wire n20602;
   wire n20603;
   wire n20604;
   wire n20605;
   wire n20606;
   wire n20607;
   wire n20608;
   wire n20609;
   wire n20610;
   wire n20611;
   wire n20612;
   wire n20613;
   wire n20614;
   wire n20615;
   wire n20616;
   wire n20617;
   wire n20618;
   wire n20619;
   wire n20620;
   wire n20621;
   wire n20622;
   wire n20623;
   wire n20624;
   wire n20625;
   wire n20626;
   wire n20627;
   wire n20628;
   wire n20629;
   wire n20630;
   wire n20631;
   wire n20632;
   wire n20633;
   wire n20634;
   wire n20635;
   wire n20636;
   wire n20637;
   wire n20638;
   wire n20639;
   wire n20640;
   wire n20641;
   wire n20642;
   wire n20643;
   wire n20644;
   wire n20645;
   wire n20646;
   wire n20647;
   wire n20648;
   wire n20649;
   wire n20650;
   wire n20651;
   wire n20652;
   wire n20653;
   wire n20654;
   wire n20655;
   wire n20656;
   wire n20657;
   wire n20658;
   wire n20659;
   wire n20660;
   wire n20661;
   wire n20662;
   wire n20663;
   wire n20664;
   wire n20665;
   wire n20666;
   wire n20667;
   wire n20668;
   wire n20669;
   wire n20670;
   wire n20671;
   wire n20672;
   wire n20673;
   wire n20674;
   wire n20675;
   wire n20676;
   wire n20677;
   wire n20678;
   wire n20679;
   wire n20680;
   wire n20681;
   wire n20682;
   wire n20683;
   wire n20684;
   wire n20685;
   wire n20686;
   wire n20687;
   wire n20688;
   wire n20689;
   wire n20690;
   wire n20691;
   wire n20692;
   wire n20693;
   wire n20694;
   wire n20695;
   wire n20696;
   wire n20697;
   wire n20698;
   wire n20699;
   wire n20700;
   wire n20701;
   wire n20702;
   wire n20703;
   wire n20704;
   wire n20705;
   wire n20706;
   wire n20707;
   wire n20708;
   wire n20709;
   wire n20710;
   wire n20711;
   wire n20712;
   wire n20713;
   wire n20714;
   wire n20715;
   wire n20717;
   wire n20718;
   wire n20719;
   wire n20720;
   wire n20721;
   wire n20722;
   wire n20723;
   wire n20724;
   wire n20725;
   wire n20726;
   wire n20727;
   wire n20728;
   wire n20729;
   wire n20730;
   wire n20731;
   wire n20732;
   wire n20733;
   wire n20734;
   wire n20735;
   wire n20736;
   wire n20737;
   wire n20738;
   wire n20739;
   wire n20740;
   wire n20741;
   wire n20742;
   wire n20743;
   wire n20744;
   wire n20745;
   wire n20746;
   wire n20747;
   wire n20748;
   wire n20749;
   wire n20750;
   wire n20751;
   wire n20752;
   wire n20753;
   wire n20754;
   wire n20755;
   wire n20756;
   wire n20757;
   wire n20758;
   wire n20759;
   wire n20760;
   wire n20761;
   wire n20762;
   wire n20763;
   wire n20764;
   wire n20765;
   wire n20766;
   wire n20767;
   wire n20768;
   wire n20769;
   wire n20770;
   wire n20771;
   wire n20772;
   wire n20773;
   wire n20774;
   wire n20775;
   wire n20776;
   wire n20777;
   wire n20778;
   wire n20779;
   wire n20780;
   wire n20781;
   wire n20782;
   wire n20783;
   wire n20784;
   wire n20785;
   wire n20786;
   wire n20787;
   wire n20788;
   wire n20789;
   wire n20790;
   wire n20791;
   wire n20792;
   wire n20793;
   wire n20794;
   wire n20795;
   wire n20796;
   wire n20797;
   wire n20798;
   wire n20799;
   wire n20800;
   wire n20801;
   wire n20802;
   wire n20803;
   wire n20804;
   wire n20805;
   wire n20806;
   wire n20809;
   wire n20810;
   wire n20811;
   wire n20812;
   wire n20813;
   wire n20814;
   wire n20815;
   wire n20816;
   wire n20817;
   wire n20818;
   wire n20819;
   wire n20820;
   wire n20821;
   wire n20822;
   wire n20823;
   wire n20824;
   wire n20825;
   wire n20826;
   wire n20827;
   wire n20828;
   wire n20829;
   wire n20830;
   wire n20831;
   wire n20832;
   wire n20833;
   wire n20834;
   wire n20835;
   wire n20836;
   wire n20837;
   wire n20838;
   wire n20839;
   wire n20840;
   wire n20841;
   wire n20842;
   wire n20843;
   wire n20844;
   wire n20845;
   wire n20846;
   wire n20847;
   wire n20848;
   wire n20849;
   wire n20850;
   wire n20851;
   wire n20852;
   wire n20853;
   wire n20854;
   wire n20855;
   wire n20856;
   wire n20857;
   wire n20858;
   wire n20859;
   wire n20860;
   wire n20861;
   wire n20862;
   wire n20863;
   wire n20864;
   wire n20865;
   wire n20866;
   wire n20867;
   wire n20868;
   wire n20870;
   wire n20871;
   wire n20872;
   wire n20873;
   wire n20874;
   wire n20875;
   wire n20876;
   wire n20877;
   wire n20878;
   wire n20879;
   wire n20880;
   wire n20881;
   wire n20882;
   wire n20883;
   wire n20884;
   wire n20885;
   wire n20887;
   wire n20888;
   wire n20889;
   wire n20890;
   wire n20891;
   wire n20892;
   wire n20893;
   wire n20894;
   wire n20895;
   wire n20896;
   wire n20897;
   wire n20898;
   wire n20899;
   wire n20900;
   wire n20901;
   wire n20902;
   wire n20903;
   wire n20904;
   wire n20905;
   wire n20907;
   wire n20908;
   wire n20909;
   wire n20910;
   wire n20911;
   wire n20912;
   wire n20913;
   wire n20914;
   wire n20915;
   wire n20916;
   wire n20917;
   wire n20918;
   wire n20919;
   wire n20920;
   wire n20921;
   wire n20922;
   wire n20923;
   wire n20924;
   wire n20925;
   wire n20926;
   wire n20927;
   wire n20928;
   wire n20929;
   wire n20930;
   wire n20931;
   wire n20932;
   wire n20933;
   wire n20934;
   wire n20935;
   wire n20936;
   wire n20937;
   wire n20938;
   wire n20939;
   wire n20940;
   wire n20941;
   wire n20942;
   wire n20943;
   wire n20944;
   wire n20945;
   wire n20946;
   wire n20947;
   wire n20948;
   wire n20949;
   wire n20950;
   wire n20951;
   wire n20952;
   wire n20953;
   wire n20954;
   wire n20955;
   wire n20956;
   wire n20957;
   wire n20958;
   wire n20959;
   wire n20960;
   wire n20961;
   wire n20962;
   wire n20963;
   wire n20964;
   wire n20965;
   wire n20966;
   wire n20967;
   wire n20968;
   wire n20969;
   wire n20970;
   wire n20971;
   wire n20972;
   wire n20973;
   wire n20974;
   wire n20975;
   wire n20976;
   wire n20977;
   wire n20978;
   wire n20979;
   wire n20980;
   wire n20981;
   wire n20982;
   wire n20983;
   wire n20984;
   wire n20985;
   wire n20986;
   wire n20987;
   wire n20988;
   wire n20989;
   wire n20990;
   wire n20991;
   wire n20992;
   wire n20993;
   wire n20994;
   wire n20995;
   wire n20996;
   wire n20997;
   wire n20998;
   wire n20999;
   wire n21000;
   wire n21001;
   wire n21002;
   wire n21003;
   wire n21004;
   wire n21005;
   wire n21006;
   wire n21007;
   wire n21008;
   wire n21009;
   wire n21010;
   wire n21011;
   wire n21012;
   wire n21013;
   wire n21014;
   wire n21015;
   wire n21016;
   wire n21017;
   wire n21018;
   wire n21019;
   wire n21020;
   wire n21021;
   wire n21022;
   wire n21023;
   wire n21024;
   wire n21025;
   wire n21026;
   wire n21027;
   wire n21029;
   wire n21030;
   wire n21031;
   wire n21032;
   wire n21033;
   wire n21034;
   wire n21035;
   wire n21037;
   wire n21038;
   wire n21039;
   wire n21040;
   wire n21041;
   wire n21042;
   wire n21043;
   wire n21044;
   wire n21045;
   wire n21046;
   wire n21047;
   wire n21048;
   wire n21049;
   wire n21050;
   wire n21051;
   wire n21052;
   wire n21053;
   wire n21054;
   wire n21055;
   wire n21056;
   wire n21058;
   wire n21059;
   wire n21060;
   wire n21061;
   wire n21062;
   wire n21063;
   wire n21064;
   wire n21065;
   wire n21066;
   wire n21067;
   wire n21068;
   wire n21069;
   wire n21070;
   wire n21071;
   wire n21072;
   wire n21073;
   wire n21074;
   wire n21076;
   wire n21077;
   wire n21078;
   wire n21079;
   wire n21080;
   wire n21081;
   wire n21082;
   wire n21083;
   wire n21084;
   wire n21085;
   wire n21086;
   wire n21087;
   wire n21088;
   wire n21089;
   wire n21090;
   wire n21091;
   wire n21092;
   wire n21093;
   wire n21094;
   wire n21095;
   wire n21096;
   wire n21097;
   wire n21098;
   wire n21099;
   wire n21100;
   wire n21101;
   wire n21102;
   wire n21103;
   wire n21104;
   wire n21105;
   wire n21106;
   wire n21107;
   wire n21108;
   wire n21109;
   wire n21110;
   wire n21111;
   wire n21112;
   wire n21113;
   wire n21114;
   wire n21115;
   wire n21116;
   wire n21117;
   wire n21118;
   wire n21119;
   wire n21120;
   wire n21121;
   wire n21122;
   wire n21123;
   wire n21124;
   wire n21125;
   wire n21126;
   wire n21127;
   wire n21128;
   wire n21129;
   wire n21130;
   wire n21131;
   wire n21132;
   wire n21133;
   wire n21134;
   wire n21135;
   wire n21136;
   wire n21137;
   wire n21138;
   wire n21140;
   wire n21141;
   wire n21143;
   wire n21144;
   wire n21145;
   wire n21146;
   wire n21147;
   wire n21148;
   wire n21149;
   wire n21150;
   wire n21151;
   wire n21152;
   wire n21153;
   wire n21154;
   wire n21155;
   wire n21156;
   wire n21157;
   wire n21158;
   wire n21159;
   wire n21160;
   wire n21161;
   wire n21162;
   wire n21163;
   wire n21164;
   wire n21165;
   wire n21166;
   wire n21167;
   wire n21168;
   wire n21169;
   wire n21170;
   wire n21171;
   wire n21172;
   wire n21173;
   wire n21174;
   wire n21175;
   wire n21176;
   wire n21177;
   wire n21178;
   wire n21179;
   wire n21180;
   wire n21181;
   wire n21182;
   wire n21183;
   wire n21184;
   wire n21185;
   wire n21186;
   wire n21187;
   wire n21188;
   wire n21189;
   wire n21190;
   wire n21191;
   wire n21192;
   wire n21193;
   wire n21194;
   wire n21195;
   wire n21196;
   wire n21197;
   wire n21198;
   wire n21199;
   wire n21200;
   wire n21201;
   wire n21202;
   wire n21203;
   wire n21204;
   wire n21205;
   wire n21206;
   wire n21207;
   wire n21208;
   wire n21209;
   wire n21210;
   wire n21212;
   wire n21213;
   wire n21214;
   wire n21215;
   wire n21216;
   wire n21217;
   wire n21218;
   wire n21219;
   wire n21220;
   wire n21221;
   wire n21222;
   wire n21223;
   wire n21224;
   wire n21225;
   wire n21226;
   wire n21227;
   wire n21228;
   wire n21229;
   wire n21230;
   wire n21231;
   wire n21232;
   wire n21233;
   wire n21234;
   wire n21235;
   wire n21236;
   wire n21237;
   wire n21238;
   wire n21239;
   wire n21240;
   wire n21241;
   wire n21242;
   wire n21243;
   wire n21244;
   wire n21245;
   wire n21246;
   wire n21247;
   wire n21248;
   wire n21249;
   wire n21250;
   wire n21251;
   wire n21252;
   wire n21253;
   wire n21254;
   wire n21255;
   wire n21256;
   wire n21257;
   wire n21258;
   wire n21259;
   wire n21260;
   wire n21261;
   wire n21262;
   wire n21263;
   wire n21264;
   wire n21265;
   wire n21266;
   wire n21267;
   wire n21268;
   wire n21269;
   wire n21270;
   wire n21271;
   wire n21272;
   wire n21273;
   wire n21274;
   wire n21275;
   wire n21276;
   wire n21277;
   wire n21278;
   wire n21279;
   wire n21280;
   wire n21281;
   wire n21282;
   wire n21283;
   wire n21284;
   wire n21285;
   wire n21286;
   wire n21287;
   wire n21288;
   wire n21289;
   wire n21290;
   wire n21291;
   wire n21292;
   wire n21293;
   wire n21294;
   wire n21295;
   wire n21296;
   wire n21297;
   wire n21298;
   wire n21299;
   wire n21300;
   wire n21301;
   wire n21302;
   wire n21303;
   wire n21304;
   wire n21305;
   wire n21306;
   wire n21307;
   wire n21308;
   wire n21309;
   wire n21310;
   wire n21311;
   wire n21312;
   wire n21313;
   wire n21314;
   wire n21315;
   wire n21316;
   wire n21317;
   wire n21318;
   wire n21319;
   wire n21320;
   wire n21321;
   wire n21322;
   wire n21323;
   wire n21324;
   wire n21325;
   wire n21326;
   wire n21327;
   wire n21328;
   wire n21329;
   wire n21330;
   wire n21331;
   wire n21332;
   wire n21333;
   wire n21334;
   wire n21335;
   wire n21336;
   wire n21337;
   wire n21338;
   wire n21339;
   wire n21340;
   wire n21341;
   wire n21342;
   wire n21343;
   wire n21344;
   wire n21345;
   wire n21346;
   wire n21347;
   wire n21348;
   wire n21349;
   wire n21350;
   wire n21351;
   wire n21352;
   wire n21353;
   wire n21354;
   wire n21355;
   wire n21356;
   wire n21357;
   wire n21358;
   wire n21359;
   wire n21360;
   wire n21361;
   wire n21362;
   wire n21363;
   wire n21364;
   wire n21365;
   wire n21366;
   wire n21367;
   wire n21368;
   wire n21369;
   wire n21370;
   wire n21371;
   wire n21372;
   wire n21373;
   wire n21374;
   wire n21375;
   wire n21376;
   wire n21377;
   wire n21378;
   wire n21379;
   wire n21380;
   wire n21381;
   wire n21382;
   wire n21383;
   wire n21384;
   wire n21385;
   wire n21386;
   wire n21387;
   wire n21388;
   wire n21389;
   wire n21390;
   wire n21391;
   wire n21393;
   wire n21394;
   wire n21395;
   wire n21396;
   wire n21397;
   wire n21398;
   wire n21399;
   wire n21400;
   wire n21401;
   wire n21402;
   wire n21403;
   wire n21404;
   wire n21405;
   wire n21406;
   wire n21407;
   wire n21408;
   wire n21409;
   wire n21410;
   wire n21411;
   wire n21412;
   wire n21413;
   wire n21414;
   wire n21415;
   wire n21416;
   wire n21417;
   wire n21418;
   wire n21419;
   wire n21420;
   wire n21421;
   wire n21422;
   wire n21423;
   wire n21424;
   wire n21425;
   wire n21426;
   wire n21427;
   wire n21428;
   wire n21429;
   wire n21430;
   wire n21431;
   wire n21432;
   wire n21433;
   wire n21434;
   wire n21435;
   wire n21436;
   wire n21437;
   wire n21438;
   wire n21439;
   wire n21440;
   wire n21441;
   wire n21442;
   wire n21443;
   wire n21444;
   wire n21445;
   wire n21446;
   wire n21447;
   wire n21448;
   wire n21449;
   wire n21450;
   wire n21451;
   wire n21452;
   wire n21453;
   wire n21454;
   wire n21455;
   wire n21457;
   wire n21458;
   wire n21459;
   wire n21460;
   wire n21461;
   wire n21462;
   wire n21463;
   wire n21464;
   wire n21465;
   wire n21466;
   wire n21467;
   wire n21468;
   wire n21469;
   wire n21471;
   wire n21472;
   wire n21473;
   wire n21474;
   wire n21475;
   wire n21476;
   wire n21477;
   wire n21478;
   wire n21479;
   wire n21480;
   wire n21482;
   wire n21483;
   wire n21484;
   wire n21485;
   wire n21486;
   wire n21487;
   wire n21488;
   wire n21489;
   wire n21490;
   wire n21491;
   wire n21492;
   wire n21493;
   wire n21494;
   wire n21495;
   wire n21496;
   wire n21497;
   wire n21498;
   wire n21499;
   wire n21500;
   wire n21501;
   wire n21502;
   wire n21503;
   wire n21504;
   wire n21505;
   wire n21506;
   wire n21507;
   wire n21508;
   wire n21509;
   wire n21510;
   wire n21511;
   wire n21513;
   wire n21514;
   wire n21516;
   wire n21517;
   wire n21518;
   wire n21519;
   wire n21520;
   wire n21521;
   wire n21522;
   wire n21523;
   wire n21524;
   wire n21525;
   wire n21526;
   wire n21527;
   wire n21528;
   wire n21529;
   wire n21530;
   wire n21531;
   wire n21532;
   wire n21533;
   wire n21534;
   wire n21535;
   wire n21536;
   wire n21537;
   wire n21538;
   wire n21539;
   wire n21540;
   wire n21541;
   wire n21542;
   wire n21543;
   wire n21544;
   wire n21545;
   wire n21546;
   wire n21547;
   wire n21548;
   wire n21549;
   wire n21550;
   wire n21551;
   wire n21552;
   wire n21553;
   wire n21554;
   wire n21556;
   wire n21557;
   wire n21558;
   wire n21559;
   wire n21560;
   wire n21561;
   wire n21562;
   wire n21563;
   wire n21564;
   wire n21565;
   wire n21566;
   wire n21567;
   wire n21568;
   wire n21569;
   wire n21570;
   wire n21571;
   wire n21572;
   wire n21573;
   wire n21574;
   wire n21575;
   wire n21576;
   wire n21577;
   wire n21578;
   wire n21579;
   wire n21580;
   wire n21581;
   wire n21582;
   wire n21583;
   wire n21584;
   wire n21585;
   wire n21586;
   wire n21587;
   wire n21588;
   wire n21589;
   wire n21590;
   wire n21591;
   wire n21592;
   wire n21593;
   wire n21594;
   wire n21595;
   wire n21596;
   wire n21597;
   wire n21598;
   wire n21599;
   wire n21600;
   wire n21601;
   wire n21602;
   wire n21603;
   wire n21604;
   wire n21605;
   wire n21606;
   wire n21607;
   wire n21608;
   wire n21609;
   wire n21611;
   wire n21613;
   wire n21615;
   wire n21616;
   wire n21617;
   wire n21618;
   wire n21619;
   wire n21620;
   wire n21621;
   wire n21622;
   wire n21623;
   wire n21624;
   wire n21625;
   wire n21626;
   wire n21627;
   wire n21628;
   wire n21629;
   wire n21630;
   wire n21631;
   wire n21632;
   wire n21633;
   wire n21634;
   wire n21635;
   wire n21636;
   wire n21637;
   wire n21638;
   wire n21639;
   wire n21640;
   wire n21641;
   wire n21642;
   wire n21643;
   wire n21644;
   wire n21645;
   wire n21646;
   wire n21647;
   wire n21648;
   wire n21649;
   wire n21650;
   wire n21651;
   wire n21652;
   wire n21653;
   wire n21654;
   wire n21655;
   wire n21656;
   wire n21657;
   wire n21658;
   wire n21659;
   wire n21660;
   wire n21661;
   wire n21662;
   wire n21663;
   wire n21664;
   wire n21665;
   wire n21666;
   wire n21667;
   wire n21668;
   wire n21669;
   wire n21670;
   wire n21671;
   wire n21672;
   wire n21673;
   wire n21674;
   wire n21675;
   wire n21676;
   wire n21677;
   wire n21678;
   wire n21679;
   wire n21680;
   wire n21681;
   wire n21682;
   wire n21683;
   wire n21684;
   wire n21685;
   wire n21686;
   wire n21687;
   wire n21688;
   wire n21689;
   wire n21690;
   wire n21691;
   wire n21692;
   wire n21693;
   wire n21694;
   wire n21695;
   wire n21696;
   wire n21697;
   wire n21698;
   wire n21699;
   wire n21700;
   wire n21701;
   wire n21703;
   wire n21704;
   wire n21705;
   wire n21706;
   wire n21707;
   wire n21708;
   wire n21709;
   wire n21710;
   wire n21711;
   wire n21712;
   wire n21713;
   wire n21714;
   wire n21715;
   wire n21716;
   wire n21717;
   wire n21718;
   wire n21719;
   wire n21720;
   wire n21721;
   wire n21722;
   wire n21724;
   wire n21725;
   wire n21726;
   wire n21727;
   wire n21728;
   wire n21729;
   wire n21730;
   wire n21731;
   wire n21732;
   wire n21733;
   wire n21734;
   wire n21735;
   wire n21736;
   wire n21737;
   wire n21738;
   wire n21739;
   wire n21740;
   wire n21742;
   wire n21743;
   wire n21744;
   wire n21745;
   wire n21746;
   wire n21747;
   wire n21748;
   wire n21749;
   wire n21750;
   wire n21751;
   wire n21752;
   wire n21753;
   wire n21754;
   wire n21755;
   wire n21756;
   wire n21757;
   wire n21758;
   wire n21759;
   wire n21760;
   wire n21761;
   wire n21762;
   wire n21763;
   wire n21764;
   wire n21765;
   wire n21766;
   wire n21767;
   wire n21768;
   wire n21769;
   wire n21770;
   wire n21771;
   wire n21772;
   wire n21773;
   wire n21774;
   wire n21775;
   wire n21776;
   wire n21777;
   wire n21778;
   wire n21779;
   wire n21780;
   wire n21781;
   wire n21782;
   wire n21783;
   wire n21784;
   wire n21785;
   wire n21786;
   wire n21787;
   wire n21788;
   wire n21789;
   wire n21790;
   wire n21791;
   wire n21792;
   wire n21793;
   wire n21794;
   wire n21795;
   wire n21796;
   wire n21797;
   wire n21798;
   wire n21799;
   wire n21800;
   wire n21801;
   wire n21802;
   wire n21803;
   wire n21804;
   wire n21805;
   wire n21806;
   wire n21807;
   wire n21808;
   wire n21809;
   wire n21810;
   wire n21811;
   wire n21812;
   wire n21813;
   wire n21814;
   wire n21815;
   wire n21816;
   wire n21817;
   wire n21818;
   wire n21819;
   wire n21820;
   wire n21821;
   wire n21822;
   wire n21823;
   wire n21824;
   wire n21825;
   wire n21826;
   wire n21827;
   wire n21828;
   wire n21829;
   wire n21830;
   wire n21831;
   wire n21832;
   wire n21833;
   wire n21834;
   wire n21835;
   wire n21836;
   wire n21837;
   wire n21838;
   wire n21839;
   wire n21840;
   wire n21841;
   wire n21842;
   wire n21843;
   wire n21844;
   wire n21845;
   wire n21846;
   wire n21847;
   wire n21848;
   wire n21849;
   wire n21850;
   wire n21851;
   wire n21852;
   wire n21853;
   wire n21854;
   wire n21855;
   wire n21856;
   wire n21857;
   wire n21858;
   wire n21859;
   wire n21860;
   wire n21861;
   wire n21862;
   wire n21863;
   wire n21864;
   wire n21865;
   wire n21866;
   wire n21867;
   wire n21868;
   wire n21869;
   wire n21870;
   wire n21872;
   wire n21873;
   wire n21874;
   wire n21875;
   wire n21876;
   wire n21877;
   wire n21878;
   wire n21879;
   wire n21880;
   wire n21881;
   wire n21882;
   wire n21883;
   wire n21884;
   wire n21885;
   wire n21886;
   wire n21887;
   wire n21888;
   wire n21889;
   wire n21890;
   wire n21891;
   wire n21892;
   wire n21893;
   wire n21894;
   wire n21895;
   wire n21896;
   wire n21897;
   wire n21898;
   wire n21899;
   wire n21900;
   wire n21901;
   wire n21902;
   wire n21903;
   wire n21904;
   wire n21905;
   wire n21906;
   wire n21907;
   wire n21908;
   wire n21909;
   wire n21910;
   wire n21911;
   wire n21912;
   wire n21913;
   wire n21914;
   wire n21915;
   wire n21916;
   wire n21917;
   wire n21918;
   wire n21919;
   wire n21920;
   wire n21921;
   wire n21922;
   wire n21923;
   wire n21924;
   wire n21925;
   wire n21926;
   wire n21927;
   wire n21928;
   wire n21929;
   wire n21930;
   wire n21931;
   wire n21932;
   wire n21933;
   wire n21934;
   wire n21935;
   wire n21936;
   wire n21937;
   wire n21938;
   wire n21939;
   wire n21940;
   wire n21941;
   wire n21942;
   wire n21943;
   wire n21944;
   wire n21945;
   wire n21946;
   wire n21947;
   wire n21948;
   wire n21949;
   wire n21950;
   wire n21951;
   wire n21952;
   wire n21953;
   wire n21954;
   wire n21955;
   wire n21956;
   wire n21957;
   wire n21958;
   wire n21959;
   wire n21960;
   wire n21961;
   wire n21962;
   wire n21963;
   wire n21964;
   wire n21965;
   wire n21966;
   wire n21967;
   wire n21968;
   wire n21969;
   wire n21970;
   wire n21971;
   wire n21972;
   wire n21974;
   wire n21975;
   wire n21977;
   wire n21978;
   wire n21979;
   wire n21980;
   wire n21981;
   wire n21982;
   wire n21983;
   wire n21984;
   wire n21985;
   wire n21986;
   wire n21987;
   wire n21988;
   wire n21989;
   wire n21990;
   wire n21991;
   wire n21992;
   wire n21993;
   wire n21994;
   wire n21995;
   wire n21996;
   wire n21997;
   wire n21998;
   wire n21999;
   wire n22000;
   wire n22001;
   wire n22002;
   wire n22003;
   wire n22004;
   wire n22005;
   wire n22006;
   wire n22007;
   wire n22008;
   wire n22009;
   wire n22010;
   wire n22011;
   wire n22012;
   wire n22013;
   wire n22014;
   wire n22015;
   wire n22016;
   wire n22018;
   wire n22019;
   wire n22020;
   wire n22021;
   wire n22022;
   wire n22024;
   wire n22025;
   wire n22026;
   wire n22027;
   wire n22028;
   wire n22029;
   wire n22030;
   wire n22031;
   wire n22032;
   wire n22033;
   wire n22034;
   wire n22035;
   wire n22036;
   wire n22038;
   wire n22039;
   wire n22040;
   wire n22041;
   wire n22042;
   wire n22043;
   wire n22044;
   wire n22045;
   wire n22046;
   wire n22047;
   wire n22048;
   wire n22049;
   wire n22050;
   wire n22051;
   wire n22052;
   wire n22053;
   wire n22054;
   wire n22055;
   wire n22056;
   wire n22057;
   wire n22058;
   wire n22059;
   wire n22060;
   wire n22061;
   wire n22062;
   wire n22063;
   wire n22064;
   wire n22065;
   wire n22066;
   wire n22067;
   wire n22068;
   wire n22069;
   wire n22070;
   wire n22071;
   wire n22072;
   wire n22073;
   wire n22074;
   wire n22075;
   wire n22076;
   wire n22077;
   wire n22078;
   wire n22079;
   wire n22081;
   wire n22082;
   wire n22083;
   wire n22084;
   wire n22085;
   wire n22086;
   wire n22087;
   wire n22088;
   wire n22089;
   wire n22090;
   wire n22091;
   wire n22092;
   wire n22093;
   wire n22094;
   wire n22095;
   wire n22096;
   wire n22098;
   wire n22099;
   wire n22100;
   wire n22101;
   wire n22102;
   wire n22103;
   wire n22104;
   wire n22105;
   wire n22106;
   wire n22107;
   wire n22108;
   wire n22109;
   wire n22110;
   wire n22111;
   wire n22112;
   wire n22113;
   wire n22114;
   wire n22115;
   wire n22116;
   wire n22117;
   wire n22118;
   wire n22119;
   wire n22120;
   wire n22121;
   wire n22122;
   wire n22123;
   wire n22124;
   wire n22125;
   wire n22126;
   wire n22127;
   wire n22128;
   wire n22129;
   wire n22130;
   wire n22131;
   wire n22132;
   wire n22133;
   wire n22134;
   wire n22135;
   wire n22136;
   wire n22137;
   wire n22138;
   wire n22139;
   wire n22140;
   wire n22141;
   wire n22142;
   wire n22143;
   wire n22144;
   wire n22145;
   wire n22146;
   wire n22147;
   wire n22148;
   wire n22149;
   wire n22150;
   wire n22151;
   wire n22152;
   wire n22153;
   wire n22154;
   wire n22155;
   wire n22156;
   wire n22157;
   wire n22158;
   wire n22159;
   wire n22160;
   wire n22161;
   wire n22162;
   wire n22163;
   wire n22164;
   wire n22165;
   wire n22166;
   wire n22167;
   wire n22168;
   wire n22169;
   wire n22170;
   wire n22171;
   wire n22172;
   wire n22173;
   wire n22174;
   wire n22175;
   wire n22176;
   wire n22177;
   wire n22178;
   wire n22179;
   wire n22180;
   wire n22181;
   wire n22182;
   wire n22183;
   wire n22184;
   wire n22185;
   wire n22186;
   wire n22187;
   wire n22188;
   wire n22189;
   wire n22190;
   wire n22191;
   wire n22192;
   wire n22193;
   wire n22194;
   wire n22195;
   wire n22196;
   wire n22197;
   wire n22198;
   wire n22199;
   wire n22200;
   wire n22201;
   wire n22202;
   wire n22203;
   wire n22204;
   wire n22205;
   wire n22206;
   wire n22207;
   wire n22208;
   wire n22209;
   wire n22210;
   wire n22211;
   wire n22212;
   wire n22214;
   wire n22215;
   wire n22216;
   wire n22217;
   wire n22218;
   wire n22219;
   wire n22220;
   wire n22221;
   wire n22222;
   wire n22223;
   wire n22224;
   wire n22225;
   wire n22226;
   wire n22227;
   wire n22228;
   wire n22229;
   wire n22230;
   wire n22231;
   wire n22232;
   wire n22233;
   wire n22234;
   wire n22235;
   wire n22236;
   wire n22237;
   wire n22238;
   wire n22239;
   wire n22240;
   wire n22241;
   wire n22242;
   wire n22243;
   wire n22244;
   wire n22245;
   wire n22246;
   wire n22247;
   wire n22248;
   wire n22249;
   wire n22250;
   wire n22251;
   wire n22252;
   wire n22253;
   wire n22254;
   wire n22255;
   wire n22256;
   wire n22257;
   wire n22258;
   wire n22259;
   wire n22260;
   wire n22261;
   wire n22262;
   wire n22263;
   wire n22264;
   wire n22265;
   wire n22266;
   wire n22267;
   wire n22268;
   wire n22269;
   wire n22270;
   wire n22271;
   wire n22272;
   wire n22273;
   wire n22274;
   wire n22275;
   wire n22276;
   wire n22277;
   wire n22278;
   wire n22279;
   wire n22280;
   wire n22281;
   wire n22282;
   wire n22283;
   wire n22284;
   wire n22285;
   wire n22286;
   wire n22287;
   wire n22288;
   wire n22289;
   wire n22290;
   wire n22291;
   wire n22292;
   wire n22293;
   wire n22294;
   wire n22295;
   wire n22296;
   wire n22297;
   wire n22298;
   wire n22299;
   wire n22300;
   wire n22301;
   wire n22302;
   wire n22303;
   wire n22304;
   wire n22305;
   wire n22306;
   wire n22307;
   wire n22308;
   wire n22309;
   wire n22310;
   wire n22311;
   wire n22312;
   wire n22313;
   wire n22314;
   wire n22315;
   wire n22316;
   wire n22317;
   wire n22318;
   wire n22319;
   wire n22320;
   wire n22321;
   wire n22322;
   wire n22323;
   wire n22324;
   wire n22325;
   wire n22326;
   wire n22327;
   wire n22328;
   wire n22329;
   wire n22330;
   wire n22331;
   wire n22332;
   wire n22333;
   wire n22334;
   wire n22335;
   wire n22336;
   wire n22337;
   wire n22338;
   wire n22339;
   wire n22340;
   wire n22341;
   wire n22342;
   wire n22343;
   wire n22344;
   wire n22345;
   wire n22346;
   wire n22347;
   wire n22348;
   wire n22349;
   wire n22350;
   wire n22351;
   wire n22352;
   wire n22353;
   wire n22354;
   wire n22355;
   wire n22356;
   wire n22357;
   wire n22358;
   wire n22359;
   wire n22360;
   wire n22361;
   wire n22362;
   wire n22363;
   wire n22364;
   wire n22365;
   wire n22366;
   wire n22367;
   wire n22368;
   wire n22369;
   wire n22370;
   wire n22371;
   wire n22372;
   wire n22373;
   wire n22374;
   wire n22375;
   wire n22376;
   wire n22377;
   wire n22378;
   wire n22379;
   wire n22380;
   wire n22381;
   wire n22382;
   wire n22383;
   wire n22384;
   wire n22385;
   wire n22386;
   wire n22387;
   wire n22388;
   wire n22389;
   wire n22390;
   wire n22391;
   wire n22392;
   wire n22393;
   wire n22394;
   wire n22395;
   wire n22396;
   wire n22397;
   wire n22398;
   wire n22399;
   wire n22400;
   wire n22401;
   wire n22402;
   wire n22403;
   wire n22405;
   wire n22406;
   wire n22407;
   wire n22409;
   wire n22410;
   wire n22411;
   wire n22412;
   wire n22414;
   wire n22415;
   wire n22416;
   wire n22417;
   wire n22418;
   wire n22419;
   wire n22420;
   wire n22421;
   wire n22422;
   wire n22423;
   wire n22424;
   wire n22425;
   wire n22426;
   wire n22427;
   wire n22428;
   wire n22429;
   wire n22430;
   wire n22431;
   wire n22432;
   wire n22433;
   wire n22434;
   wire n22435;
   wire n22436;
   wire n22437;
   wire n22438;
   wire n22439;
   wire n22442;
   wire n22443;
   wire n22444;
   wire n22445;
   wire n22446;
   wire n22447;
   wire n22448;
   wire n22449;
   wire n22450;
   wire n22451;
   wire n22452;
   wire n22453;
   wire n22455;
   wire n22456;
   wire n22457;
   wire n22458;
   wire n22459;
   wire n22460;
   wire n22461;
   wire n22462;
   wire n22463;
   wire n22464;
   wire n22467;
   wire n22468;
   wire n22469;
   wire n22470;
   wire n22471;
   wire n22472;
   wire n22473;
   wire n22474;
   wire n22475;
   wire n22476;
   wire n22477;
   wire n22478;
   wire n22479;
   wire n22480;
   wire n22481;
   wire n22482;
   wire n22483;
   wire n22484;
   wire n22485;
   wire n22486;
   wire n22487;
   wire n22488;
   wire n22489;
   wire n22490;
   wire n22491;
   wire n22492;
   wire n22493;
   wire n22494;
   wire n22495;
   wire n22496;
   wire n22497;
   wire n22498;
   wire n22499;
   wire n22500;
   wire n22501;
   wire n22502;
   wire n22503;
   wire n22504;
   wire n22505;
   wire n22506;
   wire n22507;
   wire n22508;
   wire n22509;
   wire n22510;
   wire n22511;
   wire n22512;
   wire n22513;
   wire n22514;
   wire n22515;
   wire n22516;
   wire n22517;
   wire n22518;
   wire n22519;
   wire n22520;
   wire n22521;
   wire n22522;
   wire n22523;
   wire n22524;
   wire n22526;
   wire n22527;
   wire n22528;
   wire n22529;
   wire n22530;
   wire n22531;
   wire n22532;
   wire n22533;
   wire n22534;
   wire n22535;
   wire n22536;
   wire n22537;
   wire n22538;
   wire n22539;
   wire n22540;
   wire n22541;
   wire n22542;
   wire n22543;
   wire n22544;
   wire n22545;
   wire n22546;
   wire n22547;
   wire n22548;
   wire n22549;
   wire n22550;
   wire n22551;
   wire n22552;
   wire n22553;
   wire n22554;
   wire n22555;
   wire n22556;
   wire n22557;
   wire n22558;
   wire n22559;
   wire n22560;
   wire n22561;
   wire n22562;
   wire n22563;
   wire n22564;
   wire n22565;
   wire n22566;
   wire n22567;
   wire n22568;
   wire n22569;
   wire n22570;
   wire n22571;
   wire n22572;
   wire n22573;
   wire n22574;
   wire n22575;
   wire n22576;
   wire n22577;
   wire n22578;
   wire n22579;
   wire n22580;
   wire n22581;
   wire n22582;
   wire n22583;
   wire n22584;
   wire n22585;
   wire n22586;
   wire n22587;
   wire n22588;
   wire n22589;
   wire n22590;
   wire n22591;
   wire n22592;
   wire n22593;
   wire n22594;
   wire n22595;
   wire n22596;
   wire n22597;
   wire n22598;
   wire n22599;
   wire n22600;
   wire n22601;
   wire n22602;
   wire n22603;
   wire n22604;
   wire n22605;
   wire n22606;
   wire n22607;
   wire n22608;
   wire n22609;
   wire n22610;
   wire n22611;
   wire n22612;
   wire n22613;
   wire n22614;
   wire n22615;
   wire n22616;
   wire n22617;
   wire n22618;
   wire n22619;
   wire n22620;
   wire n22621;
   wire n22622;
   wire n22623;
   wire n22624;
   wire n22625;
   wire n22626;
   wire n22627;
   wire n22628;
   wire n22629;
   wire n22630;
   wire n22631;
   wire n22632;
   wire n22633;
   wire n22634;
   wire n22635;
   wire n22636;
   wire n22637;
   wire n22638;
   wire n22639;
   wire n22640;
   wire n22641;
   wire n22642;
   wire n22643;
   wire n22644;
   wire n22645;
   wire n22646;
   wire n22647;
   wire n22648;
   wire n22649;
   wire n22650;
   wire n22651;
   wire n22652;
   wire n22653;
   wire n22654;
   wire n22655;
   wire n22656;
   wire n22657;
   wire n22658;
   wire n22659;
   wire n22660;
   wire n22661;
   wire n22662;
   wire n22663;
   wire n22664;
   wire n22665;
   wire n22666;
   wire n22667;
   wire n22668;
   wire n22669;
   wire n22670;
   wire n22671;
   wire n22672;
   wire n22673;
   wire n22674;
   wire n22675;
   wire n22676;
   wire n22677;
   wire n22678;
   wire n22679;
   wire n22681;
   wire n22682;
   wire n22683;
   wire n22684;
   wire n22685;
   wire n22686;
   wire n22687;
   wire n22688;
   wire n22689;
   wire n22690;
   wire n22692;
   wire n22693;
   wire n22694;
   wire n22695;
   wire n22696;
   wire n22697;
   wire n22698;
   wire n22699;
   wire n22700;
   wire n22701;
   wire n22702;
   wire n22703;
   wire n22704;
   wire n22705;
   wire n22706;
   wire n22707;
   wire n22708;
   wire n22709;
   wire n22710;
   wire n22711;
   wire n22712;
   wire n22713;
   wire n22714;
   wire n22715;
   wire n22716;
   wire n22717;
   wire n22718;
   wire n22719;
   wire n22720;
   wire n22721;
   wire n22722;
   wire n22723;
   wire n22724;
   wire n22725;
   wire n22726;
   wire n22727;
   wire n22728;
   wire n22730;
   wire n22731;
   wire n22732;
   wire n22733;
   wire n22734;
   wire n22735;
   wire n22736;
   wire n22737;
   wire n22738;
   wire n22739;
   wire n22740;
   wire n22741;
   wire n22742;
   wire n22743;
   wire n22744;
   wire n22745;
   wire n22746;
   wire n22747;
   wire n22748;
   wire n22749;
   wire n22750;
   wire n22751;
   wire n22752;
   wire n22753;
   wire n22754;
   wire n22755;
   wire n22756;
   wire n22757;
   wire n22758;
   wire n22759;
   wire n22760;
   wire n22761;
   wire n22762;
   wire n22763;
   wire n22764;
   wire n22765;
   wire n22766;
   wire n22767;
   wire n22768;
   wire n22769;
   wire n22770;
   wire n22771;
   wire n22772;
   wire n22773;
   wire n22774;
   wire n22775;
   wire n22776;
   wire n22777;
   wire n22778;
   wire n22779;
   wire n22780;
   wire n22781;
   wire n22782;
   wire n22783;
   wire n22784;
   wire n22785;
   wire n22786;
   wire n22787;
   wire n22788;
   wire n22789;
   wire n22790;
   wire n22791;
   wire n22792;
   wire n22793;
   wire n22794;
   wire n22795;
   wire n22796;
   wire n22797;
   wire n22798;
   wire n22799;
   wire n22800;
   wire n22801;
   wire n22802;
   wire n22803;
   wire n22804;
   wire n22805;
   wire n22806;
   wire n22807;
   wire n22808;
   wire n22809;
   wire n22810;
   wire n22811;
   wire n22812;
   wire n22813;
   wire n22814;
   wire n22815;
   wire n22816;
   wire n22817;
   wire n22819;
   wire n22820;
   wire n22821;
   wire n22822;
   wire n22823;
   wire n22824;
   wire n22825;
   wire n22826;
   wire n22827;
   wire n22828;
   wire n22829;
   wire n22830;
   wire n22831;
   wire n22832;
   wire n22833;
   wire n22834;
   wire n22835;
   wire n22836;
   wire n22837;
   wire n22838;
   wire n22839;
   wire n22840;
   wire n22841;
   wire n22842;
   wire n22843;
   wire n22844;
   wire n22845;
   wire n22846;
   wire n22847;
   wire n22848;
   wire n22849;
   wire n22850;
   wire n22851;
   wire n22852;
   wire n22853;
   wire n22854;
   wire n22855;
   wire n22856;
   wire n22857;
   wire n22858;
   wire n22859;
   wire n22860;
   wire n22861;
   wire n22862;
   wire n22863;
   wire n22864;
   wire n22865;
   wire n22866;
   wire n22867;
   wire n22868;
   wire n22869;
   wire n22870;
   wire n22871;
   wire n22872;
   wire n22873;
   wire n22874;
   wire n22875;
   wire n22876;
   wire n22877;
   wire n22878;
   wire n22879;
   wire n22880;
   wire n22881;
   wire n22882;
   wire n22883;
   wire n22884;
   wire n22885;
   wire n22886;
   wire n22888;
   wire n22889;
   wire n22890;
   wire n22891;
   wire n22892;
   wire n22893;
   wire n22894;
   wire n22895;
   wire n22896;
   wire n22897;
   wire n22898;
   wire n22899;
   wire n22900;
   wire n22901;
   wire n22902;
   wire n22903;
   wire n22904;
   wire n22905;
   wire n22906;
   wire n22907;
   wire n22908;
   wire n22909;
   wire n22910;
   wire n22911;
   wire n22912;
   wire n22913;
   wire n22914;
   wire n22915;
   wire n22916;
   wire n22917;
   wire n22918;
   wire n22919;
   wire n22920;
   wire n22921;
   wire n22922;
   wire n22923;
   wire n22924;
   wire n22925;
   wire n22926;
   wire n22927;
   wire n22928;
   wire n22929;
   wire n22930;
   wire n22931;
   wire n22932;
   wire n22933;
   wire n22934;
   wire n22935;
   wire n22936;
   wire n22937;
   wire n22938;
   wire n22939;
   wire n22940;
   wire n22941;
   wire n22942;
   wire n22943;
   wire n22944;
   wire n22945;
   wire n22946;
   wire n22947;
   wire n22948;
   wire n22949;
   wire n22950;
   wire n22951;
   wire n22952;
   wire n22953;
   wire n22954;
   wire n22955;
   wire n22956;
   wire n22957;
   wire n22958;
   wire n22959;
   wire n22960;
   wire n22961;
   wire n22962;
   wire n22963;
   wire n22964;
   wire n22965;
   wire n22966;
   wire n22967;
   wire n22968;
   wire n22969;
   wire n22970;
   wire n22971;
   wire n22972;
   wire n22973;
   wire n22974;
   wire n22975;
   wire n22976;
   wire n22977;
   wire n22978;
   wire n22979;
   wire n22980;
   wire n22981;
   wire n22982;
   wire n22983;
   wire n22984;
   wire n22985;
   wire n22986;
   wire n22987;
   wire n22988;
   wire n22989;
   wire n22990;
   wire n22992;
   wire n22993;
   wire n22994;
   wire n22995;
   wire n22996;
   wire n22997;
   wire n22998;
   wire n22999;
   wire n23000;
   wire n23001;
   wire n23002;
   wire n23003;
   wire n23004;
   wire n23005;
   wire n23006;
   wire n23007;
   wire n23008;
   wire n23009;
   wire n23010;
   wire n23012;
   wire n23013;
   wire n23014;
   wire n23015;
   wire n23016;
   wire n23017;
   wire n23018;
   wire n23020;
   wire n23021;
   wire n23022;
   wire n23024;
   wire n23025;
   wire n23026;
   wire n23027;
   wire n23028;
   wire n23029;
   wire n23030;
   wire n23031;
   wire n23032;
   wire n23033;
   wire n23034;
   wire n23035;
   wire n23036;
   wire n23037;
   wire n23038;
   wire n23039;
   wire n23040;
   wire n23041;
   wire n23042;
   wire n23043;
   wire n23044;
   wire n23046;
   wire n23048;
   wire n23050;
   wire n23051;
   wire n23052;
   wire n23053;
   wire n23054;
   wire n23055;
   wire n23056;
   wire n23057;
   wire n23058;
   wire n23059;
   wire n23060;
   wire n23061;
   wire n23062;
   wire n23063;
   wire n23064;
   wire n23065;
   wire n23066;
   wire n23067;
   wire n23068;
   wire n23069;
   wire n23071;
   wire n23072;
   wire n23073;
   wire n23074;
   wire n23075;
   wire n23076;
   wire n23077;
   wire n23078;
   wire n23079;
   wire n23080;
   wire n23081;
   wire n23082;
   wire n23083;
   wire n23084;
   wire n23085;
   wire n23086;
   wire n23087;
   wire n23088;
   wire n23089;
   wire n23090;
   wire n23091;
   wire n23092;
   wire n23093;
   wire n23094;
   wire n23095;
   wire n23096;
   wire n23097;
   wire n23099;
   wire n23100;
   wire n23101;
   wire n23102;
   wire n23103;
   wire n23104;
   wire n23105;
   wire n23106;
   wire n23107;
   wire n23108;
   wire n23109;
   wire n23110;
   wire n23111;
   wire n23112;
   wire n23113;
   wire n23114;
   wire n23115;
   wire n23116;
   wire n23117;
   wire n23118;
   wire n23119;
   wire n23120;
   wire n23121;
   wire n23122;
   wire n23123;
   wire n23124;
   wire n23125;
   wire n23126;
   wire n23127;
   wire n23128;
   wire n23129;
   wire n23130;
   wire n23131;
   wire n23132;
   wire n23133;
   wire n23134;
   wire n23135;
   wire n23136;
   wire n23137;
   wire n23138;
   wire n23139;
   wire n23140;
   wire n23141;
   wire n23143;
   wire n23144;
   wire n23145;
   wire n23147;
   wire n23148;
   wire n23149;
   wire n23150;
   wire n23151;
   wire n23152;
   wire n23153;
   wire n23154;
   wire n23155;
   wire n23156;
   wire n23157;
   wire n23158;
   wire n23159;
   wire n23160;
   wire n23161;
   wire n23162;
   wire n23164;
   wire n23165;
   wire n23166;
   wire n23167;
   wire n23168;
   wire n23169;
   wire n23170;
   wire n23171;
   wire n23172;
   wire n23173;
   wire n23174;
   wire n23175;
   wire n23176;
   wire n23177;
   wire n23178;
   wire n23179;
   wire n23180;
   wire n23181;
   wire n23182;
   wire n23183;
   wire n23184;
   wire n23185;
   wire n23186;
   wire n23187;
   wire n23188;
   wire n23189;
   wire n23190;
   wire n23191;
   wire n23192;
   wire n23193;
   wire n23194;
   wire n23195;
   wire n23196;
   wire n23197;
   wire n23198;
   wire n23199;
   wire n23200;
   wire n23201;
   wire n23202;
   wire n23203;
   wire n23204;
   wire n23205;
   wire n23206;
   wire n23207;
   wire n23208;
   wire n23209;
   wire n23210;
   wire n23211;
   wire n23212;
   wire n23213;
   wire n23214;
   wire n23215;
   wire n23216;
   wire n23217;
   wire n23218;
   wire n23219;
   wire n23220;
   wire n23221;
   wire n23222;
   wire n23223;
   wire n23224;
   wire n23225;
   wire n23226;
   wire n23227;
   wire n23228;
   wire n23229;
   wire n23230;
   wire n23231;
   wire n23232;
   wire n23233;
   wire n23234;
   wire n23235;
   wire n23236;
   wire n23237;
   wire n23238;
   wire n23239;
   wire n23240;
   wire n23241;
   wire n23242;
   wire n23243;
   wire n23244;
   wire n23245;
   wire n23246;
   wire n23247;
   wire n23248;
   wire n23249;
   wire n23250;
   wire n23251;
   wire n23252;
   wire n23253;
   wire n23254;
   wire n23255;
   wire n23256;
   wire n23257;
   wire n23258;
   wire n23259;
   wire n23260;
   wire n23261;
   wire n23262;
   wire n23263;
   wire n23264;
   wire n23265;
   wire n23266;
   wire n23267;
   wire n23268;
   wire n23269;
   wire n23270;
   wire n23271;
   wire n23272;
   wire n23273;
   wire n23274;
   wire n23275;
   wire n23276;
   wire n23277;
   wire n23278;
   wire n23279;
   wire n23280;
   wire n23281;
   wire n23282;
   wire n23283;
   wire n23284;
   wire n23285;
   wire n23286;
   wire n23287;
   wire n23288;
   wire n23289;
   wire n23290;
   wire n23291;
   wire n23292;
   wire n23293;
   wire n23294;
   wire n23295;
   wire n23296;
   wire n23297;
   wire n23298;
   wire n23299;
   wire n23300;
   wire n23301;
   wire n23302;
   wire n23303;
   wire n23304;
   wire n23305;
   wire n23306;
   wire n23307;
   wire n23308;
   wire n23309;
   wire n23310;
   wire n23311;
   wire n23312;
   wire n23313;
   wire n23314;
   wire n23315;
   wire n23316;
   wire n23317;
   wire n23318;
   wire n23319;
   wire n23320;
   wire n23321;
   wire n23322;
   wire n23323;
   wire n23324;
   wire n23325;
   wire n23326;
   wire n23327;
   wire n23328;
   wire n23329;
   wire n23330;
   wire n23331;
   wire n23332;
   wire n23333;
   wire n23334;
   wire n23335;
   wire n23336;
   wire n23337;
   wire n23338;
   wire n23339;
   wire n23340;
   wire n23341;
   wire n23342;
   wire n23343;
   wire n23344;
   wire n23345;
   wire n23346;
   wire n23347;
   wire n23348;
   wire n23349;
   wire n23350;
   wire n23351;
   wire n23352;
   wire n23353;
   wire n23354;
   wire n23355;
   wire n23356;
   wire n23357;
   wire n23358;
   wire n23359;
   wire n23360;
   wire n23361;
   wire n23362;
   wire n23363;
   wire n23364;
   wire n23365;
   wire n23366;
   wire n23367;
   wire n23368;
   wire n23369;
   wire n23370;
   wire n23371;
   wire n23372;
   wire n23373;
   wire n23374;
   wire n23375;
   wire n23376;
   wire n23377;
   wire n23378;
   wire n23379;
   wire n23380;
   wire n23381;
   wire n23382;
   wire n23383;
   wire n23384;
   wire n23385;
   wire n23386;
   wire n23387;
   wire n23388;
   wire n23389;
   wire n23390;
   wire n23391;
   wire n23392;
   wire n23393;
   wire n23394;
   wire n23395;
   wire n23396;
   wire n23397;
   wire n23398;
   wire n23399;
   wire n23400;
   wire n23401;
   wire n23402;
   wire n23403;
   wire n23404;
   wire n23405;
   wire n23406;
   wire n23407;
   wire n23408;
   wire n23409;
   wire n23410;
   wire n23411;
   wire n23412;
   wire n23413;
   wire n23414;
   wire n23415;
   wire n23416;
   wire n23417;
   wire n23418;
   wire n23419;
   wire n23420;
   wire n23421;
   wire n23422;
   wire n23423;
   wire n23424;
   wire n23425;
   wire n23426;
   wire n23427;
   wire n23428;
   wire n23429;
   wire n23430;
   wire n23431;
   wire n23432;
   wire n23433;
   wire n23435;
   wire n23436;
   wire n23437;
   wire n23438;
   wire n23439;
   wire n23440;
   wire n23441;
   wire n23442;
   wire n23443;
   wire n23444;
   wire n23446;
   wire n23447;
   wire n23448;
   wire n23449;
   wire n23450;
   wire n23451;
   wire n23452;
   wire n23453;
   wire n23454;
   wire n23455;
   wire n23456;
   wire n23457;
   wire n23458;
   wire n23459;
   wire n23460;
   wire n23461;
   wire n23462;
   wire n23463;
   wire n23464;
   wire n23465;
   wire n23466;
   wire n23467;
   wire n23468;
   wire n23469;
   wire n23470;
   wire n23471;
   wire n23472;
   wire n23473;
   wire n23474;
   wire n23475;
   wire n23476;
   wire n23477;
   wire n23478;
   wire n23479;
   wire n23480;
   wire n23481;
   wire n23482;
   wire n23483;
   wire n23484;
   wire n23485;
   wire n23486;
   wire n23487;
   wire n23488;
   wire n23489;
   wire n23490;
   wire n23491;
   wire n23492;
   wire n23493;
   wire n23494;
   wire n23495;
   wire n23496;
   wire n23497;
   wire n23498;
   wire n23499;
   wire n23500;
   wire n23501;
   wire n23502;
   wire n23503;
   wire n23504;
   wire n23505;
   wire n23506;
   wire n23507;
   wire n23508;
   wire n23509;
   wire n23510;
   wire n23511;
   wire n23512;
   wire n23513;
   wire n23514;
   wire n23515;
   wire n23516;
   wire n23517;
   wire n23518;
   wire n23519;
   wire n23520;
   wire n23521;
   wire n23522;
   wire n23523;
   wire n23524;
   wire n23525;
   wire n23526;
   wire n23527;
   wire n23528;
   wire n23529;
   wire n23530;
   wire n23531;
   wire n23532;
   wire n23533;
   wire n23534;
   wire n23535;
   wire n23536;
   wire n23537;
   wire n23538;
   wire n23539;
   wire n23540;
   wire n23541;
   wire n23542;
   wire n23543;
   wire n23544;
   wire n23545;
   wire n23546;
   wire n23547;
   wire n23548;
   wire n23549;
   wire n23550;
   wire n23551;
   wire n23552;
   wire n23553;
   wire n23554;
   wire n23555;
   wire n23556;
   wire n23557;
   wire n23558;
   wire n23559;
   wire n23560;
   wire n23561;
   wire n23562;
   wire n23563;
   wire n23564;
   wire n23565;
   wire n23566;
   wire n23567;
   wire n23568;
   wire n23569;
   wire n23570;
   wire n23571;
   wire n23572;
   wire n23573;
   wire n23574;
   wire n23575;
   wire n23576;
   wire n23577;
   wire n23578;
   wire n23579;
   wire n23580;
   wire n23581;
   wire n23582;
   wire n23583;
   wire n23584;
   wire n23585;
   wire n23586;
   wire n23587;
   wire n23588;
   wire n23589;
   wire n23590;
   wire n23592;
   wire n23593;
   wire n23594;
   wire n23595;
   wire n23596;
   wire n23597;
   wire n23598;
   wire n23599;
   wire n23600;
   wire n23601;
   wire n23602;
   wire n23603;
   wire n23604;
   wire n23605;
   wire n23606;
   wire n23607;
   wire n23608;
   wire n23609;
   wire n23610;
   wire n23611;
   wire n23612;
   wire n23613;
   wire n23614;
   wire n23615;
   wire n23616;
   wire n23617;
   wire n23618;
   wire n23619;
   wire n23620;
   wire n23621;
   wire n23622;
   wire n23623;
   wire n23624;
   wire n23625;
   wire n23626;
   wire n23627;
   wire n23628;
   wire n23630;
   wire n23631;
   wire n23632;
   wire n23633;
   wire n23634;
   wire n23635;
   wire n23636;
   wire n23637;
   wire n23638;
   wire n23639;
   wire n23640;
   wire n23641;
   wire n23642;
   wire n23643;
   wire n23644;
   wire n23645;
   wire n23646;
   wire n23647;
   wire n23648;
   wire n23649;
   wire n23650;
   wire n23651;
   wire n23652;
   wire n23653;
   wire n23654;
   wire n23655;
   wire n23656;
   wire n23657;
   wire n23658;
   wire n23659;
   wire n23660;
   wire n23661;
   wire n23662;
   wire n23663;
   wire n23664;
   wire n23665;
   wire n23666;
   wire n23667;
   wire n23668;
   wire n23669;
   wire n23670;
   wire n23671;
   wire n23672;
   wire n23673;
   wire n23674;
   wire n23675;
   wire n23676;
   wire n23677;
   wire n23678;
   wire n23679;
   wire n23680;
   wire n23681;
   wire n23682;
   wire n23683;
   wire n23684;
   wire n23685;
   wire n23686;
   wire n23687;
   wire n23688;
   wire n23689;
   wire n23690;
   wire n23691;
   wire n23692;
   wire n23693;
   wire n23694;
   wire n23695;
   wire n23696;
   wire n23697;
   wire n23698;
   wire n23699;
   wire n23700;
   wire n23701;
   wire n23702;
   wire n23703;
   wire n23704;
   wire n23705;
   wire n23706;
   wire n23707;
   wire n23708;
   wire n23709;
   wire n23710;
   wire n23711;
   wire n23712;
   wire n23713;
   wire n23714;
   wire n23715;
   wire n23716;
   wire n23717;
   wire n23718;
   wire n23719;
   wire n23720;
   wire n23721;
   wire n23722;
   wire n23723;
   wire n23724;
   wire n23725;
   wire n23726;
   wire n23727;
   wire n23728;
   wire n23729;
   wire n23730;
   wire n23731;
   wire n23732;
   wire n23733;
   wire n23734;
   wire n23735;
   wire n23736;
   wire n23737;
   wire n23738;
   wire n23739;
   wire n23740;
   wire n23741;
   wire n23743;
   wire n23744;
   wire n23745;
   wire n23746;
   wire n23747;
   wire n23748;
   wire n23749;
   wire n23750;
   wire n23751;
   wire n23752;
   wire n23753;
   wire n23754;
   wire n23755;
   wire n23757;
   wire n23758;
   wire n23759;
   wire n23760;
   wire n23761;
   wire n23762;
   wire n23763;
   wire n23764;
   wire n23765;
   wire n23766;
   wire n23767;
   wire n23768;
   wire n23769;
   wire n23770;
   wire n23771;
   wire n23773;
   wire n23774;
   wire n23775;
   wire n23776;
   wire n23777;
   wire n23778;
   wire n23779;
   wire n23780;
   wire n23781;
   wire n23782;
   wire n23783;
   wire n23784;
   wire n23785;
   wire n23786;
   wire n23787;
   wire n23788;
   wire n23789;
   wire n23790;
   wire n23791;
   wire n23792;
   wire n23793;
   wire n23794;
   wire n23795;
   wire n23796;
   wire n23797;
   wire n23798;
   wire n23799;
   wire n23800;
   wire n23801;
   wire n23802;
   wire n23803;
   wire n23804;
   wire n23805;
   wire n23806;
   wire n23807;
   wire n23808;
   wire n23809;
   wire n23810;
   wire n23811;
   wire n23812;
   wire n23813;
   wire n23814;
   wire n23815;
   wire n23816;
   wire n23817;
   wire n23818;
   wire n23819;
   wire n23821;
   wire n23822;
   wire n23823;
   wire n23824;
   wire n23825;
   wire n23826;
   wire n23827;
   wire n23828;
   wire n23829;
   wire n23830;
   wire n23831;
   wire n23832;
   wire n23833;
   wire n23834;
   wire n23835;
   wire n23836;
   wire n23837;
   wire n23838;
   wire n23839;
   wire n23840;
   wire n23841;
   wire n23842;
   wire n23843;
   wire n23844;
   wire n23845;
   wire n23846;
   wire n23847;
   wire n23848;
   wire n23849;
   wire n23850;
   wire n23851;
   wire n23852;
   wire n23853;
   wire n23854;
   wire n23855;
   wire n23856;
   wire n23857;
   wire n23858;
   wire n23859;
   wire n23860;
   wire n23861;
   wire n23862;
   wire n23863;
   wire n23864;
   wire n23865;
   wire n23866;
   wire n23867;
   wire n23868;
   wire n23869;
   wire n23870;
   wire n23871;
   wire n23872;
   wire n23873;
   wire n23874;
   wire n23875;
   wire n23876;
   wire n23877;
   wire n23878;
   wire n23879;
   wire n23880;
   wire n23882;
   wire n23883;
   wire n23884;
   wire n23885;
   wire n23886;
   wire n23887;
   wire n23888;
   wire n23889;
   wire n23890;
   wire n23891;
   wire n23892;
   wire n23893;
   wire n23894;
   wire n23895;
   wire n23896;
   wire n23897;
   wire n23898;
   wire n23899;
   wire n23900;
   wire n23901;
   wire n23902;
   wire n23903;
   wire n23904;
   wire n23905;
   wire n23906;
   wire n23907;
   wire n23908;
   wire n23909;
   wire n23910;
   wire n23911;
   wire n23913;
   wire n23914;
   wire n23915;
   wire n23916;
   wire n23917;
   wire n23918;
   wire n23919;
   wire n23920;
   wire n23921;
   wire n23922;
   wire n23923;
   wire n23924;
   wire n23925;
   wire n23926;
   wire n23927;
   wire n23928;
   wire n23929;
   wire n23930;
   wire n23931;
   wire n23932;
   wire n23933;
   wire n23934;
   wire n23935;
   wire n23936;
   wire n23937;
   wire n23938;
   wire n23939;
   wire n23940;
   wire n23941;
   wire n23942;
   wire n23943;
   wire n23944;
   wire n23945;
   wire n23946;
   wire n23948;
   wire n23949;
   wire n23950;
   wire n23951;
   wire n23952;
   wire n23953;
   wire n23954;
   wire n23955;
   wire n23956;
   wire n23957;
   wire n23958;
   wire n23959;
   wire n23960;
   wire n23961;
   wire n23962;
   wire n23963;
   wire n23964;
   wire n23965;
   wire n23966;
   wire n23967;
   wire n23968;
   wire n23969;
   wire n23970;
   wire n23971;
   wire n23972;
   wire n23973;
   wire n23974;
   wire n23975;
   wire n23976;
   wire n23977;
   wire n23978;
   wire n23979;
   wire n23980;
   wire n23981;
   wire n23982;
   wire n23983;
   wire n23984;
   wire n23985;
   wire n23986;
   wire n23987;
   wire n23988;
   wire n23989;
   wire n23990;
   wire n23991;
   wire n23992;
   wire n23993;
   wire n23994;
   wire n23995;
   wire n23996;
   wire n23997;
   wire n23998;
   wire n23999;
   wire n24000;
   wire n24001;
   wire n24002;
   wire n24003;
   wire n24004;
   wire n24005;
   wire n24006;
   wire n24007;
   wire n24008;
   wire n24009;
   wire n24010;
   wire n24011;
   wire n24012;
   wire n24013;
   wire n24014;
   wire n24015;
   wire n24016;
   wire n24017;
   wire n24018;
   wire n24019;
   wire n24020;
   wire n24021;
   wire n24022;
   wire n24023;
   wire n24024;
   wire n24025;
   wire n24027;
   wire n24028;
   wire n24029;
   wire n24030;
   wire n24031;
   wire n24032;
   wire n24033;
   wire n24034;
   wire n24035;
   wire n24037;
   wire n24038;
   wire n24040;
   wire n24041;
   wire n24042;
   wire n24043;
   wire n24044;
   wire n24045;
   wire n24046;
   wire n24047;
   wire n24048;
   wire n24049;
   wire n24050;
   wire n24051;
   wire n24052;
   wire n24053;
   wire n24054;
   wire n24055;
   wire n24056;
   wire n24057;
   wire n24058;
   wire n24059;
   wire n24060;
   wire n24061;
   wire n24062;
   wire n24063;
   wire n24064;
   wire n24065;
   wire n24066;
   wire n24067;
   wire n24068;
   wire n24069;
   wire n24070;
   wire n24071;
   wire n24072;
   wire n24073;
   wire n24074;
   wire n24075;
   wire n24076;
   wire n24077;
   wire n24078;
   wire n24079;
   wire n24080;
   wire n24081;
   wire n24082;
   wire n24083;
   wire n24084;
   wire n24085;
   wire n24086;
   wire n24087;
   wire n24088;
   wire n24089;
   wire n24090;
   wire n24091;
   wire n24092;
   wire n24093;
   wire n24094;
   wire n24095;
   wire n24096;
   wire n24097;
   wire n24098;
   wire n24099;
   wire n24100;
   wire n24101;
   wire n24102;
   wire n24103;
   wire n24104;
   wire n24105;
   wire n24106;
   wire n24107;
   wire n24108;
   wire n24109;
   wire n24110;
   wire n24111;
   wire n24112;
   wire n24113;
   wire n24114;
   wire n24115;
   wire n24116;
   wire n24117;
   wire n24118;
   wire n24119;
   wire n24120;
   wire n24121;
   wire n24122;
   wire n24123;
   wire n24124;
   wire n24125;
   wire n24126;
   wire n24127;
   wire n24128;
   wire n24129;
   wire n24130;
   wire n24131;
   wire n24132;
   wire n24133;
   wire n24134;
   wire n24135;
   wire n24136;
   wire n24137;
   wire n24138;
   wire n24139;
   wire n24140;
   wire n24141;
   wire n24142;
   wire n24143;
   wire n24144;
   wire n24145;
   wire n24146;
   wire n24147;
   wire n24148;
   wire n24149;
   wire n24150;
   wire n24151;
   wire n24152;
   wire n24153;
   wire n24154;
   wire n24155;
   wire n24156;
   wire n24157;
   wire n24158;
   wire n24159;
   wire n24160;
   wire n24161;
   wire n24162;
   wire n24163;
   wire n24164;
   wire n24165;
   wire n24166;
   wire n24167;
   wire n24168;
   wire n24169;
   wire n24170;
   wire n24171;
   wire n24172;
   wire n24173;
   wire n24174;
   wire n24175;
   wire n24176;
   wire n24177;
   wire n24178;
   wire n24179;
   wire n24180;
   wire n24181;
   wire n24182;
   wire n24183;
   wire n24184;
   wire n24185;
   wire n24186;
   wire n24187;
   wire n24188;
   wire n24189;
   wire n24190;
   wire n24191;
   wire n24192;
   wire n24193;
   wire n24194;
   wire n24195;
   wire n24196;
   wire n24197;
   wire n24198;
   wire n24199;
   wire n24200;
   wire n24201;
   wire n24202;
   wire n24203;
   wire n24204;
   wire n24205;
   wire n24206;
   wire n24207;
   wire n24208;
   wire n24209;
   wire n24210;
   wire n24211;
   wire n24212;
   wire n24213;
   wire n24214;
   wire n24216;
   wire n24217;
   wire n24218;
   wire n24219;
   wire n24220;
   wire n24221;
   wire n24222;
   wire n24223;
   wire n24224;
   wire n24225;
   wire n24226;
   wire n24227;
   wire n24228;
   wire n24229;
   wire n24230;
   wire n24231;
   wire n24232;
   wire n24233;
   wire n24235;
   wire n24236;
   wire n24237;
   wire n24238;
   wire n24239;
   wire n24240;
   wire n24241;
   wire n24243;
   wire n24244;
   wire n24245;
   wire n24246;
   wire n24247;
   wire n24248;
   wire n24249;
   wire n24250;
   wire n24251;
   wire n24252;
   wire n24253;
   wire n24254;
   wire n24255;
   wire n24256;
   wire n24257;
   wire n24258;
   wire n24259;
   wire n24260;
   wire n24261;
   wire n24262;
   wire n24263;
   wire n24264;
   wire n24265;
   wire n24266;
   wire n24267;
   wire n24268;
   wire n24269;
   wire n24270;
   wire n24271;
   wire n24272;
   wire n24273;
   wire n24274;
   wire n24275;
   wire n24276;
   wire n24277;
   wire n24278;
   wire n24279;
   wire n24280;
   wire n24281;
   wire n24282;
   wire n24283;
   wire n24284;
   wire n24285;
   wire n24286;
   wire n24287;
   wire n24288;
   wire n24289;
   wire n24290;
   wire n24291;
   wire n24293;
   wire n24294;
   wire n24295;
   wire n24296;
   wire n24297;
   wire n24298;
   wire n24299;
   wire n24300;
   wire n24301;
   wire n24302;
   wire n24303;
   wire n24304;
   wire n24305;
   wire n24306;
   wire n24307;
   wire n24308;
   wire n24309;
   wire n24310;
   wire n24311;
   wire n24312;
   wire n24313;
   wire n24314;
   wire n24315;
   wire n24318;
   wire n24319;
   wire n24320;
   wire n24321;
   wire n24322;
   wire n24323;
   wire n24324;
   wire n24325;
   wire n24326;
   wire n24327;
   wire n24328;
   wire n24329;
   wire n24330;
   wire n24331;
   wire n24333;
   wire n24334;
   wire n24335;
   wire n24336;
   wire n24337;
   wire n24338;
   wire n24339;
   wire n24340;
   wire n24341;
   wire n24342;
   wire n24343;
   wire n24344;
   wire n24345;
   wire n24346;
   wire n24347;
   wire n24348;
   wire n24349;
   wire n24350;
   wire n24351;
   wire n24352;
   wire n24353;
   wire n24354;
   wire n24355;
   wire n24356;
   wire n24357;
   wire n24358;
   wire n24359;
   wire n24360;
   wire n24361;
   wire n24362;
   wire n24363;
   wire n24364;
   wire n24365;
   wire n24366;
   wire n24367;
   wire n24368;
   wire n24369;
   wire n24370;
   wire n24371;
   wire n24372;
   wire n24373;
   wire n24374;
   wire n24375;
   wire n24376;
   wire n24377;
   wire n24378;
   wire n24379;
   wire n24380;
   wire n24381;
   wire n24382;
   wire n24383;
   wire n24384;
   wire n24385;
   wire n24386;
   wire n24387;
   wire n24388;
   wire n24389;
   wire n24390;
   wire n24391;
   wire n24392;
   wire n24393;
   wire n24394;
   wire n24395;
   wire n24396;
   wire n24397;
   wire n24398;
   wire n24399;
   wire n24400;
   wire n24401;
   wire n24402;
   wire n24403;
   wire n24404;
   wire n24405;
   wire n24406;
   wire n24407;
   wire n24408;
   wire n24409;
   wire n24410;
   wire n24411;
   wire n24412;
   wire n24413;
   wire n24414;
   wire n24415;
   wire n24416;
   wire n24417;
   wire n24418;
   wire n24419;
   wire n24420;
   wire n24421;
   wire n24422;
   wire n24423;
   wire n24424;
   wire n24426;
   wire n24427;
   wire n24428;
   wire n24429;
   wire n24430;
   wire n24431;
   wire n24432;
   wire n24433;
   wire n24434;
   wire n24435;
   wire n24436;
   wire n24437;
   wire n24438;
   wire n24439;
   wire n24440;
   wire n24441;
   wire n24442;
   wire n24444;
   wire n24445;
   wire n24446;
   wire n24447;
   wire n24448;
   wire n24449;
   wire n24450;
   wire n24451;
   wire n24452;
   wire n24453;
   wire n24454;
   wire n24455;
   wire n24456;
   wire n24457;
   wire n24458;
   wire n24459;
   wire n24460;
   wire n24461;
   wire n24462;
   wire n24463;
   wire n24464;
   wire n24465;
   wire n24466;
   wire n24467;
   wire n24468;
   wire n24469;
   wire n24470;
   wire n24471;
   wire n24472;
   wire n24473;
   wire n24474;
   wire n24475;
   wire n24476;
   wire n24477;
   wire n24478;
   wire n24479;
   wire n24480;
   wire n24481;
   wire n24482;
   wire n24483;
   wire n24484;
   wire n24485;
   wire n24486;
   wire n24487;
   wire n24488;
   wire n24489;
   wire n24490;
   wire n24491;
   wire n24492;
   wire n24493;
   wire n24494;
   wire n24495;
   wire n24496;
   wire n24497;
   wire n24498;
   wire n24499;
   wire n24500;
   wire n24501;
   wire n24502;
   wire n24503;
   wire n24504;
   wire n24505;
   wire n24506;
   wire n24507;
   wire n24508;
   wire n24509;
   wire n24510;
   wire n24511;
   wire n24512;
   wire n24513;
   wire n24514;
   wire n24515;
   wire n24516;
   wire n24517;
   wire n24518;
   wire n24519;
   wire n24520;
   wire n24521;
   wire n24522;
   wire n24523;
   wire n24524;
   wire n24525;
   wire n24526;
   wire n24527;
   wire n24528;
   wire n24529;
   wire n24530;
   wire n24531;
   wire n24532;
   wire n24533;
   wire n24534;
   wire n24535;
   wire n24537;
   wire n24538;
   wire n24539;
   wire n24540;
   wire n24541;
   wire n24542;
   wire n24543;
   wire n24544;
   wire n24545;
   wire n24546;
   wire n24547;
   wire n24548;
   wire n24549;
   wire n24550;
   wire n24551;
   wire n24552;
   wire n24553;
   wire n24554;
   wire n24555;
   wire n24556;
   wire n24557;
   wire n24558;
   wire n24559;
   wire n24560;
   wire n24561;
   wire n24562;
   wire n24563;
   wire n24564;
   wire n24565;
   wire n24566;
   wire n24567;
   wire n24568;
   wire n24569;
   wire n24570;
   wire n24571;
   wire n24572;
   wire n24573;
   wire n24574;
   wire n24575;
   wire n24576;
   wire n24577;
   wire n24578;
   wire n24579;
   wire n24580;
   wire n24581;
   wire n24582;
   wire n24583;
   wire n24584;
   wire n24585;
   wire n24586;
   wire n24587;
   wire n24588;
   wire n24589;
   wire n24590;
   wire n24591;
   wire n24592;
   wire n24593;
   wire n24594;
   wire n24595;
   wire n24596;
   wire n24597;
   wire n24598;
   wire n24599;
   wire n24600;
   wire n24601;
   wire n24602;
   wire n24603;
   wire n24604;
   wire n24605;
   wire n24606;
   wire n24607;
   wire n24608;
   wire n24609;
   wire n24610;
   wire n24611;
   wire n24612;
   wire n24613;
   wire n24614;
   wire n24615;
   wire n24616;
   wire n24617;
   wire n24618;
   wire n24619;
   wire n24620;
   wire n24622;
   wire n24623;
   wire n24624;
   wire n24625;
   wire n24626;
   wire n24627;
   wire n24628;
   wire n24629;
   wire n24630;
   wire n24631;
   wire n24632;
   wire n24633;
   wire n24634;
   wire n24635;
   wire n24636;
   wire n24637;
   wire n24638;
   wire n24639;
   wire n24640;
   wire n24641;
   wire n24642;
   wire n24643;
   wire n24644;
   wire n24645;
   wire n24646;
   wire n24647;
   wire n24648;
   wire n24649;
   wire n24650;
   wire n24651;
   wire n24652;
   wire n24653;
   wire n24654;
   wire n24655;
   wire n24656;
   wire n24657;
   wire n24658;
   wire n24659;
   wire n24660;
   wire n24661;
   wire n24662;
   wire n24663;
   wire n24664;
   wire n24665;
   wire n24666;
   wire n24667;
   wire n24668;
   wire n24669;
   wire n24670;
   wire n24671;
   wire n24673;
   wire n24674;
   wire n24675;
   wire n24676;
   wire n24677;
   wire n24678;
   wire n24679;
   wire n24680;
   wire n24681;
   wire n24682;
   wire n24683;
   wire n24684;
   wire n24685;
   wire n24686;
   wire n24687;
   wire n24688;
   wire n24689;
   wire n24690;
   wire n24691;
   wire n24692;
   wire n24693;
   wire n24694;
   wire n24695;
   wire n24696;
   wire n24697;
   wire n24698;
   wire n24699;
   wire n24700;
   wire n24701;
   wire n24702;
   wire n24703;
   wire n24704;
   wire n24705;
   wire n24706;
   wire n24707;
   wire n24708;
   wire n24709;
   wire n24710;
   wire n24711;
   wire n24712;
   wire n24713;
   wire n24714;
   wire n24715;
   wire n24716;
   wire n24717;
   wire n24718;
   wire n24719;
   wire n24720;
   wire n24721;
   wire n24722;
   wire n24723;
   wire n24724;
   wire n24725;
   wire n24726;
   wire n24727;
   wire n24728;
   wire n24729;
   wire n24730;
   wire n24731;
   wire n24732;
   wire n24733;
   wire n24734;
   wire n24735;
   wire n24736;
   wire n24737;
   wire n24738;
   wire n24739;
   wire n24740;
   wire n24741;
   wire n24742;
   wire n24743;
   wire n24744;
   wire n24745;
   wire n24746;
   wire n24747;
   wire n24748;
   wire n24749;
   wire n24750;
   wire n24751;
   wire n24752;
   wire n24753;
   wire n24754;
   wire n24755;
   wire n24756;
   wire n24757;
   wire n24758;
   wire n24759;
   wire n24760;
   wire n24761;
   wire n24762;
   wire n24763;
   wire n24765;
   wire n24766;
   wire n24767;
   wire n24768;
   wire n24769;
   wire n24770;
   wire n24771;
   wire n24772;
   wire n24773;
   wire n24774;
   wire n24775;
   wire n24776;
   wire n24777;
   wire n24778;
   wire n24779;
   wire n24780;
   wire n24781;
   wire n24782;
   wire n24783;
   wire n24784;
   wire n24785;
   wire n24786;
   wire n24787;
   wire n24788;
   wire n24789;
   wire n24790;
   wire n24791;
   wire n24792;
   wire n24793;
   wire n24794;
   wire n24795;
   wire n24796;
   wire n24797;
   wire n24798;
   wire n24799;
   wire n24800;
   wire n24801;
   wire n24802;
   wire n24803;
   wire n24805;
   wire n24806;
   wire n24807;
   wire n24809;
   wire n24810;
   wire n24811;
   wire n24812;
   wire n24813;
   wire n24814;
   wire n24815;
   wire n24816;
   wire n24817;
   wire n24818;
   wire n24819;
   wire n24820;
   wire n24821;
   wire n24822;
   wire n24823;
   wire n24824;
   wire n24825;
   wire n24826;
   wire n24827;
   wire n24828;
   wire n24829;
   wire n24830;
   wire n24831;
   wire n24832;
   wire n24833;
   wire n24834;
   wire n24835;
   wire n24837;
   wire n24838;
   wire n24839;
   wire n24841;
   wire n24842;
   wire n24843;
   wire n24844;
   wire n24845;
   wire n24846;
   wire n24847;
   wire n24848;
   wire n24849;
   wire n24850;
   wire n24851;
   wire n24852;
   wire n24853;
   wire n24854;
   wire n24855;
   wire n24856;
   wire n24858;
   wire n24859;
   wire n24860;
   wire n24861;
   wire n24862;
   wire n24863;
   wire n24864;
   wire n24865;
   wire n24866;
   wire n24867;
   wire n24868;
   wire n24869;
   wire n24870;
   wire n24871;
   wire n24872;
   wire n24873;
   wire n24874;
   wire n24875;
   wire n24876;
   wire n24877;
   wire n24878;
   wire n24879;
   wire n24880;
   wire n24881;
   wire n24883;
   wire n24884;
   wire n24885;
   wire n24886;
   wire n24887;
   wire n24888;
   wire n24889;
   wire n24890;
   wire n24891;
   wire n24892;
   wire n24893;
   wire n24894;
   wire n24895;
   wire n24896;
   wire n24897;
   wire n24898;
   wire n24899;
   wire n24900;
   wire n24901;
   wire n24902;
   wire n24903;
   wire n24904;
   wire n24905;
   wire n24906;
   wire n24907;
   wire n24909;
   wire n24910;
   wire n24911;
   wire n24912;
   wire n24913;
   wire n24914;
   wire n24915;
   wire n24916;
   wire n24917;
   wire n24918;
   wire n24919;
   wire n24920;
   wire n24921;
   wire n24922;
   wire n24923;
   wire n24924;
   wire n24925;
   wire n24926;
   wire n24927;
   wire n24928;
   wire n24929;
   wire n24930;
   wire n24931;
   wire n24932;
   wire n24933;
   wire n24934;
   wire n24935;
   wire n24936;
   wire n24937;
   wire n24938;
   wire n24939;
   wire n24941;
   wire n24942;
   wire n24943;
   wire n24944;
   wire n24945;
   wire n24946;
   wire n24947;
   wire n24948;
   wire n24949;
   wire n24950;
   wire n24951;
   wire n24952;
   wire n24953;
   wire n24954;
   wire n24955;
   wire n24956;
   wire n24957;
   wire n24958;
   wire n24959;
   wire n24960;
   wire n24961;
   wire n24962;
   wire n24963;
   wire n24964;
   wire n24965;
   wire n24966;
   wire n24967;
   wire n24968;
   wire n24969;
   wire n24970;
   wire n24971;
   wire n24972;
   wire n24973;
   wire n24974;
   wire n24975;
   wire n24976;
   wire n24977;
   wire n24978;
   wire n24979;
   wire n24980;
   wire n24981;
   wire n24982;
   wire n24983;
   wire n24985;
   wire n24986;
   wire n24987;
   wire n24988;
   wire n24989;
   wire n24991;
   wire n24992;
   wire n24993;
   wire n24994;
   wire n24995;
   wire n24996;
   wire n24997;
   wire n24998;
   wire n24999;
   wire n25000;
   wire n25001;
   wire n25002;
   wire n25003;
   wire n25004;
   wire n25005;
   wire n25006;
   wire n25007;
   wire n25008;
   wire n25009;
   wire n25010;
   wire n25011;
   wire n25012;
   wire n25013;
   wire n25014;
   wire n25015;
   wire n25017;
   wire n25018;
   wire n25019;
   wire n25020;
   wire n25021;
   wire n25022;
   wire n25023;
   wire n25024;
   wire n25025;
   wire n25026;
   wire n25027;
   wire n25028;
   wire n25029;
   wire n25030;
   wire n25031;
   wire n25032;
   wire n25033;
   wire n25034;
   wire n25035;
   wire n25036;
   wire n25037;
   wire n25038;
   wire n25039;
   wire n25040;
   wire n25041;
   wire n25042;
   wire n25043;
   wire n25044;
   wire n25045;
   wire n25046;
   wire n25047;
   wire n25048;
   wire n25049;
   wire n25050;
   wire n25051;
   wire n25052;
   wire n25053;
   wire n25054;
   wire n25055;
   wire n25056;
   wire n25057;
   wire n25058;
   wire n25059;
   wire n25060;
   wire n25061;
   wire n25062;
   wire n25063;
   wire n25064;
   wire n25065;
   wire n25066;
   wire n25067;
   wire n25068;
   wire n25069;
   wire n25070;
   wire n25071;
   wire n25072;
   wire n25073;
   wire n25074;
   wire n25075;
   wire n25076;
   wire n25077;
   wire n25078;
   wire n25079;
   wire n25080;
   wire n25081;
   wire n25082;
   wire n25083;
   wire n25084;
   wire n25085;
   wire n25086;
   wire n25087;
   wire n25088;
   wire n25089;
   wire n25090;
   wire n25091;
   wire n25092;
   wire n25093;
   wire n25094;
   wire n25095;
   wire n25096;
   wire n25097;
   wire n25098;
   wire n25099;
   wire n25100;
   wire n25101;
   wire n25102;
   wire n25103;
   wire n25104;
   wire n25105;
   wire n25106;
   wire n25107;
   wire n25108;
   wire n25109;
   wire n25110;
   wire n25111;
   wire n25112;
   wire n25113;
   wire n25114;
   wire n25115;
   wire n25116;
   wire n25117;
   wire n25118;
   wire n25119;
   wire n25120;
   wire n25121;
   wire n25122;
   wire n25123;
   wire n25124;
   wire n25125;
   wire n25126;
   wire n25127;
   wire n25128;
   wire n25129;
   wire n25130;
   wire n25131;
   wire n25132;
   wire n25133;
   wire n25134;
   wire n25136;
   wire n25137;
   wire n25138;
   wire n25139;
   wire n25140;
   wire n25141;
   wire n25142;
   wire n25143;
   wire n25144;
   wire n25145;
   wire n25146;
   wire n25147;
   wire n25148;
   wire n25149;
   wire n25150;
   wire n25151;
   wire n25152;
   wire n25153;
   wire n25154;
   wire n25155;
   wire n25156;
   wire n25158;
   wire n25159;
   wire n25160;
   wire n25161;
   wire n25162;
   wire n25163;
   wire n25164;
   wire n25165;
   wire n25166;
   wire n25167;
   wire n25168;
   wire n25169;
   wire n25170;
   wire n25171;
   wire n25172;
   wire n25173;
   wire n25174;
   wire n25176;
   wire n25177;
   wire n25178;
   wire n25179;
   wire n25180;
   wire n25181;
   wire n25182;
   wire n25183;
   wire n25184;
   wire n25185;
   wire n25186;
   wire n25187;
   wire n25188;
   wire n25189;
   wire n25190;
   wire n25191;
   wire n25192;
   wire n25193;
   wire n25194;
   wire n25195;
   wire n25196;
   wire n25197;
   wire n25198;
   wire n25199;
   wire n25200;
   wire n25201;
   wire n25202;
   wire n25203;
   wire n25204;
   wire n25205;
   wire n25206;
   wire n25207;
   wire n25208;
   wire n25210;
   wire n25211;
   wire n25212;
   wire n25213;
   wire n25214;
   wire n25215;
   wire n25216;
   wire n25217;
   wire n25218;
   wire n25219;
   wire n25220;
   wire n25221;
   wire n25222;
   wire n25223;
   wire n25224;
   wire n25225;
   wire n25226;
   wire n25227;
   wire n25228;
   wire n25229;
   wire n25230;
   wire n25231;
   wire n25232;
   wire n25233;
   wire n25234;
   wire n25235;
   wire n25236;
   wire n25237;
   wire n25238;
   wire n25239;
   wire n25240;
   wire n25241;
   wire n25242;
   wire n25243;
   wire n25244;
   wire n25245;
   wire n25246;
   wire n25247;
   wire n25248;
   wire n25249;
   wire n25250;
   wire n25251;
   wire n25252;
   wire n25253;
   wire n25254;
   wire n25255;
   wire n25256;
   wire n25257;
   wire n25258;
   wire n25259;
   wire n25260;
   wire n25261;
   wire n25262;
   wire n25263;
   wire n25264;
   wire n25265;
   wire n25266;
   wire n25267;
   wire n25268;
   wire n25269;
   wire n25270;
   wire n25271;
   wire n25272;
   wire n25273;
   wire n25274;
   wire n25275;
   wire n25276;
   wire n25277;
   wire n25278;
   wire n25279;
   wire n25280;
   wire n25281;
   wire n25282;
   wire n25283;
   wire n25284;
   wire n25285;
   wire n25286;
   wire n25287;
   wire n25288;
   wire n25289;
   wire n25290;
   wire n25291;
   wire n25292;
   wire n25293;
   wire n25294;
   wire n25295;
   wire n25296;
   wire n25297;
   wire n25298;
   wire n25299;
   wire n25300;
   wire n25301;
   wire n25302;
   wire n25303;
   wire n25304;
   wire n25305;
   wire n25306;
   wire n25307;
   wire n25308;
   wire n25309;
   wire n25310;
   wire n25311;
   wire n25312;
   wire n25313;
   wire n25314;
   wire n25315;
   wire n25316;
   wire n25317;
   wire n25318;
   wire n25319;
   wire n25320;
   wire n25321;
   wire n25322;
   wire n25323;
   wire n25324;
   wire n25325;
   wire n25326;
   wire n25327;
   wire n25328;
   wire n25329;
   wire n25330;
   wire n25331;
   wire n25332;
   wire n25333;
   wire n25334;
   wire n25335;
   wire n25336;
   wire n25337;
   wire n25338;
   wire n25339;
   wire n25340;
   wire n25341;
   wire n25342;
   wire n25343;
   wire n25344;
   wire n25345;
   wire n25346;
   wire n25347;
   wire n25348;
   wire n25349;
   wire n25350;
   wire n25351;
   wire n25352;
   wire n25353;
   wire n25354;
   wire n25355;
   wire n25356;
   wire n25357;
   wire n25358;
   wire n25359;
   wire n25360;
   wire n25361;
   wire n25362;
   wire n25363;
   wire n25364;
   wire n25365;
   wire n25366;
   wire n25367;
   wire n25368;
   wire n25369;
   wire n25370;
   wire n25371;
   wire n25372;
   wire n25373;
   wire n25375;
   wire n25376;
   wire n25377;
   wire n25378;
   wire n25379;
   wire n25380;
   wire n25381;
   wire n25382;
   wire n25383;
   wire n25384;
   wire n25385;
   wire n25386;
   wire n25387;
   wire n25388;
   wire n25389;
   wire n25390;
   wire n25391;
   wire n25392;
   wire n25393;
   wire n25394;
   wire n25395;
   wire n25396;
   wire n25397;
   wire n25398;
   wire n25399;
   wire n25400;
   wire n25401;
   wire n25402;
   wire n25403;
   wire n25404;
   wire n25405;
   wire n25406;
   wire n25407;
   wire n25408;
   wire n25409;
   wire n25410;
   wire n25411;
   wire n25412;
   wire n25413;
   wire n25414;
   wire n25417;
   wire n25418;
   wire n25419;
   wire n25420;
   wire n25421;
   wire n25422;
   wire n25423;
   wire n25424;
   wire n25425;
   wire n25426;
   wire n25427;
   wire n25428;
   wire n25429;
   wire n25430;
   wire n25431;
   wire n25432;
   wire n25434;
   wire n25435;
   wire n25436;
   wire n25437;
   wire n25438;
   wire n25439;
   wire n25440;
   wire n25441;
   wire n25442;
   wire n25443;
   wire n25444;
   wire n25445;
   wire n25446;
   wire n25447;
   wire n25449;
   wire n25450;
   wire n25451;
   wire n25452;
   wire n25453;
   wire n25454;
   wire n25455;
   wire n25456;
   wire n25457;
   wire n25459;
   wire n25460;
   wire n25461;
   wire n25462;
   wire n25463;
   wire n25464;
   wire n25465;
   wire n25466;
   wire n25467;
   wire n25468;
   wire n25469;
   wire n25470;
   wire n25471;
   wire n25472;
   wire n25473;
   wire n25474;
   wire n25475;
   wire n25476;
   wire n25478;
   wire n25479;
   wire n25480;
   wire n25481;
   wire n25482;
   wire n25483;
   wire n25484;
   wire n25485;
   wire n25486;
   wire n25487;
   wire n25488;
   wire n25489;
   wire n25490;
   wire n25491;
   wire n25492;
   wire n25493;
   wire n25494;
   wire n25495;
   wire n25496;
   wire n25497;
   wire n25498;
   wire n25499;
   wire n25500;
   wire n25501;
   wire n25502;
   wire n25503;
   wire n25504;
   wire n25505;
   wire n25506;
   wire n25507;
   wire n25508;
   wire n25509;
   wire n25510;
   wire n25511;
   wire n25512;
   wire n25513;
   wire n25514;
   wire n25515;
   wire n25516;
   wire n25517;
   wire n25518;
   wire n25519;
   wire n25520;
   wire n25521;
   wire n25522;
   wire n25523;
   wire n25524;
   wire n25525;
   wire n25526;
   wire n25527;
   wire n25528;
   wire n25529;
   wire n25530;
   wire n25531;
   wire n25532;
   wire n25533;
   wire n25534;
   wire n25535;
   wire n25536;
   wire n25537;
   wire n25538;
   wire n25539;
   wire n25540;
   wire n25541;
   wire n25542;
   wire n25543;
   wire n25544;
   wire n25545;
   wire n25546;
   wire n25547;
   wire n25548;
   wire n25549;
   wire n25550;
   wire n25551;
   wire n25552;
   wire n25553;
   wire n25554;
   wire n25555;
   wire n25556;
   wire n25557;
   wire n25558;
   wire n25559;
   wire n25560;
   wire n25561;
   wire n25562;
   wire n25563;
   wire n25564;
   wire n25565;
   wire n25566;
   wire n25567;
   wire n25568;
   wire n25569;
   wire n25570;
   wire n25571;
   wire n25572;
   wire n25573;
   wire n25574;
   wire n25575;
   wire n25576;
   wire n25577;
   wire n25578;
   wire n25579;
   wire n25580;
   wire n25581;
   wire n25582;
   wire n25583;
   wire n25584;
   wire n25585;
   wire n25586;
   wire n25587;
   wire n25588;
   wire n25589;
   wire n25590;
   wire n25591;
   wire n25592;
   wire n25593;
   wire n25594;
   wire n25595;
   wire n25596;
   wire n25597;
   wire n25598;
   wire n25599;
   wire n25600;
   wire n25601;
   wire n25602;
   wire n25603;
   wire n25604;
   wire n25605;
   wire n25606;
   wire n25607;
   wire n25608;
   wire n25609;
   wire n25610;
   wire n25611;
   wire n25612;
   wire n25613;
   wire n25614;
   wire n25615;
   wire n25616;
   wire n25617;
   wire n25618;
   wire n25619;
   wire n25620;
   wire n25621;
   wire n25622;
   wire n25623;
   wire n25624;
   wire n25625;
   wire n25626;
   wire n25627;
   wire n25628;
   wire n25629;
   wire n25630;
   wire n25631;
   wire n25632;
   wire n25633;
   wire n25634;
   wire n25635;
   wire n25636;
   wire n25637;
   wire n25638;
   wire n25639;
   wire n25640;
   wire n25641;
   wire n25642;
   wire n25643;
   wire n25644;
   wire n25645;
   wire n25646;
   wire n25647;
   wire n25648;
   wire n25649;
   wire n25650;
   wire n25651;
   wire n25652;
   wire n25654;
   wire n25655;
   wire n25657;
   wire n25658;
   wire n25659;
   wire n25660;
   wire n25661;
   wire n25662;
   wire n25663;
   wire n25664;
   wire n25665;
   wire n25666;
   wire n25667;
   wire n25669;
   wire n25670;
   wire n25671;
   wire n25672;
   wire n25673;
   wire n25674;
   wire n25675;
   wire n25676;
   wire n25677;
   wire n25678;
   wire n25679;
   wire n25680;
   wire n25681;
   wire n25682;
   wire n25683;
   wire n25684;
   wire n25685;
   wire n25686;
   wire n25687;
   wire n25688;
   wire n25689;
   wire n25690;
   wire n25691;
   wire n25692;
   wire n25693;
   wire n25694;
   wire n25695;
   wire n25696;
   wire n25697;
   wire n25698;
   wire n25699;
   wire n25700;
   wire n25701;
   wire n25702;
   wire n25703;
   wire n25704;
   wire n25705;
   wire n25706;
   wire n25707;
   wire n25708;
   wire n25709;
   wire n25710;
   wire n25711;
   wire n25712;
   wire n25713;
   wire n25714;
   wire n25715;
   wire n25716;
   wire n25717;
   wire n25718;
   wire n25719;
   wire n25721;
   wire n25722;
   wire n25723;
   wire n25724;
   wire n25725;
   wire n25726;
   wire n25727;
   wire n25728;
   wire n25729;
   wire n25730;
   wire n25731;
   wire n25732;
   wire n25733;
   wire n25734;
   wire n25735;
   wire n25736;
   wire n25737;
   wire n25738;
   wire n25739;
   wire n25740;
   wire n25741;
   wire n25742;
   wire n25743;
   wire n25744;
   wire n25745;
   wire n25746;
   wire n25747;
   wire n25748;
   wire n25749;
   wire n25750;
   wire n25751;
   wire n25752;
   wire n25753;
   wire n25754;
   wire n25755;
   wire n25756;
   wire n25757;
   wire n25758;
   wire n25759;
   wire n25760;
   wire n25761;
   wire n25762;
   wire n25763;
   wire n25764;
   wire n25765;
   wire n25766;
   wire n25767;
   wire n25768;
   wire n25769;
   wire n25770;
   wire n25771;
   wire n25772;
   wire n25773;
   wire n25774;
   wire n25775;
   wire n25776;
   wire n25777;
   wire n25778;
   wire n25779;
   wire n25780;
   wire n25781;
   wire n25782;
   wire n25783;
   wire n25784;
   wire n25785;
   wire n25786;
   wire n25787;
   wire n25788;
   wire n25789;
   wire n25790;
   wire n25791;
   wire n25792;
   wire n25793;
   wire n25794;
   wire n25795;
   wire n25796;
   wire n25797;
   wire n25798;
   wire n25799;
   wire n25800;
   wire n25801;
   wire n25802;
   wire n25803;
   wire n25804;
   wire n25805;
   wire n25806;
   wire n25807;
   wire n25808;
   wire n25809;
   wire n25810;
   wire n25811;
   wire n25812;
   wire n25813;
   wire n25814;
   wire n25815;
   wire n25816;
   wire n25817;
   wire n25818;
   wire n25819;
   wire n25820;
   wire n25821;
   wire n25822;
   wire n25823;
   wire n25824;
   wire n25825;
   wire n25826;
   wire n25827;
   wire n25828;
   wire n25829;
   wire n25830;
   wire n25831;
   wire n25832;
   wire n25833;
   wire n25834;
   wire n25835;
   wire n25836;
   wire n25837;
   wire n25838;
   wire n25839;
   wire n25840;
   wire n25841;
   wire n25842;
   wire n25843;
   wire n25844;
   wire n25845;
   wire n25846;
   wire n25847;
   wire n25848;
   wire n25849;
   wire n25850;
   wire n25851;
   wire n25852;
   wire n25853;
   wire n25854;
   wire n25855;
   wire n25856;
   wire n25857;
   wire n25858;
   wire n25859;
   wire n25860;
   wire n25861;
   wire n25862;
   wire n25863;
   wire n25864;
   wire n25866;
   wire n25867;
   wire n25868;
   wire n25869;
   wire n25870;
   wire n25872;
   wire n25873;
   wire n25874;
   wire n25875;
   wire n25876;
   wire n25877;
   wire n25878;
   wire n25879;
   wire n25880;
   wire n25881;
   wire n25882;
   wire n25883;
   wire n25884;
   wire n25885;
   wire n25886;
   wire n25887;
   wire n25888;
   wire n25889;
   wire n25890;
   wire n25891;
   wire n25892;
   wire n25893;
   wire n25894;
   wire n25895;
   wire n25896;
   wire n25897;
   wire n25898;
   wire n25899;
   wire n25900;
   wire n25901;
   wire n25902;
   wire n25903;
   wire n25904;
   wire n25905;
   wire n25906;
   wire n25907;
   wire n25908;
   wire n25909;
   wire n25910;
   wire n25911;
   wire n25912;
   wire n25913;
   wire n25914;
   wire n25915;
   wire n25916;
   wire n25917;
   wire n25918;
   wire n25919;
   wire n25920;
   wire n25921;
   wire n25922;
   wire n25923;
   wire n25924;
   wire n25925;
   wire n25926;
   wire n25927;
   wire n25928;
   wire n25929;
   wire n25930;
   wire n25931;
   wire n25932;
   wire n25933;
   wire n25934;
   wire n25935;
   wire n25936;
   wire n25937;
   wire n25938;
   wire n25939;
   wire n25940;
   wire n25941;
   wire n25942;
   wire n25943;
   wire n25944;
   wire n25946;
   wire n25947;
   wire n25948;
   wire n25949;
   wire n25950;
   wire n25951;
   wire n25952;
   wire n25953;
   wire n25954;
   wire n25956;
   wire n25957;
   wire n25958;
   wire n25959;
   wire n25960;
   wire n25961;
   wire n25962;
   wire n25963;
   wire n25964;
   wire n25965;
   wire n25966;
   wire n25967;
   wire n25968;
   wire n25969;
   wire n25970;
   wire n25971;
   wire n25972;
   wire n25973;
   wire n25974;
   wire n25975;
   wire n25976;
   wire n25977;
   wire n25978;
   wire n25979;
   wire n25980;
   wire n25981;
   wire n25982;
   wire n25983;
   wire n25984;
   wire n25985;
   wire n25986;
   wire n25987;
   wire n25988;
   wire n25989;
   wire n25990;
   wire n25991;
   wire n25992;
   wire n25993;
   wire n25994;
   wire n25995;
   wire n25996;
   wire n25997;
   wire n25998;
   wire n25999;
   wire n26000;
   wire n26001;
   wire n26002;
   wire n26003;
   wire n26004;
   wire n26005;
   wire n26006;
   wire n26007;
   wire n26008;
   wire n26009;
   wire n26010;
   wire n26011;
   wire n26012;
   wire n26013;
   wire n26014;
   wire n26015;
   wire n26016;
   wire n26017;
   wire n26018;
   wire n26019;
   wire n26020;
   wire n26021;
   wire n26022;
   wire n26023;
   wire n26024;
   wire n26025;
   wire n26026;
   wire n26027;
   wire n26028;
   wire n26029;
   wire n26030;
   wire n26031;
   wire n26032;
   wire n26033;
   wire n26034;
   wire n26035;
   wire n26036;
   wire n26037;
   wire n26038;
   wire n26039;
   wire n26040;
   wire n26041;
   wire n26042;
   wire n26043;
   wire n26044;
   wire n26045;
   wire n26046;
   wire n26047;
   wire n26048;
   wire n26049;
   wire n26050;
   wire n26051;
   wire n26052;
   wire n26053;
   wire n26054;
   wire n26055;
   wire n26056;
   wire n26057;
   wire n26058;
   wire n26059;
   wire n26060;
   wire n26061;
   wire n26062;
   wire n26063;
   wire n26064;
   wire n26065;
   wire n26066;
   wire n26067;
   wire n26068;
   wire n26069;
   wire n26070;
   wire n26071;
   wire n26072;
   wire n26073;
   wire n26074;
   wire n26075;
   wire n26076;
   wire n26077;
   wire n26078;
   wire n26079;
   wire n26080;
   wire n26081;
   wire n26082;
   wire n26083;
   wire n26084;
   wire n26085;
   wire n26086;
   wire n26087;
   wire n26088;
   wire n26089;
   wire n26090;
   wire n26091;
   wire n26092;
   wire n26093;
   wire n26094;
   wire n26095;
   wire n26096;
   wire n26097;
   wire n26098;
   wire n26099;
   wire n26100;
   wire n26101;
   wire n26102;
   wire n26103;
   wire n26104;
   wire n26105;
   wire n26106;
   wire n26107;
   wire n26108;
   wire n26109;
   wire n26110;
   wire n26111;
   wire n26112;
   wire n26113;
   wire n26114;
   wire n26115;
   wire n26116;
   wire n26117;
   wire n26118;
   wire n26119;
   wire n26120;
   wire n26121;
   wire n26122;
   wire n26123;
   wire n26124;
   wire n26125;
   wire n26126;
   wire n26127;
   wire n26128;
   wire n26129;
   wire n26130;
   wire n26131;
   wire n26132;
   wire n26133;
   wire n26134;
   wire n26135;
   wire n26136;
   wire n26137;
   wire n26138;
   wire n26139;
   wire n26140;
   wire n26141;
   wire n26142;
   wire n26143;
   wire n26144;
   wire n26145;
   wire n26146;
   wire n26147;
   wire n26148;
   wire n26149;
   wire n26150;
   wire n26151;
   wire n26152;
   wire n26153;
   wire n26154;
   wire n26155;
   wire n26156;
   wire n26157;
   wire n26158;
   wire n26159;
   wire n26160;
   wire n26161;
   wire n26162;
   wire n26163;
   wire n26164;
   wire n26165;
   wire n26166;
   wire n26167;
   wire n26168;
   wire n26169;
   wire n26170;
   wire n26171;
   wire n26172;
   wire n26173;
   wire n26174;
   wire n26175;
   wire n26176;
   wire n26177;
   wire n26178;
   wire n26179;
   wire n26180;
   wire n26181;
   wire n26182;
   wire n26183;
   wire n26184;
   wire n26185;
   wire n26186;
   wire n26187;
   wire n26188;
   wire n26189;
   wire n26190;
   wire n26192;
   wire n26193;
   wire n26194;
   wire n26195;
   wire n26196;
   wire n26197;
   wire n26198;
   wire n26199;
   wire n26200;
   wire n26201;
   wire n26202;
   wire n26203;
   wire n26204;
   wire n26205;
   wire n26206;
   wire n26207;
   wire n26208;
   wire n26209;
   wire n26210;
   wire n26211;
   wire n26212;
   wire n26213;
   wire n26214;
   wire n26215;
   wire n26216;
   wire n26217;
   wire n26218;
   wire n26219;
   wire n26220;
   wire n26221;
   wire n26222;
   wire n26223;
   wire n26224;
   wire n26225;
   wire n26226;
   wire n26227;
   wire n26228;
   wire n26229;
   wire n26230;
   wire n26231;
   wire n26232;
   wire n26233;
   wire n26234;
   wire n26235;
   wire n26236;
   wire n26237;
   wire n26238;
   wire n26239;
   wire n26240;
   wire n26241;
   wire n26242;
   wire n26243;
   wire n26245;
   wire n26246;
   wire n26247;
   wire n26248;
   wire n26249;
   wire n26250;
   wire n26251;
   wire n26252;
   wire n26253;
   wire n26254;
   wire n26255;
   wire n26256;
   wire n26257;
   wire n26258;
   wire n26259;
   wire n26260;
   wire n26261;
   wire n26262;
   wire n26263;
   wire n26264;
   wire n26265;
   wire n26266;
   wire n26267;
   wire n26268;
   wire n26269;
   wire n26270;
   wire n26271;
   wire n26272;
   wire n26273;
   wire n26274;
   wire n26276;
   wire n26277;
   wire n26279;
   wire n26280;
   wire n26281;
   wire n26282;
   wire n26283;
   wire n26284;
   wire n26285;
   wire n26286;
   wire n26287;
   wire n26288;
   wire n26289;
   wire n26290;
   wire n26291;
   wire n26292;
   wire n26293;
   wire n26294;
   wire n26295;
   wire n26296;
   wire n26297;
   wire n26298;
   wire n26299;
   wire n26300;
   wire n26301;
   wire n26302;
   wire n26303;
   wire n26304;
   wire n26305;
   wire n26306;
   wire n26307;
   wire n26308;
   wire n26309;
   wire n26310;
   wire n26311;
   wire n26312;
   wire n26313;
   wire n26314;
   wire n26315;
   wire n26317;
   wire n26318;
   wire n26319;
   wire n26320;
   wire n26321;
   wire n26322;
   wire n26323;
   wire n26324;
   wire n26325;
   wire n26326;
   wire n26327;
   wire n26328;
   wire n26329;
   wire n26330;
   wire n26331;
   wire n26332;
   wire n26333;
   wire n26334;
   wire n26335;
   wire n26336;
   wire n26337;
   wire n26338;
   wire n26339;
   wire n26340;
   wire n26342;
   wire n26343;
   wire n26344;
   wire n26345;
   wire n26346;
   wire n26347;
   wire n26348;
   wire n26349;
   wire n26350;
   wire n26351;
   wire n26352;
   wire n26353;
   wire n26354;
   wire n26355;
   wire n26356;
   wire n26357;
   wire n26358;
   wire n26359;
   wire n26360;
   wire n26361;
   wire n26362;
   wire n26363;
   wire n26364;
   wire n26365;
   wire n26366;
   wire n26367;
   wire n26368;
   wire n26369;
   wire n26370;
   wire n26371;
   wire n26372;
   wire n26373;
   wire n26374;
   wire n26375;
   wire n26376;
   wire n26377;
   wire n26378;
   wire n26379;
   wire n26380;
   wire n26381;
   wire n26382;
   wire n26383;
   wire n26384;
   wire n26385;
   wire n26386;
   wire n26387;
   wire n26388;
   wire n26389;
   wire n26390;
   wire n26391;
   wire n26392;
   wire n26393;
   wire n26394;
   wire n26395;
   wire n26396;
   wire n26397;
   wire n26398;
   wire n26399;
   wire n26400;
   wire n26401;
   wire n26402;
   wire n26403;
   wire n26404;
   wire n26405;
   wire n26406;
   wire n26407;
   wire n26408;
   wire n26409;
   wire n26410;
   wire n26412;
   wire n26413;
   wire n26414;
   wire n26415;
   wire n26416;
   wire n26417;
   wire n26418;
   wire n26419;
   wire n26420;
   wire n26421;
   wire n26422;
   wire n26423;
   wire n26424;
   wire n26425;
   wire n26426;
   wire n26427;
   wire n26428;
   wire n26429;
   wire n26430;
   wire n26431;
   wire n26432;
   wire n26433;
   wire n26434;
   wire n26435;
   wire n26436;
   wire n26437;
   wire n26438;
   wire n26439;
   wire n26440;
   wire n26441;
   wire n26442;
   wire n26443;
   wire n26444;
   wire n26445;
   wire n26446;
   wire n26447;
   wire n26448;
   wire n26449;
   wire n26450;
   wire n26451;
   wire n26452;
   wire n26453;
   wire n26454;
   wire n26455;
   wire n26456;
   wire n26457;
   wire n26458;
   wire n26459;
   wire n26460;
   wire n26461;
   wire n26462;
   wire n26463;
   wire n26464;
   wire n26465;
   wire n26466;
   wire n26467;
   wire n26468;
   wire n26469;
   wire n26470;
   wire n26471;
   wire n26472;
   wire n26473;
   wire n26474;
   wire n26475;
   wire n26476;
   wire n26477;
   wire n26478;
   wire n26479;
   wire n26480;
   wire n26481;
   wire n26482;
   wire n26483;
   wire n26484;
   wire n26485;
   wire n26486;
   wire n26487;
   wire n26488;
   wire n26491;
   wire n26492;
   wire n26493;
   wire n26494;
   wire n26495;
   wire n26496;
   wire n26497;
   wire n26498;
   wire n26499;
   wire n26500;
   wire n26501;
   wire n26502;
   wire n26503;
   wire n26504;
   wire n26505;
   wire n26506;
   wire n26507;
   wire n26508;
   wire n26509;
   wire n26510;
   wire n26511;
   wire n26512;
   wire n26513;
   wire n26514;
   wire n26515;
   wire n26516;
   wire n26517;
   wire n26518;
   wire n26519;
   wire n26520;
   wire n26521;
   wire n26522;
   wire n26523;
   wire n26524;
   wire n26527;
   wire n26528;
   wire n26529;
   wire n26530;
   wire n26531;
   wire n26532;
   wire n26533;
   wire n26534;
   wire n26535;
   wire n26536;
   wire n26537;
   wire n26538;
   wire n26539;
   wire n26540;
   wire n26541;
   wire n26542;
   wire n26543;
   wire n26544;
   wire n26545;
   wire n26546;
   wire n26547;
   wire n26548;
   wire n26549;
   wire n26550;
   wire n26551;
   wire n26552;
   wire n26553;
   wire n26554;
   wire n26555;
   wire n26556;
   wire n26557;
   wire n26558;
   wire n26559;
   wire n26560;
   wire n26561;
   wire n26562;
   wire n26563;
   wire n26564;
   wire n26565;
   wire n26566;
   wire n26567;
   wire n26568;
   wire n26569;
   wire n26570;
   wire n26571;
   wire n26572;
   wire n26573;
   wire n26574;
   wire n26575;
   wire n26576;
   wire n26577;
   wire n26578;
   wire n26579;
   wire n26580;
   wire n26581;
   wire n26582;
   wire n26583;
   wire n26584;
   wire n26585;
   wire n26586;
   wire n26587;
   wire n26588;
   wire n26589;
   wire n26590;
   wire n26591;
   wire n26592;
   wire n26593;
   wire n26594;
   wire n26595;
   wire n26596;
   wire n26597;
   wire n26598;
   wire n26599;
   wire n26600;
   wire n26601;
   wire n26603;
   wire n26604;
   wire n26605;
   wire n26606;
   wire n26607;
   wire n26608;
   wire n26609;
   wire n26610;
   wire n26611;
   wire n26612;
   wire n26613;
   wire n26615;
   wire n26616;
   wire n26617;
   wire n26618;
   wire n26619;
   wire n26620;
   wire n26621;
   wire n26622;
   wire n26623;
   wire n26624;
   wire n26625;
   wire n26626;
   wire n26627;
   wire n26628;
   wire n26629;
   wire n26630;
   wire n26631;
   wire n26632;
   wire n26633;
   wire n26634;
   wire n26635;
   wire n26636;
   wire n26637;
   wire n26638;
   wire n26639;
   wire n26640;
   wire n26641;
   wire n26642;
   wire n26643;
   wire n26644;
   wire n26645;
   wire n26646;
   wire n26647;
   wire n26648;
   wire n26649;
   wire n26651;
   wire n26652;
   wire n26653;
   wire n26654;
   wire n26655;
   wire n26656;
   wire n26657;
   wire n26658;
   wire n26659;
   wire n26660;
   wire n26661;
   wire n26662;
   wire n26663;
   wire n26664;
   wire n26665;
   wire n26666;
   wire n26667;
   wire n26668;
   wire n26669;
   wire n26670;
   wire n26671;
   wire n26672;
   wire n26673;
   wire n26674;
   wire n26675;
   wire n26676;
   wire n26677;
   wire n26678;
   wire n26679;
   wire n26680;
   wire n26681;
   wire n26682;
   wire n26683;
   wire n26684;
   wire n26685;
   wire n26686;
   wire n26687;
   wire n26688;
   wire n26689;
   wire n26690;
   wire n26691;
   wire n26692;
   wire n26693;
   wire n26694;
   wire n26695;
   wire n26696;
   wire n26697;
   wire n26698;
   wire n26699;
   wire n26700;
   wire n26701;
   wire n26702;
   wire n26703;
   wire n26704;
   wire n26705;
   wire n26706;
   wire n26707;
   wire n26708;
   wire n26709;
   wire n26710;
   wire n26711;
   wire n26712;
   wire n26713;
   wire n26714;
   wire n26715;
   wire n26716;
   wire n26717;
   wire n26718;
   wire n26719;
   wire n26721;
   wire n26722;
   wire n26723;
   wire n26724;
   wire n26725;
   wire n26726;
   wire n26727;
   wire n26728;
   wire n26729;
   wire n26730;
   wire n26731;
   wire n26732;
   wire n26734;
   wire n26735;
   wire n26736;
   wire n26737;
   wire n26738;
   wire n26739;
   wire n26740;
   wire n26741;
   wire n26742;
   wire n26743;
   wire n26744;
   wire n26745;
   wire n26746;
   wire n26747;
   wire n26748;
   wire n26749;
   wire n26750;
   wire n26751;
   wire n26752;
   wire n26753;
   wire n26754;
   wire n26755;
   wire n26756;
   wire n26757;
   wire n26758;
   wire n26759;
   wire n26760;
   wire n26761;
   wire n26762;
   wire n26764;
   wire n26765;
   wire n26766;
   wire n26767;
   wire n26768;
   wire n26769;
   wire n26770;
   wire n26771;
   wire n26772;
   wire n26773;
   wire n26774;
   wire n26775;
   wire n26776;
   wire n26777;
   wire n26778;
   wire n26779;
   wire n26780;
   wire n26781;
   wire n26782;
   wire n26783;
   wire n26784;
   wire n26785;
   wire n26786;
   wire n26787;
   wire n26788;
   wire n26789;
   wire n26790;
   wire n26791;
   wire n26792;
   wire n26793;
   wire n26794;
   wire n26795;
   wire n26796;
   wire n26797;
   wire n26798;
   wire n26799;
   wire n26800;
   wire n26801;
   wire n26802;
   wire n26803;
   wire n26804;
   wire n26805;
   wire n26806;
   wire n26807;
   wire n26808;
   wire n26809;
   wire n26810;
   wire n26811;
   wire n26812;
   wire n26813;
   wire n26814;
   wire n26815;
   wire n26816;
   wire n26817;
   wire n26818;
   wire n26819;
   wire n26820;
   wire n26821;
   wire n26822;
   wire n26823;
   wire n26824;
   wire n26825;
   wire n26826;
   wire n26827;
   wire n26828;
   wire n26829;
   wire n26830;
   wire n26831;
   wire n26832;
   wire n26833;
   wire n26834;
   wire n26835;
   wire n26836;
   wire n26837;
   wire n26838;
   wire n26839;
   wire n26840;
   wire n26841;
   wire n26842;
   wire n26843;
   wire n26844;
   wire n26845;
   wire n26846;
   wire n26848;
   wire n26849;
   wire n26850;
   wire n26851;
   wire n26852;
   wire n26853;
   wire n26854;
   wire n26855;
   wire n26856;
   wire n26857;
   wire n26858;
   wire n26859;
   wire n26860;
   wire n26861;
   wire n26863;
   wire n26864;
   wire n26866;
   wire n26867;
   wire n26868;
   wire n26869;
   wire n26870;
   wire n26871;
   wire n26872;
   wire n26873;
   wire n26874;
   wire n26875;
   wire n26876;
   wire n26877;
   wire n26878;
   wire n26879;
   wire n26880;
   wire n26881;
   wire n26882;
   wire n26883;
   wire n26884;
   wire n26885;
   wire n26886;
   wire n26887;
   wire n26888;
   wire n26889;
   wire n26890;
   wire n26891;
   wire n26892;
   wire n26893;
   wire n26894;
   wire n26895;
   wire n26896;
   wire n26897;
   wire n26898;
   wire n26899;
   wire n26900;
   wire n26901;
   wire n26902;
   wire n26903;
   wire n26904;
   wire n26905;
   wire n26906;
   wire n26907;
   wire n26910;
   wire n26911;
   wire n26912;
   wire n26913;
   wire n26914;
   wire n26915;
   wire n26916;
   wire n26917;
   wire n26918;
   wire n26919;
   wire n26920;
   wire n26921;
   wire n26922;
   wire n26923;
   wire n26924;
   wire n26925;
   wire n26926;
   wire n26927;
   wire n26928;
   wire n26929;
   wire n26930;
   wire n26931;
   wire n26932;
   wire n26933;
   wire n26934;
   wire n26935;
   wire n26936;
   wire n26937;
   wire n26938;
   wire n26939;
   wire n26940;
   wire n26941;
   wire n26942;
   wire n26943;
   wire n26944;
   wire n26945;
   wire n26946;
   wire n26947;
   wire n26948;
   wire n26950;
   wire n26951;
   wire n26952;
   wire n26953;
   wire n26954;
   wire n26955;
   wire n26956;
   wire n26957;
   wire n26958;
   wire n26959;
   wire n26960;
   wire n26961;
   wire n26962;
   wire n26963;
   wire n26964;
   wire n26965;
   wire n26966;
   wire n26967;
   wire n26968;
   wire n26969;
   wire n26970;
   wire n26971;
   wire n26972;
   wire n26973;
   wire n26974;
   wire n26975;
   wire n26976;
   wire n26978;
   wire n26979;
   wire n26980;
   wire n26981;
   wire n26982;
   wire n26983;
   wire n26984;
   wire n26985;
   wire n26986;
   wire n26987;
   wire n26988;
   wire n26989;
   wire n26990;
   wire n26991;
   wire n26992;
   wire n26993;
   wire n26994;
   wire n26995;
   wire n26996;
   wire n26997;
   wire n26998;
   wire n26999;
   wire n27000;
   wire n27001;
   wire n27002;
   wire n27003;
   wire n27004;
   wire n27005;
   wire n27006;
   wire n27007;
   wire n27008;
   wire n27009;
   wire n27010;
   wire n27011;
   wire n27012;
   wire n27013;
   wire n27014;
   wire n27015;
   wire n27016;
   wire n27017;
   wire n27018;
   wire n27019;
   wire n27020;
   wire n27022;
   wire n27023;
   wire n27024;
   wire n27025;
   wire n27027;
   wire n27028;
   wire n27029;
   wire n27030;
   wire n27031;
   wire n27033;
   wire n27034;
   wire n27036;
   wire n27037;
   wire n27038;
   wire n27039;
   wire n27040;
   wire n27041;
   wire n27042;
   wire n27044;
   wire n27045;
   wire n27046;
   wire n27049;
   wire n27050;
   wire n27051;
   wire n27052;
   wire n27053;
   wire n27054;
   wire n27055;
   wire n27056;
   wire n27057;
   wire n27058;
   wire n27059;
   wire n27060;
   wire n27061;
   wire n27062;
   wire n27063;
   wire n27064;
   wire n27065;
   wire n27066;
   wire n27067;
   wire n27068;
   wire n27069;
   wire n27070;
   wire n27071;
   wire n27072;
   wire n27073;
   wire n27074;
   wire n27075;
   wire n27076;
   wire n27077;
   wire n27078;
   wire n27079;
   wire n27080;
   wire n27081;
   wire n27082;
   wire n27083;
   wire n27084;
   wire n27085;
   wire n27086;
   wire n27087;
   wire n27088;
   wire n27089;
   wire n27090;
   wire n27091;
   wire n27093;
   wire n27094;
   wire n27095;
   wire n27096;
   wire n27097;
   wire n27098;
   wire n27099;
   wire n27100;
   wire n27101;
   wire n27102;
   wire n27103;
   wire n27105;
   wire n27106;
   wire n27107;
   wire n27108;
   wire n27109;
   wire n27110;
   wire n27113;
   wire n27114;
   wire n27115;
   wire n27116;
   wire n27117;
   wire n27118;
   wire n27119;
   wire n27120;
   wire n27121;
   wire n27122;
   wire n27123;
   wire n27124;
   wire n27125;
   wire n27126;
   wire n27127;
   wire n27128;
   wire n27129;
   wire n27130;
   wire n27131;
   wire n27132;
   wire n27133;
   wire n27135;
   wire n27136;
   wire n27137;
   wire n27138;
   wire n27139;
   wire n27140;
   wire n27141;
   wire n27142;
   wire n27143;
   wire n27144;
   wire n27145;
   wire n27146;
   wire n27147;
   wire n27148;
   wire n27149;
   wire n27150;
   wire n27151;
   wire n27152;
   wire n27153;
   wire n27155;
   wire n27156;
   wire n27157;
   wire n27158;
   wire n27159;
   wire n27160;
   wire n27161;
   wire n27162;
   wire n27163;
   wire n27164;
   wire n27165;
   wire n27166;
   wire n27167;
   wire n27168;
   wire n27169;
   wire n27170;
   wire n27171;
   wire n27172;
   wire n27173;
   wire n27174;
   wire n27175;
   wire n27176;
   wire n27177;
   wire n27178;
   wire n27179;
   wire n27180;
   wire n27181;
   wire n27182;
   wire n27183;
   wire n27184;
   wire n27185;
   wire n27186;
   wire n27187;
   wire n27188;
   wire n27189;
   wire n27190;
   wire n27191;
   wire n27192;
   wire n27194;
   wire n27195;
   wire n27196;
   wire n27197;
   wire n27198;
   wire n27199;
   wire n27200;
   wire n27201;
   wire n27202;
   wire n27203;
   wire n27204;
   wire n27205;
   wire n27206;
   wire n27207;
   wire n27208;
   wire n27209;
   wire n27210;
   wire n27211;
   wire n27212;
   wire n27213;
   wire n27214;
   wire n27215;
   wire n27216;
   wire n27218;
   wire n27219;
   wire n27220;
   wire n27221;
   wire n27222;
   wire n27223;

   HB1xp67_ASAP7_75t_L FE_PSC8338_n19791 (.Y(FE_PSN8338_n19791),
	.A(n19791));
   BUFx2_ASAP7_75t_SL FE_PSC8337_n16909 (.Y(FE_PSN8337_n16909),
	.A(n16909));
   HB1xp67_ASAP7_75t_L FE_PSC8336_n23340 (.Y(FE_PSN8336_n23340),
	.A(n23340));
   HB1xp67_ASAP7_75t_L FE_PSC8335_n17606 (.Y(FE_PSN8335_n17606),
	.A(n17606));
   BUFx3_ASAP7_75t_L FE_PSC8334_n15539 (.Y(FE_PSN8334_n15539),
	.A(n15539));
   HB1xp67_ASAP7_75t_SL FE_PSC8333_n18478 (.Y(FE_PSN8333_n18478),
	.A(n18478));
   HB1xp67_ASAP7_75t_L FE_PSC8332_n23879 (.Y(FE_PSN8332_n23879),
	.A(n23879));
   HB1xp67_ASAP7_75t_L FE_PSC8331_n24113 (.Y(FE_PSN8331_n24113),
	.A(n24113));
   HB1xp67_ASAP7_75t_L FE_PSC8330_n17761 (.Y(FE_PSN8330_n17761),
	.A(n17761));
   HB1xp67_ASAP7_75t_L FE_PSC8329_n21638 (.Y(FE_PSN8329_n21638),
	.A(n21638));
   HB1xp67_ASAP7_75t_SL FE_PSC8328_n20260 (.Y(FE_PSN8328_n20260),
	.A(n20260));
   HB1xp67_ASAP7_75t_L FE_PSC8327_n24562 (.Y(FE_PSN8327_n24562),
	.A(n24562));
   HB1xp67_ASAP7_75t_L FE_PSC8326_n21455 (.Y(FE_PSN8326_n21455),
	.A(n21455));
   HB1xp67_ASAP7_75t_SL FE_PSC8325_FE_OFN28811_n19170 (.Y(FE_PSN8325_FE_OFN28811_n19170),
	.A(FE_OFN28811_n19170));
   BUFx3_ASAP7_75t_SL FE_PSC8324_n15987 (.Y(FE_PSN8324_n15987),
	.A(n15987));
   HB1xp67_ASAP7_75t_SL FE_PSC8323_n22543 (.Y(FE_PSN8323_n22543),
	.A(n22543));
   HB1xp67_ASAP7_75t_L FE_PSC8322_n25105 (.Y(FE_PSN8322_n25105),
	.A(n25105));
   BUFx3_ASAP7_75t_SL FE_PSC8321_n26520 (.Y(FE_PSN8321_n26520),
	.A(n26520));
   BUFx2_ASAP7_75t_L FE_PSC8320_n18176 (.Y(FE_PSN8320_n18176),
	.A(n18176));
   HB1xp67_ASAP7_75t_L FE_PSC8319_n21725 (.Y(FE_PSN8319_n21725),
	.A(n21725));
   HB2xp67_ASAP7_75t_SL FE_PSC8318_n21455 (.Y(FE_PSN8318_n21455),
	.A(FE_PSN8326_n21455));
   HB1xp67_ASAP7_75t_L FE_PSC8317_n20850 (.Y(FE_PSN8317_n20850),
	.A(n20850));
   HB1xp67_ASAP7_75t_L FE_PSC8316_n23781 (.Y(FE_PSN8316_n23781),
	.A(n23781));
   BUFx3_ASAP7_75t_SL FE_PSC8315_FE_OFN16135_sa22_4 (.Y(FE_PSN8315_FE_OFN16135_sa22_4),
	.A(FE_OFN16135_sa22_4));
   HB1xp67_ASAP7_75t_L FE_PSC8314_n25722 (.Y(FE_PSN8314_n25722),
	.A(n25722));
   BUFx2_ASAP7_75t_SL FE_PSC8313_FE_OCPN29469_n17747 (.Y(FE_PSN8313_FE_OCPN29469_n17747),
	.A(FE_OCPN29469_n17747));
   HB1xp67_ASAP7_75t_L FE_PSC8312_n21442 (.Y(FE_PSN8312_n21442),
	.A(n21442));
   HB1xp67_ASAP7_75t_SL FE_PSC8311_n25105 (.Y(FE_PSN8311_n25105),
	.A(FE_PSN8322_n25105));
   HB1xp67_ASAP7_75t_SL FE_PSC8310_n17473 (.Y(FE_PSN8310_n17473),
	.A(n17473));
   HB1xp67_ASAP7_75t_L FE_PSC8309_n21372 (.Y(FE_PSN8309_n21372),
	.A(n21372));
   HB1xp67_ASAP7_75t_SL FE_PSC8308_n22624 (.Y(FE_PSN8308_n22624),
	.A(n22624));
   BUFx2_ASAP7_75t_SL FE_PSC8307_FE_OFN27207_w3_30 (.Y(FE_PSN8307_FE_OFN27207_w3_30),
	.A(FE_OFN27207_w3_30));
   HB1xp67_ASAP7_75t_L FE_PSC8306_FE_OFN28689_sa03_5 (.Y(FE_PSN8306_FE_OFN28689_sa03_5),
	.A(FE_OFN28689_sa03_5));
   HB1xp67_ASAP7_75t_L FE_PSC8305_n21217 (.Y(FE_PSN8305_n21217),
	.A(n21217));
   HB1xp67_ASAP7_75t_L FE_PSC8304_n24565 (.Y(FE_PSN8304_n24565),
	.A(n24565));
   HB1xp67_ASAP7_75t_SL FE_PSC8303_n19222 (.Y(FE_PSN8303_n19222),
	.A(n19222));
   HB1xp67_ASAP7_75t_L FE_PSC8302_n24562 (.Y(FE_PSN8302_n24562),
	.A(FE_PSN8327_n24562));
   HB1xp67_ASAP7_75t_SL FE_PSC8301_n23197 (.Y(FE_PSN8301_n23197),
	.A(n23197));
   BUFx2_ASAP7_75t_L FE_PSC8300_n26482 (.Y(FE_PSN8300_n26482),
	.A(n26482));
   HB1xp67_ASAP7_75t_L FE_PSC8299_FE_OFN4_w3_22 (.Y(FE_PSN8299_FE_OFN4_w3_22),
	.A(FE_OFN4_w3_22));
   HB1xp67_ASAP7_75t_L FE_PSC8298_FE_OFN27151_n (.Y(FE_PSN8298_FE_OFN27151_n),
	.A(FE_OFN27151_n));
   HB1xp67_ASAP7_75t_L FE_PSC8297_FE_OFN8_w3_14 (.Y(FE_PSN8297_FE_OFN8_w3_14),
	.A(FE_OFN8_w3_14));
   HB1xp67_ASAP7_75t_SL FE_PSC8296_FE_OFN26588_n24062 (.Y(FE_PSN8296_FE_OFN26588_n24062),
	.A(FE_OFN26588_n24062));
   HB1xp67_ASAP7_75t_L FE_PSC8295_FE_OFN28669_sa31_5 (.Y(FE_PSN8295_FE_OFN28669_sa31_5),
	.A(FE_OFN28669_sa31_5));
   HB1xp67_ASAP7_75t_SL FE_PSC8294_n22310 (.Y(FE_PSN8294_n22310),
	.A(n22310));
   BUFx3_ASAP7_75t_SL FE_PSC8293_n25317 (.Y(FE_PSN8293_n25317),
	.A(n25317));
   BUFx2_ASAP7_75t_L FE_PSC8292_FE_OFN26041_w3_17 (.Y(FE_PSN8292_FE_OFN26041_w3_17),
	.A(FE_OFN26041_w3_17));
   HB1xp67_ASAP7_75t_L FE_PSC8291_n26404 (.Y(FE_PSN8291_n26404),
	.A(n26404));
   HB1xp67_ASAP7_75t_SL FE_PSC8290_n21439 (.Y(FE_PSN8290_n21439),
	.A(n21439));
   HB1xp67_ASAP7_75t_L FE_PSC8289_FE_OFN28514_sa00_1 (.Y(FE_PSN8289_FE_OFN28514_sa00_1),
	.A(FE_OFN28514_sa00_1));
   HB1xp67_ASAP7_75t_L FE_PSC8288_n17275 (.Y(FE_PSN8288_n17275),
	.A(n17275));
   HB1xp67_ASAP7_75t_L FE_PSC8287_FE_OCPN27494_n26479 (.Y(FE_PSN8287_FE_OCPN27494_n26479),
	.A(FE_OCPN27494_n26479));
   HB1xp67_ASAP7_75t_L FE_PSC8286_FE_OCPN29260_sa00_5 (.Y(FE_PSN8286_FE_OCPN29260_sa00_5),
	.A(FE_OCPN29260_sa00_5));
   HB1xp67_ASAP7_75t_L FE_PSC8285_FE_OCPN29463_n (.Y(FE_PSN8285_FE_OCPN29463_n),
	.A(FE_OCPN29463_n));
   HB1xp67_ASAP7_75t_SL FE_PSC8284_n21438 (.Y(FE_PSN8284_n21438),
	.A(n21438));
   HB1xp67_ASAP7_75t_L FE_PSC8283_n22629 (.Y(FE_PSN8283_n22629),
	.A(n22629));
   BUFx2_ASAP7_75t_SL FE_PSC8282_n21154 (.Y(FE_PSN8282_n21154),
	.A(n21154));
   HB1xp67_ASAP7_75t_SL FE_PSC8281_n25118 (.Y(FE_PSN8281_n25118),
	.A(n25118));
   HB1xp67_ASAP7_75t_L FE_PSC8280_n15660 (.Y(FE_PSN8280_n15660),
	.A(n15660));
   HB1xp67_ASAP7_75t_L FE_PSC8279_FE_OCPN27292_n25389 (.Y(FE_PSN8279_FE_OCPN27292_n25389),
	.A(FE_OCPN27292_n25389));
   HB1xp67_ASAP7_75t_L FE_PSC8278_n25605 (.Y(FE_PSN8278_n25605),
	.A(n25605));
   HB1xp67_ASAP7_75t_L FE_PSC8277_n16099 (.Y(FE_PSN8277_n16099),
	.A(n16099));
   HB1xp67_ASAP7_75t_L FE_PSC8276_FE_OFN28712_n (.Y(FE_PSN8276_FE_OFN28712_n),
	.A(FE_OFN28712_n));
   BUFx6f_ASAP7_75t_SL FE_PSC8275_FE_OCPN27818_n17267 (.Y(FE_PSN8275_FE_OCPN27818_n17267),
	.A(FE_OCPN27818_n17267));
   HB1xp67_ASAP7_75t_L FE_PSC8274_n21164 (.Y(FE_PSN8274_n21164),
	.A(n21164));
   HB1xp67_ASAP7_75t_SL FE_PSC8273_n24087 (.Y(FE_PSN8273_n24087),
	.A(n24087));
   HB1xp67_ASAP7_75t_SL FE_PSC8272_n20428 (.Y(FE_PSN8272_n20428),
	.A(n20428));
   BUFx2_ASAP7_75t_L FE_PSC8271_n15924 (.Y(FE_PSN8271_n15924),
	.A(n15924));
   BUFx3_ASAP7_75t_SL FE_PSC8270_n26027 (.Y(FE_PSN8270_n26027),
	.A(n26027));
   BUFx2_ASAP7_75t_SL FE_OCPC8269_FE_OFN16136_sa02_5 (.Y(FE_OCPN8269_FE_OFN16136_sa02_5),
	.A(FE_OFN16136_sa02_5));
   HB1xp67_ASAP7_75t_L FE_OCPC8268_n26632 (.Y(FE_OCPN8268_n26632),
	.A(n26632));
   HB1xp67_ASAP7_75t_R FE_OCPC8267_n16069 (.Y(FE_OCPN8267_n16069),
	.A(n16069));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8266_sa21_2 (.Y(FE_OCPN8266_sa21_2),
	.A(sa21_2_));
   HB1xp67_ASAP7_75t_R FE_OCPC8265_n24362 (.Y(FE_OCPN8265_n24362),
	.A(n24362));
   BUFx3_ASAP7_75t_SL FE_OCPC8264_n13890 (.Y(FE_OCPN8264_n13890),
	.A(n13890));
   HB1xp67_ASAP7_75t_L FE_OCPC8263_n25039 (.Y(FE_OCPN8263_n25039),
	.A(n25039));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8262_n21726 (.Y(FE_OCPN8262_n21726),
	.A(n21726));
   HB1xp67_ASAP7_75t_R FE_OCPC8261_n26513 (.Y(FE_OCPN8261_n26513),
	.A(n26513));
   HB1xp67_ASAP7_75t_L FE_OCPC8260_n26335 (.Y(FE_OCPN8260_n26335),
	.A(n26335));
   HB1xp67_ASAP7_75t_R FE_OCPC8259_FE_OFN28686_FE_OCPN27812 (.Y(FE_OCPN8259_FE_OFN28686_FE_OCPN27812),
	.A(FE_OFN28686_FE_OCPN27812));
   HB1xp67_ASAP7_75t_L FE_OCPC8258_n26572 (.Y(FE_OCPN8258_n26572),
	.A(n26572));
   HB1xp67_ASAP7_75t_R FE_OCPC8257_n18178 (.Y(FE_OCPN8257_n18178),
	.A(n18178));
   HB1xp67_ASAP7_75t_L FE_OCPC8256_n16873 (.Y(FE_OCPN8256_n16873),
	.A(n16873));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8255_n21002 (.Y(FE_OCPN8255_n21002),
	.A(n21002));
   HB1xp67_ASAP7_75t_L FE_OCPC8254_w3_3 (.Y(FE_OCPN8254_w3_3),
	.A(FE_OCPN27978_w3_3));
   HB1xp67_ASAP7_75t_SL FE_OCPC8253_n17149 (.Y(FE_OCPN8253_n17149),
	.A(n17149));
   BUFx4f_ASAP7_75t_L FE_OCPC8252_FE_OFN28661_w3_7 (.Y(FE_OCPN8252_FE_OFN28661_w3_7),
	.A(FE_OFN28661_w3_7));
   HB1xp67_ASAP7_75t_R FE_OCPC8251_FE_OFN28672_sa01_2 (.Y(FE_OCPN8251_FE_OFN28672_sa01_2),
	.A(FE_OFN28672_sa01_2));
   HB1xp67_ASAP7_75t_L FE_OCPC8250_n22692 (.Y(FE_OCPN8250_n22692),
	.A(n22692));
   HB1xp67_ASAP7_75t_L FE_OCPC8249_n26944 (.Y(FE_OCPN8249_n26944),
	.A(n26944));
   HB1xp67_ASAP7_75t_L FE_OCPC8248_n16145 (.Y(FE_OCPN8248_n16145),
	.A(n16145));
   HB1xp67_ASAP7_75t_SL FE_OCPC8247_n21317 (.Y(FE_OCPN8247_n21317),
	.A(n21317));
   HB1xp67_ASAP7_75t_R FE_OCPC8246_n27143 (.Y(FE_OCPN8246_n27143),
	.A(n27143));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8245_n25295 (.Y(FE_OCPN8245_n25295),
	.A(n25295));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8244_n25778 (.Y(FE_OCPN8244_n25778),
	.A(n25778));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8243_n24899 (.Y(FE_OCPN8243_n24899),
	.A(n24899));
   HB1xp67_ASAP7_75t_R FE_OCPC8242_n20527 (.Y(FE_OCPN8242_n20527),
	.A(n20527));
   BUFx2_ASAP7_75t_L FE_OCPC8241_n22041 (.Y(FE_OCPN8241_n22041),
	.A(n22041));
   HB1xp67_ASAP7_75t_R FE_OCPC8240_n17618 (.Y(FE_OCPN8240_n17618),
	.A(n17618));
   HB1xp67_ASAP7_75t_R FE_OCPC8239_n24844 (.Y(FE_OCPN8239_n24844),
	.A(n24844));
   HB1xp67_ASAP7_75t_R FE_OCPC8238_n26472 (.Y(FE_OCPN8238_n26472),
	.A(n26472));
   HB1xp67_ASAP7_75t_L FE_OCPC8237_n21561 (.Y(FE_OCPN8237_n21561),
	.A(n21561));
   BUFx2_ASAP7_75t_L FE_OCPC8236_n22438 (.Y(FE_OCPN8236_n22438),
	.A(n22438));
   HB1xp67_ASAP7_75t_L FE_OCPC8235_n24589 (.Y(FE_OCPN8235_n24589),
	.A(n24589));
   HB1xp67_ASAP7_75t_L FE_OCPC8234_n25199 (.Y(FE_OCPN8234_n25199),
	.A(n25199));
   HB1xp67_ASAP7_75t_L FE_OCPC8233_n21647 (.Y(FE_OCPN8233_n21647),
	.A(n21647));
   BUFx2_ASAP7_75t_L FE_OCPC8232_FE_OFN27206_w3_30 (.Y(FE_OCPN8232_FE_OFN27206_w3_30),
	.A(FE_OFN27206_w3_30));
   BUFx2_ASAP7_75t_SL FE_OCPC8231_n20522 (.Y(FE_OCPN8231_n20522),
	.A(n20522));
   BUFx2_ASAP7_75t_R FE_OCPC8230_n20993 (.Y(FE_OCPN8230_n20993),
	.A(n20993));
   BUFx3_ASAP7_75t_SL FE_OCPC8229_n25750 (.Y(FE_OCPN8229_n25750),
	.A(n25750));
   HB1xp67_ASAP7_75t_SL FE_OCPC8228_n24165 (.Y(FE_OCPN8228_n24165),
	.A(n24165));
   BUFx3_ASAP7_75t_R FE_OCPC8227_n25950 (.Y(FE_OCPN8227_n25950),
	.A(n25950));
   OA21x2_ASAP7_75t_L FE_RC_1006_0 (.Y(n24171),
	.A1(n17176),
	.A2(n17173),
	.B(n17175));
   HB1xp67_ASAP7_75t_R FE_OCPC8226_n23113 (.Y(FE_OCPN8226_n23113),
	.A(n23113));
   HB1xp67_ASAP7_75t_R FE_OCPC8225_n26172 (.Y(FE_OCPN8225_n26172),
	.A(FE_OCPN27373_n26172));
   HB1xp67_ASAP7_75t_SL FE_OCPC8224_n22773 (.Y(FE_OCPN8224_n22773),
	.A(n22773));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8223_n16063 (.Y(FE_OCPN8223_n16063),
	.A(n16063));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8222_n27006 (.Y(FE_OCPN8222_n27006),
	.A(n27006));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8221_n26825 (.Y(FE_OCPN8221_n26825),
	.A(n26825));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8220_n26198 (.Y(FE_OCPN8220_n26198),
	.A(n26198));
   BUFx2_ASAP7_75t_SL FE_OCPC8219_n22197 (.Y(FE_OCPN8219_n22197),
	.A(n22197));
   BUFx3_ASAP7_75t_L FE_OCPC8218_n25507 (.Y(FE_OCPN8218_n25507),
	.A(n25507));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8217_n26319 (.Y(FE_OCPN8217_n26319),
	.A(n26319));
   HB1xp67_ASAP7_75t_R FE_OCPC8216_n13916 (.Y(FE_OCPN8216_n13916),
	.A(n13916));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8215_n25287 (.Y(FE_OCPN8215_n25287),
	.A(n25287));
   HB1xp67_ASAP7_75t_SL FE_OCPC8214_n27185 (.Y(FE_OCPN8214_n27185),
	.A(n27185));
   HB1xp67_ASAP7_75t_R FE_OCPC8213_FE_OFN29234_n16996 (.Y(FE_OCPN8213_FE_OFN29234_n16996),
	.A(FE_OFN29234_n16996));
   HB1xp67_ASAP7_75t_R FE_OCPC8212_n26261 (.Y(FE_OCPN8212_n26261),
	.A(n26261));
   HB1xp67_ASAP7_75t_R FE_OCPC8211_n24166 (.Y(FE_OCPN8211_n24166),
	.A(n24166));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8210_n25287 (.Y(FE_OCPN8210_n25287),
	.A(FE_OCPN8215_n25287));
   HB1xp67_ASAP7_75t_SL FE_OCPC8209_n26051 (.Y(FE_OCPN8209_n26051),
	.A(n26051));
   HB1xp67_ASAP7_75t_L FE_OCPC8208_n27094 (.Y(FE_OCPN8208_n27094),
	.A(n27094));
   BUFx6f_ASAP7_75t_SL FE_OCPC8207_n18497 (.Y(FE_OCPN8207_n18497),
	.A(n18497));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC8206_n25544 (.Y(FE_OCPN8206_n25544),
	.A(n25544));
   AOI21xp5_ASAP7_75t_L FE_RC_1005_0 (.Y(n568),
	.A1(key_36_),
	.A2(n16125),
	.B(n16079));
   OAI21x1_ASAP7_75t_L FE_RC_1004_0 (.Y(n26484),
	.A1(FE_RN_270_0),
	.A2(n26481),
	.B(n26480));
   XNOR2xp5_ASAP7_75t_SL FE_RC_1003_0 (.Y(FE_RN_247_0),
	.A(FE_OCPN29274_n26478),
	.B(n25268));
   OR3x2_ASAP7_75t_SL FE_RC_1002_0 (.Y(FE_OFN27123_n26275),
	.A(n23116),
	.B(n23115),
	.C(n23114));
   AOI31xp33_ASAP7_75t_R FE_RC_1001_0 (.Y(n17517),
	.A1(n17505),
	.A2(n24571),
	.A3(n22508),
	.B(n26078));
   AOI31xp33_ASAP7_75t_L FE_RC_1000_0 (.Y(n20777),
	.A1(n20776),
	.A2(n23189),
	.A3(n22852),
	.B(n26889));
   AO31x2_ASAP7_75t_L FE_RC_999_0 (.Y(n18868),
	.A1(n18867),
	.A2(FE_OFN27189_n),
	.A3(FE_OCPN7647_FE_OFN141_sa03_1),
	.B(n21308));
   AOI21xp5_ASAP7_75t_L FE_RC_998_0 (.Y(n21850),
	.A1(n21373),
	.A2(FE_OFN94_sa11_5),
	.B(n19200));
   AOI21xp5_ASAP7_75t_L FE_RC_997_0 (.Y(n22106),
	.A1(FE_OCPN29469_n17747),
	.A2(FE_OCPN27384_n22888),
	.B(n20208));
   AOI21xp5_ASAP7_75t_L FE_RC_996_0 (.Y(n18727),
	.A1(FE_OFN16208_n23101),
	.A2(n17382),
	.B(n23093));
   AOI21xp5_ASAP7_75t_L FE_RC_995_0 (.Y(n19445),
	.A1(n21327),
	.A2(FE_OCPN4680_n21317),
	.B(FE_OCPN27628_n23455));
   AOI21xp5_ASAP7_75t_L FE_RC_994_0 (.Y(n19095),
	.A1(FE_OCPN28021_n21445),
	.A2(n12998),
	.B(n19129));
   AOI21xp5_ASAP7_75t_SL FE_RC_993_0 (.Y(n15478),
	.A1(FE_OFN26053_n25415),
	.A2(FE_OFN28706_n),
	.B(FE_OFN5_w3_22));
   AOI31xp33_ASAP7_75t_SL FE_RC_992_0 (.Y(n22254),
	.A1(FE_OCPN27729_n24362),
	.A2(FE_OCPN28386_n17899),
	.A3(FE_OFN28764_n17928),
	.B(n22750));
   AOI31xp33_ASAP7_75t_SL FE_RC_991_0 (.Y(n24677),
	.A1(n19803),
	.A2(n19804),
	.A3(n19802),
	.B(n24978));
   BUFx2_ASAP7_75t_SL FE_OCPC8205_n449 (.Y(FE_OCPN29590_n449),
	.A(n449));
   BUFx2_ASAP7_75t_SL FE_OCPC8204_n426 (.Y(FE_OCPN29589_n426),
	.A(n426));
   BUFx2_ASAP7_75t_SL FE_OCPC8203_n457 (.Y(FE_OCPN29588_n457),
	.A(n457));
   AOI31xp33_ASAP7_75t_SL FE_RC_990_0 (.Y(n16484),
	.A1(n16482),
	.A2(n16483),
	.A3(n16710),
	.B(n23548));
   NOR3x2_ASAP7_75t_SL FE_RC_989_0 (.Y(n26149),
	.A(FE_OCPN28071_n25092),
	.B(FE_OCPN28107_n23504),
	.C(FE_OCPN29374_FE_OFN29191_sa23_2));
   HB1xp67_ASAP7_75t_L FE_OCPC8202_n26857 (.Y(FE_OCPN29587_n26857),
	.A(FE_OCPN29586_n26857));
   HB1xp67_ASAP7_75t_L FE_OCPC8201_n26857 (.Y(FE_OCPN29586_n26857),
	.A(n26857));
   OAI21xp33_ASAP7_75t_L FE_RC_988_0 (.Y(n17469),
	.A1(FE_OCPN28175_n21818),
	.A2(FE_OCPN27757_n21819),
	.B(n21858));
   INVx2_ASAP7_75t_SL FE_RC_987_0 (.Y(n27028),
	.A(FE_RN_286_0));
   OR2x2_ASAP7_75t_SRAM FE_RC_986_0 (.Y(FE_RN_287_0),
	.A(n27027),
	.B(FE_RN_213_0));
   AO21x1_ASAP7_75t_L FE_RC_985_0 (.Y(FE_RN_286_0),
	.A1(FE_RN_287_0),
	.A2(n27025),
	.B(n27024));
   INVx3_ASAP7_75t_SL FE_RC_984_0 (.Y(n18166),
	.A(FE_RN_285_0));
   AND2x2_ASAP7_75t_L FE_RC_983_0 (.Y(FE_RN_285_0),
	.A(FE_OFN16135_sa22_4),
	.B(n18165));
   XOR2xp5_ASAP7_75t_L FE_RC_982_0 (.Y(FE_RN_284_0),
	.A(FE_OCPN27234_n26837),
	.B(n24753));
   INVx1_ASAP7_75t_SL FE_RC_981_0 (.Y(FE_RN_283_0),
	.A(FE_RN_284_0));
   XOR2x1_ASAP7_75t_L FE_RC_980_0 (.Y(n24758),
	.A(FE_RN_283_0),
	.B(FE_OCPN7637_n25422));
   BUFx2_ASAP7_75t_SL FE_OCPC8200_n22281 (.Y(FE_OCPN29585_n22281),
	.A(n22281));
   NAND2xp5_ASAP7_75t_L FE_RC_979_0 (.Y(n21467),
	.A(FE_OCPN27679_n18631),
	.B(n17245));
   INVxp67_ASAP7_75t_L FE_RC_978_0 (.Y(FE_RN_282_0),
	.A(FE_OCPN27818_n17267));
   AND3x4_ASAP7_75t_SL FE_RC_977_0 (.Y(n19845),
	.A(FE_RN_282_0),
	.B(FE_OCPN27679_n18631),
	.C(n17245));
   BUFx2_ASAP7_75t_SL FE_OCPC8199_sa20_1 (.Y(FE_OCPN29584_n),
	.A(FE_OCPN29380_sa20_1));
   NAND3x1_ASAP7_75t_L FE_RC_976_0 (.Y(n24142),
	.A(n20385),
	.B(FE_OCPN28427_n25064),
	.C(n25063));
   BUFx2_ASAP7_75t_SL FE_OCPC8198_n15422 (.Y(FE_OCPN29583_n15422),
	.A(n15422));
   NOR3x1_ASAP7_75t_L FE_RC_975_0 (.Y(n15080),
	.A(FE_OFN28732_n),
	.B(FE_OCPN29537_FE_OFN28699_w3_6),
	.C(n25140));
   NOR3x1_ASAP7_75t_R FE_RC_974_0 (.Y(n26258),
	.A(n25087),
	.B(n25089),
	.C(FE_OFN28511_n25088));
   INVxp67_ASAP7_75t_L FE_RC_973_0 (.Y(FE_RN_278_0),
	.A(n24556));
   INVxp33_ASAP7_75t_L FE_RC_972_0 (.Y(FE_RN_279_0),
	.A(n17463));
   NAND2xp5_ASAP7_75t_L FE_RC_971_0 (.Y(FE_RN_280_0),
	.A(FE_RN_278_0),
	.B(FE_RN_279_0));
   NAND2xp5_ASAP7_75t_R FE_RC_970_0 (.Y(FE_RN_281_0),
	.A(FE_RN_129_0),
	.B(n24553));
   AOI22xp5_ASAP7_75t_SL FE_RC_969_0 (.Y(n26389),
	.A1(FE_RN_281_0),
	.A2(n24315),
	.B1(FE_RN_280_0),
	.B2(n24318));
   BUFx2_ASAP7_75t_SL FE_OCPC8196_n16097 (.Y(FE_OCPN29581_n16097),
	.A(n16097));
   HB1xp67_ASAP7_75t_SL FE_OCPC8195_sa21_2 (.Y(FE_OCPN29580_n),
	.A(FE_OCPN27328_sa21_2));
   OAI21x1_ASAP7_75t_SL FE_RC_968_0 (.Y(n16156),
	.A1(n16152),
	.A2(w2_7_),
	.B(n16151));
   BUFx2_ASAP7_75t_L FE_OCPC8194_n18837 (.Y(FE_OCPN29579_n18837),
	.A(n18837));
   HB1xp67_ASAP7_75t_SL FE_OCPC8193_FE_OFN27214_w3_17 (.Y(FE_OCPN29578_FE_OFN27214_w3_17),
	.A(FE_OFN27214_w3_17));
   BUFx2_ASAP7_75t_SL FE_OCPC8192_n24298 (.Y(FE_OCPN29577_n24298),
	.A(n24298));
   AOI21x1_ASAP7_75t_SL FE_RC_967_0 (.Y(n416),
	.A1(n25944),
	.A2(FE_RN_114_0),
	.B(n25943));
   BUFx2_ASAP7_75t_SL FE_OCPC8191_n26930 (.Y(FE_OCPN29576_n26930),
	.A(n26930));
   OAI222xp33_ASAP7_75t_SL FE_RC_966_0 (.Y(n18233),
	.A1(n18232),
	.A2(n23345),
	.B1(n20745),
	.B2(n23345),
	.C1(n22806),
	.C2(n23345));
   OAI22xp33_ASAP7_75t_SL FE_RC_965_0 (.Y(n589),
	.A1(FE_OFN26646_n16159),
	.A2(ld),
	.B1(FE_OFN26646_n16159),
	.B2(key_58_));
   BUFx3_ASAP7_75t_SL FE_OCPC8189_n484 (.Y(FE_OCPN29574_n484),
	.A(n484));
   AOI31xp33_ASAP7_75t_SL FE_RC_964_0 (.Y(n21574),
	.A1(n24205),
	.A2(n21573),
	.A3(n21572),
	.B(n27004));
   BUFx2_ASAP7_75t_L FE_OCPC8188_n15184 (.Y(FE_OCPN29573_n15184),
	.A(n15184));
   HB1xp67_ASAP7_75t_L FE_OCPC8187_n24468 (.Y(FE_OCPN29572_n24468),
	.A(n24468));
   BUFx2_ASAP7_75t_L FE_OCPC8186_n26355 (.Y(FE_OCPN29571_n26355),
	.A(n26355));
   BUFx3_ASAP7_75t_SL FE_OCPC8185_n15423 (.Y(FE_OCPN29570_n15423),
	.A(n15423));
   NAND3x1_ASAP7_75t_L FE_RC_963_0 (.Y(n23127),
	.A(n19787),
	.B(FE_OCPN28040_n19766),
	.C(FE_OFN27196_n));
   OAI222xp33_ASAP7_75t_L FE_RC_962_0 (.Y(n18436),
	.A1(n18429),
	.A2(n23548),
	.B1(n23548),
	.B2(n18446),
	.C1(n23548),
	.C2(n18445));
   OAI22x1_ASAP7_75t_SL FE_RC_961_0 (.Y(n15901),
	.A1(n25648),
	.A2(FE_OFN21_n16125),
	.B1(n15902),
	.B2(FE_OFN21_n16125));
   OAI22xp33_ASAP7_75t_L FE_RC_960_0 (.Y(n13961),
	.A1(FE_OCPN29536_FE_OFN8_w3_14),
	.A2(n14098),
	.B1(FE_OFN28856_n15450),
	.B2(n14098));
   BUFx2_ASAP7_75t_L FE_OCPC8184_n18947 (.Y(FE_OCPN29569_n18947),
	.A(n18947));
   OAI21xp5_ASAP7_75t_SL FE_RC_959_0 (.Y(n17154),
	.A1(FE_OCPN27836_n16976),
	.A2(FE_OFN28775_n16992),
	.B(n27089));
   INVx2_ASAP7_75t_SL FE_RC_958_0 (.Y(n26418),
	.A(FE_RN_276_0));
   AND2x2_ASAP7_75t_L FE_RC_957_0 (.Y(FE_RN_277_0),
	.A(FE_OCPN7625_n26501),
	.B(FE_OFN16215_ld_r));
   OA21x2_ASAP7_75t_SL FE_RC_956_0 (.Y(FE_RN_276_0),
	.A1(FE_RN_277_0),
	.A2(n26414),
	.B(n26413));
   AOI31xp33_ASAP7_75t_SL FE_RC_955_0 (.Y(n22570),
	.A1(n22558),
	.A2(n22557),
	.A3(n22559),
	.B(n26976));
   BUFx2_ASAP7_75t_SL FE_OCPC8183_n18257 (.Y(FE_OCPN29568_n18257),
	.A(n18257));
   OAI21xp5_ASAP7_75t_SL FE_RC_954_0 (.Y(n23522),
	.A1(FE_OCPN29488_FE_OFN25883_n22945),
	.A2(FE_OFN28841_n22980),
	.B(n22036));
   BUFx3_ASAP7_75t_SL FE_OCPC8182_n23806 (.Y(FE_OCPN29567_n23806),
	.A(n23806));
   BUFx2_ASAP7_75t_SL FE_OCPC8180_n432 (.Y(FE_OCPN29565_n432),
	.A(n432));
   HB1xp67_ASAP7_75t_L FE_OCPC8179_n16012 (.Y(FE_OCPN29564_n16012),
	.A(n16012));
   OAI21x1_ASAP7_75t_SL FE_RC_953_0 (.Y(n15776),
	.A1(n15367),
	.A2(n24200),
	.B(n15366));
   BUFx2_ASAP7_75t_L FE_OCPC8178_n18602 (.Y(FE_OCPN29563_n18602),
	.A(n18602));
   NAND3x1_ASAP7_75t_L FE_RC_952_0 (.Y(n20153),
	.A(FE_OCPN27570_n17791),
	.B(FE_OFN28730_FE_OCPN28416_sa02_3),
	.C(FE_OFN28703_FE_OCPN27740_sa02_4));
   NOR2xp33_ASAP7_75t_L FE_RC_951_0 (.Y(FE_RN_271_0),
	.A(FE_OFN26072_n26720),
	.B(text_in_r_20_));
   INVxp67_ASAP7_75t_L FE_RC_950_0 (.Y(FE_RN_272_0),
	.A(n26734));
   NOR2xp33_ASAP7_75t_L FE_RC_949_0 (.Y(FE_RN_273_0),
	.A(FE_RN_271_0),
	.B(FE_RN_272_0));
   OAI21xp33_ASAP7_75t_SL FE_RC_948_0 (.Y(FE_RN_274_0),
	.A1(n26732),
	.A2(FE_OFN16214_ld_r),
	.B(n26731));
   INVxp67_ASAP7_75t_SL FE_RC_947_0 (.Y(FE_RN_275_0),
	.A(n26730));
   AOI21x1_ASAP7_75t_L FE_RC_946_0 (.Y(n517),
	.A1(FE_RN_275_0),
	.A2(FE_RN_274_0),
	.B(FE_RN_273_0));
   HB1xp67_ASAP7_75t_SL FE_OCPC8177_n25138 (.Y(FE_OCPN29562_n25138),
	.A(n25138));
   OAI21xp33_ASAP7_75t_SL FE_RC_945_0 (.Y(n17414),
	.A1(FE_OCPN28127_n16872),
	.A2(n16874),
	.B(n16959));
   NAND3x1_ASAP7_75t_SL FE_RC_944_0 (.Y(n24182),
	.A(n16299),
	.B(FE_OFN16415_sa31_2),
	.C(n16295));
   NAND3x1_ASAP7_75t_L FE_RC_943_0 (.Y(n23172),
	.A(n18161),
	.B(FE_OCPN27979_FE_OFN16147_sa22_1),
	.C(FE_PSN8320_n18176));
   BUFx2_ASAP7_75t_SL FE_OCPC8176_n23532 (.Y(FE_OCPN29561_n23532),
	.A(n23532));
   OAI21xp5_ASAP7_75t_SL FE_RC_941_0 (.Y(n27066),
	.A1(n27067),
	.A2(n27068),
	.B(FE_OFN15_FE_DBTN0_ld_r));
   OAI21x1_ASAP7_75t_SL FE_RC_940_0 (.Y(n24306),
	.A1(n24305),
	.A2(FE_RN_118_0),
	.B(n24304));
   BUFx3_ASAP7_75t_SL FE_OCPC8174_n17900 (.Y(FE_OCPN29559_n17900),
	.A(n17900));
   BUFx2_ASAP7_75t_L FE_OCPC8172_n18161 (.Y(FE_OCPN29557_n18161),
	.A(n18161));
   AOI31xp33_ASAP7_75t_SL FE_RC_939_0 (.Y(n24167),
	.A1(n17141),
	.A2(n17140),
	.A3(n18262),
	.B(n27095));
   BUFx3_ASAP7_75t_SL FE_OCPC8171_n383 (.Y(FE_OCPN29556_n383),
	.A(n383));
   AOI31xp33_ASAP7_75t_SL FE_RC_938_0 (.Y(n23005),
	.A1(n23003),
	.A2(n23004),
	.A3(n23002),
	.B(n26710));
   NAND3x1_ASAP7_75t_L FE_RC_937_0 (.Y(n25220),
	.A(n17048),
	.B(n17049),
	.C(FE_OCPN8228_n24165));
   AOI21xp5_ASAP7_75t_L FE_RC_936_0 (.Y(n23786),
	.A1(n23784),
	.A2(n26323),
	.B(n23785));
   NAND3x1_ASAP7_75t_R FE_RC_935_0 (.Y(n23950),
	.A(n24955),
	.B(FE_OCPN28052_sa10_1),
	.C(n23035));
   AOI21xp5_ASAP7_75t_SL FE_RC_934_0 (.Y(n26274),
	.A1(FE_OFN2_ld_r),
	.A2(text_in_r_111_),
	.B(n26269));
   AOI31xp33_ASAP7_75t_SL FE_RC_933_0 (.Y(n26074),
	.A1(n21387),
	.A2(n24081),
	.A3(FE_OCPN29416_n22516),
	.B(n17463));
   HB1xp67_ASAP7_75t_L FE_OCPC8170_n20593 (.Y(FE_OCPN29555_n20593),
	.A(n20593));
   HB1xp67_ASAP7_75t_L FE_OCPC8169_n22507 (.Y(FE_OCPN29554_n22507),
	.A(n22507));
   BUFx2_ASAP7_75t_L FE_OCPC8168_n19602 (.Y(FE_OCPN29553_n19602),
	.A(n19602));
   BUFx2_ASAP7_75t_SL FE_OCPC8167_n393 (.Y(FE_OCPN29552_n393),
	.A(n393));
   HB1xp67_ASAP7_75t_L FE_OCPC8166_sa23_3 (.Y(FE_OCPN29551_n),
	.A(FE_OCPN29489_sa23_3));
   AND2x2_ASAP7_75t_SRAM FE_RC_931_0 (.Y(FE_RN_270_0),
	.A(n27117),
	.B(FE_PSN8300_n26482));
   AOI31xp33_ASAP7_75t_SL FE_RC_929_0 (.Y(n22863),
	.A1(n22861),
	.A2(n22862),
	.A3(n22860),
	.B(n26889));
   BUFx2_ASAP7_75t_SL FE_OCPC8165_n16114 (.Y(FE_OCPN29550_n16114),
	.A(n16114));
   AOI31xp33_ASAP7_75t_SL FE_RC_928_0 (.Y(n21184),
	.A1(n21182),
	.A2(n21183),
	.A3(n21181),
	.B(n21493));
   BUFx2_ASAP7_75t_L FE_OCPC8163_n25717 (.Y(FE_OCPN29548_n25717),
	.A(n25717));
   NAND3x2_ASAP7_75t_SL FE_RC_927_0 (.Y(n20527),
	.A(FE_OFN27186_sa13_4),
	.B(FE_OFN16181_sa13_5),
	.C(FE_OFN16268_sa13_3));
   OAI222xp33_ASAP7_75t_L FE_RC_926_0 (.Y(n26235),
	.A1(n17151),
	.A2(n26959),
	.B1(n26959),
	.B2(n25549),
	.C1(n26959),
	.C2(n25197));
   BUFx2_ASAP7_75t_SL FE_OCPC8162_n15183 (.Y(FE_OCPN29547_n15183),
	.A(n15183));
   OAI21xp33_ASAP7_75t_SL FE_RC_925_0 (.Y(n25677),
	.A1(FE_OCPN27362_n25679),
	.A2(n25678),
	.B(FE_OFN28490_ld_r));
   AOI31xp33_ASAP7_75t_SL FE_RC_924_0 (.Y(n25295),
	.A1(n19427),
	.A2(n27088),
	.A3(FE_RN_231_0),
	.B(n27095));
   OAI21xp33_ASAP7_75t_L FE_RC_923_0 (.Y(n21464),
	.A1(sa00_5_),
	.A2(n21152),
	.B(n21451));
   INVx2_ASAP7_75t_SL FE_RC_922_0 (.Y(n26431),
	.A(FE_RN_268_0));
   OR3x1_ASAP7_75t_SL FE_RC_921_0 (.Y(FE_RN_268_0),
	.A(n16926),
	.B(FE_OFN28936_n18104),
	.C(n18135));
   HB1xp67_ASAP7_75t_SL FE_OCPC8161_n19275 (.Y(FE_OCPN29546_n),
	.A(FE_OCPN27771_n19275));
   BUFx3_ASAP7_75t_SL FE_OCPC8160_n22529 (.Y(FE_OCPN29545_n22529),
	.A(n22529));
   NAND3x2_ASAP7_75t_SL FE_RC_920_0 (.Y(n23259),
	.A(FE_OFN29054_n17453),
	.B(FE_OCPN28321_n21341),
	.C(FE_OFN94_sa11_5));
   BUFx6f_ASAP7_75t_SL FE_OCPC8159_n20527 (.Y(FE_OCPN29544_n20527),
	.A(n20527));
   AOI21x1_ASAP7_75t_SL FE_RC_919_0 (.Y(FE_OCPN27419_n26602),
	.A1(FE_RN_126_0),
	.A2(n24806),
	.B(n24805));
   BUFx2_ASAP7_75t_L FE_OCPC8158_FE_OFN28862_n (.Y(FE_OCPN29543_FE_OFN28862_n),
	.A(FE_OFN28862_n));
   BUFx3_ASAP7_75t_SL FE_OCPC8157_n21151 (.Y(FE_OCPN29542_n21151),
	.A(n21151));
   BUFx3_ASAP7_75t_SL FE_OCPC8156_n25870 (.Y(FE_OCPN29541_n25870),
	.A(n25870));
   AND2x2_ASAP7_75t_R FE_RC_918_0 (.Y(FE_RN_267_0),
	.A(n18764),
	.B(FE_OCPN7640_n18765));
   NAND2xp5_ASAP7_75t_SL FE_RC_917_0 (.Y(n18769),
	.A(FE_RN_267_0),
	.B(n18763));
   AOI31xp33_ASAP7_75t_SL FE_RC_916_0 (.Y(n19155),
	.A1(n19153),
	.A2(n19154),
	.A3(n19152),
	.B(n21493));
   NOR3x1_ASAP7_75t_R FE_RC_915_0 (.Y(n24155),
	.A(n17065),
	.B(n17115),
	.C(FE_OFN28725_n16982));
   HB1xp67_ASAP7_75t_L FE_OCPC8155_FE_OFN25927_n26527 (.Y(FE_OCPN29540_FE_OFN25927_n26527),
	.A(FE_OFN25927_n26527));
   INVx1_ASAP7_75t_SL FE_OCPC8154_n24927 (.Y(FE_OCPN29539_n24927),
	.A(FE_OFN16260_n24927));
   INVx1_ASAP7_75t_L FE_OCPC8153_n24927 (.Y(FE_OCPN29538_n24927),
	.A(n24925));
   INVxp67_ASAP7_75t_L FE_OCPC8152_n24927 (.Y(FE_OFN16260_n24927),
	.A(n24925));
   INVx2_ASAP7_75t_SL FE_OCPC8151_n24927 (.Y(n24925),
	.A(n24927));
   INVx3_ASAP7_75t_SL FE_OCPC8150_n16534 (.Y(FE_OCPN28157_n16534),
	.A(FE_OFN28911_n16534));
   INVx1_ASAP7_75t_SL FE_OCPC8149_n16534 (.Y(FE_OFN28911_n16534),
	.A(n16534));
   BUFx3_ASAP7_75t_SL FE_OCPC8148_n18177 (.Y(FE_OCPN27947_n18177),
	.A(n18177));
   INVx2_ASAP7_75t_L FE_OCPC8147_FE_OFN28699_w3_6 (.Y(FE_OCPN29537_FE_OFN28699_w3_6),
	.A(FE_OFN28734_n));
   INVxp67_ASAP7_75t_L FE_OCPC8145_FE_OFN28699_w3_6 (.Y(FE_OFN28734_n),
	.A(FE_OFN28699_w3_6));
   INVxp67_ASAP7_75t_L FE_OCPC8144_n16263 (.Y(FE_OFN16361_n16263),
	.A(FE_OFN25892_n16264));
   BUFx3_ASAP7_75t_SL FE_OCPC8143_n16263 (.Y(FE_OFN25892_n16264),
	.A(n16263));
   INVx3_ASAP7_75t_SL FE_OCPC8142_FE_OFN8_w3_14 (.Y(FE_OCPN29536_FE_OFN8_w3_14),
	.A(FE_OFN28894_n));
   INVx4_ASAP7_75t_SL FE_OCPC8141_FE_OFN8_w3_14 (.Y(FE_OCPN29535_FE_OFN8_w3_14),
	.A(FE_OFN28894_n));
   INVx2_ASAP7_75t_SL FE_OCPC8140_FE_OFN8_w3_14 (.Y(FE_OCPN29534_FE_OFN8_w3_14),
	.A(FE_OFN28894_n));
   BUFx3_ASAP7_75t_SL FE_OCPC8139_FE_OFN8_w3_14 (.Y(FE_OFN28894_n),
	.A(FE_OFN8_w3_14));
   INVx4_ASAP7_75t_SL FE_OCPC8138_n17993 (.Y(FE_OFN29158_n18860),
	.A(n17993));
   BUFx3_ASAP7_75t_SL FE_OCPC8137_n14091 (.Y(n14090),
	.A(n14091));
   INVx1_ASAP7_75t_SL FE_OCPC8136_n14091 (.Y(FE_OFN27216_n14091),
	.A(n14091));
   BUFx2_ASAP7_75t_L FE_OCPC8135_n26971 (.Y(FE_OCPN29533_n26971),
	.A(FE_OCPN27624_n26971));
   BUFx3_ASAP7_75t_SL FE_OCPC8134_n26971 (.Y(FE_OCPN27624_n26971),
	.A(n26971));
   INVxp67_ASAP7_75t_SL FE_OCPC8133_n25697 (.Y(FE_OCPN29532_n25697),
	.A(n25697));
   INVx1_ASAP7_75t_SL FE_OCPC8131_FE_OFN25926_n26922 (.Y(FE_OCPN29531_FE_OFN25926_n26922),
	.A(FE_OFN25926_n26922));
   INVx1_ASAP7_75t_SL FE_OCPC8129_FE_OFN25926_n26922 (.Y(n26923),
	.A(FE_OFN25926_n26922));
   INVxp67_ASAP7_75t_SL FE_OCPC8128_n27033 (.Y(FE_RN_151_0),
	.A(n27033));
   INVxp67_ASAP7_75t_L FE_OCPC8127_n23125 (.Y(FE_OCPN29529_n23125),
	.A(n24725));
   INVx1_ASAP7_75t_SL FE_OCPC8126_n23125 (.Y(n24725),
	.A(n23125));
   INVxp67_ASAP7_75t_SL FE_OCPC8124_n25721 (.Y(n25719),
	.A(n25721));
   INVxp67_ASAP7_75t_SL FE_OCPC8123_n16751 (.Y(FE_OCPN27367_sa21_0),
	.A(n16751));
   BUFx2_ASAP7_75t_SL FE_OCPC8122_n22850 (.Y(FE_OFN29195_n22850),
	.A(n22850));
   BUFx2_ASAP7_75t_SL FE_OCPC8120_n16581 (.Y(FE_OCPN29498_n16581),
	.A(n16581));
   BUFx3_ASAP7_75t_SL FE_OCPC8119_n25389 (.Y(FE_OCPN27292_n25389),
	.A(n25389));
   INVx3_ASAP7_75t_SL FE_OCPC8117_n16923 (.Y(FE_OFN28998_n16923),
	.A(n16923));
   INVxp67_ASAP7_75t_SL FE_OCPC8116_n24138 (.Y(FE_OCPN29528_n24138),
	.A(n24139));
   INVxp33_ASAP7_75t_L FE_OCPC8115_n24138 (.Y(FE_OCPN29527_n24138),
	.A(n24139));
   INVx2_ASAP7_75t_SL FE_OCPC8114_n24138 (.Y(n24139),
	.A(n24138));
   INVx3_ASAP7_75t_SL FE_OCPC8113_sa31_4 (.Y(FE_OCPN29526_sa31_4),
	.A(FE_OFN26595_sa31_4));
   INVx1_ASAP7_75t_SL FE_OCPC8112_sa31_4 (.Y(n16298),
	.A(FE_OFN26595_sa31_4));
   INVx3_ASAP7_75t_SL FE_OCPC8111_sa31_4 (.Y(FE_OFN26595_sa31_4),
	.A(sa31_4_));
   BUFx2_ASAP7_75t_L FE_OCPC8110_n18947 (.Y(FE_OCPN29525_n18947),
	.A(n25991));
   INVx2_ASAP7_75t_SL FE_OCPC8109_n18947 (.Y(n25991),
	.A(n18947));
   INVx1_ASAP7_75t_SL FE_OCPC8108_n25029 (.Y(FE_OCPN29524_n25029),
	.A(FE_OFN26577_n));
   BUFx3_ASAP7_75t_SL FE_OCPC8107_n25029 (.Y(FE_OFN26577_n),
	.A(n25029));
   BUFx2_ASAP7_75t_SL FE_OCPC8106_n25029 (.Y(n19920),
	.A(n25029));
   INVxp67_ASAP7_75t_SL FE_OCPC8105_n25544 (.Y(FE_OCPN29523_n25544),
	.A(n25544));
   HB1xp67_ASAP7_75t_SL FE_OCPC8103_n23558 (.Y(FE_OFN29005_n23558),
	.A(n23558));
   INVxp67_ASAP7_75t_SL FE_OCPC8102_n23558 (.Y(FE_OFN27089_n23558),
	.A(n23558));
   INVx1_ASAP7_75t_L FE_OCPC8100_n24755 (.Y(FE_OCPN29521_n24755),
	.A(FE_OFN101_w3_12));
   INVx1_ASAP7_75t_SL FE_OCPC8099_n24755 (.Y(FE_OCPN29520_n24755),
	.A(n24755));
   INVxp67_ASAP7_75t_L FE_OCPC8098_n24755 (.Y(FE_OFN101_w3_12),
	.A(n24755));
   INVxp67_ASAP7_75t_L FE_OCPC8097_n18871 (.Y(n18051),
	.A(FE_OCPN27975_n18871));
   BUFx2_ASAP7_75t_SL FE_OCPC8096_n20064 (.Y(FE_OCPN27444_n20064),
	.A(n20064));
   INVxp67_ASAP7_75t_SL FE_OCPC8095_n20007 (.Y(FE_OCPN29519_n),
	.A(FE_OCPN27554_n20007));
   HB1xp67_ASAP7_75t_L FE_OCPC8094_n20007 (.Y(FE_OFN27140_n20007),
	.A(FE_OCPN27554_n20007));
   INVxp67_ASAP7_75t_L FE_OCPC8092_FE_OFN25874_sa03_2 (.Y(FE_OCPN29517_n),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2));
   HB1xp67_ASAP7_75t_L FE_OCPC8090_FE_OFN25874_sa03_2 (.Y(FE_OFN27189_n),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2));
   BUFx6f_ASAP7_75t_SL FE_OCPC8089_n17475 (.Y(FE_OCPN27601_n17475),
	.A(n17475));
   HB1xp67_ASAP7_75t_L FE_OCPC8088_n27136 (.Y(FE_OCPN29515_n27136),
	.A(FE_OCPN29514_n27136));
   INVx1_ASAP7_75t_SL FE_OCPC8087_n27136 (.Y(FE_OCPN29514_n27136),
	.A(n27136));
   INVx1_ASAP7_75t_SL FE_OCPC8085_n17429 (.Y(n17430),
	.A(n17429));
   BUFx2_ASAP7_75t_SL FE_OCPC8084_n17447 (.Y(FE_OCPN29513_n17447),
	.A(n17447));
   BUFx2_ASAP7_75t_SL FE_OCPC8083_n17447 (.Y(FE_OCPN29439_n17447),
	.A(n17447));
   INVx1_ASAP7_75t_L FE_OCPC8082_n16750 (.Y(FE_OCPN29512_n16750),
	.A(FE_OCPN27735_n16750));
   INVx3_ASAP7_75t_SL FE_OCPC8081_n16750 (.Y(FE_OFN29023_n16750),
	.A(FE_OCPN27735_n16750));
   INVx2_ASAP7_75t_SL FE_OCPC8080_n16750 (.Y(FE_OCPN27735_n16750),
	.A(n16750));
   INVxp67_ASAP7_75t_SL FE_OCPC8079_n20395 (.Y(n20396),
	.A(n20395));
   INVxp67_ASAP7_75t_SL FE_OCPC8078_n22226 (.Y(FE_OCPN29511_n22226),
	.A(n22226));
   HB1xp67_ASAP7_75t_SL FE_OCPC8076_n23357 (.Y(FE_OCPN27605_n23357),
	.A(n23357));
   BUFx2_ASAP7_75t_SL FE_OCPC8075_n25444 (.Y(n25710),
	.A(FE_OFN29143_n25444));
   INVx1_ASAP7_75t_SL FE_OCPC8074_n25444 (.Y(FE_OFN29143_n25444),
	.A(n25444));
   INVxp67_ASAP7_75t_SL FE_OCPC8073_n26363 (.Y(n26361),
	.A(n26363));
   BUFx6f_ASAP7_75t_SL FE_OCPC8072_sa30_1 (.Y(FE_OFN16247_sa30_1),
	.A(sa30_1_));
   BUFx6f_ASAP7_75t_SL FE_OCPC8071_n21845 (.Y(FE_OCPN27313_n21845),
	.A(n21845));
   INVxp67_ASAP7_75t_SL FE_OCPC8070_n15776 (.Y(n15777),
	.A(n15776));
   INVx1_ASAP7_75t_L FE_OCPC8069_n14745 (.Y(n14744),
	.A(n14745));
   BUFx2_ASAP7_75t_SL FE_OCPC8068_n14745 (.Y(FE_OFN27218_n14745),
	.A(n14745));
   BUFx4f_ASAP7_75t_SL FE_OCPC8067_n16189 (.Y(FE_OFN16253_n16189),
	.A(n16189));
   HB1xp67_ASAP7_75t_SL FE_OCPC8066_n16996 (.Y(FE_OCPN29510_n16996),
	.A(FE_OFN29234_n16996));
   BUFx3_ASAP7_75t_SL FE_OCPC8065_n16996 (.Y(FE_OFN29234_n16996),
	.A(n16996));
   BUFx2_ASAP7_75t_L FE_OCPC8063_FE_OFN16184_w3_9 (.Y(FE_OCPN29509_FE_OFN16184_w3_9),
	.A(FE_OCPN29506_FE_OFN16184_w3_9));
   INVx6_ASAP7_75t_SL FE_OCPC8062_FE_OFN16184_w3_9 (.Y(FE_OCPN29508_FE_OFN16184_w3_9),
	.A(FE_OCPN7616_FE_OFN16184_w3_9));
   BUFx5_ASAP7_75t_SL FE_OCPC8060_FE_OFN16184_w3_9 (.Y(FE_OCPN29506_FE_OFN16184_w3_9),
	.A(FE_OFN16184_w3_9));
   INVx2_ASAP7_75t_SL FE_OCPC8059_FE_OFN16184_w3_9 (.Y(FE_OCPN7616_FE_OFN16184_w3_9),
	.A(FE_OFN16184_w3_9));
   BUFx2_ASAP7_75t_SL FE_OCPC8058_n22380 (.Y(FE_OCPN28392_n22380),
	.A(n22380));
   BUFx3_ASAP7_75t_SL FE_OCPC8057_n22448 (.Y(FE_OCPN28301_n22448),
	.A(n22448));
   INVx1_ASAP7_75t_SL FE_OCPC8056_n16534 (.Y(FE_OFN28910_n16534),
	.A(FE_OFN28912_n16534));
   INVx1_ASAP7_75t_SL FE_OCPC8054_n16534 (.Y(FE_OFN28912_n16534),
	.A(FE_OFN28911_n16534));
   INVxp67_ASAP7_75t_L FE_OCPC8053_n22457 (.Y(FE_OCPN29505_n22457),
	.A(FE_OFN78_n22457));
   INVx1_ASAP7_75t_SL FE_OCPC8052_n22457 (.Y(FE_OFN78_n22457),
	.A(n22457));
   BUFx4f_ASAP7_75t_SL FE_OCPC8051_n18206 (.Y(FE_OFN26548_n18206),
	.A(n18206));
   INVx3_ASAP7_75t_SL FE_OCPC8050_sa11_4 (.Y(FE_OCPN29504_sa11_4),
	.A(FE_OCPN27365_sa11_4));
   INVx2_ASAP7_75t_SL FE_OCPC8048_sa11_4 (.Y(FE_OCPN27365_sa11_4),
	.A(sa11_4_));
   INVx1_ASAP7_75t_R FE_OCPC8047_n24627 (.Y(FE_OCPN29503_n24627),
	.A(n24630));
   INVx1_ASAP7_75t_SL FE_OCPC8046_n24627 (.Y(n24630),
	.A(n24627));
   BUFx2_ASAP7_75t_SL FE_OCPC8044_n26103 (.Y(FE_OFN28767_n26103),
	.A(n26103));
   HB1xp67_ASAP7_75t_L FE_OCPC8043_w3_23 (.Y(FE_OCPN29502_w3_23),
	.A(FE_OFN37_w3_23));
   INVxp67_ASAP7_75t_L FE_OCPC8042_w3_23 (.Y(FE_OFN28908_w3_23),
	.A(FE_OFN37_w3_23));
   BUFx3_ASAP7_75t_SL FE_OCPC8041_w3_23 (.Y(FE_OFN28_w3_23),
	.A(w3_23_));
   INVx3_ASAP7_75t_SL FE_OCPC8040_w3_23 (.Y(FE_OFN37_w3_23),
	.A(w3_23_));
   HB1xp67_ASAP7_75t_L FE_OCPC8039_FE_OFN28662_w3_7 (.Y(FE_OCPN29501_FE_OFN28662_w3_7),
	.A(FE_OCPN29500_FE_OFN28662_w3_7));
   INVx2_ASAP7_75t_SL FE_OCPC8038_FE_OFN28662_w3_7 (.Y(FE_OCPN29500_FE_OFN28662_w3_7),
	.A(FE_OFN28662_w3_7));
   INVx1_ASAP7_75t_SL FE_OCPC8036_FE_OFN16131_sa12_1 (.Y(FE_OCPN29499_FE_OFN16131_sa12_1),
	.A(FE_OFN16131_sa12_1));
   INVx3_ASAP7_75t_SL FE_OCPC8035_FE_OFN16131_sa12_1 (.Y(FE_OFN28764_n17928),
	.A(FE_OFN16131_sa12_1));
   INVxp67_ASAP7_75t_SL FE_OCPC8034_FE_OFN16131_sa12_1 (.Y(n17928),
	.A(FE_OFN16131_sa12_1));
   BUFx2_ASAP7_75t_SL FE_OCPC8031_n20195 (.Y(FE_OCPN27503_n20195),
	.A(n20195));
   BUFx2_ASAP7_75t_R FE_OCPC8030_FE_OFN27148_sa32_3 (.Y(FE_OCPN27230_sa32_3),
	.A(FE_OFN27148_sa32_3));
   BUFx2_ASAP7_75t_L FE_OCPC8026_sa21_1 (.Y(FE_OCPN29497_sa21_1),
	.A(FE_OFN28698_sa21_1));
   BUFx6f_ASAP7_75t_SL FE_OCPC8025_sa21_1 (.Y(FE_OFN28698_sa21_1),
	.A(sa21_1_));
   INVxp67_ASAP7_75t_L FE_OCPC8024_n24789 (.Y(FE_OCPN29496_n24789),
	.A(n21592));
   INVx2_ASAP7_75t_SL FE_OCPC8022_n24789 (.Y(n21592),
	.A(n24789));
   INVxp67_ASAP7_75t_SL FE_OCPC8021_n25168 (.Y(n25166),
	.A(n25168));
   INVx3_ASAP7_75t_L FE_OCPC8020_sa30_0 (.Y(n17601),
	.A(FE_OFN28925_sa30_0));
   INVx3_ASAP7_75t_SL FE_OCPC8019_sa30_0 (.Y(FE_OCPN28049_sa30_0),
	.A(FE_OFN28925_sa30_0));
   INVx4_ASAP7_75t_SL FE_OCPC8018_sa30_0 (.Y(FE_OFN28925_sa30_0),
	.A(sa30_0_));
   BUFx2_ASAP7_75t_SL FE_OCPC8017_n25524 (.Y(FE_OCPN29318_n25524),
	.A(n25524));
   BUFx2_ASAP7_75t_SL FE_OCPC8016_n27049 (.Y(FE_OFN29142_n27049),
	.A(n27049));
   INVx1_ASAP7_75t_SL FE_OCPC8015_n25414 (.Y(FE_OFN28902_n25414),
	.A(FE_OCPN27682_n25414));
   INVx2_ASAP7_75t_SL FE_OCPC8014_n25414 (.Y(FE_OCPN27682_n25414),
	.A(n25414));
   INVx2_ASAP7_75t_L FE_OCPC8013_sa12_4 (.Y(FE_OCPN29494_sa12_4),
	.A(FE_OCPN29491_sa12_4));
   INVx2_ASAP7_75t_L FE_OCPC8012_sa12_4 (.Y(FE_OCPN29493_sa12_4),
	.A(FE_OCPN29491_sa12_4));
   INVx2_ASAP7_75t_SL FE_OCPC8011_sa12_4 (.Y(FE_OCPN29492_sa12_4),
	.A(FE_OCPN29491_sa12_4));
   INVx2_ASAP7_75t_SL FE_OCPC8010_sa12_4 (.Y(FE_OCPN29491_sa12_4),
	.A(sa12_4_));
   BUFx2_ASAP7_75t_SL FE_OCPC8009_sa12_4 (.Y(FE_OCPN29453_sa12_4),
	.A(sa12_4_));
   BUFx2_ASAP7_75t_L FE_OCPC8007_n17001 (.Y(FE_OCPN29490_n17001),
	.A(FE_OFN28583_n17001));
   INVx1_ASAP7_75t_L FE_OCPC8006_n17001 (.Y(FE_OFN28583_n17001),
	.A(n17001));
   INVx1_ASAP7_75t_SL FE_OCPC8005_sa10_1 (.Y(FE_OFN29042_n),
	.A(FE_OCPN28053_sa10_1));
   BUFx6f_ASAP7_75t_SL FE_OCPC8004_sa10_1 (.Y(FE_OCPN28053_sa10_1),
	.A(sa10_1_));
   INVx1_ASAP7_75t_L FE_OCPC8003_n26579 (.Y(n26580),
	.A(FE_OFN29029_n26579));
   INVx2_ASAP7_75t_SL FE_OCPC8002_n26579 (.Y(FE_OFN29029_n26579),
	.A(n26579));
   INVx2_ASAP7_75t_SL FE_OCPC8001_sa11_1 (.Y(FE_OCPN27241_sa11_1),
	.A(FE_OCPN27242_sa11_1));
   BUFx6f_ASAP7_75t_SL FE_OCPC8000_sa11_1 (.Y(FE_OCPN27242_sa11_1),
	.A(sa11_1_));
   INVx2_ASAP7_75t_SL FE_OCPC7999_sa23_3 (.Y(FE_OCPN29489_sa23_3),
	.A(FE_OFN27128_sa23_3));
   INVx2_ASAP7_75t_SL FE_OCPC7998_sa23_3 (.Y(FE_OFN27126_sa23_3),
	.A(FE_OFN27128_sa23_3));
   BUFx2_ASAP7_75t_SL FE_OCPC7996_sa23_3 (.Y(FE_OFN27127_sa23_3),
	.A(FE_OFN27128_sa23_3));
   INVx2_ASAP7_75t_SL FE_OCPC7995_sa23_3 (.Y(FE_OFN27128_sa23_3),
	.A(sa23_3_));
   BUFx3_ASAP7_75t_L FE_OCPC7994_n18640 (.Y(FE_OCPN29292_n18640),
	.A(n18640));
   BUFx3_ASAP7_75t_SL FE_OCPC7993_FE_OFN25883_n22945 (.Y(FE_OCPN29488_FE_OFN25883_n22945),
	.A(FE_OFN25883_n22945));
   BUFx2_ASAP7_75t_SL FE_OCPC7992_FE_OFN25883_n22945 (.Y(FE_OCPN27954_n22945),
	.A(FE_OFN25883_n22945));
   BUFx2_ASAP7_75t_SL FE_OCPC7990_n26712 (.Y(FE_OCPN27922_n26712),
	.A(n26712));
   INVx1_ASAP7_75t_L FE_OCPC7989_sa01_4 (.Y(FE_OCPN27712_sa01_4),
	.A(sa01_4_));
   BUFx6f_ASAP7_75t_SL FE_OCPC7988_sa01_4 (.Y(n17326),
	.A(sa01_4_));
   BUFx2_ASAP7_75t_SL FE_OCPC7986_n22414 (.Y(FE_OCPN5188_n22414),
	.A(n22414));
   BUFx3_ASAP7_75t_SL FE_OCPC7984_n27157 (.Y(FE_OCPN28122_n27157),
	.A(n27157));
   BUFx2_ASAP7_75t_SL FE_OCPC7983_FE_OFN28694_sa33_4 (.Y(FE_OCPN29487_FE_OFN28694_sa33_4),
	.A(FE_OFN28694_sa33_4));
   INVx2_ASAP7_75t_SL FE_OCPC7981_FE_OFN28694_sa33_4 (.Y(FE_OCPN27544_sa33_4),
	.A(FE_OFN28694_sa33_4));
   INVx4_ASAP7_75t_SL FE_OCPC7980_FE_OFN28689_sa03_5 (.Y(n17992),
	.A(FE_OFN28689_sa03_5));
   INVx1_ASAP7_75t_L FE_OCPC7979_sa12_3 (.Y(FE_OCPN29486_sa12_3),
	.A(FE_OCPN28135_sa12_3));
   INVx3_ASAP7_75t_SL FE_OCPC7978_sa12_3 (.Y(FE_OCPN29485_sa12_3),
	.A(FE_OCPN28135_sa12_3));
   INVx1_ASAP7_75t_L FE_OCPC7977_sa12_3 (.Y(FE_OCPN29484_sa12_3),
	.A(FE_OCPN28135_sa12_3));
   INVx1_ASAP7_75t_SL FE_OCPC7976_sa12_3 (.Y(n19538),
	.A(FE_OCPN28135_sa12_3));
   INVx2_ASAP7_75t_SL FE_OCPC7975_sa12_3 (.Y(FE_OCPN28135_sa12_3),
	.A(sa12_3_));
   BUFx3_ASAP7_75t_SL FE_OCPC7972_n20514 (.Y(FE_OCPN27902_n20514),
	.A(n20514));
   INVx1_ASAP7_75t_SL FE_OCPC7971_n16222 (.Y(n16223),
	.A(n16222));
   BUFx3_ASAP7_75t_SL FE_OCPC7970_sa32_5 (.Y(FE_OCPN27499_FE_OFN16151_sa32_5),
	.A(sa32_5_));
   INVx1_ASAP7_75t_L FE_OCPC7969_FE_OFN26014_sa31_3 (.Y(FE_OCPN29483_FE_OFN26014_sa31_3),
	.A(FE_OFN26014_sa31_3));
   INVx3_ASAP7_75t_SL FE_OCPC7968_FE_OFN26014_sa31_3 (.Y(FE_OCPN29482_FE_OFN26014_sa31_3),
	.A(FE_OFN26014_sa31_3));
   INVx3_ASAP7_75t_SL FE_OCPC7966_FE_OFN26014_sa31_3 (.Y(n16493),
	.A(FE_OFN26014_sa31_3));
   INVx2_ASAP7_75t_L FE_OCPC7965_FE_OFN26014_sa31_3 (.Y(FE_OFN28840_n),
	.A(FE_OFN26014_sa31_3));
   INVxp67_ASAP7_75t_SL FE_OCPC7964_n25799 (.Y(n25798),
	.A(n25799));
   BUFx2_ASAP7_75t_L FE_OCPC7963_sa31_2 (.Y(FE_OFN16415_sa31_2),
	.A(FE_OFN28516_FE_OFN27192_sa31_2));
   BUFx4f_ASAP7_75t_SL FE_OCPC7962_sa31_2 (.Y(FE_OFN28753_sa31_2),
	.A(sa31_2_));
   BUFx3_ASAP7_75t_SL FE_OCPC7961_sa31_2 (.Y(FE_OFN28516_FE_OFN27192_sa31_2),
	.A(sa31_2_));
   BUFx3_ASAP7_75t_SL FE_OCPC7960_n26537 (.Y(FE_OCPN29481_n26537),
	.A(n26537));
   INVxp67_ASAP7_75t_L FE_OCPC7958_n24936 (.Y(n24935),
	.A(n24936));
   INVx1_ASAP7_75t_SL FE_OCPC7957_n20913 (.Y(FE_OCPN29480_n20913),
	.A(FE_OFN25889_n20913));
   BUFx2_ASAP7_75t_SL FE_OCPC7955_n20913 (.Y(FE_OFN25889_n20913),
	.A(n20913));
   INVx3_ASAP7_75t_SL FE_OCPC7954_n23306 (.Y(FE_OCPN29478_n23306),
	.A(FE_OCPN27720_n23306));
   INVx2_ASAP7_75t_SL FE_OCPC7952_n23306 (.Y(FE_OCPN27719_n23306),
	.A(FE_OCPN27720_n23306));
   INVx2_ASAP7_75t_SL FE_OCPC7951_n23306 (.Y(FE_OCPN27720_n23306),
	.A(n23306));
   INVx1_ASAP7_75t_L FE_OCPC7950_sa12_5 (.Y(FE_OCPN29477_sa12_5),
	.A(FE_OFN28947_sa12_5));
   INVx1_ASAP7_75t_SL FE_OCPC7949_sa12_5 (.Y(FE_OCPN29476_sa12_5),
	.A(FE_OFN28947_sa12_5));
   BUFx3_ASAP7_75t_SL FE_OCPC7948_sa12_5 (.Y(FE_OFN73_sa12_5),
	.A(sa12_5_));
   INVx1_ASAP7_75t_SL FE_OCPC7947_sa12_5 (.Y(FE_OFN28676_sa12_5),
	.A(sa12_5_));
   INVx1_ASAP7_75t_SL FE_OCPC7946_sa12_5 (.Y(FE_OFN28947_sa12_5),
	.A(sa12_5_));
   HB1xp67_ASAP7_75t_SL FE_OCPC7945_sa02_4 (.Y(FE_OFN27202_n),
	.A(n17760));
   INVx2_ASAP7_75t_L FE_OCPC7944_sa02_4 (.Y(FE_OFN26077_n),
	.A(FE_OCPN27740_sa02_4));
   BUFx3_ASAP7_75t_SL FE_OCPC7943_sa02_4 (.Y(n17760),
	.A(sa02_4_));
   INVx1_ASAP7_75t_SL FE_OCPC7942_sa02_4 (.Y(FE_OCPN27740_sa02_4),
	.A(sa02_4_));
   INVx1_ASAP7_75t_L FE_OCPC7941_sa11_5 (.Y(n17451),
	.A(FE_OCPN27625_sa11_5));
   BUFx6f_ASAP7_75t_SL FE_OCPC7940_sa11_5 (.Y(FE_OCPN27625_sa11_5),
	.A(sa11_5_));
   INVx1_ASAP7_75t_L FE_OCPC7938_n25054 (.Y(FE_OCPN29475_n25054),
	.A(n26456));
   INVx2_ASAP7_75t_SL FE_OCPC7937_n25054 (.Y(n26456),
	.A(n25054));
   INVx2_ASAP7_75t_SL FE_OCPC7935_n25696 (.Y(n25697),
	.A(n25696));
   INVx2_ASAP7_75t_SL FE_OCPC7934_n19119 (.Y(FE_OCPN29474_n19119),
	.A(FE_OFN16130_n19119));
   INVx3_ASAP7_75t_SL FE_OCPC7933_n19119 (.Y(FE_OFN28835_n),
	.A(FE_OFN16130_n19119));
   INVx1_ASAP7_75t_SL FE_OCPC7932_n19119 (.Y(FE_OFN16130_n19119),
	.A(n19119));
   INVxp67_ASAP7_75t_L FE_OCPC7931_n26579 (.Y(FE_OCPN29473_n26579),
	.A(n26580));
   BUFx2_ASAP7_75t_L FE_OCPC7927_n24175 (.Y(FE_OCPN29471_n24175),
	.A(FE_OCPN29470_n24175));
   INVx1_ASAP7_75t_SL FE_OCPC7926_n24175 (.Y(FE_OCPN29470_n24175),
	.A(n24175));
   INVx3_ASAP7_75t_SL FE_OCPC7924_n17747 (.Y(FE_OCPN29469_n17747),
	.A(FE_OCPN27838_n17747));
   BUFx2_ASAP7_75t_SL FE_OCPC7923_n17747 (.Y(FE_OFN29144_n17747),
	.A(FE_OCPN27838_n17747));
   INVx2_ASAP7_75t_SL FE_OCPC7922_n17747 (.Y(FE_OCPN27838_n17747),
	.A(n17747));
   INVx2_ASAP7_75t_SL FE_OCPC7921_n15919 (.Y(FE_OCPN29468_n15919),
	.A(n15918));
   INVx2_ASAP7_75t_SL FE_OCPC7919_n15919 (.Y(n15918),
	.A(n15919));
   INVx2_ASAP7_75t_L FE_OCPC7918_n25102 (.Y(FE_OCPN29467_n25102),
	.A(n21605));
   INVx2_ASAP7_75t_SL FE_OCPC7916_n25102 (.Y(FE_OCPN27829_n25102),
	.A(n25102));
   INVx2_ASAP7_75t_L FE_OCPC7915_n25102 (.Y(n21605),
	.A(n25102));
   BUFx3_ASAP7_75t_SL FE_OCPC7913_n16989 (.Y(FE_OFN28738_n16989),
	.A(n16989));
   BUFx3_ASAP7_75t_SL FE_OCPC7911_n16230 (.Y(FE_OFN16287_n16230),
	.A(n16230));
   INVx1_ASAP7_75t_L FE_OCPC7910_n16230 (.Y(FE_OFN25975_n16217),
	.A(n16230));
   INVxp67_ASAP7_75t_SL FE_OCPC7909_n16751 (.Y(FE_OCPN29450_sa21_0),
	.A(n16751));
   INVx1_ASAP7_75t_SL FE_OCPC7907_n16751 (.Y(FE_OCPN29418_n),
	.A(n16751));
   INVxp67_ASAP7_75t_L FE_OCPC7906_n19149 (.Y(FE_OCPN29464_n),
	.A(n19149));
   INVx2_ASAP7_75t_SL FE_OCPC7905_n19149 (.Y(FE_OCPN29463_n),
	.A(FE_OCPN27337_n19149));
   INVx2_ASAP7_75t_SL FE_OCPC7904_n19149 (.Y(FE_OFN29249_n),
	.A(FE_OCPN27337_n19149));
   INVx1_ASAP7_75t_SL FE_OCPC7903_n19149 (.Y(n19149),
	.A(FE_OCPN27337_n19149));
   BUFx6f_ASAP7_75t_L FE_OCPC7901_n15233 (.Y(FE_OFN25893_n15214),
	.A(n15233));
   BUFx2_ASAP7_75t_SL FE_OCPC7900_sa01_5 (.Y(FE_OFN28736_FE_OCPN28216_sa01_5),
	.A(FE_OCPN28217_sa01_5));
   INVxp67_ASAP7_75t_L FE_OCPC7898_n22197 (.Y(FE_OCPN29461_n22197),
	.A(FE_OFN26648_n22197));
   INVx3_ASAP7_75t_L FE_OCPC7897_n22197 (.Y(FE_OFN26648_n22197),
	.A(n22197));
   INVx1_ASAP7_75t_SL FE_OCPC7896_n22499 (.Y(FE_OFN26031_n22499),
	.A(n22499));
   BUFx2_ASAP7_75t_R FE_OCPC7895_n26227 (.Y(FE_OCPN29460_n26227),
	.A(FE_OCPN27678_n26227));
   BUFx3_ASAP7_75t_SL FE_OCPC7894_n26227 (.Y(FE_OCPN27678_n26227),
	.A(n26227));
   BUFx3_ASAP7_75t_SL FE_OCPC7893_FE_OFN16151_sa32_5 (.Y(FE_OCPN29459_n),
	.A(FE_OCPN27499_FE_OFN16151_sa32_5));
   INVxp67_ASAP7_75t_SL FE_OCPC7892_FE_OFN16151_sa32_5 (.Y(FE_OFN28707_n),
	.A(FE_OCPN27499_FE_OFN16151_sa32_5));
   BUFx2_ASAP7_75t_SL FE_OCPC7890_n26982 (.Y(FE_OCPN27354_n26982),
	.A(n26982));
   HB1xp67_ASAP7_75t_L FE_OCPC7889_n26442 (.Y(FE_OCPN29458_n26442),
	.A(n26442));
   INVxp67_ASAP7_75t_L FE_OCPC7887_n25722 (.Y(FE_OCPN29457_n25722),
	.A(n25722));
   INVxp67_ASAP7_75t_L FE_OCPC7883_n18671 (.Y(FE_OCPN29455_n18671),
	.A(FE_OFN27072_n18671));
   INVxp67_ASAP7_75t_SL FE_OCPC7882_n18671 (.Y(FE_OCPN29454_n18671),
	.A(FE_OFN27072_n18671));
   INVx4_ASAP7_75t_SL FE_OCPC7881_n18671 (.Y(FE_OFN27072_n18671),
	.A(n18671));
   BUFx2_ASAP7_75t_SL FE_OCPC7880_n24847 (.Y(FE_OCPN27446_n24847),
	.A(n24847));
   INVx2_ASAP7_75t_SL FE_OCPC7879_sa33_5 (.Y(FE_OFN26628_n),
	.A(FE_OFN28679_sa33_5));
   BUFx6f_ASAP7_75t_SL FE_OCPC7878_sa33_5 (.Y(FE_OFN28679_sa33_5),
	.A(sa33_5_));
   BUFx6f_ASAP7_75t_SL FE_OCPC7877_sa10_2 (.Y(FE_OFN28749_n),
	.A(sa10_2_));
   INVxp67_ASAP7_75t_L FE_OCPC7876_n25599 (.Y(n24478),
	.A(n25599));
   BUFx2_ASAP7_75t_SL FE_OCPC7875_n17001 (.Y(n19376),
	.A(n17001));
   BUFx2_ASAP7_75t_SL FE_OCPC7873_FE_OFN28689_sa03_5 (.Y(FE_OFN29179_n),
	.A(FE_OFN28689_sa03_5));
   INVxp67_ASAP7_75t_SL FE_OCPC7870_sa12_4 (.Y(n23220),
	.A(FE_OCPN29492_sa12_4));
   BUFx6f_ASAP7_75t_SL FE_OCPC7866_sa02_2 (.Y(FE_OFN16234_sa02_2),
	.A(sa02_2_));
   INVxp67_ASAP7_75t_SL FE_OCPC7864_n16240 (.Y(FE_OCPN29452_n16240),
	.A(n16240));
   HB1xp67_ASAP7_75t_L FE_OCPC7862_n (.Y(FE_OCPN29451_n),
	.A(FE_OCPN27726_n));
   BUFx2_ASAP7_75t_SL FE_OCPC7861_n (.Y(FE_OCPN27393_sa03_0),
	.A(FE_OCPN27726_n));
   INVx2_ASAP7_75t_SL FE_OCPC7860_n (.Y(FE_OCPN27726_n),
	.A(FE_OCPN27800_n));
   BUFx3_ASAP7_75t_SL FE_OCPC7859_n (.Y(FE_OFN29199_FE_OCPN27726_n),
	.A(FE_OCPN27800_n));
   BUFx3_ASAP7_75t_SL FE_OCPC7858_n24099 (.Y(FE_OCPN29376_n24099),
	.A(n24099));
   INVx2_ASAP7_75t_SL FE_OCPC7854_sa21_0 (.Y(n16751),
	.A(sa21_0_));
   INVx2_ASAP7_75t_SL FE_OCPC7853_n17441 (.Y(n24310),
	.A(n17441));
   BUFx3_ASAP7_75t_L FE_OCPC7852_n17521 (.Y(FE_OCPN29449_n17521),
	.A(n17521));
   INVx3_ASAP7_75t_SL FE_OCPC7850_sa11_0 (.Y(FE_OFN28507_sa11_0),
	.A(FE_OFN25879_sa11_0));
   INVx2_ASAP7_75t_SL FE_OCPC7849_sa11_0 (.Y(n21844),
	.A(FE_OFN25879_sa11_0));
   INVx2_ASAP7_75t_SL FE_OCPC7848_sa11_0 (.Y(FE_OFN25879_sa11_0),
	.A(sa11_0_));
   INVx4_ASAP7_75t_SL FE_OCPC7847_sa30_4 (.Y(FE_OFN28901_sa30_4),
	.A(FE_OFN29067_n));
   BUFx3_ASAP7_75t_SL FE_OCPC7846_sa30_4 (.Y(FE_OFN16333_sa30_4),
	.A(FE_OFN29067_n));
   INVx2_ASAP7_75t_SL FE_OCPC7845_sa30_4 (.Y(FE_OFN29067_n),
	.A(sa30_4_));
   INVx1_ASAP7_75t_R FE_OCPC7843_n27189 (.Y(FE_OCPN29448_n27189),
	.A(n27188));
   INVxp67_ASAP7_75t_SL FE_OCPC7842_n27189 (.Y(FE_OCPN29447_n27189),
	.A(FE_OCPN27456_n27189));
   INVx1_ASAP7_75t_R FE_OCPC7841_n27189 (.Y(n27188),
	.A(FE_OCPN27456_n27189));
   INVx2_ASAP7_75t_SL FE_OCPC7840_n27189 (.Y(FE_OCPN27456_n27189),
	.A(n27189));
   INVx1_ASAP7_75t_SL FE_OCPC7839_n26789 (.Y(FE_OFN155_n26788),
	.A(FE_OCPN28311_n26789));
   INVx1_ASAP7_75t_L FE_OCPC7838_n26789 (.Y(FE_OCPN28311_n26789),
	.A(n26789));
   BUFx3_ASAP7_75t_SL FE_OCPC7837_n27203 (.Y(FE_OCPN29445_n27203),
	.A(n27203));
   BUFx4f_ASAP7_75t_SL FE_OCPC7836_n17115 (.Y(FE_OCPN29446_n17115),
	.A(n17115));
   INVxp67_ASAP7_75t_L FE_OCPC7834_n25507 (.Y(FE_OCPN29444_n25507),
	.A(FE_OCPN29443_n25507));
   INVx2_ASAP7_75t_SL FE_OCPC7833_n25507 (.Y(FE_OCPN29443_n25507),
	.A(FE_OCPN8218_n25507));
   BUFx2_ASAP7_75t_L FE_OCPC7831_n17261 (.Y(FE_OFN28958_n17261),
	.A(n19594));
   INVx1_ASAP7_75t_SL FE_OCPC7830_n17261 (.Y(n19594),
	.A(n17261));
   INVxp67_ASAP7_75t_SL FE_OCPC7829_n26369 (.Y(n26368),
	.A(FE_OCPN27357_n26369));
   HB1xp67_ASAP7_75t_SL FE_OCPC7828_n26369 (.Y(FE_OCPN27357_n26369),
	.A(n26369));
   BUFx2_ASAP7_75t_SL FE_OCPC7827_n458 (.Y(FE_OCPN29442_n458),
	.A(n458));
   BUFx2_ASAP7_75t_L FE_OCPC7826_sa23_4 (.Y(FE_OCPN29441_sa23_4),
	.A(FE_OCPN27803_sa23_4));
   INVxp67_ASAP7_75t_SL FE_OCPC7825_sa23_4 (.Y(FE_OCPN29440_sa23_4),
	.A(FE_OCPN27577_sa23_4));
   BUFx4f_ASAP7_75t_SL FE_OCPC7824_sa23_4 (.Y(FE_OCPN27803_sa23_4),
	.A(sa23_4_));
   INVx1_ASAP7_75t_SL FE_OCPC7823_sa23_4 (.Y(FE_OCPN27577_sa23_4),
	.A(sa23_4_));
   BUFx2_ASAP7_75t_SL FE_OCPC7821_n17447 (.Y(FE_OCPN27562_n17447),
	.A(n17447));
   BUFx2_ASAP7_75t_SL FE_OCPC7820_n23255 (.Y(FE_OCPN27848_n23255),
	.A(n23255));
   INVx2_ASAP7_75t_SL FE_OCPC7819_n18443 (.Y(n16701),
	.A(n18443));
   BUFx2_ASAP7_75t_SL FE_OCPC7818_sa33_2 (.Y(FE_OCPN29438_sa33_2),
	.A(FE_OFN26062_n16435));
   INVx3_ASAP7_75t_SL FE_OCPC7817_sa33_2 (.Y(FE_OCPN29391_FE_OFN29162_sa33_2),
	.A(FE_OFN26062_n16435));
   INVxp67_ASAP7_75t_L FE_OCPC7816_sa33_2 (.Y(FE_OFN29162_sa33_2),
	.A(FE_OFN26062_n16435));
   INVx1_ASAP7_75t_SL FE_OCPC7815_sa33_2 (.Y(FE_OFN29163_sa33_2),
	.A(FE_OFN26062_n16435));
   INVx4_ASAP7_75t_SL FE_OCPC7814_sa33_2 (.Y(FE_OFN26062_n16435),
	.A(sa33_2_));
   BUFx2_ASAP7_75t_L FE_OCPC7813_sa33_2 (.Y(FE_OFN26078_sa33_2),
	.A(sa33_2_));
   BUFx2_ASAP7_75t_SL FE_OCPC7812_n16143 (.Y(FE_OFN25904_n16143),
	.A(n16143));
   INVxp67_ASAP7_75t_L FE_OCPC7811_n16143 (.Y(FE_OFN26154_n16132),
	.A(n16143));
   BUFx3_ASAP7_75t_SL FE_OCPC7810_n14008 (.Y(n14007),
	.A(n14008));
   INVx1_ASAP7_75t_SL FE_OCPC7809_n14008 (.Y(FE_OFN16254_n14008),
	.A(n14008));
   INVx1_ASAP7_75t_SL FE_OCPC7808_n25935 (.Y(FE_OCPN29267_n25935),
	.A(n25935));
   HB1xp67_ASAP7_75t_L FE_OCPC7807_n25422 (.Y(FE_OCPN7637_n25422),
	.A(n25422));
   INVx1_ASAP7_75t_SL FE_OCPC7806_n25864 (.Y(FE_OCPN29437_n25864),
	.A(n25864));
   HB1xp67_ASAP7_75t_L FE_OCPC7805_n25864 (.Y(n25997),
	.A(n25864));
   INVx2_ASAP7_75t_R FE_OCPC7804_n22080 (.Y(FE_OCPN29436_n22080),
	.A(FE_OFN16234_sa02_2));
   HB1xp67_ASAP7_75t_L FE_OCPC7803_n22080 (.Y(FE_OFN26159_n22080),
	.A(FE_OFN16234_sa02_2));
   BUFx2_ASAP7_75t_SL FE_OCPC7800_n17445 (.Y(FE_OCPN29435_n17445),
	.A(n17445));
   BUFx2_ASAP7_75t_SL FE_OCPC7798_n408 (.Y(FE_OCPN29434_n408),
	.A(n408));
   INVxp67_ASAP7_75t_SL FE_OCPC7797_n25040 (.Y(FE_OCPN29433_n25040),
	.A(n25041));
   BUFx2_ASAP7_75t_SL FE_OCPC7796_n25040 (.Y(n25041),
	.A(n25040));
   INVxp67_ASAP7_75t_L FE_OCPC7795_n25040 (.Y(FE_OFN29015_n25040),
	.A(n25040));
   HB1xp67_ASAP7_75t_L FE_OCPC7794_sa30_3 (.Y(FE_OCPN29432_sa30_3),
	.A(FE_OCPN29431_sa30_3));
   INVx5_ASAP7_75t_SL FE_OCPC7793_sa30_3 (.Y(FE_OCPN29431_sa30_3),
	.A(FE_OFN25958_sa30_3));
   INVx2_ASAP7_75t_SL FE_OCPC7791_sa30_3 (.Y(FE_OFN25958_sa30_3),
	.A(sa30_3_));
   BUFx2_ASAP7_75t_SL FE_OCPC7790_FE_OFN31_sa20_0 (.Y(FE_OCPN29430_FE_OFN31_sa20_0),
	.A(n18522));
   INVx2_ASAP7_75t_SL FE_OCPC7789_FE_OFN31_sa20_0 (.Y(n18522),
	.A(FE_OFN31_sa20_0));
   INVx4_ASAP7_75t_SL FE_OCPC7788_FE_OFN31_sa20_0 (.Y(FE_OCPN28223_FE_OFN27219_n18522),
	.A(FE_OFN31_sa20_0));
   INVx1_ASAP7_75t_SL FE_OCPC7787_FE_OFN31_sa20_0 (.Y(FE_OFN29223_sa20_0),
	.A(FE_OFN31_sa20_0));
   BUFx4f_ASAP7_75t_SL FE_OCPC7786_FE_OFN16141_sa01_3 (.Y(FE_OCPN29429_FE_OFN16141_sa01_3),
	.A(FE_OFN16141_sa01_3));
   BUFx6f_ASAP7_75t_L FE_OCPC7785_FE_OFN27131_w3_29 (.Y(FE_OCPN29428_FE_OFN27131_w3_29),
	.A(FE_OFN27131_w3_29));
   INVxp67_ASAP7_75t_L FE_OCPC7784_FE_OFN27131_w3_29 (.Y(FE_OFN28663_n),
	.A(FE_OFN27131_w3_29));
   INVx2_ASAP7_75t_SL FE_OCPC7783_FE_OFN27131_w3_29 (.Y(FE_OFN28452_w3_29),
	.A(FE_OFN27131_w3_29));
   BUFx3_ASAP7_75t_SL FE_OCPC7782_w3_15 (.Y(FE_OCPN29427_w3_15),
	.A(FE_OFN27200_n));
   BUFx4f_ASAP7_75t_SL FE_OCPC7781_w3_15 (.Y(FE_OFN27200_n),
	.A(w3_15_));
   BUFx2_ASAP7_75t_SL FE_OCPC7780_FE_OFN16444_sa13_1 (.Y(FE_OCPN29426_FE_OFN16444_sa13_1),
	.A(FE_OFN16444_sa13_1));
   INVxp67_ASAP7_75t_SL FE_OCPC7778_sa11_5 (.Y(FE_OFN26005_n17451),
	.A(FE_OCPN27625_sa11_5));
   HB1xp67_ASAP7_75t_L FE_OCPC7776_n24172 (.Y(FE_OCPN29425_n24172),
	.A(n24172));
   HB1xp67_ASAP7_75t_L FE_OCPC7775_FE_OFN26039_sa10_2 (.Y(FE_OCPN29424_FE_OFN26039_sa10_2),
	.A(FE_OFN26039_sa10_2));
   HB1xp67_ASAP7_75t_SL FE_OCPC7774_n26970 (.Y(FE_OCPN29423_n26970),
	.A(n26970));
   BUFx2_ASAP7_75t_SL FE_OCPC7773_n23397 (.Y(FE_OCPN29422_n23397),
	.A(n23397));
   BUFx2_ASAP7_75t_R FE_OCPC7772_FE_OFN16128_sa32_2 (.Y(FE_OCPN29421_FE_OFN16128_sa32_2),
	.A(FE_OCPN29420_FE_OFN16128_sa32_2));
   BUFx3_ASAP7_75t_SL FE_OCPC7771_FE_OFN16128_sa32_2 (.Y(FE_OCPN29420_FE_OFN16128_sa32_2),
	.A(FE_OFN28892_n));
   HB1xp67_ASAP7_75t_L FE_OCPC7770_FE_OFN16128_sa32_2 (.Y(FE_OCPN29419_FE_OFN16128_sa32_2),
	.A(FE_OFN28892_n));
   BUFx2_ASAP7_75t_SL FE_OCPC7769_FE_OFN16128_sa32_2 (.Y(FE_OFN28893_n),
	.A(FE_OFN28892_n));
   INVx3_ASAP7_75t_L FE_OCPC7768_FE_OFN16128_sa32_2 (.Y(n17564),
	.A(FE_OFN28892_n));
   INVx5_ASAP7_75t_SL FE_OCPC7767_FE_OFN16128_sa32_2 (.Y(FE_OFN28892_n),
	.A(FE_OFN16128_sa32_2));
   INVx2_ASAP7_75t_L FE_OCPC7763_sa21_0 (.Y(FE_OFN28903_sa21_0),
	.A(n16751));
   BUFx2_ASAP7_75t_SL FE_OCPC7761_n455 (.Y(FE_OCPN29417_n455),
	.A(n455));
   BUFx2_ASAP7_75t_L FE_OCPC7760_n22516 (.Y(FE_OCPN29416_n22516),
	.A(n22516));
   HB1xp67_ASAP7_75t_SL FE_OCPC7759_n17237 (.Y(FE_OCPN29415_n17237),
	.A(n17237));
   BUFx4f_ASAP7_75t_SL FE_OCPC7758_FE_OFN25990_sa21_4 (.Y(FE_OCPN29414_n),
	.A(FE_OFN25989_sa21_4));
   INVx1_ASAP7_75t_R FE_OCPC7757_FE_OFN25990_sa21_4 (.Y(FE_OFN27155_sa21_4),
	.A(FE_OFN25989_sa21_4));
   INVx4_ASAP7_75t_SL FE_OCPC7756_FE_OFN25990_sa21_4 (.Y(FE_OFN25989_sa21_4),
	.A(FE_OCPN27388_FE_OFN25990_sa21_4));
   BUFx2_ASAP7_75t_SL FE_OCPC7754_FE_OFN25990_sa21_4 (.Y(FE_OCPN29307_FE_OFN25989_sa21_4),
	.A(FE_OCPN27388_FE_OFN25990_sa21_4));
   INVx1_ASAP7_75t_SL FE_OCPC7753_n26955 (.Y(n26954),
	.A(n26955));
   BUFx2_ASAP7_75t_SL FE_OCPC7752_n26955 (.Y(FE_OCPN28119_n26955),
	.A(n26955));
   BUFx2_ASAP7_75t_SL FE_OCPC7751_sa30_5 (.Y(FE_OCPN29413_sa30_5),
	.A(n17618));
   INVx1_ASAP7_75t_SL FE_OCPC7750_sa30_5 (.Y(FE_OCPN29412_sa30_5),
	.A(sa30_5_));
   BUFx6f_ASAP7_75t_SL FE_OCPC7749_sa30_5 (.Y(n17618),
	.A(sa30_5_));
   BUFx3_ASAP7_75t_SL FE_OCPC7747_sa12_0 (.Y(FE_OFN28476_sa12_0),
	.A(FE_OFN29225_sa12_0));
   BUFx3_ASAP7_75t_SL FE_OCPC7746_sa12_0 (.Y(FE_OFN29225_sa12_0),
	.A(sa12_0_));
   BUFx2_ASAP7_75t_SL FE_OCPC7745_sa00_5 (.Y(FE_OCPN29411_n),
	.A(FE_OCPN27227_sa00_5));
   INVx1_ASAP7_75t_L FE_OCPC7743_n22461 (.Y(FE_OCPN29409_n22461),
	.A(n22461));
   INVx1_ASAP7_75t_SL FE_OCPC7742_n22461 (.Y(FE_OCPN29408_n22461),
	.A(n22461));
   INVx1_ASAP7_75t_L FE_OCPC7741_n22461 (.Y(FE_OCPN29388_n22461),
	.A(n22461));
   BUFx3_ASAP7_75t_SL FE_OCPC7740_n22461 (.Y(FE_OCPN29320_n22461),
	.A(n22461));
   OAI222xp33_ASAP7_75t_SL FE_RC_914_0 (.Y(n26441),
	.A1(n24580),
	.A2(n24800),
	.B1(n24581),
	.B2(n24800),
	.C1(n24579),
	.C2(n24800));
   INVx1_ASAP7_75t_L FE_RC_913_0 (.Y(n20985),
	.A(FE_RN_266_0));
   OR3x1_ASAP7_75t_L FE_RC_912_0 (.Y(FE_RN_266_0),
	.A(FE_OCPN29341_FE_OFN29148_n),
	.B(FE_OFN28800_n22526),
	.C(FE_OFN28812_FE_OCPN27261_sa02_0));
   HB1xp67_ASAP7_75t_L FE_OCPC7735_FE_OFN142_sa10_0 (.Y(FE_OCPN29407_FE_OFN142_sa10_0),
	.A(FE_OFN142_sa10_0));
   AND2x2_ASAP7_75t_R FE_RC_911_0 (.Y(FE_RN_265_0),
	.A(n22487),
	.B(n22495));
   NAND2x1p5_ASAP7_75t_SL FE_RC_910_0 (.Y(n17459),
	.A(FE_RN_265_0),
	.B(n26071));
   AOI31xp33_ASAP7_75t_SL FE_RC_909_0 (.Y(n23732),
	.A1(n23729),
	.A2(n23730),
	.A3(n23731),
	.B(n25641));
   INVx1_ASAP7_75t_L FE_RC_908_0 (.Y(n19774),
	.A(FE_RN_264_0));
   OR3x1_ASAP7_75t_L FE_RC_907_0 (.Y(FE_RN_264_0),
	.A(n16533),
	.B(FE_OCPN29498_n16581),
	.C(FE_OFN26160_sa10_4));
   BUFx2_ASAP7_75t_SL FE_OCPC7734_n26145 (.Y(FE_OCPN7609_n26145),
	.A(n26145));
   AOI31xp33_ASAP7_75t_SL FE_RC_906_0 (.Y(n19495),
	.A1(n19494),
	.A2(n19493),
	.A3(n21292),
	.B(n25420));
   AOI21xp5_ASAP7_75t_L FE_RC_905_0 (.Y(n19595),
	.A1(n17254),
	.A2(FE_PSN8282_n21154),
	.B(FE_OFN26644_n19599));
   INVx1_ASAP7_75t_SL FE_RC_904_0 (.Y(n16653),
	.A(FE_RN_263_0));
   OR3x1_ASAP7_75t_L FE_RC_903_0 (.Y(FE_RN_263_0),
	.A(n16581),
	.B(n17191),
	.C(FE_OFN26161_sa10_4));
   BUFx3_ASAP7_75t_SL FE_OCPC7733_n15899 (.Y(FE_OCPN28327_n15899),
	.A(n15899));
   INVx1_ASAP7_75t_SL FE_OCPC7732_n15899 (.Y(n15898),
	.A(n15899));
   BUFx2_ASAP7_75t_SL FE_OCPC7731_n26093 (.Y(FE_OCPN27941_n),
	.A(n26093));
   BUFx6f_ASAP7_75t_SL FE_OCPC7730_n18710 (.Y(FE_OCPN29406_n18710),
	.A(n18710));
   OAI21xp5_ASAP7_75t_SL FE_RC_902_0 (.Y(n26921),
	.A1(n26917),
	.A2(FE_RN_250_0),
	.B(n26916));
   OAI21x1_ASAP7_75t_SL FE_RC_901_0 (.Y(n26339),
	.A1(FE_RN_107_0),
	.A2(n25365),
	.B(n25364));
   AOI31xp33_ASAP7_75t_SL FE_RC_900_0 (.Y(n24706),
	.A1(n24704),
	.A2(FE_RN_2_0),
	.A3(n26874),
	.B(n26889));
   BUFx2_ASAP7_75t_SL FE_OCPC7729_FE_OFN27148_sa32_3 (.Y(FE_OCPN29405_FE_OFN27148_sa32_3),
	.A(FE_OFN27148_sa32_3));
   HB1xp67_ASAP7_75t_L FE_OCPC7728_FE_OFN27148_sa32_3 (.Y(FE_OCPN29404_FE_OFN27148_sa32_3),
	.A(FE_OFN27148_sa32_3));
   INVx3_ASAP7_75t_SL FE_OCPC7723_sa31_3 (.Y(FE_OFN26014_sa31_3),
	.A(sa31_3_));
   BUFx2_ASAP7_75t_L FE_OCPC7719_sa30_3 (.Y(FE_OCPN29400_sa30_3),
	.A(FE_OCPN29431_sa30_3));
   BUFx2_ASAP7_75t_SL FE_OCPC7718_sa30_3 (.Y(FE_OCPN29399_sa30_3),
	.A(FE_OCPN29431_sa30_3));
   BUFx2_ASAP7_75t_SL FE_OCPC7717_sa30_3 (.Y(FE_OCPN29398_sa30_3),
	.A(FE_OFN25958_sa30_3));
   BUFx2_ASAP7_75t_SL FE_OCPC7711_n26502 (.Y(FE_OCPN29397_n26502),
	.A(n26502));
   BUFx2_ASAP7_75t_SL FE_OCPC7710_n19149 (.Y(FE_OCPN29396_n19149),
	.A(FE_OFN29249_n));
   AOI31xp33_ASAP7_75t_SL FE_RC_899_0 (.Y(n24270),
	.A1(n23674),
	.A2(n20017),
	.A3(n20016),
	.B(n25585));
   BUFx2_ASAP7_75t_SL FE_OCPC7708_n479 (.Y(FE_OCPN29394_n479),
	.A(n479));
   BUFx3_ASAP7_75t_SL FE_OCPC7707_n26420 (.Y(FE_OCPN7589_n26420),
	.A(n26420));
   BUFx2_ASAP7_75t_SL FE_OCPC7706_n483 (.Y(FE_OCPN29393_n483),
	.A(n483));
   BUFx3_ASAP7_75t_SL FE_OCPC7705_n26334 (.Y(FE_OCPN27430_n26334),
	.A(n26334));
   BUFx2_ASAP7_75t_SL FE_OCPC7704_n16117 (.Y(FE_OFN16405_n16117),
	.A(n16117));
   NAND3x2_ASAP7_75t_L FE_RC_898_0 (.Y(n22529),
	.A(FE_OCPN27585_sa02_1),
	.B(FE_OCPN27261_sa02_0),
	.C(FE_OFN16234_sa02_2));
   BUFx6f_ASAP7_75t_SL FE_OCPC7703_sa13_3 (.Y(FE_OFN16268_sa13_3),
	.A(sa13_3_));
   INVx1_ASAP7_75t_L FE_OCPC7702_n16078 (.Y(n16079),
	.A(n16078));
   BUFx3_ASAP7_75t_SL FE_OCPC7700_n26528 (.Y(FE_OCPN29389_n26528),
	.A(n26528));
   OAI22xp33_ASAP7_75t_L FE_RC_897_0 (.Y(n19584),
	.A1(FE_OCPN28389_n21479),
	.A2(n19139),
	.B1(FE_OCPN28021_n21445),
	.B2(n19139));
   INVx2_ASAP7_75t_L FE_OCPC7698_n26528 (.Y(FE_OCPN29390_n26528),
	.A(FE_OCPN29389_n26528));
   BUFx6f_ASAP7_75t_SL FE_OCPC7694_n17237 (.Y(FE_OCPN28270_n17237),
	.A(n17237));
   INVxp67_ASAP7_75t_SL FE_RC_896_0 (.Y(FE_RN_260_0),
	.A(n25521));
   INVxp67_ASAP7_75t_SL FE_RC_895_0 (.Y(FE_RN_261_0),
	.A(n25522));
   INVxp67_ASAP7_75t_L FE_RC_894_0 (.Y(FE_RN_262_0),
	.A(FE_RN_86_0));
   AO21x2_ASAP7_75t_SL FE_RC_893_0 (.Y(n26520),
	.A1(FE_RN_262_0),
	.A2(FE_RN_261_0),
	.B(FE_RN_260_0));
   BUFx2_ASAP7_75t_SL FE_OCPC7690_n25273 (.Y(FE_OCPN29387_n25273),
	.A(n25273));
   INVx2_ASAP7_75t_SL FE_OCPC7689_n16073 (.Y(FE_OCPN29386_n16073),
	.A(FE_OFN25929_n16073));
   BUFx3_ASAP7_75t_SL FE_OCPC7688_n16073 (.Y(FE_OFN25929_n16073),
	.A(n16073));
   BUFx2_ASAP7_75t_SL FE_OCPC7687_n26193 (.Y(FE_OCPN27583_n26193),
	.A(n26193));
   BUFx6f_ASAP7_75t_SL FE_OCPC7686_n17267 (.Y(FE_OCPN29385_n),
	.A(FE_OCPN27818_n17267));
   INVx1_ASAP7_75t_L FE_OCPC7684_n26674 (.Y(FE_OCPN29383_n26674),
	.A(n26672));
   INVx1_ASAP7_75t_R FE_OCPC7683_n26674 (.Y(FE_OCPN29382_n26674),
	.A(n26672));
   INVxp67_ASAP7_75t_SL FE_OCPC7682_n26674 (.Y(FE_OFN86_n26674),
	.A(n26674));
   INVx1_ASAP7_75t_SL FE_OCPC7681_n26674 (.Y(n26672),
	.A(n26674));
   INVx1_ASAP7_75t_SL FE_OCPC7680_n26938 (.Y(FE_OCPN27809_n26938),
	.A(n26936));
   INVx2_ASAP7_75t_SL FE_OCPC7679_n26938 (.Y(n26936),
	.A(n26938));
   BUFx2_ASAP7_75t_L FE_OCPC7678_n26215 (.Y(FE_OCPN27462_n26215),
	.A(n26215));
   BUFx2_ASAP7_75t_SL FE_OCPC7677_n26380 (.Y(FE_OCPN27321_n26380),
	.A(n26380));
   BUFx2_ASAP7_75t_L FE_OCPC7674_n26796 (.Y(FE_OCPN29381_n26796),
	.A(FE_OCPN28131_n26796));
   BUFx2_ASAP7_75t_SL FE_OCPC7673_n26796 (.Y(FE_OCPN28131_n26796),
	.A(n26796));
   BUFx3_ASAP7_75t_SL FE_OCPC7672_n26809 (.Y(FE_OCPN27379_n26809),
	.A(n26809));
   AOI22xp5_ASAP7_75t_SL FE_RC_892_0 (.Y(n16175),
	.A1(w1_19_),
	.A2(n16063),
	.B1(n25732),
	.B2(n16062));
   BUFx6f_ASAP7_75t_SL FE_OCPC7671_n26434 (.Y(FE_OCPN27525_n26434),
	.A(n26434));
   INVx4_ASAP7_75t_SL FE_OCPC7670_sa20_1 (.Y(FE_OCPN29380_sa20_1),
	.A(FE_OFN28720_sa20_1));
   BUFx2_ASAP7_75t_L FE_OCPC7669_sa20_1 (.Y(FE_OCPN29379_sa20_1),
	.A(FE_OFN28720_sa20_1));
   INVxp67_ASAP7_75t_SL FE_OCPC7668_sa20_1 (.Y(FE_OFN16385_n18525),
	.A(FE_OFN28720_sa20_1));
   INVx2_ASAP7_75t_SL FE_OCPC7667_sa20_1 (.Y(FE_OFN28720_sa20_1),
	.A(sa20_1_));
   BUFx6f_ASAP7_75t_SL FE_OCPC7666_n23266 (.Y(FE_OCPN29378_n23266),
	.A(n23266));
   BUFx2_ASAP7_75t_SL FE_OCPC7664_n26716 (.Y(FE_OCPN5022_n26716),
	.A(n26716));
   BUFx2_ASAP7_75t_SL FE_OCPC7663_n26659 (.Y(FE_OCPN27796_n26659),
	.A(n26659));
   INVx2_ASAP7_75t_SL FE_OCPC7662_n23409 (.Y(n25606),
	.A(n23409));
   AOI31xp33_ASAP7_75t_SL FE_RC_891_0 (.Y(n26267),
	.A1(n24568),
	.A2(n24566),
	.A3(n24567),
	.B(n26078));
   OAI21xp5_ASAP7_75t_SL FE_RC_890_0 (.Y(n26470),
	.A1(FE_OFN16213_ld_r),
	.A2(n26472),
	.B(n26471));
   NAND3x1_ASAP7_75t_R FE_RC_889_0 (.Y(n24422),
	.A(n22620),
	.B(n22622),
	.C(n22621));
   INVxp67_ASAP7_75t_SL FE_OCPC7661_n26910 (.Y(FE_OCPN27302_n26910),
	.A(n26910));
   INVx2_ASAP7_75t_L FE_OCPC7660_n26910 (.Y(FE_OCPN27741_n),
	.A(n26910));
   BUFx3_ASAP7_75t_SL FE_OCPC7659_n25868 (.Y(FE_OCPN27859_n25868),
	.A(n25868));
   INVx2_ASAP7_75t_SL FE_OCPC7655_FE_OFN29191_sa23_2 (.Y(FE_OCPN29374_FE_OFN29191_sa23_2),
	.A(FE_OCPN27498_sa23_2));
   BUFx3_ASAP7_75t_SL FE_OCPC7654_FE_OFN29191_sa23_2 (.Y(FE_OCPN29373_FE_OFN29191_sa23_2),
	.A(FE_OFN29191_sa23_2));
   INVx1_ASAP7_75t_SL FE_OCPC7652_FE_OFN29191_sa23_2 (.Y(n22951),
	.A(FE_OFN29191_sa23_2));
   INVx1_ASAP7_75t_L FE_OCPC7651_FE_OFN29191_sa23_2 (.Y(FE_OCPN27498_sa23_2),
	.A(FE_OFN29191_sa23_2));
   INVxp67_ASAP7_75t_L FE_OCPC7650_n26317 (.Y(n26318),
	.A(FE_OFN16340_n26317));
   INVx2_ASAP7_75t_SL FE_OCPC7649_n26317 (.Y(FE_OFN16340_n26317),
	.A(n26317));
   BUFx2_ASAP7_75t_SL FE_OCPC7648_n16191 (.Y(FE_OCPN29371_n16191),
	.A(n16191));
   BUFx2_ASAP7_75t_L FE_OCPC7647_FE_OFN28744_FE_OCPN27908 (.Y(FE_OCPN29370_FE_OFN28744),
	.A(FE_OFN28744_FE_OCPN27908));
   BUFx2_ASAP7_75t_SL FE_OCPC7646_n16982 (.Y(FE_OCPN29369_n16982),
	.A(FE_OFN28725_n16982));
   BUFx6f_ASAP7_75t_SL FE_OCPC7645_n16982 (.Y(FE_OFN28725_n16982),
	.A(n16982));
   BUFx2_ASAP7_75t_L FE_OCPC7644_FE_OFN16247_sa30_1 (.Y(FE_OCPN29368_FE_OFN16247_sa30_1),
	.A(FE_OFN16247_sa30_1));
   INVx1_ASAP7_75t_L FE_OCPC7643_sa22_0 (.Y(FE_OCPN29281_sa22_0),
	.A(n23183));
   INVx3_ASAP7_75t_SL FE_OCPC7642_sa22_0 (.Y(n23183),
	.A(sa22_0_));
   BUFx3_ASAP7_75t_SL FE_OCPC7641_sa22_0 (.Y(FE_OFN29152_sa22_0),
	.A(sa22_0_));
   BUFx2_ASAP7_75t_SL FE_OCPC7640_n26944 (.Y(n25621),
	.A(FE_OCPN27778_n25621));
   INVx1_ASAP7_75t_SL FE_OCPC7639_n26944 (.Y(FE_OCPN27778_n25621),
	.A(n26944));
   INVxp67_ASAP7_75t_SL FE_OCPC7637_n26773 (.Y(n26771),
	.A(FE_OCPN27935_n26773));
   BUFx2_ASAP7_75t_SL FE_OCPC7636_n26773 (.Y(FE_OCPN27935_n26773),
	.A(n26773));
   OAI21xp33_ASAP7_75t_SL FE_RC_888_0 (.Y(n637),
	.A1(n23937),
	.A2(n15915),
	.B(n15914));
   BUFx2_ASAP7_75t_SL FE_OCPC7635_n24639 (.Y(FE_OCPN29365_n24639),
	.A(n24639));
   INVx1_ASAP7_75t_L FE_RC_887_0 (.Y(n23725),
	.A(FE_RN_259_0));
   OR3x1_ASAP7_75t_L FE_RC_886_0 (.Y(FE_RN_259_0),
	.A(n23819),
	.B(n18571),
	.C(FE_OFN29250_FE_OCPN27371_sa20_2));
   BUFx3_ASAP7_75t_SL FE_OCPC7632_n25981 (.Y(FE_OCPN27514_n25981),
	.A(n25981));
   BUFx3_ASAP7_75t_SL FE_OCPC7631_n448 (.Y(FE_OCPN29364_n448),
	.A(n448));
   INVx1_ASAP7_75t_L FE_OCPC7630_n14011 (.Y(FE_OCPN29363_n14011),
	.A(FE_OFN28501_FE_OFN26020_n14010));
   BUFx2_ASAP7_75t_SL FE_OCPC7629_n14011 (.Y(FE_OFN26020_n14010),
	.A(FE_OFN28501_FE_OFN26020_n14010));
   INVx1_ASAP7_75t_SL FE_OCPC7628_n14011 (.Y(FE_OFN28501_FE_OFN26020_n14010),
	.A(n14011));
   INVxp33_ASAP7_75t_L FE_OCPC7626_n25696 (.Y(FE_OCPN29361_n25696),
	.A(n25697));
   BUFx2_ASAP7_75t_SL FE_OCPC7624_n26780 (.Y(FE_OFN28968_n26780),
	.A(n26780));
   AOI31xp33_ASAP7_75t_SL FE_RC_885_0 (.Y(n22214),
	.A1(n22212),
	.A2(n22474),
	.A3(FE_RN_4_0),
	.B(n27004));
   INVx2_ASAP7_75t_L FE_OCPC7622_n26990 (.Y(FE_OFN28451_n26990),
	.A(n26992));
   INVx2_ASAP7_75t_SL FE_OCPC7621_n26990 (.Y(n26992),
	.A(n26990));
   BUFx2_ASAP7_75t_SL FE_OCPC7620_n26586 (.Y(FE_OCPN29359_n26586),
	.A(FE_OCPN27358_n26586));
   BUFx2_ASAP7_75t_SL FE_OCPC7619_n26586 (.Y(FE_OCPN27358_n26586),
	.A(n26586));
   OAI22x1_ASAP7_75t_SL FE_RC_884_0 (.Y(n26632),
	.A1(n26082),
	.A2(n25606),
	.B1(n25606),
	.B2(n25605));
   INVx3_ASAP7_75t_SL FE_OCPC7618_n26115 (.Y(FE_OFN26024_n26115),
	.A(n26784));
   BUFx3_ASAP7_75t_SL FE_OCPC7617_n26115 (.Y(n26784),
	.A(n26115));
   INVx1_ASAP7_75t_SL FE_OCPC7616_n14664 (.Y(FE_OFN16273_n14664),
	.A(n14664));
   BUFx2_ASAP7_75t_SL FE_OCPC7615_n14664 (.Y(n14663),
	.A(n14664));
   BUFx6f_ASAP7_75t_SL FE_OCPC7614_sa13_1 (.Y(FE_OFN16444_sa13_1),
	.A(sa13_1_));
   OAI21xp33_ASAP7_75t_L FE_RC_883_0 (.Y(n18146),
	.A1(FE_OCPN27460_n16913),
	.A2(n16874),
	.B(n16945));
   INVx2_ASAP7_75t_SL FE_OCPC7613_n25132 (.Y(FE_OCPN5112_n25135),
	.A(n25132));
   INVxp67_ASAP7_75t_SL FE_OCPC7612_n17159 (.Y(FE_OCPN29358_n17159),
	.A(n17103));
   INVx2_ASAP7_75t_SL FE_OCPC7610_n17159 (.Y(n17103),
	.A(n17159));
   INVxp67_ASAP7_75t_SL FE_OCPC7609_n27110 (.Y(FE_OCPN29356_n27110),
	.A(n27110));
   INVx1_ASAP7_75t_SL FE_OCPC7608_n27110 (.Y(n26754),
	.A(n27110));
   BUFx2_ASAP7_75t_SL FE_OCPC7607_n492 (.Y(FE_OCPN29355_n492),
	.A(n492));
   AOI31xp33_ASAP7_75t_SL FE_RC_882_0 (.Y(n22172),
	.A1(n22171),
	.A2(n24795),
	.A3(n22170),
	.B(n26926));
   INVxp67_ASAP7_75t_L FE_OCPC7606_n26853 (.Y(n26850),
	.A(FE_OCPN27377_n26853));
   HB1xp67_ASAP7_75t_SL FE_OCPC7605_n26853 (.Y(FE_OCPN27377_n26853),
	.A(n26853));
   INVx2_ASAP7_75t_SL FE_OCPC7604_sa00_1 (.Y(FE_OFN148_sa00_1),
	.A(sa00_1_));
   BUFx4f_ASAP7_75t_SL FE_OCPC7603_sa00_1 (.Y(FE_OFN28514_sa00_1),
	.A(sa00_1_));
   BUFx2_ASAP7_75t_L FE_OCPC7601_n26586 (.Y(FE_OCPN29353_n26586),
	.A(FE_OCPN27358_n26586));
   BUFx2_ASAP7_75t_L FE_OCPC7599_n25173 (.Y(FE_OCPN29352_n25173),
	.A(n25173));
   BUFx3_ASAP7_75t_SL FE_OCPC7598_FE_OFN26116_sa13_1 (.Y(FE_OCPN29351_FE_OFN26116_sa13_1),
	.A(FE_OFN16444_sa13_1));
   INVx3_ASAP7_75t_SL FE_OCPC7597_FE_OFN26116_sa13_1 (.Y(FE_OFN26061_n),
	.A(FE_OFN16444_sa13_1));
   INVx2_ASAP7_75t_SL FE_OCPC7593_n27158 (.Y(n27162),
	.A(n27158));
   HB1xp67_ASAP7_75t_SL FE_OCPC7592_w3_25 (.Y(FE_OCPN29350_w3_25),
	.A(w3_25_));
   INVxp67_ASAP7_75t_R FE_OCPC7591_n26113 (.Y(n24540),
	.A(FE_OCPN27314_n26113));
   HB1xp67_ASAP7_75t_L FE_OCPC7590_n26113 (.Y(FE_OCPN27314_n26113),
	.A(n26113));
   BUFx2_ASAP7_75t_SL FE_OCPC7589_n26098 (.Y(FE_OCPN5045_n26098),
	.A(n26098));
   NAND3xp33_ASAP7_75t_SL FE_RC_881_0 (.Y(n15195),
	.A(FE_OFN27129_w3_28),
	.B(FE_OCPN28096_w3_31),
	.C(FE_OFN28452_w3_29));
   BUFx12f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_8 (.Y(CTS_39),
	.A(CTS_40));
   BUFx12f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_7 (.Y(CTS_38),
	.A(CTS_40));
   BUFx12f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_6 (.Y(CTS_37),
	.A(CTS_40));
   BUFx16f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_5 (.Y(CTS_36),
	.A(CTS_40));
   BUFx6f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L1_2 (.Y(CTS_40),
	.A(clk));
   BUFx16f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_4 (.Y(CTS_34),
	.A(CTS_35));
   BUFx16f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_3 (.Y(CTS_33),
	.A(CTS_35));
   BUFx10_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_2 (.Y(CTS_32),
	.A(CTS_35));
   BUFx12f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L2_1 (.Y(CTS_31),
	.A(CTS_35));
   BUFx6f_ASAP7_75t_SL CTS_ccl_a_BUF_clk_G0_L1_1 (.Y(CTS_35),
	.A(clk));
   HB1xp67_ASAP7_75t_R FE_OCPC7662_n26633 (.Y(FE_OCPN7662_n26633),
	.A(FE_OCPN27284_n26633));
   BUFx6f_ASAP7_75t_L FE_OCPC7584_n27113 (.Y(FE_OFN29010_n27113),
	.A(n27113));
   BUFx6f_ASAP7_75t_L FE_OCPC7583_FE_OCPN27405_sa03_4 (.Y(FE_OCPN29349_FE_OCPN27405_sa03_4),
	.A(FE_OCPN27405_sa03_4));
   BUFx2_ASAP7_75t_SRAM FE_OCPC7582_FE_OCPN27405_sa03_4 (.Y(FE_OFN28997_sa03_4),
	.A(FE_OCPN27405_sa03_4));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7660_FE_OFN28720_sa20_1 (.Y(FE_OCPN7660_FE_OFN28720_sa20_1),
	.A(FE_OCPN29380_sa20_1));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7658_n27056 (.Y(FE_OCPN7658_n27056),
	.A(n27056));
   BUFx2_ASAP7_75t_L FE_OCPC7657_n26213 (.Y(FE_OCPN7657_n26213),
	.A(n26213));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7656_n24301 (.Y(FE_OCPN7656_n24301),
	.A(n24301));
   HB1xp67_ASAP7_75t_L FE_OCPC7653_n24270 (.Y(FE_OCPN7653_n24270),
	.A(n24270));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7650_n27110 (.Y(FE_OCPN7650_n27110),
	.A(n27110));
   HB1xp67_ASAP7_75t_SL FE_OCPC7649_n23259 (.Y(FE_OCPN7649_n23259),
	.A(n23259));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7647_FE_OFN141_sa03_1 (.Y(FE_OCPN7647_FE_OFN141_sa03_1),
	.A(FE_OFN141_sa03_1));
   HB1xp67_ASAP7_75t_SL FE_OCPC7645_n20962 (.Y(FE_OCPN7645_n20962),
	.A(n20962));
   BUFx2_ASAP7_75t_SL FE_OCPC7644_n21523 (.Y(FE_OCPN7644_n21523),
	.A(n21523));
   HB1xp67_ASAP7_75t_R FE_OCPC7643_n17646 (.Y(FE_OCPN7643_n17646),
	.A(n17646));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7642_n26319 (.Y(FE_OCPN7642_n26319),
	.A(FE_OCPN8217_n26319));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7641_n25778 (.Y(FE_OCPN7641_n25778),
	.A(n25778));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7640_n18765 (.Y(FE_OCPN7640_n18765),
	.A(n18765));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7638_n26183 (.Y(FE_OCPN7638_n26183),
	.A(n26183));
   BUFx2_ASAP7_75t_L FE_OCPC7636_n25940 (.Y(FE_OCPN7636_n25940),
	.A(n25940));
   HB1xp67_ASAP7_75t_R FE_OCPC7633_n26815 (.Y(FE_OCPN7633_n26815),
	.A(n26815));
   HB1xp67_ASAP7_75t_R FE_OCPC7631_n24750 (.Y(FE_OCPN7631_n24750),
	.A(FE_OCPN29262_n24750));
   HB1xp67_ASAP7_75t_R FE_OCPC7629_FE_OFN105_n27178 (.Y(FE_OCPN7629_FE_OFN105_n27178),
	.A(FE_OFN105_n27178));
   HB1xp67_ASAP7_75t_L FE_OCPC7626_n18582 (.Y(FE_OCPN7626_n18582),
	.A(n18582));
   HB1xp67_ASAP7_75t_L FE_OCPC7625_n26501 (.Y(FE_OCPN7625_n26501),
	.A(FE_OCPN28054_n26501));
   HB1xp67_ASAP7_75t_R FE_OCPC7623_FE_OFN4_w3_22 (.Y(FE_OCPN7623_FE_OFN4_w3_22),
	.A(FE_OFN4_w3_22));
   BUFx2_ASAP7_75t_SL FE_OCPC7622_n24526 (.Y(FE_OCPN7622_n24526),
	.A(n24526));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7621_n26898 (.Y(FE_OCPN7621_n26898),
	.A(n26898));
   HB1xp67_ASAP7_75t_R FE_OCPC7620_n25761 (.Y(FE_OCPN7620_n25761),
	.A(n25761));
   HB1xp67_ASAP7_75t_R FE_OCPC7619_FE_OFN28689_sa03_5 (.Y(FE_OCPN7619_FE_OFN28689_sa03_5),
	.A(FE_OFN29179_n));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7618_n21027 (.Y(FE_OCPN7618_n21027),
	.A(n21027));
   HB1xp67_ASAP7_75t_L FE_OCPC7617_n26009 (.Y(FE_OCPN7617_n26009),
	.A(n26009));
   HB1xp67_ASAP7_75t_R FE_OCPC7613_n24166 (.Y(FE_OCPN7613_n24166),
	.A(FE_OCPN8211_n24166));
   HB1xp67_ASAP7_75t_R FE_OCPC7612_n25229 (.Y(FE_OCPN7612_n25229),
	.A(n25229));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7610_n25861 (.Y(FE_OCPN7610_n25861),
	.A(n25861));
   HB1xp67_ASAP7_75t_L FE_OCPC7607_n23539 (.Y(FE_OCPN7607_n23539),
	.A(n23539));
   HB1xp67_ASAP7_75t_R FE_OCPC7605_n26234 (.Y(FE_OCPN7605_n26234),
	.A(n26234));
   HB1xp67_ASAP7_75t_SL FE_OCPC7599_n26721 (.Y(FE_OCPN7599_n26721),
	.A(n26721));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7598_n25174 (.Y(FE_OCPN7598_n25174),
	.A(n25174));
   BUFx2_ASAP7_75t_SL FE_OCPC7597_n21981 (.Y(FE_OCPN7597_n21981),
	.A(n21981));
   HB1xp67_ASAP7_75t_R FE_OCPC7596_n24647 (.Y(FE_OCPN7596_n24647),
	.A(n24647));
   HB1xp67_ASAP7_75t_L FE_OCPC7595_n17426 (.Y(FE_OCPN7595_n17426),
	.A(n17426));
   BUFx2_ASAP7_75t_L FE_OCPC7586_n17693 (.Y(FE_OCPN7586_n17693),
	.A(n17693));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7585_FE_OFN25926_n26922 (.Y(FE_OCPN7585_FE_OFN25926_n26922),
	.A(FE_OFN25926_n26922));
   HB1xp67_ASAP7_75t_L FE_OCPC7584_n23447 (.Y(FE_OCPN7584_n23447),
	.A(n23447));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC7583_n26983 (.Y(FE_OCPN7583_n26983),
	.A(n26983));
   BUFx2_ASAP7_75t_SL FE_OCPC7581_n17592 (.Y(FE_OCPN29348_n17592),
	.A(n17592));
   INVx2_ASAP7_75t_L FE_RC_880_0 (.Y(n25149),
	.A(FE_RN_258_0));
   OR3x1_ASAP7_75t_L FE_RC_879_0 (.Y(FE_RN_258_0),
	.A(n18305),
	.B(FE_OFN28928_n22374),
	.C(n20112));
   BUFx3_ASAP7_75t_SL FE_OCPC7579_n12998 (.Y(FE_OCPN29346_n12998),
	.A(n12998));
   NAND3x1_ASAP7_75t_L FE_RC_878_0 (.Y(n23762),
	.A(n20658),
	.B(n20659),
	.C(n23870));
   AOI22x1_ASAP7_75t_SL FE_RC_877_0 (.Y(n16127),
	.A1(n25411),
	.A2(n15898),
	.B1(w1_15_),
	.B2(FE_OCPN28327_n15899));
   NOR3xp33_ASAP7_75t_SL FE_RC_876_0 (.Y(n24000),
	.A(n24943),
	.B(n21900),
	.C(n19675));
   NOR3x1_ASAP7_75t_L FE_RC_875_0 (.Y(n27078),
	.A(FE_OCPN27391_n27079),
	.B(n27081),
	.C(FE_OCPN28438_n27080));
   AOI21xp5_ASAP7_75t_SL FE_RC_874_0 (.Y(n14080),
	.A1(n14078),
	.A2(n15757),
	.B(n14079));
   BUFx2_ASAP7_75t_SL FE_OCPC7575_n25357 (.Y(FE_OCPN29342_n25357),
	.A(n25357));
   BUFx2_ASAP7_75t_SL FE_OCPC7574_FE_OFN29148_n (.Y(FE_OCPN29341_FE_OFN29148_n),
	.A(FE_OFN29148_n));
   BUFx2_ASAP7_75t_L FE_OCPC7573_n17079 (.Y(FE_OCPN29340_n17079),
	.A(n17079));
   AOI31xp33_ASAP7_75t_SL FE_RC_873_0 (.Y(n18782),
	.A1(n19141),
	.A2(n18781),
	.A3(n18780),
	.B(n26777));
   NOR3x1_ASAP7_75t_L FE_RC_872_0 (.Y(n24887),
	.A(n22672),
	.B(n22671),
	.C(n22673));
   OAI21xp5_ASAP7_75t_SL FE_RC_871_0 (.Y(n27108),
	.A1(FE_OFN26559_n26754),
	.A2(n27109),
	.B(FE_OFN16215_ld_r));
   HB1xp67_ASAP7_75t_SL FE_OCPC7556_n26504 (.Y(FE_OCPN7556_n26504),
	.A(n26504));
   BUFx3_ASAP7_75t_SL FE_OCPC7568_n26602 (.Y(FE_OCPN29335_n),
	.A(FE_OCPN27419_n26602));
   NAND3x1_ASAP7_75t_L FE_RC_870_0 (.Y(n21268),
	.A(n19457),
	.B(n23416),
	.C(n19456));
   BUFx2_ASAP7_75t_L FE_OCPC7567_n17330 (.Y(FE_OCPN29334_n17330),
	.A(n17330));
   HB1xp67_ASAP7_75t_SL FE_OCPC7566_n17330 (.Y(FE_OCPN29333_n17330),
	.A(n17330));
   INVx1_ASAP7_75t_L FE_RC_869_0 (.Y(n20265),
	.A(FE_RN_257_0));
   OR3x1_ASAP7_75t_L FE_RC_868_0 (.Y(FE_RN_257_0),
	.A(n22979),
	.B(FE_OCPN27710_n19011),
	.C(FE_OCPN27881_FE_OFN27126_sa23_3));
   HB1xp67_ASAP7_75t_L FE_OCPC7564_n20933 (.Y(FE_OCPN29331_n20933),
	.A(n20933));
   BUFx2_ASAP7_75t_L FE_OCPC7563_n26459 (.Y(FE_OCPN29330_n26459),
	.A(n26459));
   NAND3x1_ASAP7_75t_SL FE_RC_867_0 (.Y(n26395),
	.A(n26398),
	.B(n26397),
	.C(n26396));
   HB1xp67_ASAP7_75t_SL FE_OCPC7562_n15517 (.Y(FE_OCPN29329_n15517),
	.A(n15517));
   NAND3x1_ASAP7_75t_L FE_RC_866_0 (.Y(n24485),
	.A(n16686),
	.B(n18128),
	.C(n16840));
   AOI31xp33_ASAP7_75t_SL FE_RC_865_0 (.Y(n24265),
	.A1(n24264),
	.A2(n24261),
	.A3(FE_OFN29215_n24262),
	.B(n24263));
   INVx2_ASAP7_75t_L FE_RC_864_0 (.Y(n15779),
	.A(FE_RN_256_0));
   OR3x1_ASAP7_75t_L FE_RC_863_0 (.Y(FE_RN_256_0),
	.A(FE_OFN25899_w3_4),
	.B(FE_OFN29052_w3_5),
	.C(FE_OFN28661_w3_7));
   OAI21xp33_ASAP7_75t_R FE_RC_862_0 (.Y(n13428),
	.A1(FE_OCPN29547_n15183),
	.A2(FE_OFN27212_w3_30),
	.B(FE_OFN28817_n));
   INVxp67_ASAP7_75t_L FE_RC_861_0 (.Y(FE_RN_253_0),
	.A(n21477));
   INVxp67_ASAP7_75t_L FE_RC_860_0 (.Y(FE_RN_254_0),
	.A(n21478));
   NAND2xp5_ASAP7_75t_L FE_RC_859_0 (.Y(FE_RN_255_0),
	.A(FE_RN_253_0),
	.B(FE_RN_254_0));
   NOR2xp33_ASAP7_75t_SL FE_RC_858_0 (.Y(n21487),
	.A(FE_RN_255_0),
	.B(FE_OFN25949_n21475));
   NAND3x1_ASAP7_75t_SL FE_RC_857_0 (.Y(n21799),
	.A(n18208),
	.B(n21085),
	.C(n20702));
   AOI31xp33_ASAP7_75t_SL FE_RC_856_0 (.Y(n21489),
	.A1(n21487),
	.A2(n21488),
	.A3(n21486),
	.B(n26777));
   BUFx2_ASAP7_75t_SL FE_OCPC7560_n21017 (.Y(FE_OCPN29327_n21017),
	.A(n21017));
   AOI22x1_ASAP7_75t_SL FE_RC_854_0 (.Y(n16134),
	.A1(n24073),
	.A2(n15773),
	.B1(w1_22_),
	.B2(FE_OCPN28065_n15774));
   OAI21xp5_ASAP7_75t_SL FE_RC_853_0 (.Y(n25572),
	.A1(FE_OCPN29356_n27110),
	.A2(n25573),
	.B(FE_OFN16215_ld_r));
   OAI21xp5_ASAP7_75t_L FE_RC_852_0 (.Y(n23139),
	.A1(n16533),
	.A2(FE_OFN28910_n16534),
	.B(n16637));
   OAI21x1_ASAP7_75t_SL FE_RC_851_0 (.Y(n26694),
	.A1(n26695),
	.A2(n26696),
	.B(FE_OFN14_FE_DBTN0_ld_r));
   BUFx4f_ASAP7_75t_SL FE_OCPC7557_n23216 (.Y(FE_OCPN29324_n23216),
	.A(n23216));
   BUFx3_ASAP7_75t_SL FE_OCPC7556_n19721 (.Y(FE_OCPN29323_n19721),
	.A(n19721));
   AOI31xp33_ASAP7_75t_SL FE_RC_850_0 (.Y(n25883),
	.A1(n19370),
	.A2(n18962),
	.A3(n26001),
	.B(n27095));
   AND2x2_ASAP7_75t_R FE_RC_849_0 (.Y(FE_RN_252_0),
	.A(n26942),
	.B(n26907));
   OAI21x1_ASAP7_75t_SL FE_RC_848_0 (.Y(n27202),
	.A1(FE_RN_252_0),
	.A2(n26906),
	.B(n26905));
   OAI211xp5_ASAP7_75t_SL FE_RC_847_0 (.Y(n24114),
	.A1(n23345),
	.A2(FE_RN_158_0),
	.B(FE_RN_154_0),
	.C(FE_RN_155_0));
   AND2x2_ASAP7_75t_L FE_RC_846_0 (.Y(FE_RN_251_0),
	.A(n27117),
	.B(FE_PSN8300_n26482));
   OAI21xp5_ASAP7_75t_SL FE_RC_845_0 (.Y(n26434),
	.A1(FE_RN_251_0),
	.A2(n25973),
	.B(n25972));
   NOR3x1_ASAP7_75t_L FE_RC_844_0 (.Y(n21806),
	.A(n22320),
	.B(n21802),
	.C(n22838));
   AND2x2_ASAP7_75t_SRAM FE_RC_843_0 (.Y(FE_RN_250_0),
	.A(FE_OCPN27442_n27202),
	.B(FE_OFN16215_ld_r));
   AND2x2_ASAP7_75t_SL FE_RC_841_0 (.Y(FE_RN_249_0),
	.A(n25652),
	.B(n25651));
   OAI21x1_ASAP7_75t_SL FE_RC_840_0 (.Y(n465),
	.A1(FE_RN_249_0),
	.A2(n25650),
	.B(n25649));
   INVx1_ASAP7_75t_SL FE_RC_835_0 (.Y(FE_RN_248_0),
	.A(FE_RN_247_0));
   OAI22xp5_ASAP7_75t_SL FE_RC_834_0 (.Y(n25270),
	.A1(FE_OCPN27310_n26389),
	.A2(FE_RN_248_0),
	.B1(n26388),
	.B2(FE_RN_247_0));
   AO21x1_ASAP7_75t_SL FE_RC_833_0 (.Y(FE_RN_243_0),
	.A1(FE_OCPN27274_n26394),
	.A2(FE_OFN28484_ld_r),
	.B(n26393));
   NAND2x1p5_ASAP7_75t_SL FE_RC_832_0 (.Y(n26398),
	.A(FE_RN_243_0),
	.B(n26392));
   OA21x2_ASAP7_75t_L FE_RC_831_0 (.Y(FE_RN_242_0),
	.A1(n25359),
	.A2(n25358),
	.B(n26829));
   NOR2x1p5_ASAP7_75t_SL FE_RC_830_0 (.Y(n25362),
	.A(FE_RN_242_0),
	.B(FE_OCPN29342_n25357));
   BUFx2_ASAP7_75t_SL FE_OCPC7554_n17876 (.Y(FE_OCPN29321_n17876),
	.A(n17876));
   HB1xp67_ASAP7_75t_R FE_OCPC7547_sa03_4 (.Y(FE_OCPN29314_n),
	.A(FE_OCPN27405_sa03_4));
   BUFx2_ASAP7_75t_SL FE_OCPC7542_n26452 (.Y(FE_OCPN29309_n26452),
	.A(n26452));
   HB1xp67_ASAP7_75t_L FE_OCPC7541_sa22_1 (.Y(FE_OCPN29308_n),
	.A(FE_OCPN29269_sa22_1));
   BUFx3_ASAP7_75t_SL FE_OCPC7538_n23302 (.Y(FE_OCPN29305_n23302),
	.A(n23302));
   BUFx2_ASAP7_75t_L FE_OCPC7537_n17526 (.Y(FE_OCPN29304_n17526),
	.A(n17526));
   BUFx6f_ASAP7_75t_SL FE_OCPC7535_sa00_4 (.Y(FE_OCPN29302_sa00_4),
	.A(sa00_4_));
   BUFx2_ASAP7_75t_L FE_OCPC7532_FE_OFN29232_n16875 (.Y(FE_OCPN29299_FE_OFN29232_n16875),
	.A(n16875));
   BUFx3_ASAP7_75t_SL FE_OCPC7531_n25028 (.Y(FE_OCPN29298_n25028),
	.A(n25028));
   HB1xp67_ASAP7_75t_SL FE_OCPC7528_n18739 (.Y(FE_OCPN29295_n18739),
	.A(n18739));
   BUFx2_ASAP7_75t_L FE_OCPC7527_n23925 (.Y(FE_OCPN29294_n23925),
	.A(n23925));
   BUFx3_ASAP7_75t_SL FE_OCPC7526_FE_OFN28678_sa21_3 (.Y(FE_OCPN29293_FE_OFN28678_sa21_3),
	.A(FE_OFN28678_sa21_3));
   BUFx4f_ASAP7_75t_SL FE_OCPC7524_n17282 (.Y(FE_OCPN29291_n17282),
	.A(n17282));
   BUFx2_ASAP7_75t_SL FE_OCPC7522_n22162 (.Y(FE_OCPN29289_n22162),
	.A(n22162));
   BUFx3_ASAP7_75t_SL FE_OCPC7520_n27210 (.Y(FE_OCPN29287_n27210),
	.A(n27210));
   BUFx2_ASAP7_75t_SL FE_OCPC7517_n19821 (.Y(FE_OCPN29284_n19821),
	.A(n19821));
   BUFx6f_ASAP7_75t_SL FE_OCPC7516_n23439 (.Y(FE_OCPN29283_n23439),
	.A(n23439));
   BUFx2_ASAP7_75t_SL FE_OCPC7512_n25353 (.Y(FE_OCPN29279_n25353),
	.A(n25353));
   BUFx2_ASAP7_75t_SL FE_OCPC7510_n26713 (.Y(FE_OCPN29277_n26713),
	.A(n26713));
   BUFx3_ASAP7_75t_SL FE_OCPC7507_n26478 (.Y(FE_OCPN29274_n26478),
	.A(n26478));
   BUFx4f_ASAP7_75t_SL FE_OCPC7502_sa22_1 (.Y(FE_OCPN29269_sa22_1),
	.A(sa22_1_));
   BUFx2_ASAP7_75t_L FE_OCPC7498_FE_OFN28698_sa21_1 (.Y(FE_OCPN29265_FE_OFN28698_sa21_1),
	.A(FE_OFN28698_sa21_1));
   BUFx2_ASAP7_75t_SL FE_OCPC7496_n24537 (.Y(FE_OCPN29263_n24537),
	.A(n24537));
   BUFx3_ASAP7_75t_SL FE_OCPC7495_n24750 (.Y(FE_OCPN29262_n24750),
	.A(n24750));
   BUFx4f_ASAP7_75t_SL FE_OCPC7493_sa00_5 (.Y(FE_OCPN29260_sa00_5),
	.A(sa00_5_));
   BUFx2_ASAP7_75t_L FE_OCPC7491_n27171 (.Y(FE_OCPN29258_n27171),
	.A(n27171));
   OAI21x1_ASAP7_75t_SL FE_RC_829_0 (.Y(n27171),
	.A1(n25918),
	.A2(FE_RN_110_0),
	.B(n25917));
   NOR3xp33_ASAP7_75t_SL FE_RC_828_0 (.Y(n25929),
	.A(n25927),
	.B(FE_OCPN7636_n25940),
	.C(FE_OFN13_FE_DBTN0_ld_r));
   INVx1_ASAP7_75t_L FE_RC_827_0 (.Y(FE_RN_238_0),
	.A(n25423));
   NAND2xp5_ASAP7_75t_SL FE_RC_826_0 (.Y(FE_RN_239_0),
	.A(n25422),
	.B(n25421));
   OAI21xp5_ASAP7_75t_SL FE_RC_825_0 (.Y(FE_RN_240_0),
	.A1(n25422),
	.A2(n25421),
	.B(FE_RN_239_0));
   INVx1_ASAP7_75t_SL FE_RC_824_0 (.Y(FE_RN_241_0),
	.A(FE_RN_240_0));
   OAI22xp5_ASAP7_75t_SL FE_RC_823_0 (.Y(n25425),
	.A1(n25423),
	.A2(FE_RN_241_0),
	.B1(FE_RN_238_0),
	.B2(FE_RN_240_0));
   BUFx2_ASAP7_75t_SL FE_OCPC7490_n474 (.Y(FE_OCPN29257_n474),
	.A(n474));
   BUFx3_ASAP7_75t_SL FE_OCPC7489_n418 (.Y(FE_OCPN29256_n418),
	.A(n418));
   AOI21xp5_ASAP7_75t_L FE_RC_822_0 (.Y(n580),
	.A1(key_34_),
	.A2(ld),
	.B(n15903));
   AOI21xp33_ASAP7_75t_L FE_RC_821_0 (.Y(n23174),
	.A1(FE_OFN26141_n23307),
	.A2(n18161),
	.B(n21122));
   AOI21x1_ASAP7_75t_SL FE_RC_819_0 (.Y(n16058),
	.A1(n26202),
	.A2(n16059),
	.B(n16125));
   INVxp67_ASAP7_75t_L FE_RC_818_0 (.Y(FE_RN_237_0),
	.A(n16172));
   AOI21xp5_ASAP7_75t_SRAM FE_RC_817_0 (.Y(n610),
	.A1(key_49_),
	.A2(FE_OFN0_ld),
	.B(FE_RN_237_0));
   XOR2xp5_ASAP7_75t_SL FE_RC_816_0 (.Y(n26133),
	.A(FE_OCPN28140_FE_OFN133_n24306),
	.B(FE_RN_24_0));
   AOI21xp33_ASAP7_75t_L FE_RC_815_0 (.Y(n622),
	.A1(key_48_),
	.A2(ld),
	.B(FE_OFN26021_n16253));
   AOI21xp5_ASAP7_75t_L FE_RC_814_0 (.Y(n547),
	.A1(key_43_),
	.A2(FE_OFN21_n16125),
	.B(n16266));
   XOR2xp5_ASAP7_75t_SL FE_RC_813_0 (.Y(n25154),
	.A(FE_OCPN5041_n26726),
	.B(FE_RN_74_0));
   XOR2xp5_ASAP7_75t_SL FE_RC_812_0 (.Y(FE_RN_26_0),
	.A(n27143),
	.B(n27141));
   AOI21xp5_ASAP7_75t_SL FE_RC_811_0 (.Y(n16224),
	.A1(n26963),
	.A2(n16225),
	.B(n16125));
   AOI21xp5_ASAP7_75t_SL FE_RC_810_0 (.Y(n16126),
	.A1(n27085),
	.A2(n16127),
	.B(FE_OFN21_n16125));
   AOI21xp5_ASAP7_75t_SL FE_RC_809_0 (.Y(n16218),
	.A1(n26951),
	.A2(n16219),
	.B(FE_OFN21_n16125));
   OR2x2_ASAP7_75t_SL FE_RC_808_0 (.Y(n25447),
	.A(FE_RN_204_0),
	.B(FE_RN_205_0));
   AOI21xp5_ASAP7_75t_L FE_RC_807_0 (.Y(n23291),
	.A1(n23289),
	.A2(n26082),
	.B(n23290));
   OR2x2_ASAP7_75t_L FE_RC_806_0 (.Y(n27022),
	.A(n27019),
	.B(n27018));
   AND2x2_ASAP7_75t_SL FE_RC_805_0 (.Y(n26765),
	.A(n26882),
	.B(n24707));
   OR3x1_ASAP7_75t_SL FE_RC_804_0 (.Y(FE_OFN16316_n24840),
	.A(n23904),
	.B(n23906),
	.C(n23911));
   AOI21xp5_ASAP7_75t_L FE_RC_803_0 (.Y(n27074),
	.A1(n26046),
	.A2(n26407),
	.B(n26047));
   OR3x1_ASAP7_75t_SL FE_RC_802_0 (.Y(FE_OFN16235_n15055),
	.A(n15054),
	.B(n15053),
	.C(n15052));
   OR2x2_ASAP7_75t_SL FE_RC_801_0 (.Y(n25038),
	.A(n19459),
	.B(n18057));
   AOI31xp33_ASAP7_75t_SL FE_RC_800_0 (.Y(n20484),
	.A1(n20448),
	.A2(n20447),
	.A3(FE_OCPN28172_n20449),
	.B(n26687));
   AOI31xp33_ASAP7_75t_R FE_RC_799_0 (.Y(n24730),
	.A1(n24728),
	.A2(n24964),
	.A3(n24729),
	.B(n25139));
   OR3x1_ASAP7_75t_SL FE_RC_798_0 (.Y(n24440),
	.A(n19458),
	.B(n23450),
	.C(n21268));
   AND2x2_ASAP7_75t_L FE_RC_797_0 (.Y(n19419),
	.A(n18941),
	.B(n17101));
   AOI21x1_ASAP7_75t_SL FE_RC_796_0 (.Y(n20417),
	.A1(n25069),
	.A2(n26457),
	.B(n27004));
   INVxp33_ASAP7_75t_R FE_RC_795_0 (.Y(FE_RN_236_0),
	.A(FE_PSN8296_FE_OFN26588_n24062));
   AOI31xp33_ASAP7_75t_SL FE_RC_794_0 (.Y(n24063),
	.A1(FE_RN_236_0),
	.A2(n24061),
	.A3(n24060),
	.B(n24377));
   AOI21xp33_ASAP7_75t_R FE_RC_793_0 (.Y(n23116),
	.A1(n23084),
	.A2(n23085),
	.B(n27015));
   A2O1A1Ixp33_ASAP7_75t_L FE_RC_792_0 (.Y(n19496),
	.A1(n19484),
	.A2(n21506),
	.B(n23467),
	.C(FE_RN_40_0));
   AOI31xp33_ASAP7_75t_L FE_RC_791_0 (.Y(n24132),
	.A1(n24130),
	.A2(n24137),
	.A3(n24131),
	.B(n26687));
   AOI31xp33_ASAP7_75t_L FE_RC_790_0 (.Y(n25626),
	.A1(n20216),
	.A2(n25275),
	.A3(n25274),
	.B(n27140));
   AOI31xp33_ASAP7_75t_SL FE_RC_789_0 (.Y(n27120),
	.A1(n26359),
	.A2(n26358),
	.A3(n26360),
	.B(n26542));
   AOI31xp33_ASAP7_75t_L FE_RC_788_0 (.Y(n24049),
	.A1(n20604),
	.A2(n20603),
	.A3(n25163),
	.B(n26607));
   NOR3xp33_ASAP7_75t_L FE_RC_787_0 (.Y(n20283),
	.A(n20236),
	.B(n22929),
	.C(n22002));
   AOI21xp5_ASAP7_75t_SL FE_RC_786_0 (.Y(n14958),
	.A1(n14955),
	.A2(n14957),
	.B(n14956));
   OR3x1_ASAP7_75t_SL FE_RC_785_0 (.Y(n25996),
	.A(n18287),
	.B(n20490),
	.C(n18286));
   AOI21xp33_ASAP7_75t_L FE_RC_784_0 (.Y(n26073),
	.A1(n21349),
	.A2(FE_PSN8310_n17473),
	.B(n21346));
   AOI31xp33_ASAP7_75t_SL FE_RC_783_0 (.Y(n13694),
	.A1(n13692),
	.A2(n13691),
	.A3(FE_OFN28717_n15158),
	.B(n13693));
   INVx1_ASAP7_75t_L FE_RC_782_0 (.Y(FE_RN_235_0),
	.A(n21442));
   NOR2x1_ASAP7_75t_SL FE_RC_781_0 (.Y(n18653),
	.A(FE_RN_235_0),
	.B(n26101));
   AND2x2_ASAP7_75t_SL FE_RC_780_0 (.Y(n24669),
	.A(n19665),
	.B(n19664));
   AOI31xp33_ASAP7_75t_L FE_RC_779_0 (.Y(n14082),
	.A1(FE_OFN28623_n13874),
	.A2(FE_OFN27066_n13869),
	.A3(FE_OFN5_w3_22),
	.B(n14029));
   AOI31xp33_ASAP7_75t_SL FE_RC_778_0 (.Y(n20210),
	.A1(FE_OCPN27579_FE_OFN16138_sa02_5),
	.A2(FE_OFN28730_FE_OCPN28416_sa02_3),
	.A3(FE_OCPN27384_n22888),
	.B(n20209));
   OA21x2_ASAP7_75t_R FE_RC_777_0 (.Y(n20865),
	.A1(n16397),
	.A2(FE_OCPN28394_FE_OFN27043_n),
	.B(n16519));
   OA21x2_ASAP7_75t_L FE_RC_776_0 (.Y(n16544),
	.A1(FE_OFN28751_n),
	.A2(n16616),
	.B(n17222));
   AOI21xp5_ASAP7_75t_L FE_RC_775_0 (.Y(n23034),
	.A1(FE_OCPN28157_n16534),
	.A2(FE_OFN28807_n24944),
	.B(FE_OFN29159_n21892));
   AOI21x1_ASAP7_75t_L FE_RC_774_0 (.Y(n23370),
	.A1(FE_OCPN29435_n17445),
	.A2(FE_OCPN5021_n17446),
	.B(n21854));
   AOI31xp33_ASAP7_75t_L FE_RC_773_0 (.Y(n15971),
	.A1(n15959),
	.A2(FE_OFN26131_n15376),
	.A3(n15948),
	.B(n15947));
   INVxp33_ASAP7_75t_L FE_RC_772_0 (.Y(FE_RN_234_0),
	.A(n15616));
   AOI21xp33_ASAP7_75t_R FE_RC_771_0 (.Y(n15620),
	.A1(n15617),
	.A2(n15619),
	.B(FE_RN_234_0));
   AOI21xp33_ASAP7_75t_L FE_RC_770_0 (.Y(n23333),
	.A1(FE_OFN27173_n),
	.A2(n22828),
	.B(n22825));
   AOI21xp5_ASAP7_75t_L FE_RC_769_0 (.Y(n17417),
	.A1(n16417),
	.A2(n17416),
	.B(n17415));
   AOI21xp5_ASAP7_75t_SL FE_RC_768_0 (.Y(n17807),
	.A1(FE_OCPN27570_n17791),
	.A2(FE_OFN108_n26971),
	.B(n25524));
   AOI31xp33_ASAP7_75t_L FE_RC_767_0 (.Y(n16761),
	.A1(FE_OFN28779_n24257),
	.A2(FE_OCPN27616_n16760),
	.A3(FE_OCPN29265_FE_OFN28698_sa21_1),
	.B(n20345));
   OR2x2_ASAP7_75t_SL FE_RC_766_0 (.Y(n18742),
	.A(FE_OFN29062_n18651),
	.B(n17300));
   AOI21x1_ASAP7_75t_L FE_RC_765_0 (.Y(n22021),
	.A1(FE_OFN16248_n20235),
	.A2(n19000),
	.B(n18988));
   AOI21xp5_ASAP7_75t_L FE_RC_764_0 (.Y(n18009),
	.A1(FE_OCPN28001_n21310),
	.A2(n21708),
	.B(n18008));
   AOI21xp5_ASAP7_75t_L FE_RC_763_0 (.Y(n18191),
	.A1(n18176),
	.A2(FE_OFN26528_n23302),
	.B(FE_OFN29195_n22850));
   AOI21xp33_ASAP7_75t_L FE_RC_762_0 (.Y(n19114),
	.A1(FE_PSN8282_n21154),
	.A2(n17254),
	.B(n18746));
   AOI21xp5_ASAP7_75t_SL FE_RC_761_0 (.Y(n20395),
	.A1(FE_OFN16208_n23101),
	.A2(n17382),
	.B(n22601));
   AOI21xp5_ASAP7_75t_L FE_RC_760_0 (.Y(n22280),
	.A1(n18162),
	.A2(FE_RN_0_0),
	.B(n24694));
   AOI21xp5_ASAP7_75t_SL FE_RC_759_0 (.Y(n23716),
	.A1(n23869),
	.A2(FE_OCPN27715_n23875),
	.B(n21649));
   AOI21xp5_ASAP7_75t_SL FE_RC_758_0 (.Y(n22877),
	.A1(FE_PSN8330_n17761),
	.A2(FE_OFN28844_FE_OCPN27570_n17791),
	.B(n20978));
   AOI21xp33_ASAP7_75t_L FE_RC_757_0 (.Y(n20237),
	.A1(n19019),
	.A2(FE_OFN28752_n),
	.B(n19013));
   AOI21xp5_ASAP7_75t_L FE_RC_756_0 (.Y(n23852),
	.A1(FE_OCPN27896_n18583),
	.A2(n20617),
	.B(n21676));
   AOI21x1_ASAP7_75t_SL FE_RC_755_0 (.Y(n19894),
	.A1(n16771),
	.A2(FE_OFN28529_n16774),
	.B(FE_OCPN27508_n20339));
   AOI21x1_ASAP7_75t_L FE_RC_754_0 (.Y(n20098),
	.A1(FE_OCPN28229_n17529),
	.A2(n17560),
	.B(n20107));
   AOI31xp33_ASAP7_75t_SL FE_RC_753_0 (.Y(n22270),
	.A1(FE_OCPN27947_n18177),
	.A2(FE_OCPN27750_n22293),
	.A3(FE_OFN28688_sa22_2),
	.B(n22807));
   AOI31xp67_ASAP7_75t_SL FE_RC_752_0 (.Y(n19591),
	.A1(FE_OFN28835_n),
	.A2(n17245),
	.A3(FE_OCPN29370_FE_OFN28744),
	.B(n21453));
   OR2x2_ASAP7_75t_SL FE_RC_751_0 (.Y(n17284),
	.A(n17237),
	.B(n17236));
   INVx5_ASAP7_75t_SL FE_OFC7488_sa02_5 (.Y(FE_OCPN27566_FE_OFN16138_sa02_5),
	.A(FE_OFN16136_sa02_5));
   INVx3_ASAP7_75t_SL FE_OFC7487_sa02_5 (.Y(FE_OFN16136_sa02_5),
	.A(sa02_5_));
   INVx3_ASAP7_75t_SL FE_OFC7485_sa10_0 (.Y(FE_OFN29161_n),
	.A(FE_OCPN28145_n16535));
   INVx5_ASAP7_75t_SL FE_OFC7484_sa10_0 (.Y(FE_OCPN28145_n16535),
	.A(FE_OCPN28179_n16535));
   INVx2_ASAP7_75t_SL FE_OFC7482_sa10_0 (.Y(FE_OCPN28179_n16535),
	.A(sa10_0_));
   BUFx2_ASAP7_75t_SL FE_OFC7481_sa10_2 (.Y(FE_OFN29255_n),
	.A(FE_OFN28749_n));
   BUFx2_ASAP7_75t_SL FE_OFC7480_sa01_2 (.Y(FE_OFN29254_n),
	.A(FE_OFN28672_sa01_2));
   BUFx4f_ASAP7_75t_SL FE_OFC7477_n18536 (.Y(FE_OFN29251_n18536),
	.A(n18536));
   BUFx2_ASAP7_75t_SL FE_OFC7476_FE_OCPN27371_sa20_2 (.Y(FE_OFN29250_FE_OCPN27371_sa20_2),
	.A(FE_OCPN27371_sa20_2));
   BUFx2_ASAP7_75t_L FE_OFC7472_sa20_0 (.Y(FE_OFN29246_n),
	.A(n18522));
   BUFx2_ASAP7_75t_L FE_OFC7469_n17065 (.Y(FE_OFN29243_n17065),
	.A(n17065));
   HB1xp67_ASAP7_75t_SL FE_OFC7468_n26856 (.Y(FE_OFN29242_n26856),
	.A(n26856));
   INVx1_ASAP7_75t_L FE_OFC7467_FE_OCPN27399_n22598 (.Y(n17335),
	.A(FE_OCPN27399_n22598));
   INVx1_ASAP7_75t_R FE_OFC7466_n22811 (.Y(FE_OFN29241_n22811),
	.A(FE_OFN29237_n22811));
   INVx1_ASAP7_75t_SL FE_OFC7463_n22811 (.Y(FE_OFN29238_n22811),
	.A(FE_OFN29237_n22811));
   INVx2_ASAP7_75t_L FE_OFC7462_n22811 (.Y(FE_OFN29237_n22811),
	.A(n22811));
   HB1xp67_ASAP7_75t_R FE_OFC7460_n26631 (.Y(FE_OCPN28235_n26631),
	.A(n26631));
   INVx1_ASAP7_75t_SL FE_OFC7457_n19361 (.Y(FE_OFN26170_n19361),
	.A(FE_OCPN5143_n19361));
   BUFx6f_ASAP7_75t_L FE_OFC7456_n19361 (.Y(FE_OCPN5143_n19361),
	.A(n19361));
   INVx2_ASAP7_75t_SL FE_OFC7455_sa32_4 (.Y(FE_OFN29235_n),
	.A(FE_OFN28696_sa32_4));
   INVxp67_ASAP7_75t_SL FE_OFC7450_n16996 (.Y(n16997),
	.A(n16996));
   HB1xp67_ASAP7_75t_SL FE_OFC7446_n16875 (.Y(FE_OCPN27539_n16875),
	.A(n16875));
   INVx1_ASAP7_75t_SL FE_OFC7445_FE_RN_65_0 (.Y(n26753),
	.A(FE_RN_65_0));
   BUFx2_ASAP7_75t_L FE_OFC7444_n18631 (.Y(FE_OCPN27679_n18631),
	.A(n18631));
   INVx2_ASAP7_75t_SL FE_OFC7443_n22585 (.Y(FE_OCPN28310_n22585),
	.A(n22585));
   BUFx3_ASAP7_75t_SL FE_OFC7440_n27030 (.Y(FE_OCPN27439_n27030),
	.A(n27030));
   BUFx2_ASAP7_75t_L FE_OFC7435_n19975 (.Y(FE_OCPN27553_n19975),
	.A(n19975));
   INVx1_ASAP7_75t_L FE_OFC7434_n23999 (.Y(n16558),
	.A(n23999));
   BUFx2_ASAP7_75t_SL FE_OFC7433_n17501 (.Y(FE_OCPN27592_n17501),
	.A(n17501));
   INVx1_ASAP7_75t_R FE_OFC7431_n20345 (.Y(n24918),
	.A(n20345));
   INVx2_ASAP7_75t_SL FE_OFC7430_n18750 (.Y(FE_OCPN27843_n18750),
	.A(n18750));
   INVxp67_ASAP7_75t_SL FE_OFC7429_n26339 (.Y(FE_OCPN27535_n),
	.A(n26339));
   INVx1_ASAP7_75t_R FE_OFC7428_n25218 (.Y(FE_OFN29228_n25218),
	.A(n19366));
   INVx1_ASAP7_75t_L FE_OFC7427_n25218 (.Y(n19366),
	.A(n25218));
   INVxp67_ASAP7_75t_SL FE_OFC7426_n24510 (.Y(FE_OFN29227_n24510),
	.A(FE_OFN106_n24511));
   INVx1_ASAP7_75t_L FE_OFC7425_n24510 (.Y(FE_OFN106_n24511),
	.A(n24510));
   BUFx6f_ASAP7_75t_SL FE_OFC7422_sa23_2 (.Y(FE_OFN29191_sa23_2),
	.A(sa23_2_));
   INVxp33_ASAP7_75t_L FE_OFC7421_n22208 (.Y(FE_OFN26649_n22206),
	.A(n22208));
   INVxp67_ASAP7_75t_SL FE_OFC7417_n16793 (.Y(FE_OFN29226_n16793),
	.A(FE_OCPN27327_sa21_2));
   INVx2_ASAP7_75t_SL FE_OFC7416_n16793 (.Y(FE_OCPN27327_sa21_2),
	.A(n16793));
   BUFx6f_ASAP7_75t_SL FE_OFC7415_sa20_5 (.Y(FE_OFN29150_sa20_5),
	.A(FE_OCPN27633_sa20_5));
   BUFx6f_ASAP7_75t_SL FE_OFC7414_sa20_5 (.Y(FE_OCPN27633_sa20_5),
	.A(sa20_5_));
   INVx2_ASAP7_75t_L FE_OFC7413_n16438 (.Y(FE_OFN16430_sa33_3),
	.A(FE_OFN27062_n16438));
   BUFx3_ASAP7_75t_SL FE_OFC7408_n21479 (.Y(FE_OCPN28389_n21479),
	.A(n21479));
   HB1xp67_ASAP7_75t_SL FE_OFC7406_n23829 (.Y(FE_OCPN28432_n23829),
	.A(n23829));
   INVx1_ASAP7_75t_L FE_OFC7401_FE_OCPN28074_n27049 (.Y(FE_OFN29224_FE_OCPN28074_n27049),
	.A(FE_OFN29142_n27049));
   BUFx6f_ASAP7_75t_SL FE_OFC7399_n16748 (.Y(FE_OFN28778_FE_OCPN28352_n16748),
	.A(n16748));
   INVx1_ASAP7_75t_SL FE_OFC7398_n26632 (.Y(n26630),
	.A(n26632));
   INVx3_ASAP7_75t_SL FE_OFC7394_sa20_0 (.Y(FE_OFN31_sa20_0),
	.A(sa20_0_));
   INVx4_ASAP7_75t_SL FE_OFC7393_n17510 (.Y(n21366),
	.A(n17510));
   INVx2_ASAP7_75t_L FE_OFC7392_n16774 (.Y(FE_OFN28529_n16774),
	.A(FE_OCPN27632_n16774));
   INVx2_ASAP7_75t_SL FE_OFC7391_n16774 (.Y(FE_OCPN27632_n16774),
	.A(n16774));
   INVx1_ASAP7_75t_SL FE_OFC7390_n25751 (.Y(FE_OFN28525_n25751),
	.A(n26251));
   INVx2_ASAP7_75t_SL FE_OFC7389_n25751 (.Y(n26251),
	.A(n25751));
   INVx2_ASAP7_75t_SL FE_OFC7385_sa10_2 (.Y(FE_OFN28751_n),
	.A(FE_OFN29207_n));
   INVx1_ASAP7_75t_SL FE_OFC7384_sa10_2 (.Y(FE_OFN29207_n),
	.A(FE_OFN28749_n));
   BUFx4f_ASAP7_75t_SL FE_OFC7378_sa20_3 (.Y(n18536),
	.A(sa20_3_));
   BUFx3_ASAP7_75t_SL FE_OFC7370_n24262 (.Y(FE_OFN29215_n24262),
	.A(n24262));
   HB1xp67_ASAP7_75t_SL FE_OFC7366_n23587 (.Y(FE_OFN29211_n23587),
	.A(n23587));
   BUFx2_ASAP7_75t_L FE_OFC7365_FE_OCPN27261_sa02_0 (.Y(FE_OFN29210_FE_OCPN27261_sa02_0),
	.A(FE_OCPN27261_sa02_0));
   HB1xp67_ASAP7_75t_L FE_OFC7364_FE_OCPN27978_w3_3 (.Y(FE_OFN29209_FE_OCPN27978_w3_3),
	.A(FE_OCPN27978_w3_3));
   BUFx3_ASAP7_75t_SL FE_OFC7363_n16436 (.Y(FE_OFN29208_n16436),
	.A(n16436));
   HB1xp67_ASAP7_75t_R FE_OFC7359_sa10_2 (.Y(FE_OFN29204_sa10_2),
	.A(FE_OFN28749_n));
   BUFx2_ASAP7_75t_SL FE_OFC7355_n18521 (.Y(FE_OFN29200_n18521),
	.A(n18521));
   BUFx2_ASAP7_75t_SL FE_OFC7347_n13870 (.Y(FE_OFN29192_n13870),
	.A(n13870));
   BUFx6f_ASAP7_75t_SL FE_OFC7344_sa23_0 (.Y(FE_OFN29189_sa23_0),
	.A(sa23_0_));
   INVx1_ASAP7_75t_L FE_OFC7343_n22313 (.Y(n22812),
	.A(n22313));
   INVx1_ASAP7_75t_SL FE_OFC7341_n16783 (.Y(FE_OFN28985_sa21_5),
	.A(n16783));
   INVx1_ASAP7_75t_L FE_OFC7339_FE_OCPN27571_n20235 (.Y(FE_OFN29187_FE_OCPN27571_n20235),
	.A(FE_OFN16248_n20235));
   INVx2_ASAP7_75t_SL FE_OFC7337_FE_OCPN27571_n20235 (.Y(FE_OFN16248_n20235),
	.A(n20235));
   INVxp33_ASAP7_75t_L FE_OFC7336_FE_RN_14_0 (.Y(FE_OFN28933_n16321),
	.A(n16321));
   INVx2_ASAP7_75t_L FE_OFC7333_n17744 (.Y(FE_OFN29184_n17744),
	.A(FE_OFN28962_n17744));
   INVx2_ASAP7_75t_SL FE_OFC7330_n17744 (.Y(FE_OFN28962_n17744),
	.A(n17744));
   BUFx2_ASAP7_75t_L FE_OFC7329_n21310 (.Y(FE_OCPN28001_n21310),
	.A(n21310));
   INVxp33_ASAP7_75t_L FE_OFC7328_n25627 (.Y(n25629),
	.A(n25627));
   INVx1_ASAP7_75t_SL FE_OFC7327_n21708 (.Y(FE_OFN29182_n21708),
	.A(n21708));
   BUFx3_ASAP7_75t_SL FE_OFC7322_n16872 (.Y(FE_OCPN28127_n16872),
	.A(n16872));
   INVx1_ASAP7_75t_SL FE_OFC7319_n26165 (.Y(FE_OFN16250_n26165),
	.A(n26165));
   INVx1_ASAP7_75t_R FE_OFC7317_n24479 (.Y(FE_OFN29181_n24479),
	.A(FE_OFN28963_n24480));
   INVx2_ASAP7_75t_L FE_OFC7316_n24479 (.Y(FE_OFN28963_n24480),
	.A(n24479));
   INVx2_ASAP7_75t_SL FE_OFC7315_FE_OCPN28237_n17970 (.Y(n23587),
	.A(n17970));
   INVxp33_ASAP7_75t_R FE_OFC7313_n26222 (.Y(FE_OFN29180_n26222),
	.A(FE_OCPN27394_n26223));
   INVx1_ASAP7_75t_SL FE_OFC7312_n26222 (.Y(FE_OCPN27394_n26223),
	.A(n26222));
   INVx1_ASAP7_75t_SL FE_OFC7308_sa20_4 (.Y(FE_OFN29178_sa20_4),
	.A(FE_OFN16229_sa20_4));
   INVxp67_ASAP7_75t_SL FE_OFC7307_sa20_4 (.Y(FE_OFN29177_sa20_4),
	.A(FE_OFN16229_sa20_4));
   INVx1_ASAP7_75t_R FE_OFC7306_sa20_4 (.Y(FE_OCPN27557_sa20_4),
	.A(FE_OFN16229_sa20_4));
   INVx3_ASAP7_75t_SL FE_OFC7305_sa20_4 (.Y(FE_OFN16229_sa20_4),
	.A(sa20_4_));
   INVx1_ASAP7_75t_L FE_OFC7301_FE_OCPN28425_n18597 (.Y(FE_OFN28987_n18597),
	.A(FE_OCPN28425_n18597));
   INVx1_ASAP7_75t_L FE_OFC7300_n22024 (.Y(n26163),
	.A(n22024));
   BUFx3_ASAP7_75t_SL FE_OFC7299_n26351 (.Y(FE_OCPN27491_n26351),
	.A(n26351));
   INVx1_ASAP7_75t_L FE_OFC7298_n21755 (.Y(FE_OFN29175_n21755),
	.A(FE_RN_230_0));
   INVx1_ASAP7_75t_SL FE_OFC7296_n21755 (.Y(FE_RN_230_0),
	.A(n21755));
   INVx1_ASAP7_75t_L FE_OFC7295_n21129 (.Y(n21115),
	.A(n21129));
   INVx1_ASAP7_75t_L FE_OFC7294_sa13_2 (.Y(FE_OFN29173_n),
	.A(FE_OFN28479_sa13_2));
   INVx4_ASAP7_75t_SL FE_OFC7293_sa13_2 (.Y(FE_OFN28478_sa13_2),
	.A(FE_OFN16298_sa13_2));
   BUFx2_ASAP7_75t_L FE_OFC7291_sa13_2 (.Y(FE_OFN28479_sa13_2),
	.A(FE_OFN16298_sa13_2));
   BUFx3_ASAP7_75t_SL FE_OFC7290_sa00_4 (.Y(FE_OFN29172_sa00_4),
	.A(FE_OCPN29302_sa00_4));
   INVx1_ASAP7_75t_L FE_OFC7289_sa00_4 (.Y(n17248),
	.A(FE_OCPN29302_sa00_4));
   HB1xp67_ASAP7_75t_L FE_OFC7287_n17510 (.Y(FE_OFN29171_n17510),
	.A(n21366));
   INVxp67_ASAP7_75t_L FE_OFC7286_n17510 (.Y(FE_OFN29170_n17510),
	.A(n21366));
   INVx1_ASAP7_75t_SL FE_OFC7285_n17510 (.Y(FE_OFN29169_n17510),
	.A(n21366));
   INVx1_ASAP7_75t_L FE_OFC7283_n22585 (.Y(n18698),
	.A(FE_OCPN28310_n22585));
   INVx1_ASAP7_75t_L FE_OFC7280_n23701 (.Y(n20619),
	.A(n23701));
   INVx2_ASAP7_75t_L FE_OFC7278_n17274 (.Y(n21152),
	.A(n17274));
   INVx1_ASAP7_75t_SL FE_OFC7276_n16949 (.Y(n18133),
	.A(n16949));
   INVx1_ASAP7_75t_SL FE_OFC7274_n18536 (.Y(FE_OFN29021_sa20_3),
	.A(FE_OFN29251_n18536));
   BUFx6f_ASAP7_75t_SL FE_OFC7270_n23928 (.Y(n23633),
	.A(n23928));
   BUFx2_ASAP7_75t_SL FE_OFC7269_n18425 (.Y(FE_OCPN28141_n),
	.A(n18425));
   INVx2_ASAP7_75t_SL FE_OFC7267_n25256 (.Y(n26101),
	.A(n25256));
   INVx1_ASAP7_75t_L FE_OFC7266_n25967 (.Y(n25966),
	.A(n25967));
   INVx2_ASAP7_75t_SL FE_OFC7265_FE_OCPN27978_w3_3 (.Y(FE_OFN25886_w3_3),
	.A(FE_OCPN27978_w3_3));
   HB1xp67_ASAP7_75t_SL FE_OFC7264_n23082 (.Y(FE_OCPN28397_n23082),
	.A(n23082));
   INVx1_ASAP7_75t_SL FE_OFC7263_n23160 (.Y(FE_OFN25952_n22312),
	.A(n23160));
   BUFx3_ASAP7_75t_SL FE_OFC7262_sa33_2 (.Y(FE_OFN29164_sa33_2),
	.A(FE_OCPN29391_FE_OFN29162_sa33_2));
   INVxp67_ASAP7_75t_L FE_OFC7257_n23853 (.Y(n20623),
	.A(n23853));
   INVx3_ASAP7_75t_L FE_OFC7255_n16767 (.Y(FE_OFN28820_n),
	.A(FE_OFN25993_n16767));
   INVx2_ASAP7_75t_SL FE_OFC7254_n16767 (.Y(FE_OFN25993_n16767),
	.A(n16767));
   INVxp33_ASAP7_75t_R FE_OFC7251_n25363 (.Y(FE_OFN29160_n25363),
	.A(n25361));
   INVx1_ASAP7_75t_SL FE_OFC7250_n25363 (.Y(n25361),
	.A(n25363));
   INVx1_ASAP7_75t_L FE_OFC7249_n21892 (.Y(FE_OFN29159_n21892),
	.A(n16642));
   INVx2_ASAP7_75t_L FE_OFC7248_n21892 (.Y(n16642),
	.A(n21892));
   INVx3_ASAP7_75t_SL FE_OFC7244_n18860 (.Y(n17993),
	.A(n18860));
   BUFx2_ASAP7_75t_SL FE_OFC7243_n20841 (.Y(FE_OFN28710_n20841),
	.A(n20841));
   BUFx3_ASAP7_75t_SL FE_OFC7241_n18875 (.Y(FE_OCPN27599_n18875),
	.A(n18875));
   INVx2_ASAP7_75t_L FE_OFC7240_n19753 (.Y(FE_OFN29154_n19753),
	.A(FE_OFN29153_n19753));
   INVx1_ASAP7_75t_L FE_OFC7239_n19753 (.Y(FE_OFN29153_n19753),
	.A(n19753));
   INVx1_ASAP7_75t_L FE_OFC7236_n20327 (.Y(FE_OFN27179_n20327),
	.A(n20327));
   INVx1_ASAP7_75t_SL FE_OFC7234_n21921 (.Y(n25322),
	.A(n21921));
   INVxp67_ASAP7_75t_L FE_OFC7231_sa12_0 (.Y(FE_OFN28931_n17897),
	.A(FE_OFN29225_sa12_0));
   INVx1_ASAP7_75t_SL FE_OFC7227_n25390 (.Y(n26732),
	.A(n25390));
   INVx1_ASAP7_75t_L FE_OFC7225_n22988 (.Y(FE_OFN29151_n22988),
	.A(n20274));
   INVx1_ASAP7_75t_L FE_OFC7224_n22988 (.Y(n20274),
	.A(n22988));
   BUFx3_ASAP7_75t_SL FE_OFC7221_n17418 (.Y(FE_OCPN27666_n17418),
	.A(n17418));
   INVx2_ASAP7_75t_SL FE_OFC7219_n15376 (.Y(FE_OFN28574_n16016),
	.A(n15376));
   INVxp67_ASAP7_75t_L FE_OFC7218_n23726 (.Y(n23727),
	.A(n23726));
   INVxp67_ASAP7_75t_L FE_OFC7215_n20994 (.Y(FE_OFN97_n20994),
	.A(n20994));
   INVx1_ASAP7_75t_SL FE_OFC7214_n17756 (.Y(FE_OFN29148_n),
	.A(FE_OFN29048_n17756));
   INVx1_ASAP7_75t_SL FE_OFC7213_n17756 (.Y(FE_OFN29049_n17756),
	.A(FE_OFN29048_n17756));
   INVxp67_ASAP7_75t_L FE_OFC7210_n18969 (.Y(FE_OFN28850_FE_OCPN27840),
	.A(FE_OFN27078_sa23_5));
   INVx2_ASAP7_75t_SL FE_OFC7209_sa31_1 (.Y(FE_OFN29147_sa31_1),
	.A(FE_OFN26096_n16294));
   INVx1_ASAP7_75t_L FE_OFC7207_sa31_1 (.Y(FE_OFN29145_sa31_1),
	.A(FE_OFN26096_n16294));
   INVx2_ASAP7_75t_SL FE_OFC7206_sa31_1 (.Y(FE_OFN100_sa31_1),
	.A(FE_OFN26096_n16294));
   INVx3_ASAP7_75t_SL FE_OFC7205_sa31_1 (.Y(FE_OFN26096_n16294),
	.A(sa31_1_));
   HB1xp67_ASAP7_75t_R FE_OFC7203_n21472 (.Y(FE_OCPN28167_n21472),
	.A(n21472));
   INVxp67_ASAP7_75t_SL FE_OFC7195_n26574 (.Y(FE_OFN29141_n26574),
	.A(n26574));
   INVxp67_ASAP7_75t_L FE_OFC7194_n26574 (.Y(n26575),
	.A(n26574));
   INVx2_ASAP7_75t_SL FE_OFC7193_n18479 (.Y(FE_OFN26597_n),
	.A(n18479));
   BUFx2_ASAP7_75t_SL FE_OFC7192_n18479 (.Y(FE_OFN16200_sa30_2),
	.A(n18479));
   INVx2_ASAP7_75t_SL FE_OFC7191_n18479 (.Y(FE_OFN28895_sa30_2),
	.A(n18479));
   INVxp33_ASAP7_75t_L FE_OFC7190_n20237 (.Y(n20240),
	.A(n20237));
   BUFx6f_ASAP7_75t_SL FE_OFC7188_sa01_2 (.Y(FE_OFN28672_sa01_2),
	.A(sa01_2_));
   INVx1_ASAP7_75t_L FE_OFC7187_n23322 (.Y(n21769),
	.A(n23322));
   BUFx3_ASAP7_75t_SL FE_OFC7184_n16747 (.Y(FE_OFN16153_n16747),
	.A(n16747));
   INVx1_ASAP7_75t_L FE_OFC7183_n25384 (.Y(FE_OCPN27538_n25383),
	.A(n25384));
   INVx2_ASAP7_75t_SL FE_OFC7182_sa10_4 (.Y(FE_OCPN27636_sa10_4),
	.A(FE_OFN16150_sa10_4));
   INVx2_ASAP7_75t_SL FE_OFC7181_n20189 (.Y(n22903),
	.A(n20189));
   INVx2_ASAP7_75t_L FE_OFC7180_n19479 (.Y(FE_OFN28588_n21048),
	.A(n19479));
   BUFx2_ASAP7_75t_L FE_OFC7178_n26788 (.Y(FE_OFN154_n26788),
	.A(FE_OFN16283_n26788));
   INVx1_ASAP7_75t_L FE_OFC7177_n26178 (.Y(FE_OFN28904_n25733),
	.A(n26178));
   BUFx3_ASAP7_75t_L FE_OFC7176_n20854 (.Y(FE_OCPN28394_FE_OFN27043_n),
	.A(n20854));
   INVx1_ASAP7_75t_SL FE_OFC7175_n20854 (.Y(FE_OFN27043_n),
	.A(n20854));
   BUFx3_ASAP7_75t_SL FE_OFC7174_n26440 (.Y(FE_OFN160_n26440),
	.A(n26440));
   INVxp33_ASAP7_75t_L FE_OFC7173_n26883 (.Y(n26885),
	.A(n26883));
   INVxp67_ASAP7_75t_SL FE_OFC7172_n26172 (.Y(FE_OFN135_n26172),
	.A(FE_OCPN27373_n26172));
   BUFx3_ASAP7_75t_SL FE_OFC7171_n26172 (.Y(FE_OCPN27373_n26172),
	.A(n26172));
   INVx3_ASAP7_75t_SL FE_OFC7169_n23875 (.Y(n21639),
	.A(FE_OCPN27715_n23875));
   BUFx5_ASAP7_75t_SL FE_OFC7168_n23875 (.Y(FE_OCPN27715_n23875),
	.A(n23875));
   BUFx6f_ASAP7_75t_SL FE_OFC7167_n16758 (.Y(FE_OCPN27642_n16758),
	.A(n16758));
   BUFx2_ASAP7_75t_L FE_OFC7165_n19011 (.Y(FE_OCPN27710_n19011),
	.A(n19011));
   INVx2_ASAP7_75t_SL FE_OFC7164_n18527 (.Y(FE_OFN29140_n18527),
	.A(FE_OCPN27870_n18527));
   INVx2_ASAP7_75t_SL FE_OFC7163_n18527 (.Y(FE_OFN29139_n18527),
	.A(FE_OCPN27870_n18527));
   INVx2_ASAP7_75t_SL FE_OFC7160_n18527 (.Y(FE_OCPN27870_n18527),
	.A(n18527));
   INVx1_ASAP7_75t_L FE_OFC7159_n26362 (.Y(n26364),
	.A(FE_OCPN27744_n26362));
   INVx3_ASAP7_75t_SL FE_OFC7158_n26362 (.Y(FE_OCPN27744_n26362),
	.A(n26362));
   INVx2_ASAP7_75t_L FE_OFC7157_n21317 (.Y(FE_OFN26581_n21317),
	.A(n21317));
   INVxp67_ASAP7_75t_L FE_OFC7156_n24765 (.Y(n24766),
	.A(n24765));
   INVx2_ASAP7_75t_SL FE_OFC7155_n23359 (.Y(FE_OFN29033_FE_OCPN27414_n23359),
	.A(FE_OCPN27414_n23359));
   BUFx2_ASAP7_75t_SL FE_OFC7154_n23359 (.Y(FE_OCPN27414_n23359),
	.A(n23359));
   INVx3_ASAP7_75t_SL FE_OFC7153_FE_OCPN27228_sa11_2 (.Y(FE_OFN29137_FE_OCPN27228_sa11_2),
	.A(FE_OCPN27228_sa11_2));
   INVx3_ASAP7_75t_SL FE_OFC7150_n18164 (.Y(FE_OFN55_sa22_5),
	.A(n18164));
   INVxp67_ASAP7_75t_SL FE_OFC7149_n23968 (.Y(n23965),
	.A(n23968));
   INVx1_ASAP7_75t_L FE_OFC7148_n26427 (.Y(FE_OCPN27637_n26428),
	.A(FE_OCPN28024_n26427));
   BUFx2_ASAP7_75t_L FE_OFC7147_n26427 (.Y(FE_OCPN28024_n26427),
	.A(n26427));
   INVx1_ASAP7_75t_SL FE_OFC7142_n23884 (.Y(n18564),
	.A(n23884));
   INVx2_ASAP7_75t_SL FE_OFC7141_sa31_2 (.Y(FE_OFN29136_n),
	.A(FE_OFN28753_sa31_2));
   INVx2_ASAP7_75t_SL FE_OFC7136_n22009 (.Y(n22970),
	.A(n22009));
   INVx3_ASAP7_75t_L FE_OFC7134_n21551 (.Y(FE_OFN29135_n21551),
	.A(FE_OFN87_n21551));
   INVx1_ASAP7_75t_SL FE_OFC7133_n21551 (.Y(FE_OFN87_n21551),
	.A(n21551));
   INVx1_ASAP7_75t_SL FE_OFC7132_n21551 (.Y(FE_OFN27052_n21551),
	.A(n21551));
   INVx1_ASAP7_75t_SL FE_OFC7131_n21980 (.Y(FE_OCPN27877_n21980),
	.A(n21980));
   INVx2_ASAP7_75t_SL FE_OFC7130_n25545 (.Y(FE_OFN27065_n17059),
	.A(n25545));
   HB1xp67_ASAP7_75t_L FE_OFC7128_n26339 (.Y(FE_OCPN27534_n),
	.A(n26339));
   INVx2_ASAP7_75t_L FE_OFC7127_n24552 (.Y(FE_OFN28934_n24552),
	.A(n24553));
   INVx2_ASAP7_75t_SL FE_OFC7126_n24552 (.Y(n24553),
	.A(n24552));
   INVx2_ASAP7_75t_SL FE_OFC7121_n22206 (.Y(n22208),
	.A(n22206));
   INVx2_ASAP7_75t_SL FE_OFC7110_n19142 (.Y(n19145),
	.A(FE_OCPN4686_n19142));
   INVx2_ASAP7_75t_SL FE_OFC7109_n19142 (.Y(FE_OCPN4686_n19142),
	.A(n19142));
   INVx3_ASAP7_75t_SL FE_OFC7108_sa33_0 (.Y(FE_OFN29134_sa33_0),
	.A(FE_OFN28643_sa33_0));
   INVx2_ASAP7_75t_SL FE_OFC7103_sa33_0 (.Y(FE_OFN28643_sa33_0),
	.A(sa33_0_));
   INVx4_ASAP7_75t_SL FE_OFC7101_sa00_2 (.Y(FE_OFN28744_FE_OCPN27908),
	.A(n19821));
   INVx4_ASAP7_75t_SL FE_OFC7100_sa00_2 (.Y(FE_OCPN27908_FE_OFN16156_sa00_2),
	.A(FE_OCPN29284_n19821));
   INVx2_ASAP7_75t_SL FE_OFC7098_sa00_2 (.Y(n19821),
	.A(sa00_2_));
   HB1xp67_ASAP7_75t_R FE_OFC7097_sa03_3 (.Y(FE_OFN29122_n),
	.A(FE_OFN21730_sa03_3));
   HB1xp67_ASAP7_75t_L FE_OFC7096_sa03_3 (.Y(FE_OFN29124_n),
	.A(FE_OFN21730_sa03_3));
   INVx1_ASAP7_75t_L FE_OFC7094_n16850 (.Y(FE_OFN28995_n16850),
	.A(n18415));
   INVx1_ASAP7_75t_SL FE_OFC7093_n16850 (.Y(n18415),
	.A(n16850));
   BUFx2_ASAP7_75t_SL FE_OFC7092_n23329 (.Y(FE_OFN28966_n23329),
	.A(n23329));
   INVx3_ASAP7_75t_SL FE_OFC7091_n24767 (.Y(n22010),
	.A(FE_OFN16272_n24767));
   INVx2_ASAP7_75t_SL FE_OFC7090_n24767 (.Y(FE_OFN16272_n24767),
	.A(n24767));
   BUFx4_ASAP7_75t_SL FE_OFC7089_n21591 (.Y(FE_OFN25917_n21591),
	.A(n21591));
   INVx1_ASAP7_75t_L FE_OFC7088_n21591 (.Y(FE_OFN28790_n),
	.A(n21591));
   BUFx3_ASAP7_75t_SL FE_OFC7087_n16421 (.Y(FE_OCPN27604_n16421),
	.A(n16421));
   INVx1_ASAP7_75t_SL FE_OFC7084_sa03_0 (.Y(FE_OCPN27800_n),
	.A(sa03_0_));
   INVx1_ASAP7_75t_SL FE_OFC7078_sa10_2 (.Y(FE_OFN26039_sa10_2),
	.A(FE_OFN28749_n));
   BUFx3_ASAP7_75t_SL FE_OFC7077_FE_OCPN27371_sa20_2 (.Y(FE_OFN29131_FE_OCPN27371_sa20_2),
	.A(FE_OFN29250_FE_OCPN27371_sa20_2));
   HB1xp67_ASAP7_75t_SL FE_OFC7071_n (.Y(FE_OFN29125_n),
	.A(FE_OFN27115_n));
   BUFx4f_ASAP7_75t_SL FE_OFC7069_sa03_3 (.Y(FE_OFN29123_n),
	.A(FE_OFN21730_sa03_3));
   BUFx4f_ASAP7_75t_SL FE_OFC7067_n26026 (.Y(FE_OFN29121_n26026),
	.A(n26026));
   BUFx2_ASAP7_75t_L FE_OFC7063_n21980 (.Y(FE_OFN29117_n),
	.A(n21980));
   BUFx2_ASAP7_75t_SL FE_OFC7058_FE_OCPN27870_n18527 (.Y(FE_OFN29112_FE_OCPN27870_n18527),
	.A(FE_OFN29139_n18527));
   HB1xp67_ASAP7_75t_SL FE_OFC7055_sa03_2 (.Y(FE_OFN29109_n),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2));
   HB1xp67_ASAP7_75t_L FE_OFC7048_FE_OCPN27261_sa02_0 (.Y(FE_OFN29102_FE_OCPN27261_sa02_0),
	.A(FE_OCPN27261_sa02_0));
   BUFx2_ASAP7_75t_SL FE_OFC7047_n16418 (.Y(FE_OFN29101_n16418),
	.A(n16418));
   BUFx2_ASAP7_75t_L FE_OFC7042_n25188 (.Y(FE_OFN29096_n25188),
	.A(n25188));
   BUFx2_ASAP7_75t_SL FE_OFC7040_n21607 (.Y(FE_OFN29094_n21607),
	.A(n21607));
   HB1xp67_ASAP7_75t_L FE_OFC7037_n18525 (.Y(FE_OFN29091_n),
	.A(FE_OCPN29380_sa20_1));
   BUFx3_ASAP7_75t_SL FE_OFC7033_n25415 (.Y(FE_OFN29087_n),
	.A(FE_OFN26053_n25415));
   BUFx6f_ASAP7_75t_SL FE_OFC7027_n18526 (.Y(FE_OFN29081_n18526),
	.A(n18526));
   BUFx2_ASAP7_75t_L FE_OFC7026_n22310 (.Y(FE_OFN29080_n22310),
	.A(n22310));
   BUFx3_ASAP7_75t_SL FE_OFC7025_FE_OCPN27518_n17251 (.Y(FE_OFN29079_FE_OCPN27518_n17251),
	.A(FE_OCPN27518_n17251));
   BUFx2_ASAP7_75t_SL FE_OFC7022_n18540 (.Y(FE_OFN29076_n18540),
	.A(n18540));
   BUFx2_ASAP7_75t_SL FE_OFC7021_n22745 (.Y(FE_OFN29075_n22745),
	.A(n22745));
   HB1xp67_ASAP7_75t_SL FE_OFC7020_n17170 (.Y(FE_OFN29074_n17170),
	.A(n17170));
   HB1xp67_ASAP7_75t_R FE_OFC7012_FE_OCPN27328_sa21_2 (.Y(FE_OFN29066_FE_OCPN27328_sa21_2),
	.A(FE_OCPN27328_sa21_2));
   BUFx2_ASAP7_75t_L FE_OFC7009_n25433 (.Y(FE_OFN29063_n25433),
	.A(FE_OFN27115_n));
   BUFx3_ASAP7_75t_SL FE_OFC7008_n18651 (.Y(FE_OFN29062_n18651),
	.A(n18651));
   BUFx4f_ASAP7_75t_SL FE_OFC7007_n22505 (.Y(FE_OFN29061_n22505),
	.A(n22505));
   BUFx6f_ASAP7_75t_SL FE_OFC7000_n17453 (.Y(FE_OFN29054_n17453),
	.A(n17453));
   BUFx3_ASAP7_75t_SL FE_OFC6998_w3_5 (.Y(FE_OFN29052_w3_5),
	.A(w3_5_));
   HB1xp67_ASAP7_75t_SL FE_OFC6997_n25465 (.Y(FE_OFN29051_n25465),
	.A(n25465));
   INVx1_ASAP7_75t_SL FE_OFC6994_n17756 (.Y(FE_OFN29048_n17756),
	.A(n17756));
   INVx1_ASAP7_75t_SL FE_OFC6993_n21980 (.Y(FE_OFN29047_n21980),
	.A(FE_OCPN27877_n21980));
   INVxp67_ASAP7_75t_R FE_OFC6987_n19967 (.Y(FE_OFN29044_n19967),
	.A(n17863));
   INVx1_ASAP7_75t_L FE_OFC6986_n19967 (.Y(n17863),
	.A(n19967));
   BUFx3_ASAP7_75t_SL FE_OFC6985_FE_OCPN27696_n26027 (.Y(FE_OCPN27428_n26027),
	.A(n26027));
   INVx1_ASAP7_75t_L FE_OFC6984_n24787 (.Y(n17609),
	.A(n24787));
   HB1xp67_ASAP7_75t_SL FE_OFC6982_n25121 (.Y(FE_OCPN28169_n25121),
	.A(n25121));
   BUFx2_ASAP7_75t_SL FE_OFC6981_n19834 (.Y(FE_OCPN27500_n19834),
	.A(n19834));
   BUFx3_ASAP7_75t_SL FE_OFC6979_n17446 (.Y(FE_OCPN5021_n17446),
	.A(n17446));
   INVx1_ASAP7_75t_L FE_OFC6978_n25956 (.Y(FE_OFN28504_n25956),
	.A(FE_OFN16249_n25956));
   INVx1_ASAP7_75t_L FE_OFC6975_n25531 (.Y(n19242),
	.A(n25531));
   INVxp67_ASAP7_75t_SL FE_OFC6974_sa10_1 (.Y(FE_OFN29043_n),
	.A(FE_OFN29042_n));
   BUFx2_ASAP7_75t_L FE_OFC6972_sa10_1 (.Y(FE_OCPN28052_sa10_1),
	.A(FE_OCPN28053_sa10_1));
   INVxp33_ASAP7_75t_L FE_OFC6970_n21415 (.Y(FE_OFN29041_n21415),
	.A(n19202));
   INVx1_ASAP7_75t_SL FE_OFC6969_n21415 (.Y(n19202),
	.A(n21415));
   INVxp67_ASAP7_75t_L FE_OFC6968_n16935 (.Y(n16968),
	.A(n16935));
   INVx2_ASAP7_75t_L FE_OFC6967_n26443 (.Y(n26714),
	.A(n26443));
   INVxp33_ASAP7_75t_R FE_OFC6966_n17404 (.Y(FE_OFN29040_n17404),
	.A(FE_OFN16400_n17404));
   INVx1_ASAP7_75t_SL FE_OFC6965_n17404 (.Y(FE_OFN16400_n17404),
	.A(n17404));
   INVx1_ASAP7_75t_L FE_OFC6963_n26763 (.Y(FE_OFN29039_n26763),
	.A(n26765));
   INVx1_ASAP7_75t_SL FE_OFC6960_FE_OCPN27510_n27203 (.Y(n27201),
	.A(FE_OCPN29445_n27203));
   HB1xp67_ASAP7_75t_L FE_OFC6959_n26968 (.Y(FE_OCPN27685_n26968),
	.A(n26968));
   INVxp67_ASAP7_75t_L FE_OFC6958_n26440 (.Y(FE_OFN29037_n),
	.A(FE_OFN161_n26440));
   INVxp67_ASAP7_75t_L FE_OFC6957_n26440 (.Y(FE_OFN161_n26440),
	.A(FE_OFN160_n26440));
   BUFx2_ASAP7_75t_L FE_OFC6956_n20907 (.Y(FE_OCPN28098_n20907),
	.A(n20907));
   INVx1_ASAP7_75t_L FE_OFC6955_n27041 (.Y(FE_OFN16306_n27041),
	.A(n27041));
   INVx1_ASAP7_75t_L FE_OFC6954_n20806 (.Y(FE_OFN29036_n20806),
	.A(n20806));
   INVx1_ASAP7_75t_SL FE_OFC6952_n17116 (.Y(FE_OFN29035_n17116),
	.A(n17116));
   INVxp67_ASAP7_75t_R FE_OFC6949_FE_OCPN27414_n23359 (.Y(FE_OFN29034_FE_OCPN27414_n23359),
	.A(FE_OFN29033_FE_OCPN27414_n23359));
   BUFx2_ASAP7_75t_SL FE_OFC6947_FE_OCPN27414_n23359 (.Y(n19162),
	.A(FE_OCPN27414_n23359));
   INVx1_ASAP7_75t_SL FE_OFC6946_FE_OCPN27728_n21981 (.Y(FE_OFN29032_FE_OCPN27728_n21981),
	.A(n21981));
   INVxp33_ASAP7_75t_R FE_OFC6944_n23968 (.Y(FE_OFN29031_n23968),
	.A(n23965));
   INVxp67_ASAP7_75t_L FE_OFC6938_n19135 (.Y(FE_OFN29027_n19135),
	.A(n18653));
   INVxp67_ASAP7_75t_SL FE_OFC6936_n17077 (.Y(n17078),
	.A(n17077));
   INVx2_ASAP7_75t_L FE_OFC6935_n20911 (.Y(FE_OFN29026_n20911),
	.A(n20911));
   INVx1_ASAP7_75t_L FE_OFC6932_n27123 (.Y(FE_OFN29024_n),
	.A(n27122));
   INVx2_ASAP7_75t_L FE_OFC6930_n27123 (.Y(n27122),
	.A(FE_OFN25963_n27123));
   BUFx2_ASAP7_75t_L FE_OFC6922_sa20_3 (.Y(FE_OCPN27542_sa20_3),
	.A(FE_OFN29251_n18536));
   BUFx3_ASAP7_75t_SL FE_OFC6920_sa20_3 (.Y(FE_OCPN27580_n),
	.A(n18536));
   INVxp67_ASAP7_75t_R FE_OFC6919_n22282 (.Y(n21108),
	.A(n22282));
   INVxp33_ASAP7_75t_L FE_OFC6918_n25146 (.Y(FE_OFN29020_n25146),
	.A(n25143));
   INVxp67_ASAP7_75t_L FE_OFC6916_n25146 (.Y(n25143),
	.A(n25146));
   INVx1_ASAP7_75t_L FE_OFC6915_n15921 (.Y(FE_OFN29018_n15921),
	.A(FE_OFN29017_n15921));
   INVx2_ASAP7_75t_L FE_OFC6914_n15921 (.Y(FE_OFN29017_n15921),
	.A(n15921));
   INVx3_ASAP7_75t_L FE_OFC6912_FE_OCPN28120_n16975 (.Y(FE_OCPN28121_n16975),
	.A(FE_OCPN28120_n16975));
   INVx1_ASAP7_75t_L FE_OFC6911_n22874 (.Y(n25504),
	.A(n22874));
   INVxp67_ASAP7_75t_SL FE_OFC6909_FE_OCPN5182_n21090 (.Y(n20747),
	.A(FE_OCPN5182_n21090));
   BUFx2_ASAP7_75t_SL FE_OFC6908_n16512 (.Y(FE_OFN29016_n16512),
	.A(n16512));
   INVxp67_ASAP7_75t_L FE_OFC6906_n21246 (.Y(n21247),
	.A(n21246));
   INVxp67_ASAP7_75t_L FE_OFC6905_n26400 (.Y(FE_OFN26584_n20059),
	.A(n20059));
   INVx2_ASAP7_75t_SL FE_OFC6904_n26400 (.Y(n20059),
	.A(n26400));
   INVx1_ASAP7_75t_L FE_OFC6896_n27113 (.Y(FE_OFN29011_n27113),
	.A(FE_OFN29010_n27113));
   INVx1_ASAP7_75t_SL FE_OFC6891_n27003 (.Y(n21545),
	.A(n27003));
   INVxp67_ASAP7_75t_L FE_OFC6890_n20303 (.Y(n22677),
	.A(n20303));
   BUFx2_ASAP7_75t_L FE_OFC6888_n25351 (.Y(FE_OCPN27774_n25351),
	.A(n25351));
   INVx5_ASAP7_75t_SL FE_OFC6884_n16981 (.Y(FE_OFN16181_sa13_5),
	.A(n16981));
   INVx1_ASAP7_75t_SL FE_OFC6880_n16521 (.Y(n26045),
	.A(n16521));
   INVx1_ASAP7_75t_SL FE_OFC6879_n21225 (.Y(FE_OCPN27532_n21643),
	.A(n21225));
   INVxp33_ASAP7_75t_SL FE_OFC6878_n19733 (.Y(FE_OFN28609_n19730),
	.A(n19733));
   INVx1_ASAP7_75t_L FE_OFC6877_n23491 (.Y(FE_OFN29003_n23491),
	.A(FE_OFN28579_n23491));
   INVx1_ASAP7_75t_L FE_OFC6875_n23491 (.Y(FE_OFN29001_n23491),
	.A(FE_OFN28579_n23491));
   INVx1_ASAP7_75t_SL FE_OFC6872_n23491 (.Y(FE_OFN28579_n23491),
	.A(n23491));
   INVx1_ASAP7_75t_L FE_OFC6871_n26495 (.Y(n26496),
	.A(n26495));
   INVx1_ASAP7_75t_L FE_OFC6870_n26585 (.Y(n26587),
	.A(n26585));
   INVxp33_ASAP7_75t_L FE_OFC6869_n21395 (.Y(n19211),
	.A(n21395));
   BUFx2_ASAP7_75t_L FE_OFC6868_n18841 (.Y(FE_OCPN27937_n18841),
	.A(n18841));
   HB1xp67_ASAP7_75t_R FE_OFC6867_n18698 (.Y(FE_OFN29000_n18698),
	.A(FE_OCPN28310_n22585));
   INVx2_ASAP7_75t_L FE_OFC6865_n16923 (.Y(FE_OFN28999_n16923),
	.A(n16923));
   HB1xp67_ASAP7_75t_SL FE_OFC6863_n16923 (.Y(FE_OFN25960_n),
	.A(n16923));
   BUFx6f_ASAP7_75t_SL FE_OFC6861_sa03_4 (.Y(FE_OCPN27405_sa03_4),
	.A(sa03_4_));
   INVx1_ASAP7_75t_L FE_OFC6860_n16635 (.Y(n24967),
	.A(n16635));
   INVxp67_ASAP7_75t_L FE_OFC6857_n17464 (.Y(FE_OFN28996_n17464),
	.A(n17464));
   INVxp67_ASAP7_75t_L FE_OFC6852_n19841 (.Y(n19842),
	.A(n19841));
   INVx1_ASAP7_75t_L FE_OFC6851_FE_OCPN5176_n25870 (.Y(FE_OFN28994_FE_OCPN5176_n25870),
	.A(FE_OCPN29541_n25870));
   INVx1_ASAP7_75t_SL FE_OFC6847_FE_RN_60_0 (.Y(n26296),
	.A(FE_RN_60_0));
   INVx1_ASAP7_75t_L FE_OFC6846_n26904 (.Y(n26902),
	.A(n26904));
   INVx1_ASAP7_75t_L FE_OFC6843_n19938 (.Y(FE_OFN28991_n19938),
	.A(n18298));
   BUFx2_ASAP7_75t_SL FE_OFC6842_n19938 (.Y(n18298),
	.A(n19938));
   INVxp67_ASAP7_75t_L FE_OFC6840_n26276 (.Y(FE_OFN28990_n26276),
	.A(n26277));
   INVx1_ASAP7_75t_SL FE_OFC6838_n26276 (.Y(n26277),
	.A(n26276));
   INVx1_ASAP7_75t_SL FE_OFC6837_n26697 (.Y(n26699),
	.A(n26697));
   INVx2_ASAP7_75t_R FE_OFC6836_n18597 (.Y(FE_OFN28988_n18597),
	.A(FE_OCPN28425_n18597));
   INVx2_ASAP7_75t_L FE_OFC6834_n18597 (.Y(FE_OFN28986_n18597),
	.A(FE_OCPN28425_n18597));
   INVx2_ASAP7_75t_SL FE_OFC6833_n18597 (.Y(FE_OCPN28425_n18597),
	.A(n18597));
   BUFx4f_ASAP7_75t_SL FE_OFC6831_sa21_5 (.Y(n16783),
	.A(sa21_5_));
   INVxp67_ASAP7_75t_L FE_OFC6830_n20851 (.Y(FE_OFN28984_n20851),
	.A(n26302));
   INVx1_ASAP7_75t_SL FE_OFC6828_n20851 (.Y(n26302),
	.A(n20851));
   BUFx2_ASAP7_75t_L FE_OFC6825_n16767 (.Y(FE_OFN28981_n16767),
	.A(FE_OFN25993_n16767));
   INVxp67_ASAP7_75t_L FE_OFC6820_n18771 (.Y(n18645),
	.A(n18771));
   INVx1_ASAP7_75t_SL FE_OFC6819_n26198 (.Y(n26197),
	.A(n26198));
   INVxp67_ASAP7_75t_SL FE_OFC6818_n18169 (.Y(FE_OFN28980_n18169),
	.A(n18199));
   INVx2_ASAP7_75t_L FE_OFC6817_n18169 (.Y(n18199),
	.A(n18169));
   BUFx2_ASAP7_75t_SL FE_OFC6816_n (.Y(FE_OFN28979_n),
	.A(FE_OFN16268_sa13_3));
   INVx1_ASAP7_75t_SL FE_OFC6814_n21253 (.Y(n18570),
	.A(n21253));
   INVx2_ASAP7_75t_R FE_OFC6812_n17329 (.Y(n17382),
	.A(FE_OFN25878_n17329));
   INVxp67_ASAP7_75t_L FE_OFC6810_n15711 (.Y(n15728),
	.A(n15711));
   INVx1_ASAP7_75t_L FE_OFC6808_n15409 (.Y(FE_OFN28659_n15934),
	.A(n15409));
   BUFx2_ASAP7_75t_SL FE_OFC6806_w3_17 (.Y(FE_OFN28977_n),
	.A(FE_OFN27214_w3_17));
   HB1xp67_ASAP7_75t_L FE_OFC6805_w3_17 (.Y(FE_OFN28976_n),
	.A(FE_OFN27214_w3_17));
   BUFx2_ASAP7_75t_L FE_OFC6804_w3_17 (.Y(FE_OFN26045_n25377),
	.A(FE_OFN27214_w3_17));
   INVx1_ASAP7_75t_L FE_OFC6798_n25273 (.Y(FE_OFN28973_n25273),
	.A(FE_OCPN29387_n25273));
   INVxp67_ASAP7_75t_SL FE_OFC6796_n27021 (.Y(FE_OFN28972_n27021),
	.A(n27022));
   INVxp33_ASAP7_75t_R FE_OFC6794_n23947 (.Y(FE_OFN28971_n23947),
	.A(n25038));
   INVx1_ASAP7_75t_L FE_OFC6792_n19890 (.Y(FE_OFN28970_n19890),
	.A(FE_OFN28969_n19890));
   INVx1_ASAP7_75t_L FE_OFC6791_n19890 (.Y(FE_OFN28969_n19890),
	.A(n19890));
   INVx1_ASAP7_75t_SL FE_OFC6787_sa10_0 (.Y(FE_OFN142_sa10_0),
	.A(FE_OFN29161_n));
   INVxp67_ASAP7_75t_L FE_OFC6783_n22490 (.Y(FE_OFN28627_n21377),
	.A(FE_OFN16391_n22490));
   BUFx3_ASAP7_75t_SL FE_OFC6782_n26961 (.Y(FE_OCPN27271_n26961),
	.A(n26961));
   INVx1_ASAP7_75t_SL FE_OFC6779_n16640 (.Y(n16584),
	.A(n16640));
   BUFx2_ASAP7_75t_SL FE_OFC6777_n16497 (.Y(FE_OCPN28334_n16497),
	.A(n16497));
   INVxp67_ASAP7_75t_L FE_OFC6776_n20454 (.Y(n17641),
	.A(n20454));
   HB1xp67_ASAP7_75t_L FE_OFC6775_n25762 (.Y(FE_OCPN5119_n25762),
	.A(n25762));
   INVxp33_ASAP7_75t_L FE_OFC6774_n16248 (.Y(FE_OFN26549_n16248),
	.A(n16250));
   INVx1_ASAP7_75t_SL FE_OFC6773_n16248 (.Y(n16250),
	.A(n16248));
   INVx1_ASAP7_75t_SL FE_OFC6772_FE_OCPN5129_sa32_3 (.Y(FE_OCPN28245_n),
	.A(FE_OFN27148_sa32_3));
   INVx5_ASAP7_75t_SL FE_OFC6771_FE_OCPN5129_sa32_3 (.Y(FE_OFN27148_sa32_3),
	.A(FE_OCPN5129_sa32_3));
   INVxp67_ASAP7_75t_L FE_OFC6770_n23131 (.Y(FE_OCPN27906_n23131),
	.A(n23131));
   INVx1_ASAP7_75t_SL FE_OFC6768_n20437 (.Y(n24131),
	.A(n20437));
   INVx1_ASAP7_75t_SL FE_OFC6765_n24869 (.Y(FE_OFN28965_n24869),
	.A(n24869));
   INVxp67_ASAP7_75t_SL FE_OFC6763_n16273 (.Y(FE_OFN28964_n16273),
	.A(n16273));
   INVxp67_ASAP7_75t_SL FE_OFC6762_n16273 (.Y(n16276),
	.A(n16273));
   BUFx3_ASAP7_75t_SL FE_OFC6761_n25755 (.Y(FE_OCPN27322_n25755),
	.A(n25755));
   INVx1_ASAP7_75t_SL FE_OFC6759_n24480 (.Y(n24479),
	.A(n24480));
   INVx2_ASAP7_75t_SL FE_OFC6757_n17744 (.Y(FE_OFN28961_n17744),
	.A(FE_OFN28962_n17744));
   INVx1_ASAP7_75t_SL FE_OFC6753_n21426 (.Y(n19218),
	.A(n21426));
   INVx1_ASAP7_75t_L FE_OFC6752_n24941 (.Y(n24945),
	.A(n24941));
   INVxp67_ASAP7_75t_L FE_OFC6751_n22593 (.Y(n22186),
	.A(n22593));
   INVx1_ASAP7_75t_R FE_OFC6750_n25379 (.Y(FE_OFN28960_n25379),
	.A(n25378));
   INVx1_ASAP7_75t_L FE_OFC6748_n25379 (.Y(n25378),
	.A(n25379));
   INVx1_ASAP7_75t_SL FE_OFC6744_n22125 (.Y(FE_OCPN28027_n22125),
	.A(n22125));
   INVxp33_ASAP7_75t_R FE_OFC6743_n18011 (.Y(FE_OFN28956_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp67_ASAP7_75t_L FE_OFC6742_n18011 (.Y(FE_OFN28955_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp33_ASAP7_75t_R FE_OFC6741_n18011 (.Y(FE_OFN28954_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp33_ASAP7_75t_L FE_OFC6740_n18011 (.Y(FE_OFN28953_n18011),
	.A(FE_OCPN27285_n18011));
   INVx1_ASAP7_75t_L FE_OFC6739_n18011 (.Y(FE_OFN28952_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp67_ASAP7_75t_L FE_OFC6738_n18011 (.Y(FE_OFN28951_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp33_ASAP7_75t_L FE_OFC6737_n18011 (.Y(FE_OFN28950_n18011),
	.A(FE_OCPN27285_n18011));
   INVx1_ASAP7_75t_R FE_OFC6736_n18011 (.Y(FE_OFN28949_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp33_ASAP7_75t_R FE_OFC6735_n18011 (.Y(FE_OFN28948_n18011),
	.A(FE_OCPN27285_n18011));
   INVxp67_ASAP7_75t_L FE_OFC6734_n18011 (.Y(n21067),
	.A(FE_OCPN27285_n18011));
   INVx3_ASAP7_75t_SL FE_OFC6733_n18011 (.Y(FE_OCPN27285_n18011),
	.A(n18011));
   INVx1_ASAP7_75t_L FE_OFC6732_n26155 (.Y(n23511),
	.A(n26155));
   HB1xp67_ASAP7_75t_L FE_OFC6731_n21549 (.Y(FE_OCPN28365_n21549),
	.A(n21549));
   INVx1_ASAP7_75t_R FE_OFC6728_n23135 (.Y(FE_OFN28946_n23135),
	.A(n24958));
   INVx1_ASAP7_75t_L FE_OFC6727_n23135 (.Y(n24958),
	.A(n23135));
   INVxp67_ASAP7_75t_R FE_OFC6724_n16191 (.Y(n16192),
	.A(n16191));
   INVx1_ASAP7_75t_SL FE_OFC6723_n23498 (.Y(n20261),
	.A(n23498));
   INVx1_ASAP7_75t_L FE_OFC6722_n23265 (.Y(n24078),
	.A(n23265));
   INVx1_ASAP7_75t_SL FE_OFC6721_n19461 (.Y(n18879),
	.A(FE_OFN16294_n19461));
   INVx1_ASAP7_75t_SL FE_OFC6720_n19461 (.Y(FE_OFN16294_n19461),
	.A(n19461));
   BUFx2_ASAP7_75t_SL FE_OFC6719_n14472 (.Y(n13723),
	.A(n14472));
   INVx2_ASAP7_75t_SL FE_OFC6711_n26245 (.Y(FE_OFN26149_n26245),
	.A(FE_OFN26148_n26245));
   INVx2_ASAP7_75t_SL FE_OFC6710_n26245 (.Y(FE_OFN26148_n26245),
	.A(n26245));
   INVx2_ASAP7_75t_SL FE_OFC6709_n21456 (.Y(FE_OFN28942_n21456),
	.A(n18742));
   INVx1_ASAP7_75t_SL FE_OFC6707_n17876 (.Y(n23625),
	.A(FE_OCPN29321_n17876));
   INVx1_ASAP7_75t_SL FE_OFC6705_n26351 (.Y(n24826),
	.A(FE_OCPN27491_n26351));
   INVxp67_ASAP7_75t_R FE_OFC6703_sa02_2 (.Y(FE_OFN28941_sa02_2),
	.A(FE_OCPN29436_n22080));
   INVx1_ASAP7_75t_L FE_OFC6694_n21129 (.Y(FE_OFN28939_n21129),
	.A(n21115));
   INVx1_ASAP7_75t_L FE_OFC6691_n21015 (.Y(n21018),
	.A(n21015));
   INVx2_ASAP7_75t_SL FE_OFC6689_FE_OCPN27512_sa11_2 (.Y(FE_OCPN27229_sa11_2),
	.A(FE_OCPN27228_sa11_2));
   BUFx2_ASAP7_75t_SL FE_OFC6688_FE_OCPN27512_sa11_2 (.Y(n17473),
	.A(FE_OCPN27512_sa11_2));
   INVx4_ASAP7_75t_SL FE_OFC6687_FE_OCPN27512_sa11_2 (.Y(FE_OCPN27228_sa11_2),
	.A(FE_OCPN27512_sa11_2));
   INVx1_ASAP7_75t_L FE_OFC6686_n18104 (.Y(FE_OFN28936_n18104),
	.A(FE_OFN28935_n18104));
   INVxp67_ASAP7_75t_L FE_OFC6685_n18104 (.Y(FE_OFN28935_n18104),
	.A(n18104));
   INVx2_ASAP7_75t_SL FE_OFC6680_n26911 (.Y(FE_OFN26558_n26911),
	.A(FE_OFN28473_n26911));
   BUFx3_ASAP7_75t_SL FE_OFC6679_n26911 (.Y(FE_OFN28473_n26911),
	.A(n26911));
   INVx1_ASAP7_75t_SL FE_OFC6678_n16088 (.Y(n16087),
	.A(n16088));
   INVxp67_ASAP7_75t_SL FE_OFC6677_n20486 (.Y(FE_RN_204_0),
	.A(n20486));
   INVxp67_ASAP7_75t_L FE_OFC6675_n20563 (.Y(n17901),
	.A(n20563));
   INVx1_ASAP7_75t_L FE_OFC6672_n24713 (.Y(n24714),
	.A(n24713));
   INVx1_ASAP7_75t_SL FE_OFC6671_n19679 (.Y(n19680),
	.A(n19679));
   INVxp67_ASAP7_75t_L FE_OFC6667_n17475 (.Y(n22489),
	.A(FE_OCPN27601_n17475));
   INVxp33_ASAP7_75t_L FE_OFC6665_n22836 (.Y(FE_OFN28930_n22836),
	.A(n22839));
   INVxp67_ASAP7_75t_L FE_OFC6664_n22836 (.Y(n22839),
	.A(n22836));
   INVx1_ASAP7_75t_SL FE_OFC6663_n23677 (.Y(FE_OFN16295_n23837),
	.A(n23677));
   INVxp67_ASAP7_75t_L FE_OFC6662_n23451 (.Y(n21320),
	.A(n23451));
   INVxp33_ASAP7_75t_R FE_OFC6661_FE_OCPN27519_n25407 (.Y(n27034),
	.A(FE_OCPN27519_n25407));
   BUFx2_ASAP7_75t_SL FE_OFC6660_n20272 (.Y(FE_OCPN5191_n20272),
	.A(n20272));
   INVx1_ASAP7_75t_L FE_OFC6658_n15182 (.Y(FE_OFN28929_n15182),
	.A(FE_OFN26112_n13288));
   INVx2_ASAP7_75t_SL FE_OFC6657_n15182 (.Y(FE_OFN26111_n13288),
	.A(FE_OFN26112_n13288));
   BUFx2_ASAP7_75t_SL FE_OFC6656_n15182 (.Y(FE_OFN26112_n13288),
	.A(n15182));
   INVx1_ASAP7_75t_R FE_OFC6655_n22374 (.Y(FE_OFN28928_n22374),
	.A(FE_OFN28927_n22374));
   INVx1_ASAP7_75t_L FE_OFC6654_n22374 (.Y(FE_OFN28927_n22374),
	.A(n22374));
   BUFx2_ASAP7_75t_SL FE_OFC6647_n20449 (.Y(FE_OCPN28172_n20449),
	.A(n20449));
   INVxp67_ASAP7_75t_SL FE_OFC6644_n24877 (.Y(n24876),
	.A(n24877));
   INVx1_ASAP7_75t_L FE_OFC6639_n25912 (.Y(FE_OFN28924_n25912),
	.A(n22062));
   INVxp67_ASAP7_75t_L FE_OFC6638_n25912 (.Y(n22062),
	.A(n25912));
   BUFx3_ASAP7_75t_SL FE_OFC6637_n19573 (.Y(FE_OFN26651_n19573),
	.A(n19573));
   BUFx3_ASAP7_75t_SL FE_OFC6636_n15994 (.Y(FE_OFN109_n15994),
	.A(n15994));
   INVx1_ASAP7_75t_L FE_OFC6635_n16717 (.Y(n17398),
	.A(n16717));
   INVxp67_ASAP7_75t_L FE_OFC6634_n22095 (.Y(n22098),
	.A(n22095));
   INVx1_ASAP7_75t_R FE_OFC6633_n21873 (.Y(FE_OFN28923_n21873),
	.A(n16566));
   INVx1_ASAP7_75t_L FE_OFC6631_n21873 (.Y(n16566),
	.A(n21873));
   INVx1_ASAP7_75t_L FE_OFC6630_n20265 (.Y(n22953),
	.A(n20265));
   BUFx2_ASAP7_75t_L FE_OFC6629_w3_13 (.Y(FE_OCPN28402_w3_13),
	.A(w3_13_));
   INVx1_ASAP7_75t_SL FE_OFC6627_n25971 (.Y(n25970),
	.A(n25971));
   INVx1_ASAP7_75t_SRAM FE_OFC6626_n25284 (.Y(FE_OFN27147_n25284),
	.A(n20523));
   INVx1_ASAP7_75t_SL FE_OFC6625_n25284 (.Y(n20523),
	.A(n25284));
   INVx1_ASAP7_75t_SL FE_OFC6623_n24249 (.Y(FE_OFN28922_n24249),
	.A(n21285));
   INVx1_ASAP7_75t_L FE_OFC6622_n24249 (.Y(n21285),
	.A(n24249));
   INVxp67_ASAP7_75t_SL FE_OFC6621_n24926 (.Y(n24924),
	.A(n24926));
   INVx1_ASAP7_75t_L FE_OFC6620_n21301 (.Y(n19452),
	.A(n21301));
   INVx2_ASAP7_75t_SL FE_OFC6619_n13348 (.Y(FE_OFN28456_n13348),
	.A(n14535));
   INVx2_ASAP7_75t_SL FE_OFC6618_n13348 (.Y(n14535),
	.A(FE_OFN28454_n13348));
   INVx1_ASAP7_75t_SL FE_OFC6617_n13348 (.Y(FE_OFN28454_n13348),
	.A(n13348));
   INVxp33_ASAP7_75t_L FE_OFC6613_n20660 (.Y(FE_OFN28921_n20660),
	.A(n20662));
   INVxp67_ASAP7_75t_L FE_OFC6612_n20660 (.Y(n20662),
	.A(n20660));
   BUFx2_ASAP7_75t_SL FE_OFC6611_n27121 (.Y(FE_OCPN27641_n27121),
	.A(n27121));
   INVxp67_ASAP7_75t_L FE_OFC6610_n24254 (.Y(FE_OFN28920_n24254),
	.A(n24883));
   INVx1_ASAP7_75t_L FE_OFC6609_n24254 (.Y(n24883),
	.A(n24254));
   INVx1_ASAP7_75t_R FE_OFC6608_n24155 (.Y(FE_OFN28919_n24155),
	.A(n25872));
   INVxp67_ASAP7_75t_L FE_OFC6607_n24155 (.Y(n25872),
	.A(n24155));
   INVx1_ASAP7_75t_L FE_OFC6606_n25236 (.Y(n25235),
	.A(n25236));
   INVxp67_ASAP7_75t_L FE_OFC6605_n16949 (.Y(FE_OFN28918_n16949),
	.A(n18133));
   INVx3_ASAP7_75t_SL FE_OFC6601_sa10_4 (.Y(FE_OFN28916_sa10_4),
	.A(FE_OFN26160_sa10_4));
   INVx2_ASAP7_75t_L FE_OFC6599_sa10_4 (.Y(FE_OCPN27635_sa10_4),
	.A(FE_OFN16150_sa10_4));
   INVx3_ASAP7_75t_SL FE_OFC6598_sa10_4 (.Y(FE_OFN26160_sa10_4),
	.A(FE_OFN16150_sa10_4));
   INVx2_ASAP7_75t_SL FE_OFC6597_sa10_4 (.Y(FE_OFN26161_sa10_4),
	.A(FE_OFN16150_sa10_4));
   INVx3_ASAP7_75t_SL FE_OFC6596_sa10_4 (.Y(FE_OFN16150_sa10_4),
	.A(sa10_4_));
   INVx2_ASAP7_75t_L FE_OFC6595_sa12_2 (.Y(FE_OFN27070_n),
	.A(n22721));
   INVx1_ASAP7_75t_SL FE_OFC6594_sa12_2 (.Y(n22721),
	.A(FE_OFN25906_sa12_2));
   BUFx3_ASAP7_75t_SL FE_OFC6593_n25091 (.Y(FE_OCPN27288_n25091),
	.A(n25091));
   INVx2_ASAP7_75t_SL FE_OFC6592_FE_OCPN27633_sa20_5 (.Y(FE_OFN16368_n18545),
	.A(FE_OFN29150_sa20_5));
   INVxp67_ASAP7_75t_SL FE_OFC6591_n14245 (.Y(n14244),
	.A(n14245));
   INVx2_ASAP7_75t_SL FE_OFC6589_sa01_3 (.Y(FE_OFN26132_sa01_3),
	.A(sa01_3_));
   INVxp67_ASAP7_75t_L FE_OFC6588_n26603 (.Y(n26600),
	.A(n26603));
   INVxp33_ASAP7_75t_L FE_OFC6587_sa03_7 (.Y(FE_OFN118_sa03_7),
	.A(sa03_7_));
   INVx1_ASAP7_75t_L FE_OFC6586_FE_OCPN27241_sa11_1 (.Y(FE_OFN28915_FE_OCPN27241_sa11_1),
	.A(FE_OCPN27241_sa11_1));
   HB1xp67_ASAP7_75t_L FE_OFC6584_FE_OCPN27241_sa11_1 (.Y(FE_OCPN27866_n),
	.A(FE_OCPN27242_sa11_1));
   INVxp67_ASAP7_75t_SL FE_OFC6583_n27187 (.Y(n25237),
	.A(FE_OFN115_n27187));
   INVx1_ASAP7_75t_SL FE_OFC6582_n27187 (.Y(FE_OFN115_n27187),
	.A(n27187));
   HB1xp67_ASAP7_75t_SL FE_OFC6581_n26638 (.Y(FE_OCPN27447_n26638),
	.A(n26638));
   INVx1_ASAP7_75t_L FE_OFC6580_n26638 (.Y(n26639),
	.A(n26638));
   BUFx2_ASAP7_75t_SL FE_OFC6579_n15376 (.Y(FE_OFN26624_n15376),
	.A(FE_OFN28574_n16016));
   BUFx2_ASAP7_75t_L FE_OFC6578_n15376 (.Y(FE_OFN26131_n15376),
	.A(FE_OFN28574_n16016));
   INVx3_ASAP7_75t_L FE_OFC6577_n15376 (.Y(n16016),
	.A(FE_OFN28574_n16016));
   INVxp67_ASAP7_75t_R FE_OFC6571_n26431 (.Y(n16974),
	.A(n26431));
   BUFx3_ASAP7_75t_SL FE_OFC6570_n22293 (.Y(FE_OCPN27750_n22293),
	.A(n22293));
   INVx4_ASAP7_75t_SL FE_OFC6568_sa02_3 (.Y(n17763),
	.A(FE_OCPN27273_sa02_3));
   INVx2_ASAP7_75t_SL FE_OFC6566_sa02_3 (.Y(FE_OCPN27273_sa02_3),
	.A(sa02_3_));
   INVxp33_ASAP7_75t_L FE_OFC6565_n20007 (.Y(FE_OFN28914_n20007),
	.A(FE_OFN27140_n20007));
   INVx2_ASAP7_75t_L FE_OFC6563_n20007 (.Y(FE_OCPN27554_n20007),
	.A(n20007));
   INVx3_ASAP7_75t_L FE_OFC6562_n24292 (.Y(FE_OFN16459_n),
	.A(FE_OFN16184_w3_9));
   INVx1_ASAP7_75t_SL FE_OFC6561_n18247 (.Y(FE_OFN28913_n18247),
	.A(FE_OFN132_n18247));
   INVx1_ASAP7_75t_SL FE_OFC6559_n18247 (.Y(FE_OFN132_n18247),
	.A(n18247));
   INVx2_ASAP7_75t_L FE_OFC6557_n18015 (.Y(n23431),
	.A(n18015));
   INVx1_ASAP7_75t_L FE_OFC6552_n24229 (.Y(n24230),
	.A(n24229));
   INVxp67_ASAP7_75t_L FE_OFC6551_n18719 (.Y(n22447),
	.A(n18719));
   HB1xp67_ASAP7_75t_SL FE_OFC6550_n18767 (.Y(FE_OCPN27968_n21154),
	.A(n18767));
   INVx3_ASAP7_75t_SL FE_OFC6549_n18767 (.Y(n21154),
	.A(n18767));
   INVx1_ASAP7_75t_SL FE_OFC6544_n21475 (.Y(FE_OFN25949_n21475),
	.A(n21475));
   INVx2_ASAP7_75t_SL FE_OFC6543_n18206 (.Y(n22795),
	.A(n18206));
   INVx1_ASAP7_75t_L FE_OFC6541_n17284 (.Y(FE_OFN26644_n19599),
	.A(n17284));
   INVx4_ASAP7_75t_L FE_OFC6540_sa32_0 (.Y(FE_OFN16463_sa32_0),
	.A(FE_OCPN27812_FE_OFN16463_sa32_0));
   INVx2_ASAP7_75t_SL FE_OFC6539_sa32_0 (.Y(FE_OFN28686_FE_OCPN27812),
	.A(FE_OCPN27812_FE_OFN16463_sa32_0));
   INVx3_ASAP7_75t_SL FE_OFC6538_sa32_0 (.Y(FE_OCPN27812_FE_OFN16463_sa32_0),
	.A(sa32_0_));
   INVx1_ASAP7_75t_R FE_OFC6537_w3_23 (.Y(FE_OFN28909_w3_23),
	.A(FE_OFN37_w3_23));
   INVx1_ASAP7_75t_L FE_OFC6533_n26049 (.Y(FE_OFN28907_n26049),
	.A(FE_OCPN27770_n26049));
   INVx1_ASAP7_75t_L FE_OFC6531_n26049 (.Y(n25506),
	.A(FE_OCPN27770_n26049));
   INVx2_ASAP7_75t_SL FE_OFC6530_n26049 (.Y(FE_OCPN27770_n26049),
	.A(n26049));
   INVx2_ASAP7_75t_SL FE_OFC6528_n26922 (.Y(FE_OFN25926_n26922),
	.A(n26922));
   BUFx2_ASAP7_75t_SL FE_OFC6527_n15386 (.Y(FE_OCPN28296_n15386),
	.A(n15386));
   INVx1_ASAP7_75t_R FE_OFC6525_FE_OCPN27337_n19149 (.Y(FE_OCPN27338_n19149),
	.A(FE_OCPN29463_n));
   INVx3_ASAP7_75t_SL FE_OFC6520_sa32_4 (.Y(FE_OFN69_sa32_4),
	.A(FE_OFN16192_n17524));
   INVx4_ASAP7_75t_SL FE_OFC6519_sa32_4 (.Y(FE_OFN28696_sa32_4),
	.A(FE_OFN16192_n17524));
   INVx2_ASAP7_75t_SL FE_OFC6518_sa32_4 (.Y(FE_OFN16192_n17524),
	.A(sa32_4_));
   BUFx2_ASAP7_75t_SL FE_OFC6517_n23127 (.Y(FE_OCPN5153_n23127),
	.A(n23127));
   BUFx2_ASAP7_75t_SL FE_OFC6516_FE_OCPN27557_sa20_4 (.Y(FE_OFN28791_n),
	.A(FE_OFN29177_sa20_4));
   INVx2_ASAP7_75t_SL FE_OFC6513_n25733 (.Y(n26178),
	.A(n25733));
   INVx1_ASAP7_75t_L FE_OFC6512_n21571 (.Y(n20391),
	.A(FE_OCPN27433_n21571));
   INVx1_ASAP7_75t_L FE_OFC6511_n21571 (.Y(FE_OCPN27433_n21571),
	.A(n21571));
   BUFx2_ASAP7_75t_SL FE_OFC6510_n23252 (.Y(FE_OCPN28038_n23252),
	.A(n23252));
   INVx1_ASAP7_75t_L FE_OFC6509_n14289 (.Y(FE_OFN28600_n14289),
	.A(n14289));
   INVx1_ASAP7_75t_L FE_OFC6507_n23932 (.Y(n23933),
	.A(FE_OCPN28437_n23932));
   INVx1_ASAP7_75t_SL FE_OFC6506_n23932 (.Y(FE_OCPN28437_n23932),
	.A(n23932));
   BUFx6f_ASAP7_75t_SL FE_OFC6505_sa13_4 (.Y(FE_OFN27186_sa13_4),
	.A(sa13_4_));
   INVx1_ASAP7_75t_SL FE_OFC6504_n18666 (.Y(n22595),
	.A(n18666));
   INVx1_ASAP7_75t_SL FE_OFC6503_n13874 (.Y(FE_OCPN28404_n13874),
	.A(n13874));
   INVxp33_ASAP7_75t_L FE_OFC6500_w3_15 (.Y(FE_OFN28741_n),
	.A(FE_OFN27200_n));
   INVx4_ASAP7_75t_SL FE_OFC6496_n23322 (.Y(FE_OFN25987_n23322),
	.A(n23322));
   BUFx2_ASAP7_75t_L FE_OFC6492_sa11_5 (.Y(FE_OFN94_sa11_5),
	.A(FE_OCPN27625_sa11_5));
   HB1xp67_ASAP7_75t_L FE_OFC6488_n23417 (.Y(FE_OCPN28297_n23417),
	.A(n23417));
   BUFx3_ASAP7_75t_SL FE_OFC6487_n16980 (.Y(FE_OCPN28212_n16980),
	.A(n16980));
   INVx1_ASAP7_75t_SL FE_OFC6486_n22013 (.Y(n24218),
	.A(n22013));
   INVxp33_ASAP7_75t_L FE_OFC6485_n24836 (.Y(FE_OFN26001_n24836),
	.A(n24440));
   BUFx6f_ASAP7_75t_SL FE_OFC6473_sa31_5 (.Y(FE_OFN28669_sa31_5),
	.A(sa31_5_));
   INVxp33_ASAP7_75t_R FE_OFC6472_sa21_2 (.Y(FE_OCPN5083_sa21_2),
	.A(FE_OCPN27328_sa21_2));
   INVx2_ASAP7_75t_L FE_OFC6470_sa21_2 (.Y(FE_OCPN5126_sa21_2),
	.A(FE_OFN29226_n16793));
   BUFx4f_ASAP7_75t_SL FE_OFC6469_sa21_2 (.Y(FE_OCPN27328_sa21_2),
	.A(sa21_2_));
   INVx1_ASAP7_75t_SL FE_OFC6468_sa21_2 (.Y(n16793),
	.A(sa21_2_));
   INVx5_ASAP7_75t_SL FE_OFC6466_sa23_5 (.Y(FE_OFN27078_sa23_5),
	.A(FE_OCPN27840_FE_OFN27078_sa23_5));
   INVx2_ASAP7_75t_SL FE_OFC6463_sa23_5 (.Y(FE_OCPN27840_FE_OFN27078_sa23_5),
	.A(sa23_5_));
   INVx2_ASAP7_75t_SL FE_OFC6462_n16493 (.Y(FE_OFN26015_sa31_3),
	.A(n16493));
   INVx5_ASAP7_75t_SL FE_OFC6455_w3_11 (.Y(FE_OFN27115_n),
	.A(FE_OFN16436_w3_11));
   INVx2_ASAP7_75t_SL FE_OFC6453_w3_11 (.Y(FE_OCPN28407_FE_OFN16433_w3_11),
	.A(FE_OFN16436_w3_11));
   INVx2_ASAP7_75t_SL FE_OFC6452_w3_11 (.Y(FE_OFN16436_w3_11),
	.A(w3_11_));
   BUFx2_ASAP7_75t_L FE_OFC6450_w3_19 (.Y(FE_OFN26535_w3_19),
	.A(FE_OFN27096_n));
   BUFx2_ASAP7_75t_SL FE_OFC6449_w3_19 (.Y(FE_OFN26538_w3_19),
	.A(FE_OFN27096_n));
   INVx6_ASAP7_75t_SL FE_OFC6448_w3_19 (.Y(FE_OFN27096_n),
	.A(FE_OFN26534_w3_19));
   INVx2_ASAP7_75t_SL FE_OFC6446_w3_19 (.Y(FE_OFN26534_w3_19),
	.A(w3_19_));
   BUFx2_ASAP7_75t_L FE_OFC6444_n17603 (.Y(FE_OCPN28057_n17603),
	.A(n17603));
   INVx3_ASAP7_75t_L FE_OFC6443_n21012 (.Y(n21706),
	.A(FE_OFN28655_FE_OFN25986_n21012));
   INVx1_ASAP7_75t_L FE_OFC6442_n21012 (.Y(FE_OFN25986_n21012),
	.A(n21012));
   INVx2_ASAP7_75t_SL FE_OFC6441_n21012 (.Y(FE_OFN28655_FE_OFN25986_n21012),
	.A(n21012));
   INVx1_ASAP7_75t_L FE_OFC6438_sa30_4 (.Y(n18463),
	.A(FE_OFN16333_sa30_4));
   INVx1_ASAP7_75t_L FE_OFC6436_n23644 (.Y(FE_OCPN28299_n),
	.A(FE_OCPN28230_n23644));
   INVx3_ASAP7_75t_L FE_OFC6435_n23644 (.Y(FE_OCPN28298_n),
	.A(FE_OCPN28230_n23644));
   INVx1_ASAP7_75t_SL FE_OFC6434_n23644 (.Y(FE_OCPN28230_n23644),
	.A(n23644));
   INVx2_ASAP7_75t_R FE_OFC6433_sa01_2 (.Y(FE_OFN27152_n17315),
	.A(FE_OFN25950_sa01_2));
   INVx2_ASAP7_75t_R FE_OFC6431_sa02_5 (.Y(FE_OFN28665_FE_OCPN27566),
	.A(FE_OFN16136_sa02_5));
   INVx1_ASAP7_75t_L FE_OFC6427_n13805 (.Y(FE_OFN28898_n13805),
	.A(n14112));
   INVx2_ASAP7_75t_R FE_OFC6425_n13805 (.Y(n14112),
	.A(n13805));
   INVxp67_ASAP7_75t_L FE_OFC6423_n20132 (.Y(FE_OFN28897_n20132),
	.A(n20198));
   INVx1_ASAP7_75t_L FE_OFC6422_n20132 (.Y(n20198),
	.A(n20132));
   INVx1_ASAP7_75t_L FE_OFC6420_n23802 (.Y(FE_OFN28650_n23802),
	.A(n23802));
   INVx2_ASAP7_75t_SL FE_OFC6418_n23216 (.Y(n20796),
	.A(FE_OCPN29324_n23216));
   BUFx2_ASAP7_75t_SL FE_OFC6417_n23216 (.Y(FE_OFN27145_n23216),
	.A(FE_OCPN29324_n23216));
   INVxp67_ASAP7_75t_L FE_OFC6416_n23225 (.Y(n20575),
	.A(n23225));
   BUFx12f_ASAP7_75t_SL FE_OFC6415_sa10_3 (.Y(FE_OFN27196_n),
	.A(FE_OFN28722_sa10_3));
   INVx1_ASAP7_75t_SL FE_OFC6414_sa10_3 (.Y(FE_OCPN28323_FE_OFN16427_sa10_3),
	.A(FE_OFN28722_sa10_3));
   BUFx2_ASAP7_75t_SL FE_OFC6411_sa13_2 (.Y(FE_OFN28809_n),
	.A(FE_OFN28478_sa13_2));
   BUFx3_ASAP7_75t_SL FE_OFC6408_n26292 (.Y(FE_OCPN27516_n26292),
	.A(n26292));
   BUFx3_ASAP7_75t_SL FE_OFC6405_n22312 (.Y(n23160),
	.A(n22312));
   INVx2_ASAP7_75t_L FE_OFC6402_n14514 (.Y(FE_OFN28817_n),
	.A(n14514));
   BUFx2_ASAP7_75t_R FE_OFC6399_sa30_2 (.Y(FE_OFN28896_sa30_2),
	.A(FE_OFN28895_sa30_2));
   INVx2_ASAP7_75t_SL FE_OFC6394_sa30_2 (.Y(n18479),
	.A(sa30_2_));
   INVx1_ASAP7_75t_L FE_OFC6393_w3_22 (.Y(FE_OFN26114_n),
	.A(n24663));
   INVx4_ASAP7_75t_SL FE_OFC6392_w3_22 (.Y(FE_OFN27151_n),
	.A(n24663));
   INVx3_ASAP7_75t_SL FE_OFC6391_w3_22 (.Y(FE_OFN5_w3_22),
	.A(n24663));
   INVx5_ASAP7_75t_SL FE_OFC6390_w3_22 (.Y(n24663),
	.A(FE_OFN4_w3_22));
   BUFx2_ASAP7_75t_SL FE_OFC6389_w3_22 (.Y(FE_OFN6_w3_22),
	.A(FE_OFN4_w3_22));
   BUFx2_ASAP7_75t_R FE_OFC6388_w3_22 (.Y(FE_OCPN27987_FE_OFN4_w3_22),
	.A(FE_OFN4_w3_22));
   INVx1_ASAP7_75t_L FE_OFC6387_sa11_0 (.Y(FE_OFN28508_sa11_0),
	.A(FE_OFN28507_sa11_0));
   INVx1_ASAP7_75t_R FE_OFC6386_sa11_0 (.Y(FE_OFN138_sa11_0),
	.A(FE_OFN25879_sa11_0));
   INVx1_ASAP7_75t_R FE_OFC6383_n22945 (.Y(FE_OCPN27955_n22945),
	.A(FE_OCPN29488_FE_OFN25883_n22945));
   INVxp33_ASAP7_75t_L FE_OFC6381_n22945 (.Y(FE_OCPN27953_n22945),
	.A(FE_OFN25883_n22945));
   INVx1_ASAP7_75t_L FE_OFC6380_n19302 (.Y(FE_OFN26557_n19302),
	.A(n19302));
   INVx3_ASAP7_75t_SL FE_OFC6378_n21166 (.Y(n19609),
	.A(FE_OFN26172_n19609));
   INVx2_ASAP7_75t_L FE_OFC6377_n21166 (.Y(FE_OFN26172_n19609),
	.A(n21166));
   BUFx2_ASAP7_75t_SL FE_OFC6376_w3_6 (.Y(FE_OFN28695_n),
	.A(FE_OFN28699_w3_6));
   BUFx2_ASAP7_75t_SL FE_OFC6373_w3_14 (.Y(FE_OFN26635_w3_14),
	.A(FE_OFN8_w3_14));
   INVx1_ASAP7_75t_SL FE_OFC6372_w3_14 (.Y(FE_OFN16417_n),
	.A(FE_OFN8_w3_14));
   INVx1_ASAP7_75t_SL FE_OFC6371_sa03_1 (.Y(FE_OFN28523_sa03_1),
	.A(FE_OFN141_sa03_1));
   BUFx6f_ASAP7_75t_SL FE_OFC6370_sa03_1 (.Y(FE_OFN141_sa03_1),
	.A(sa03_1_));
   INVx5_ASAP7_75t_SL FE_OFC6369_n17526 (.Y(FE_OFN26035_n),
	.A(n17526));
   INVx1_ASAP7_75t_L FE_OFC6366_n15667 (.Y(n15301),
	.A(n15667));
   INVxp67_ASAP7_75t_L FE_OFC6365_n23328 (.Y(n20733),
	.A(FE_OCPN27933_n23328));
   INVx1_ASAP7_75t_L FE_OFC6364_n23328 (.Y(FE_OCPN27933_n23328),
	.A(n23328));
   INVx1_ASAP7_75t_L FE_OFC6358_w3_27 (.Y(FE_OFN28891_n),
	.A(FE_OFN27100_n25675));
   INVx1_ASAP7_75t_L FE_OFC6357_w3_27 (.Y(FE_OFN28890_n),
	.A(FE_OFN27100_n25675));
   INVxp67_ASAP7_75t_R FE_OFC6356_w3_27 (.Y(FE_OFN26120_n),
	.A(FE_OFN27100_n25675));
   INVx1_ASAP7_75t_SL FE_OFC6355_w3_27 (.Y(FE_OFN27100_n25675),
	.A(FE_OFN26048_w3_27));
   BUFx4f_ASAP7_75t_SL FE_OFC6354_sa31_2 (.Y(FE_OFN28719_n20025),
	.A(FE_OFN28753_sa31_2));
   INVx2_ASAP7_75t_SL FE_OFC6353_sa23_0 (.Y(n22950),
	.A(FE_OFN29189_sa23_0));
   INVx1_ASAP7_75t_SL FE_OFC6352_n15845 (.Y(FE_OFN28889_n15845),
	.A(n15787));
   INVx1_ASAP7_75t_L FE_OFC6351_n15845 (.Y(FE_OFN28792_n15787),
	.A(n15787));
   BUFx2_ASAP7_75t_SL FE_OFC6350_n15845 (.Y(n15787),
	.A(n15845));
   BUFx4f_ASAP7_75t_SL FE_OFC6347_sa03_2 (.Y(FE_OCPN5195_FE_OFN25874_sa03_2),
	.A(sa03_2_));
   INVxp33_ASAP7_75t_L FE_OFC6346_FE_OCPN27655_w3_25 (.Y(FE_OCPN27664_w3_25),
	.A(FE_OCPN27655_w3_25));
   HB1xp67_ASAP7_75t_SL FE_OFC6343_FE_OCPN27675_n17986 (.Y(FE_OFN28886_FE_OCPN27675_n17986),
	.A(FE_OCPN27675_n17986));
   BUFx2_ASAP7_75t_L FE_OFC6341_w3_14 (.Y(FE_OFN28884_n),
	.A(FE_OFN26642_w3_14));
   HB1xp67_ASAP7_75t_L FE_OFC6340_w3_14 (.Y(FE_OFN28883_n),
	.A(FE_OFN26642_w3_14));
   BUFx2_ASAP7_75t_SL FE_OFC6339_FE_OCPN27356_sa12_0 (.Y(FE_OFN28882_FE_OCPN27356_sa12_0),
	.A(FE_OFN28476_sa12_0));
   HB1xp67_ASAP7_75t_R FE_OFC6334_FE_OCPN27730_n17464 (.Y(FE_OFN28877_FE_OCPN27730_n17464),
	.A(FE_OCPN27730_n17464));
   BUFx6f_ASAP7_75t_SL FE_OFC6331_FE_OCPN27551_sa11_4 (.Y(FE_OFN28874_FE_OCPN27551_sa11_4),
	.A(FE_OCPN29504_sa11_4));
   BUFx2_ASAP7_75t_R FE_OFC6326_FE_OCPN27715_n23875 (.Y(FE_OFN28869_FE_OCPN27715_n23875),
	.A(FE_OCPN27715_n23875));
   HB1xp67_ASAP7_75t_L FE_OFC6325_FE_OCPN27715_n23875 (.Y(FE_OFN28868_FE_OCPN27715_n23875),
	.A(FE_OCPN27715_n23875));
   BUFx6f_ASAP7_75t_SL FE_OFC6319_sa13_4 (.Y(FE_OFN28862_n),
	.A(FE_OFN27186_sa13_4));
   HB1xp67_ASAP7_75t_R FE_OFC6316_FE_OCPN27664_w3_25 (.Y(FE_OFN28859_FE_OCPN27664_w3_25),
	.A(FE_OCPN27655_w3_25));
   HB1xp67_ASAP7_75t_R FE_OFC6315_FE_OCPN27664_w3_25 (.Y(FE_OFN28858_FE_OCPN27664_w3_25),
	.A(FE_OCPN27655_w3_25));
   BUFx2_ASAP7_75t_SL FE_OFC6313_n15450 (.Y(FE_OFN28856_n15450),
	.A(n15450));
   HB1xp67_ASAP7_75t_R FE_OFC6310_FE_OCPN28408_FE_OFN16433_w3_11 (.Y(FE_OFN28853_FE_OCPN28408),
	.A(FE_OCPN28408_FE_OFN16433_w3_11));
   HB1xp67_ASAP7_75t_SL FE_OFC6305_n14912 (.Y(FE_OFN28848_n14912),
	.A(n14912));
   BUFx2_ASAP7_75t_L FE_OFC6303_n26367 (.Y(FE_OFN28846_n26367),
	.A(n26367));
   BUFx2_ASAP7_75t_SL FE_OFC6301_FE_OCPN27570_n17791 (.Y(FE_OFN28844_FE_OCPN27570_n17791),
	.A(FE_OCPN27570_n17791));
   HB1xp67_ASAP7_75t_SL FE_OFC6298_n22980 (.Y(FE_OFN28841_n22980),
	.A(n22980));
   HB1xp67_ASAP7_75t_L FE_OFC6293_FE_OCPN27631_n16774 (.Y(FE_OFN28836_FE_OCPN27631_n16774),
	.A(FE_OCPN27631_n16774));
   HB1xp67_ASAP7_75t_SL FE_OFC6291_FE_OCPN28371_n17900 (.Y(FE_OFN28834_FE_OCPN28371_n17900),
	.A(FE_OCPN29559_n17900));
   BUFx2_ASAP7_75t_SL FE_OFC6289_n19789 (.Y(FE_OFN28832_n19789),
	.A(n19789));
   HB1xp67_ASAP7_75t_L FE_OFC6288_n15838 (.Y(FE_OFN28831_n15838),
	.A(n15838));
   BUFx2_ASAP7_75t_SL FE_OFC6286_n (.Y(FE_OFN28829_n),
	.A(FE_OFN26531_n));
   HB1xp67_ASAP7_75t_SL FE_OFC6284_n15683 (.Y(FE_OFN28827_n15683),
	.A(n15683));
   BUFx2_ASAP7_75t_L FE_OFC6280_n17860 (.Y(FE_OFN28823_n17860),
	.A(n17860));
   HB1xp67_ASAP7_75t_SL FE_OFC6275_n17602 (.Y(FE_OFN28818_n17602),
	.A(n17602));
   BUFx4f_ASAP7_75t_SL FE_OFC6272_n18523 (.Y(FE_OFN28815_n18523),
	.A(n18523));
   HB1xp67_ASAP7_75t_L FE_OFC6270_n15414 (.Y(FE_OFN28813_n15414),
	.A(n15414));
   HB1xp67_ASAP7_75t_L FE_OFC6269_FE_OCPN27261_sa02_0 (.Y(FE_OFN28812_FE_OCPN27261_sa02_0),
	.A(FE_OCPN27261_sa02_0));
   BUFx2_ASAP7_75t_L FE_OFC6268_n19170 (.Y(FE_OFN28811_n19170),
	.A(n19170));
   HB1xp67_ASAP7_75t_L FE_OFC6265_n26291 (.Y(FE_OFN28808_n26291),
	.A(n26291));
   INVx1_ASAP7_75t_SL FE_OFC6264_n24944 (.Y(FE_OFN28807_n24944),
	.A(FE_OFN28806_n24944));
   INVx1_ASAP7_75t_L FE_OFC6263_n24944 (.Y(FE_OFN28806_n24944),
	.A(n24944));
   BUFx6f_ASAP7_75t_SL FE_OFC6258_n16978 (.Y(FE_OFN28801_n16978),
	.A(n16978));
   BUFx3_ASAP7_75t_SL FE_OFC6257_n22526 (.Y(FE_OFN28800_n22526),
	.A(n22526));
   HB1xp67_ASAP7_75t_L FE_OFC6255_FE_OCPN27947_n18177 (.Y(FE_OFN28798_FE_OCPN27947_n18177),
	.A(FE_OCPN27947_n18177));
   BUFx2_ASAP7_75t_L FE_OFC6253_n17301 (.Y(FE_OFN28796_n17301),
	.A(n17301));
   HB1xp67_ASAP7_75t_R FE_OFC6244_n19000 (.Y(FE_OFN28787_n19000),
	.A(n19000));
   HB1xp67_ASAP7_75t_L FE_OFC6240_n26099 (.Y(FE_OFN28783_n26099),
	.A(n26099));
   BUFx6f_ASAP7_75t_SL FE_OFC6236_n24257 (.Y(FE_OFN28779_n24257),
	.A(n24257));
   HB1xp67_ASAP7_75t_L FE_OFC6233_n18532 (.Y(FE_OFN28776_n18532),
	.A(n18532));
   BUFx2_ASAP7_75t_L FE_OFC6232_n16992 (.Y(FE_OFN28775_n16992),
	.A(n16992));
   HB1xp67_ASAP7_75t_L FE_OFC6228_sa33_3 (.Y(FE_OFN28771_n),
	.A(FE_OFN25938_sa33_3));
   BUFx2_ASAP7_75t_SL FE_OFC6226_n15478 (.Y(FE_OFN28769_n15478),
	.A(n15478));
   BUFx2_ASAP7_75t_R FE_OFC6215_n15422 (.Y(FE_OFN28758_n15422),
	.A(n15422));
   BUFx3_ASAP7_75t_L FE_OFC6209_n22995 (.Y(FE_OFN28752_n),
	.A(FE_OFN27056_n22995));
   BUFx2_ASAP7_75t_R FE_OFC6204_w3_6 (.Y(FE_OFN28747_n),
	.A(FE_OCPN29537_FE_OFN28699_w3_6));
   BUFx3_ASAP7_75t_SL FE_OFC6196_n17898 (.Y(FE_OFN28739_n17898),
	.A(n17898));
   BUFx3_ASAP7_75t_SL FE_OFC6189_w3_1 (.Y(FE_OFN28732_n),
	.A(FE_OFN26058_w3_1));
   BUFx3_ASAP7_75t_SL FE_OFC6187_FE_OCPN28416_sa02_3 (.Y(FE_OFN28730_FE_OCPN28416_sa02_3),
	.A(n17763));
   HB1xp67_ASAP7_75t_L FE_OFC6186_n20617 (.Y(FE_OFN28729_n20617),
	.A(n20617));
   BUFx6f_ASAP7_75t_SL FE_OFC6184_sa33_1 (.Y(FE_OFN28727_sa33_1),
	.A(sa33_1_));
   HB1xp67_ASAP7_75t_SL FE_OFC6180_n22750 (.Y(FE_OFN28723_n22750),
	.A(n22750));
   BUFx6f_ASAP7_75t_SL FE_OFC6179_sa10_3 (.Y(FE_OFN28722_sa10_3),
	.A(sa10_3_));
   BUFx2_ASAP7_75t_SRAM FE_OFC6178_n (.Y(FE_OFN28721_n),
	.A(FE_OFN28699_w3_6));
   BUFx3_ASAP7_75t_SL FE_OFC6175_sa01_1 (.Y(FE_OFN28718_sa01_1),
	.A(sa01_1_));
   HB1xp67_ASAP7_75t_L FE_OFC6174_n15158 (.Y(FE_OFN28717_n15158),
	.A(n15158));
   INVxp67_ASAP7_75t_L FE_OFC6172_w3_15 (.Y(FE_OFN28715_w3_15),
	.A(FE_OFN28741_n));
   INVxp67_ASAP7_75t_R FE_OFC6170_w3_20 (.Y(FE_OFN28713_n),
	.A(FE_OFN28711_n));
   INVx3_ASAP7_75t_SL FE_OFC6169_w3_20 (.Y(FE_OFN28712_n),
	.A(FE_OFN28711_n));
   INVx1_ASAP7_75t_L FE_OFC6168_w3_20 (.Y(FE_OFN28711_n),
	.A(FE_OFN25909_w3_20));
   BUFx4_ASAP7_75t_SL FE_OFC6163_n25377 (.Y(FE_OFN28706_n),
	.A(FE_OFN26041_w3_17));
   HB1xp67_ASAP7_75t_L FE_OFC6161_FE_OCPN27740_sa02_4 (.Y(FE_OFN28704_FE_OCPN27740_sa02_4),
	.A(n17760));
   BUFx2_ASAP7_75t_L FE_OFC6160_FE_OCPN27740_sa02_4 (.Y(FE_OFN28703_FE_OCPN27740_sa02_4),
	.A(n17760));
   BUFx2_ASAP7_75t_SL FE_OFC6158_w3_16 (.Y(FE_OFN28701_w3_16),
	.A(w3_16_));
   BUFx4f_ASAP7_75t_SL FE_OFC6156_w3_6 (.Y(FE_OFN28699_w3_6),
	.A(w3_6_));
   BUFx6f_ASAP7_75t_SL FE_OFC6151_sa33_4 (.Y(FE_OFN28694_sa33_4),
	.A(sa33_4_));
   BUFx2_ASAP7_75t_L FE_OFC6148_n13725 (.Y(FE_OFN28691_n13725),
	.A(n13725));
   BUFx2_ASAP7_75t_L FE_OFC6147_n25979 (.Y(FE_OFN28690_n25979),
	.A(n25979));
   BUFx6f_ASAP7_75t_SL FE_OFC6146_sa03_5 (.Y(FE_OFN28689_sa03_5),
	.A(sa03_5_));
   BUFx6f_ASAP7_75t_SL FE_OFC6145_sa22_2 (.Y(FE_OFN28688_sa22_2),
	.A(sa22_2_));
   BUFx3_ASAP7_75t_SL FE_OFC6140_w3_21 (.Y(FE_OFN28683_w3_21),
	.A(w3_21_));
   HB1xp67_ASAP7_75t_SL FE_OFC6139_n15888 (.Y(FE_OFN28682_n15888),
	.A(n15888));
   BUFx3_ASAP7_75t_SL FE_OFC6137_sa22_5 (.Y(FE_OFN28680_n),
	.A(FE_OFN55_sa22_5));
   BUFx6f_ASAP7_75t_SL FE_OFC6135_sa21_3 (.Y(FE_OFN28678_sa21_3),
	.A(sa21_3_));
   BUFx2_ASAP7_75t_SL FE_OFC6134_n17998 (.Y(FE_OFN28677_n17998),
	.A(n17998));
   INVxp67_ASAP7_75t_L FE_OFC6131_n25377 (.Y(FE_OFN28674_n),
	.A(FE_OFN28673_n));
   INVxp67_ASAP7_75t_R FE_OFC6130_n25377 (.Y(FE_OFN28673_n),
	.A(FE_OFN28706_n));
   BUFx2_ASAP7_75t_L FE_OFC6128_FE_OCPN28076_FE_OFN9_w3_6 (.Y(FE_OFN28671_FE_OCPN28076),
	.A(FE_OCPN28076_FE_OFN9_w3_6));
   INVx2_ASAP7_75t_SL FE_OFC6119_w3_7 (.Y(FE_OFN28662_w3_7),
	.A(FE_OFN28660_w3_7));
   INVx2_ASAP7_75t_L FE_OFC6118_w3_7 (.Y(FE_OFN28661_w3_7),
	.A(FE_OFN28660_w3_7));
   INVx1_ASAP7_75t_SL FE_OFC6117_w3_7 (.Y(FE_OFN28660_w3_7),
	.A(w3_7_));
   INVxp67_ASAP7_75t_L FE_OFC6116_n23311 (.Y(FE_OFN25941_n22857),
	.A(n23311));
   INVxp67_ASAP7_75t_L FE_OFC6115_n25200 (.Y(n25203),
	.A(n25200));
   INVxp33_ASAP7_75t_R FE_OFC6114_FE_OCPN28321_n21341 (.Y(n26068),
	.A(FE_OCPN28321_n21341));
   INVx1_ASAP7_75t_SL FE_OFC6113_n21731 (.Y(n19466),
	.A(n21731));
   HB1xp67_ASAP7_75t_R FE_OFC6112_n25769 (.Y(FE_OCPN27815_n25769),
	.A(n25769));
   INVx1_ASAP7_75t_L FE_OFC6111_n25438 (.Y(n23604),
	.A(n25438));
   INVxp67_ASAP7_75t_R FE_OFC6110_n23298 (.Y(n21780),
	.A(n23298));
   INVxp33_ASAP7_75t_L FE_OFC6109_n19806 (.Y(FE_OFN16202_n19806),
	.A(n24669));
   INVxp33_ASAP7_75t_R FE_OFC6106_n15934 (.Y(FE_OFN28658_n15934),
	.A(n15934));
   INVx1_ASAP7_75t_L FE_OFC6104_n15934 (.Y(n15409),
	.A(n15934));
   INVxp67_ASAP7_75t_L FE_OFC6102_FE_OFN25986_n21012 (.Y(FE_OFN28656_FE_OFN25986_n21012),
	.A(n21706));
   INVx1_ASAP7_75t_L FE_OFC6098_n22751 (.Y(FE_OFN28654_n22751),
	.A(FE_OFN122_n22751));
   INVx1_ASAP7_75t_L FE_OFC6096_n22751 (.Y(FE_OFN122_n22751),
	.A(n22751));
   INVxp33_ASAP7_75t_L FE_OFC6094_n21642 (.Y(FE_OFN28652_n21642),
	.A(n18605));
   INVx1_ASAP7_75t_R FE_OFC6093_n21642 (.Y(n18605),
	.A(n21642));
   INVxp67_ASAP7_75t_R FE_OFC6092_FE_OFN26140_n23585 (.Y(FE_OFN28651_FE_OFN26140_n23585),
	.A(FE_OFN26140_n23585));
   INVxp33_ASAP7_75t_L FE_OFC6089_n23802 (.Y(FE_OFN28649_n23802),
	.A(FE_OFN28650_n23802));
   INVxp33_ASAP7_75t_R FE_OFC6086_n23549 (.Y(FE_OFN28648_n23549),
	.A(n16727));
   INVx1_ASAP7_75t_L FE_OFC6085_n23549 (.Y(n16727),
	.A(n23549));
   INVxp67_ASAP7_75t_R FE_OFC6084_n21764 (.Y(FE_OFN28647_n21764),
	.A(n21764));
   INVx1_ASAP7_75t_R FE_OFC6078_n15950 (.Y(FE_OFN16348_n15949),
	.A(n15950));
   INVxp67_ASAP7_75t_L FE_OFC6077_n17398 (.Y(FE_OFN16369_n16717),
	.A(n17398));
   HB1xp67_ASAP7_75t_SL FE_OFC6066_n15240 (.Y(FE_OFN16206_n15240),
	.A(n15240));
   INVx2_ASAP7_75t_SL FE_OFC6065_n15240 (.Y(n14504),
	.A(n15240));
   INVx1_ASAP7_75t_L FE_OFC6063_n25102 (.Y(FE_OFN28637_n25102),
	.A(FE_OCPN27829_n25102));
   INVxp33_ASAP7_75t_R FE_OFC6059_n24010 (.Y(n24011),
	.A(n24010));
   INVx1_ASAP7_75t_L FE_OFC6058_n21034 (.Y(FE_OFN28635_n21034),
	.A(n19492));
   INVx1_ASAP7_75t_R FE_OFC6056_n21034 (.Y(n19492),
	.A(n21034));
   INVxp33_ASAP7_75t_L FE_OFC6055_n17716 (.Y(FE_OFN28633_n17716),
	.A(n17723));
   INVx1_ASAP7_75t_R FE_OFC6054_n17716 (.Y(n17723),
	.A(n17716));
   BUFx2_ASAP7_75t_L FE_OFC6052_n20988 (.Y(FE_OCPN27972_n20988),
	.A(n20988));
   INVx1_ASAP7_75t_L FE_OFC6049_n20460 (.Y(n20462),
	.A(n20460));
   INVxp33_ASAP7_75t_L FE_OFC6048_n19087 (.Y(FE_OFN25980_n19087),
	.A(n21167));
   INVx1_ASAP7_75t_SL FE_OFC6047_n19087 (.Y(n21167),
	.A(n19087));
   INVxp33_ASAP7_75t_L FE_OFC6046_n18437 (.Y(FE_RN_191_0),
	.A(n18437));
   BUFx2_ASAP7_75t_SL FE_OFC6045_n26860 (.Y(FE_OCPN27375_n26860),
	.A(n26860));
   INVxp67_ASAP7_75t_R FE_OFC6044_n23385 (.Y(FE_OFN28630_n23385),
	.A(n23386));
   INVx1_ASAP7_75t_L FE_OFC6042_n23385 (.Y(n23386),
	.A(n23385));
   INVx1_ASAP7_75t_L FE_OFC6041_n15667 (.Y(FE_OFN28628_n15667),
	.A(n15301));
   INVx1_ASAP7_75t_R FE_OFC6037_n21377 (.Y(FE_OFN16391_n22490),
	.A(n21377));
   INVxp33_ASAP7_75t_R FE_OFC6036_n22094 (.Y(FE_OFN28626_n22094),
	.A(FE_OFN27058_n22094));
   INVx1_ASAP7_75t_SL FE_OFC6035_n22094 (.Y(FE_OFN25998_n17781),
	.A(FE_OFN27058_n22094));
   INVx5_ASAP7_75t_SL FE_OFC6034_n22094 (.Y(FE_OFN27058_n22094),
	.A(n22094));
   INVxp33_ASAP7_75t_L FE_OFC6033_n26101 (.Y(FE_OFN28625_n26101),
	.A(FE_OFN30_n25256));
   INVx1_ASAP7_75t_R FE_OFC6032_n26101 (.Y(FE_OFN30_n25256),
	.A(n26101));
   INVx1_ASAP7_75t_L FE_OFC6031_n13874 (.Y(FE_OFN28624_n13874),
	.A(FE_OCPN28404_n13874));
   BUFx2_ASAP7_75t_L FE_OFC6030_n13874 (.Y(FE_OFN28623_n13874),
	.A(n13874));
   INVx1_ASAP7_75t_L FE_OFC6027_n25870 (.Y(FE_OFN28622_n25870),
	.A(FE_OFN28994_FE_OCPN5176_n25870));
   INVxp33_ASAP7_75t_R FE_OFC6021_n20437 (.Y(FE_OFN28619_n20437),
	.A(n24131));
   INVx1_ASAP7_75t_R FE_OFC6018_n25322 (.Y(FE_OFN28618_n25322),
	.A(FE_OCPN27817_n21921));
   INVxp67_ASAP7_75t_L FE_OFC6016_n25322 (.Y(FE_OCPN27817_n21921),
	.A(n25322));
   BUFx2_ASAP7_75t_L FE_OFC6015_n21396 (.Y(FE_OCPN28417_n21396),
	.A(n21396));
   INVxp33_ASAP7_75t_R FE_OFC6013_n26191 (.Y(FE_OFN28616_n26191),
	.A(FE_OCPN27583_n26193));
   INVx1_ASAP7_75t_SL FE_OFC6012_n26191 (.Y(FE_OFN28615_n26191),
	.A(FE_OCPN27583_n26193));
   BUFx2_ASAP7_75t_SL FE_OFC6010_n20169 (.Y(FE_OCPN27634_n20169),
	.A(n20169));
   INVx1_ASAP7_75t_R FE_OFC6009_n21715 (.Y(FE_OFN28614_n21715),
	.A(n19450));
   INVx1_ASAP7_75t_L FE_OFC6005_n21715 (.Y(n19450),
	.A(n21715));
   INVx1_ASAP7_75t_SL FE_OFC6004_FE_RN_53_0 (.Y(n26294),
	.A(FE_RN_53_0));
   INVx1_ASAP7_75t_SL FE_OFC6003_n22125 (.Y(FE_OFN28610_n22125),
	.A(FE_OCPN28027_n22125));
   INVxp33_ASAP7_75t_L FE_OFC6000_n21204 (.Y(n18528),
	.A(n21204));
   INVxp67_ASAP7_75t_R FE_OFC5999_n22838 (.Y(n23337),
	.A(n22838));
   INVx1_ASAP7_75t_SL FE_OFC5997_n16761 (.Y(n23926),
	.A(n16761));
   INVx1_ASAP7_75t_SL FE_OFC5994_n19730 (.Y(n19733),
	.A(n19730));
   INVx1_ASAP7_75t_L FE_OFC5993_n21027 (.Y(FE_OFN28608_n21027),
	.A(n21027));
   INVxp33_ASAP7_75t_L FE_OFC5991_n24220 (.Y(n17343),
	.A(n24220));
   INVx1_ASAP7_75t_R FE_OFC5990_FE_RN_54_0 (.Y(n17272),
	.A(n18656));
   INVx2_ASAP7_75t_SL FE_OFC5989_FE_RN_54_0 (.Y(n18656),
	.A(FE_RN_54_0));
   INVxp67_ASAP7_75t_R FE_OFC5988_n23884 (.Y(FE_OFN28607_n23884),
	.A(n18564));
   INVxp67_ASAP7_75t_L FE_OFC5985_n21107 (.Y(n21782),
	.A(n21107));
   INVxp33_ASAP7_75t_L FE_OFC5984_n17854 (.Y(n17859),
	.A(n17854));
   INVxp33_ASAP7_75t_L FE_OFC5983_n25737 (.Y(n25747),
	.A(n25737));
   INVxp67_ASAP7_75t_SL FE_OFC5982_n23949 (.Y(FE_OFN28605_n23949),
	.A(n16646));
   INVx1_ASAP7_75t_SL FE_OFC5981_n23949 (.Y(FE_OCPN27900_n23949),
	.A(n16646));
   INVx1_ASAP7_75t_SL FE_OFC5980_n23949 (.Y(n16646),
	.A(n23949));
   INVx1_ASAP7_75t_L FE_OFC5979_n27010 (.Y(FE_OFN16307_n27010),
	.A(n22579));
   INVx1_ASAP7_75t_L FE_OFC5978_n27010 (.Y(n22579),
	.A(n27010));
   BUFx2_ASAP7_75t_SL FE_OFC5975_n14534 (.Y(FE_OFN28604_n14534),
	.A(FE_OFN28602_n14534));
   INVx1_ASAP7_75t_SL FE_OFC5974_n14534 (.Y(FE_OFN28603_n14534),
	.A(FE_OFN28602_n14534));
   INVx1_ASAP7_75t_L FE_OFC5973_n14534 (.Y(FE_OFN28602_n14534),
	.A(n14534));
   INVx1_ASAP7_75t_SL FE_OFC5969_n21090 (.Y(FE_OCPN5182_n21090),
	.A(n21090));
   INVx1_ASAP7_75t_R FE_OFC5967_n23588 (.Y(FE_OFN85_n23588),
	.A(n23588));
   INVx2_ASAP7_75t_SL FE_OFC5965_n16773 (.Y(n23668),
	.A(n16773));
   INVxp33_ASAP7_75t_L FE_OFC5964_n20497 (.Y(FE_RN_63_0),
	.A(n20497));
   INVxp67_ASAP7_75t_L FE_OFC5963_n20212 (.Y(n20213),
	.A(n20212));
   INVxp33_ASAP7_75t_L FE_OFC5962_n22704 (.Y(n22705),
	.A(n22704));
   INVx1_ASAP7_75t_R FE_OFC5960_n25082 (.Y(n21620),
	.A(n25082));
   INVxp33_ASAP7_75t_L FE_OFC5959_n22631 (.Y(n22651),
	.A(n22631));
   INVxp67_ASAP7_75t_L FE_OFC5958_n13596 (.Y(FE_OFN27044_n15236),
	.A(n13596));
   BUFx2_ASAP7_75t_SL FE_OFC5955_n14289 (.Y(FE_OFN16352_n14289),
	.A(n14289));
   INVxp67_ASAP7_75t_L FE_OFC5951_n22156 (.Y(n17659),
	.A(n22156));
   INVx1_ASAP7_75t_SL FE_OFC5950_n23018 (.Y(n23989),
	.A(n23018));
   INVx2_ASAP7_75t_L FE_OFC5949_n19817 (.Y(FE_OFN26146_n18774),
	.A(n19817));
   INVxp33_ASAP7_75t_R FE_OFC5948_n20933 (.Y(FE_OFN28598_n20933),
	.A(FE_OCPN29331_n20933));
   INVx1_ASAP7_75t_SL FE_OFC5946_n23583 (.Y(n19555),
	.A(n23583));
   INVx3_ASAP7_75t_SL FE_OFC5943_FE_RN_222_0 (.Y(n15729),
	.A(FE_RN_222_0));
   INVxp67_ASAP7_75t_R FE_OFC5942_n23948 (.Y(FE_OFN28596_n23948),
	.A(n23948));
   INVx1_ASAP7_75t_L FE_OFC5940_n16361 (.Y(FE_OFN27168_n16334),
	.A(n16361));
   BUFx2_ASAP7_75t_SL FE_OFC5938_n22776 (.Y(FE_OCPN28198_n22776),
	.A(n22776));
   INVxp33_ASAP7_75t_L FE_OFC5937_n20189 (.Y(FE_OFN28595_n20189),
	.A(n22903));
   INVxp67_ASAP7_75t_R FE_OFC5935_n24102 (.Y(FE_OFN16392_n24102),
	.A(n24517));
   INVx1_ASAP7_75t_L FE_OFC5934_n24102 (.Y(n24517),
	.A(n24102));
   BUFx2_ASAP7_75t_SL FE_OFC5933_n26454 (.Y(FE_OFN28594_n26454),
	.A(n26454));
   BUFx3_ASAP7_75t_SL FE_OFC5932_n26454 (.Y(FE_OCPN27988_n26454),
	.A(n26454));
   INVxp33_ASAP7_75t_R FE_OFC5931_n18627 (.Y(FE_OFN28593_n18627),
	.A(n24084));
   INVx1_ASAP7_75t_L FE_OFC5930_n18627 (.Y(n24084),
	.A(n18627));
   HB1xp67_ASAP7_75t_SL FE_OFC5929_n16427 (.Y(FE_OFN28592_n16427),
	.A(n16427));
   INVx1_ASAP7_75t_SL FE_OFC5926_n24062 (.Y(FE_OFN26588_n24062),
	.A(n24062));
   BUFx2_ASAP7_75t_L FE_OFC5925_n20176 (.Y(FE_OCPN27652_n20176),
	.A(n20176));
   INVx2_ASAP7_75t_SL FE_OFC5924_FE_RN_229_0 (.Y(n25395),
	.A(FE_RN_229_0));
   INVx1_ASAP7_75t_R FE_OFC5922_n21557 (.Y(n18696),
	.A(n21557));
   INVxp67_ASAP7_75t_R FE_OFC5921_n24391 (.Y(FE_OFN28590_n24391),
	.A(n18722));
   INVx1_ASAP7_75t_SL FE_OFC5920_n24391 (.Y(n18722),
	.A(n24391));
   INVx1_ASAP7_75t_L FE_OFC5919_n15239 (.Y(FE_OFN27061_n15239),
	.A(n15239));
   HB1xp67_ASAP7_75t_R FE_OFC5918_n15239 (.Y(n14516),
	.A(n15239));
   INVx1_ASAP7_75t_SL FE_OFC5917_n23761 (.Y(n21197),
	.A(n23761));
   INVxp67_ASAP7_75t_L FE_OFC5916_n15002 (.Y(n15004),
	.A(n15002));
   INVxp67_ASAP7_75t_L FE_OFC5915_n20096 (.Y(n17578),
	.A(n20096));
   INVxp67_ASAP7_75t_R FE_OFC5914_n24368 (.Y(n24371),
	.A(n24368));
   INVxp33_ASAP7_75t_R FE_OFC5913_n27041 (.Y(FE_OFN26147_n27041),
	.A(FE_OFN16306_n27041));
   INVxp67_ASAP7_75t_R FE_OFC5910_n23490 (.Y(n22936),
	.A(n23490));
   INVxp67_ASAP7_75t_L FE_OFC5909_n25750 (.Y(FE_OFN16375_n25750),
	.A(FE_OCPN8229_n25750));
   BUFx2_ASAP7_75t_L FE_OFC5906_n21042 (.Y(FE_OCPN27918_n21042),
	.A(n21042));
   INVx1_ASAP7_75t_L FE_OFC5905_FE_OCPN27274_n26394 (.Y(n24514),
	.A(FE_OCPN27274_n26394));
   INVxp33_ASAP7_75t_L FE_OFC5904_n26084 (.Y(n21417),
	.A(FE_OFN16351_n26084));
   INVx1_ASAP7_75t_SL FE_OFC5903_n26084 (.Y(FE_OFN16351_n26084),
	.A(n26084));
   INVx2_ASAP7_75t_L FE_OFC5902_n21048 (.Y(FE_OFN28589_n21048),
	.A(FE_OFN28588_n21048));
   INVx1_ASAP7_75t_L FE_OFC5898_n21048 (.Y(n19479),
	.A(n21048));
   INVxp33_ASAP7_75t_R FE_OFC5897_FE_OCPN28230_n23644 (.Y(n22706),
	.A(FE_OCPN28299_n));
   INVx1_ASAP7_75t_R FE_OFC5896_n24692 (.Y(n24695),
	.A(n24692));
   INVxp33_ASAP7_75t_L FE_OFC5895_n24736 (.Y(FE_OFN28586_n24736),
	.A(n24737));
   INVxp67_ASAP7_75t_L FE_OFC5893_n24736 (.Y(n24737),
	.A(n24736));
   INVx1_ASAP7_75t_L FE_OFC5892_n17001 (.Y(FE_OFN28584_n17001),
	.A(FE_OCPN29490_n17001));
   INVxp33_ASAP7_75t_L FE_OFC5889_n22453 (.Y(FE_RN_232_0),
	.A(n22453));
   INVx1_ASAP7_75t_R FE_OFC5888_n23449 (.Y(n21024),
	.A(n23449));
   INVxp67_ASAP7_75t_L FE_OFC5887_n25657 (.Y(FE_OFN28582_n25657),
	.A(n25657));
   INVx1_ASAP7_75t_L FE_OFC5885_n19044 (.Y(n17619),
	.A(n19044));
   INVx1_ASAP7_75t_L FE_OFC5881_n19893 (.Y(n23662),
	.A(n19893));
   INVxp33_ASAP7_75t_L FE_OFC5880_n23451 (.Y(FE_OCPN5072_n23451),
	.A(n21320));
   BUFx2_ASAP7_75t_L FE_OFC5878_n15106 (.Y(FE_OFN26084_n15106),
	.A(n15813));
   INVxp67_ASAP7_75t_SL FE_OFC5877_n15106 (.Y(FE_OFN25918_n15813),
	.A(n15813));
   INVxp67_ASAP7_75t_L FE_OFC5876_FE_OFN16246_n16113 (.Y(FE_OFN26121_n16107),
	.A(FE_OFN16246_n16113));
   INVxp33_ASAP7_75t_R FE_OFC5873_n23491 (.Y(FE_OFN28581_n23491),
	.A(FE_OFN29001_n23491));
   INVx1_ASAP7_75t_L FE_OFC5872_n23491 (.Y(FE_OFN28580_n23491),
	.A(FE_OFN28579_n23491));
   INVxp67_ASAP7_75t_SL FE_OFC5868_n15218 (.Y(n13656),
	.A(n15218));
   INVx1_ASAP7_75t_R FE_OFC5867_n23691 (.Y(FE_OFN16221_n21234),
	.A(n23691));
   INVxp67_ASAP7_75t_SL FE_OFC5866_FE_OFN16316_n24840 (.Y(FE_OFN28578_FE_OFN16316_n24840),
	.A(n24841));
   INVxp67_ASAP7_75t_L FE_OFC5864_FE_OFN16316_n24840 (.Y(n24841),
	.A(FE_OFN16316_n24840));
   INVxp67_ASAP7_75t_L FE_OFC5863_n23821 (.Y(n23841),
	.A(FE_OFN16328_n23821));
   INVx1_ASAP7_75t_SL FE_OFC5862_n23821 (.Y(FE_OFN16328_n23821),
	.A(n23821));
   INVx1_ASAP7_75t_L FE_OFC5861_n22709 (.Y(n17884),
	.A(n22709));
   INVx1_ASAP7_75t_L FE_OFC5860_FE_OFN16231_n17691 (.Y(FE_OFN16232_n17691),
	.A(FE_OFN16231_n17691));
   INVx1_ASAP7_75t_R FE_OFC5859_n27003 (.Y(FE_OFN28576_n27003),
	.A(FE_OFN16252_n27003));
   BUFx2_ASAP7_75t_SL FE_OFC5858_n27003 (.Y(FE_OFN16252_n27003),
	.A(n21545));
   INVxp67_ASAP7_75t_L FE_OFC5856_n15746 (.Y(n14054),
	.A(n15746));
   INVxp33_ASAP7_75t_L FE_OFC5851_n26748 (.Y(FE_OFN28573_n26748),
	.A(FE_OCPN27541_n26748));
   INVx1_ASAP7_75t_SL FE_OFC5850_n26748 (.Y(FE_OCPN27541_n26748),
	.A(n26750));
   INVx1_ASAP7_75t_SL FE_OFC5849_n26748 (.Y(n26750),
	.A(n26748));
   INVxp33_ASAP7_75t_L FE_OFC5847_n26165 (.Y(n22917),
	.A(FE_OFN16250_n26165));
   INVx2_ASAP7_75t_R FE_OFC5844_n13359 (.Y(n14514),
	.A(n13359));
   INVx1_ASAP7_75t_L FE_OFC5843_n23830 (.Y(n21692),
	.A(n23830));
   INVxp67_ASAP7_75t_R FE_OFC5841_n20446 (.Y(n20447),
	.A(n20446));
   INVxp33_ASAP7_75t_L FE_OFC5840_n16544 (.Y(FE_OFN27048_n23045),
	.A(n16544));
   INVxp67_ASAP7_75t_R FE_OFC5839_n15997 (.Y(FE_OFN25985_n15997),
	.A(n14098));
   INVx1_ASAP7_75t_SL FE_OFC5838_n15997 (.Y(n14098),
	.A(n15997));
   INVxp67_ASAP7_75t_L FE_OFC5837_n15637 (.Y(n15640),
	.A(n15637));
   INVxp33_ASAP7_75t_L FE_OFC5836_n20477 (.Y(n20451),
	.A(n20477));
   INVxp67_ASAP7_75t_L FE_OFC5834_n16345 (.Y(n18079),
	.A(n16345));
   INVxp33_ASAP7_75t_L FE_OFC5833_n21922 (.Y(FE_OFN26533_n21922),
	.A(n25323));
   INVx1_ASAP7_75t_L FE_OFC5832_n21922 (.Y(n25323),
	.A(n21922));
   INVxp67_ASAP7_75t_L FE_OFC5828_n18369 (.Y(n18354),
	.A(n18369));
   INVxp33_ASAP7_75t_R FE_OFC5827_n24153 (.Y(n21705),
	.A(n24153));
   INVxp33_ASAP7_75t_R FE_OFC5826_n24077 (.Y(n24080),
	.A(n24077));
   INVxp33_ASAP7_75t_L FE_OFC5825_n21723 (.Y(FE_OFN28572_n21723),
	.A(n18868));
   INVx2_ASAP7_75t_L FE_OFC5821_w3_28 (.Y(FE_OFN28571_w3_28),
	.A(FE_OFN27130_w3_28));
   INVx1_ASAP7_75t_SL FE_OFC5820_w3_28 (.Y(FE_OFN27129_w3_28),
	.A(FE_OFN27130_w3_28));
   BUFx4f_ASAP7_75t_SL FE_OFC5819_w3_28 (.Y(FE_OFN27130_w3_28),
	.A(w3_28_));
   INVx1_ASAP7_75t_R FE_OFC5818_n19172 (.Y(FE_OFN28570_n19172),
	.A(n21815));
   BUFx3_ASAP7_75t_SL FE_OFC5817_n19172 (.Y(n21815),
	.A(n19172));
   BUFx3_ASAP7_75t_SL FE_OFC5816_n26501 (.Y(FE_OCPN28054_n26501),
	.A(n26501));
   INVxp33_ASAP7_75t_L FE_OFC5815_n18755 (.Y(FE_OFN28569_n18755),
	.A(n24092));
   INVx1_ASAP7_75t_L FE_OFC5814_n18755 (.Y(n24092),
	.A(n18755));
   INVxp67_ASAP7_75t_R FE_OFC5813_n24523 (.Y(n24522),
	.A(FE_OCPN27402_n24523));
   BUFx3_ASAP7_75t_SL FE_OFC5812_n24523 (.Y(FE_OCPN27402_n24523),
	.A(n24523));
   INVx1_ASAP7_75t_SL FE_OFC5809_FE_OCPN28279_n (.Y(n26673),
	.A(FE_OCPN28279_n));
   INVxp67_ASAP7_75t_L FE_OFC5808_n15747 (.Y(n15751),
	.A(n15747));
   INVxp67_ASAP7_75t_L FE_OFC5807_n19514 (.Y(FE_OFN28567_n19514),
	.A(n24056));
   INVx2_ASAP7_75t_SL FE_OFC5806_n19514 (.Y(n24056),
	.A(n19514));
   INVx1_ASAP7_75t_L FE_OFC5805_n26275 (.Y(FE_OFN25939_n26275),
	.A(FE_OFN27123_n26275));
   INVxp33_ASAP7_75t_R FE_OFC5802_n21491 (.Y(FE_OFN28566_n21491),
	.A(n19579));
   INVx1_ASAP7_75t_L FE_OFC5801_n21491 (.Y(n19579),
	.A(n21491));
   INVxp67_ASAP7_75t_L FE_OFC5800_n21475 (.Y(n21476),
	.A(FE_OFN25949_n21475));
   INVxp67_ASAP7_75t_L FE_OFC5798_n21667 (.Y(n21192),
	.A(n21667));
   BUFx2_ASAP7_75t_SL FE_OFC5797_n26845 (.Y(FE_OFN28565_n26845),
	.A(n26845));
   INVxp67_ASAP7_75t_L FE_OFC5794_n18308 (.Y(FE_OFN28564_n18308),
	.A(n17712));
   INVx1_ASAP7_75t_SL FE_OFC5793_n18308 (.Y(n17712),
	.A(n18308));
   INVxp33_ASAP7_75t_L FE_OFC5792_n24277 (.Y(n19870),
	.A(n24277));
   INVx1_ASAP7_75t_L FE_OFC5791_FE_OCPN28322_n18141 (.Y(n16686),
	.A(FE_OCPN28322_n18141));
   INVxp67_ASAP7_75t_L FE_OFC5790_n22189 (.Y(FE_OFN27150_n22175),
	.A(n22189));
   INVxp33_ASAP7_75t_L FE_OFC5789_n21159 (.Y(FE_RN_3_0),
	.A(n21159));
   INVxp67_ASAP7_75t_R FE_OFC5788_n22313 (.Y(FE_OFN16203_n22313),
	.A(n22812));
   INVxp67_ASAP7_75t_L FE_OFC5786_n26875 (.Y(FE_RN_2_0),
	.A(n26875));
   INVxp67_ASAP7_75t_L FE_OFC5784_n22447 (.Y(FE_OFN25954_n18719),
	.A(n22447));
   BUFx4f_ASAP7_75t_SL FE_OFC5783_n18020 (.Y(FE_OCPN28184_n18020),
	.A(n18020));
   INVx1_ASAP7_75t_L FE_OFC5782_n20480 (.Y(FE_OFN28563_n20480),
	.A(n17632));
   INVxp67_ASAP7_75t_L FE_OFC5781_n20480 (.Y(n17632),
	.A(n20480));
   INVxp67_ASAP7_75t_L FE_OFC5780_FE_RN_175_0 (.Y(FE_RN_171_0),
	.A(FE_RN_175_0));
   INVx1_ASAP7_75t_L FE_OFC5779_n19342 (.Y(FE_OFN28562_n19342),
	.A(n22019));
   INVx1_ASAP7_75t_L FE_OFC5778_n19342 (.Y(n22019),
	.A(n19342));
   INVx1_ASAP7_75t_L FE_OFC5776_n24122 (.Y(n24123),
	.A(n24122));
   INVx1_ASAP7_75t_L FE_OFC5775_n25419 (.Y(FE_OFN28561_n25419),
	.A(n18914));
   INVx1_ASAP7_75t_L FE_OFC5774_n25419 (.Y(n18914),
	.A(n25419));
   INVxp33_ASAP7_75t_L FE_OFC5773_n22749 (.Y(FE_OFN28560_n22749),
	.A(n25740));
   INVx1_ASAP7_75t_SL FE_OFC5772_n22749 (.Y(n25740),
	.A(n22749));
   INVxp67_ASAP7_75t_L FE_OFC5771_n18278 (.Y(FE_OFN28559_n18278),
	.A(n17070));
   INVx1_ASAP7_75t_SL FE_OFC5770_n18278 (.Y(n17070),
	.A(n18278));
   INVxp67_ASAP7_75t_L FE_OFC5769_n23073 (.Y(FE_OFN28558_n23073),
	.A(n18724));
   INVx1_ASAP7_75t_L FE_OFC5768_n23073 (.Y(n18724),
	.A(n23073));
   INVxp33_ASAP7_75t_L FE_OFC5763_n23955 (.Y(n19638),
	.A(n23955));
   INVxp67_ASAP7_75t_R FE_OFC5762_n24960 (.Y(FE_OFN27094_n24956),
	.A(n24960));
   INVxp67_ASAP7_75t_L FE_OFC5760_n15688 (.Y(n14043),
	.A(n15688));
   INVxp67_ASAP7_75t_L FE_OFC5759_n25073 (.Y(n25072),
	.A(n25073));
   INVxp33_ASAP7_75t_L FE_OFC5758_n25031 (.Y(FE_OFN28557_n25031),
	.A(n24646));
   INVx1_ASAP7_75t_SL FE_OFC5757_n25031 (.Y(n24646),
	.A(n25031));
   INVx1_ASAP7_75t_L FE_OFC5756_n23236 (.Y(FE_OFN26556_n23236),
	.A(n23236));
   INVxp67_ASAP7_75t_R FE_OFC5755_n19784 (.Y(n19785),
	.A(n19784));
   INVx1_ASAP7_75t_L FE_OFC5754_n24516 (.Y(FE_OFN28556_n24516),
	.A(n24101));
   INVx1_ASAP7_75t_L FE_OFC5752_n24516 (.Y(n24101),
	.A(n24516));
   INVxp67_ASAP7_75t_L FE_OFC5749_n23552 (.Y(FE_OFN16241_n23552),
	.A(n16694));
   INVx1_ASAP7_75t_L FE_OFC5748_n23552 (.Y(n16694),
	.A(n23552));
   INVx1_ASAP7_75t_L FE_OFC5747_n15253 (.Y(FE_OFN75_n15253),
	.A(n15253));
   INVxp67_ASAP7_75t_R FE_OFC5746_n25875 (.Y(FE_OFN25999_n25875),
	.A(n25875));
   INVxp67_ASAP7_75t_L FE_OFC5745_n19498 (.Y(n24837),
	.A(n19498));
   INVx1_ASAP7_75t_SL FE_OFC5744_n19498 (.Y(FE_OFN95_n19498),
	.A(n19498));
   INVxp67_ASAP7_75t_R FE_OFC5743_n21876 (.Y(FE_OFN28554_n21876),
	.A(n16538));
   INVx1_ASAP7_75t_L FE_OFC5742_n21876 (.Y(n16538),
	.A(n21876));
   BUFx2_ASAP7_75t_SL FE_OFC5741_n24491 (.Y(FE_OCPN27412_n24491),
	.A(n24491));
   INVxp33_ASAP7_75t_L FE_OFC5740_n25599 (.Y(FE_OFN28553_n25599),
	.A(FE_OFN27069_n24478));
   INVxp67_ASAP7_75t_R FE_OFC5739_n25599 (.Y(FE_OFN27069_n24478),
	.A(n24478));
   INVxp67_ASAP7_75t_L FE_OFC5737_n23943 (.Y(FE_OFN25937_n23943),
	.A(n21077));
   INVx1_ASAP7_75t_L FE_OFC5736_n23943 (.Y(n21077),
	.A(n23943));
   INVxp33_ASAP7_75t_L FE_OFC5735_n20105 (.Y(FE_OFN28552_n20105),
	.A(n19945));
   INVxp67_ASAP7_75t_L FE_OFC5734_n20105 (.Y(n19945),
	.A(n20105));
   BUFx3_ASAP7_75t_SL FE_OFC5733_FE_OFN26114_n (.Y(FE_OFN28551_FE_OFN26114_n),
	.A(FE_OFN27151_n));
   INVxp67_ASAP7_75t_L FE_OFC5729_n18805 (.Y(n18807),
	.A(n18805));
   BUFx2_ASAP7_75t_L FE_OFC5728_n20339 (.Y(FE_OCPN27508_n20339),
	.A(n20339));
   INVxp33_ASAP7_75t_L FE_OFC5727_n22386 (.Y(n22388),
	.A(n22386));
   INVxp33_ASAP7_75t_R FE_OFC5726_n25149 (.Y(n18349),
	.A(n25149));
   INVxp67_ASAP7_75t_SL FE_OFC5725_n15763 (.Y(n15764),
	.A(n15763));
   INVxp67_ASAP7_75t_R FE_OFC5723_n21934 (.Y(FE_OFN28549_n21934),
	.A(n16330));
   INVx1_ASAP7_75t_R FE_OFC5722_n21934 (.Y(n16330),
	.A(n21934));
   INVxp33_ASAP7_75t_L FE_OFC5721_n22499 (.Y(n17485),
	.A(FE_OFN26031_n22499));
   INVxp67_ASAP7_75t_L FE_OFC5719_n27092 (.Y(FE_OFN28548_n27092),
	.A(n19419));
   INVxp67_ASAP7_75t_L FE_OFC5716_n20876 (.Y(n20878),
	.A(n20876));
   BUFx2_ASAP7_75t_L FE_OFC5715_n27178 (.Y(n27176),
	.A(n27178));
   INVx2_ASAP7_75t_SL FE_OFC5714_n27178 (.Y(FE_OFN105_n27178),
	.A(n27178));
   INVxp67_ASAP7_75t_L FE_OFC5712_n23176 (.Y(n22843),
	.A(n23176));
   INVxp67_ASAP7_75t_R FE_OFC5711_n23015 (.Y(n23979),
	.A(n23015));
   INVxp33_ASAP7_75t_R FE_OFC5710_n26091 (.Y(FE_OFN28546_n26091),
	.A(n18158));
   HB1xp67_ASAP7_75t_SL FE_OFC5709_n26091 (.Y(n18158),
	.A(n26091));
   INVxp33_ASAP7_75t_R FE_OFC5708_FE_OCPN28448_n27048 (.Y(FE_OCPN28073_n27049),
	.A(FE_OFN29224_FE_OCPN28074_n27049));
   INVxp33_ASAP7_75t_L FE_OFC5707_n26685 (.Y(n26686),
	.A(FE_OCPN27753_n26685));
   BUFx2_ASAP7_75t_SL FE_OFC5706_n26685 (.Y(FE_OCPN27753_n26685),
	.A(n26685));
   INVxp67_ASAP7_75t_L FE_OFC5704_n24861 (.Y(n24862),
	.A(n24861));
   INVx1_ASAP7_75t_SL FE_OFC5703_n25002 (.Y(n25000),
	.A(n25002));
   INVx1_ASAP7_75t_R FE_OFC5701_n21587 (.Y(n20423),
	.A(n21587));
   HB1xp67_ASAP7_75t_L FE_OFC5699_n13805 (.Y(FE_OFN28544_n13805),
	.A(n13805));
   INVxp67_ASAP7_75t_R FE_OFC5697_n21368 (.Y(FE_OFN65_n21412),
	.A(n21368));
   INVxp67_ASAP7_75t_L FE_OFC5696_n25987 (.Y(n25989),
	.A(FE_OCPN27589_n25987));
   BUFx2_ASAP7_75t_SL FE_OFC5695_n25987 (.Y(FE_OCPN27589_n25987),
	.A(n25987));
   INVxp67_ASAP7_75t_R FE_OFC5694_FE_OFN109_n15994 (.Y(FE_OFN28543_FE_OFN109_n15994),
	.A(FE_OFN112_n15994));
   BUFx2_ASAP7_75t_SL FE_OFC5693_FE_OFN109_n15994 (.Y(FE_OFN112_n15994),
	.A(FE_OFN109_n15994));
   INVxp33_ASAP7_75t_R FE_OFC5691_n22874 (.Y(FE_OFN16356_n22874),
	.A(n25504));
   INVxp33_ASAP7_75t_L FE_OFC5689_sa02_6 (.Y(n17815),
	.A(sa02_6_));
   INVx1_ASAP7_75t_L FE_OFC5687_FE_OFN25901_n22133 (.Y(FE_OFN27176_n),
	.A(FE_OFN25901_n22133));
   INVxp67_ASAP7_75t_R FE_OFC5686_n15433 (.Y(FE_OFN28542_n15433),
	.A(n14159));
   INVx2_ASAP7_75t_SL FE_OFC5685_n15433 (.Y(n14159),
	.A(n15433));
   INVxp33_ASAP7_75t_R FE_OFC5684_n16476 (.Y(FE_OFN28541_n16476),
	.A(n24487));
   INVx2_ASAP7_75t_L FE_OFC5683_n16476 (.Y(n24487),
	.A(n16476));
   INVxp33_ASAP7_75t_L FE_OFC5682_n23145 (.Y(FE_OFN16291_n23142),
	.A(n23145));
   INVxp67_ASAP7_75t_L FE_OFC5681_n25219 (.Y(FE_OFN16220_n25219),
	.A(n27090));
   INVx1_ASAP7_75t_L FE_OFC5680_n25219 (.Y(n27090),
	.A(n25219));
   INVx1_ASAP7_75t_SL FE_OFC5679_n26839 (.Y(n26836),
	.A(n26839));
   INVxp67_ASAP7_75t_L FE_OFC5678_n27097 (.Y(n27098),
	.A(n27097));
   INVxp67_ASAP7_75t_R FE_OFC5676_n21599 (.Y(FE_OFN28540_n21599),
	.A(n22148));
   INVx1_ASAP7_75t_L FE_OFC5675_n21599 (.Y(n22148),
	.A(n21599));
   INVxp33_ASAP7_75t_L FE_OFC5674_n22336 (.Y(FE_OFN28539_n22336),
	.A(FE_OCPN5167_n22336));
   INVx1_ASAP7_75t_SL FE_OFC5673_n22336 (.Y(n19968),
	.A(FE_OCPN5167_n22336));
   INVx2_ASAP7_75t_SL FE_OFC5672_n22336 (.Y(FE_OCPN5167_n22336),
	.A(n22336));
   INVx1_ASAP7_75t_R FE_OFC5671_n23027 (.Y(n23029),
	.A(n23027));
   INVx1_ASAP7_75t_L FE_OFC5670_n18922 (.Y(n17021),
	.A(FE_OFN25977_n18922));
   INVx1_ASAP7_75t_L FE_OFC5669_n18922 (.Y(FE_OFN25977_n18922),
	.A(n18922));
   INVx1_ASAP7_75t_L FE_OFC5668_n14667 (.Y(n14714),
	.A(n14667));
   INVx2_ASAP7_75t_L FE_OFC5667_n16166 (.Y(FE_OFN28538_n16166),
	.A(n16166));
   INVxp67_ASAP7_75t_L FE_OFC5665_n20205 (.Y(FE_RN_201_0),
	.A(n20205));
   INVx2_ASAP7_75t_SL FE_OFC5662_n25462 (.Y(FE_OCPN28106_FE_OFN25876_n25462),
	.A(n24903));
   INVx2_ASAP7_75t_SL FE_OFC5661_n25462 (.Y(n24903),
	.A(n25462));
   INVxp67_ASAP7_75t_L FE_OFC5658_sa20_2 (.Y(FE_OFN28537_sa20_2),
	.A(FE_OFN28536_sa20_2));
   INVx1_ASAP7_75t_L FE_OFC5657_sa20_2 (.Y(FE_OFN28536_sa20_2),
	.A(n18533));
   INVxp67_ASAP7_75t_SL FE_OFC5656_sa20_2 (.Y(FE_RN_168_0),
	.A(n18533));
   INVx2_ASAP7_75t_L FE_OFC5655_sa20_2 (.Y(n18533),
	.A(FE_OCPN27371_sa20_2));
   INVx5_ASAP7_75t_SL FE_OFC5653_sa20_2 (.Y(FE_OCPN27371_sa20_2),
	.A(FE_RN_165_0));
   INVx2_ASAP7_75t_SL FE_OFC5651_sa20_2 (.Y(FE_RN_165_0),
	.A(sa20_2_));
   INVxp33_ASAP7_75t_R FE_OFC5650_n24046 (.Y(n20552),
	.A(n24046));
   INVxp33_ASAP7_75t_L FE_OFC5649_n24835 (.Y(n24441),
	.A(n24835));
   INVxp33_ASAP7_75t_L FE_OFC5648_n19738 (.Y(FE_OFN28535_n19738),
	.A(n18797));
   INVx1_ASAP7_75t_L FE_OFC5647_n19738 (.Y(n18797),
	.A(n19738));
   INVx1_ASAP7_75t_SL FE_OFC5646_FE_OCPN27333_n25250 (.Y(n25252),
	.A(FE_OCPN27333_n25250));
   INVxp67_ASAP7_75t_R FE_OFC5645_n21462 (.Y(FE_OFN28534_n21462),
	.A(n19593));
   INVx1_ASAP7_75t_L FE_OFC5644_n21462 (.Y(n19593),
	.A(n21462));
   INVx1_ASAP7_75t_R FE_OFC5643_n24995 (.Y(FE_OFN28533_n24995),
	.A(FE_OFN27138_n24012));
   INVx1_ASAP7_75t_L FE_OFC5642_n24995 (.Y(FE_OFN27138_n24012),
	.A(n24995));
   INVx1_ASAP7_75t_SL FE_OFC5640_FE_OFN56_n14826 (.Y(FE_OFN28531_FE_OFN56_n14826),
	.A(FE_OFN16300_n14826));
   INVx2_ASAP7_75t_L FE_OFC5639_FE_OFN56_n14826 (.Y(FE_OFN16300_n14826),
	.A(FE_OFN56_n14826));
   INVx1_ASAP7_75t_SL FE_OFC5638_n14593 (.Y(FE_OFN28530_n14593),
	.A(FE_OFN27222_n14593));
   INVx1_ASAP7_75t_L FE_OFC5637_n14593 (.Y(FE_OFN27222_n14593),
	.A(n14593));
   INVx1_ASAP7_75t_L FE_OFC5635_n14593 (.Y(FE_OFN26104_n13659),
	.A(n14593));
   INVx1_ASAP7_75t_SL FE_OFC5634_n22966 (.Y(n24812),
	.A(n22966));
   INVxp67_ASAP7_75t_L FE_OFC5633_n23724 (.Y(n20638),
	.A(n23724));
   INVxp33_ASAP7_75t_R FE_OFC5632_FE_OCPN5067_n24089 (.Y(n24090),
	.A(n24089));
   INVx1_ASAP7_75t_L FE_OFC5630_n22024 (.Y(FE_OFN27046_n22024),
	.A(n26163));
   INVxp33_ASAP7_75t_R FE_OFC5628_n15683 (.Y(FE_OFN16211_n13876),
	.A(n15683));
   INVxp67_ASAP7_75t_L FE_OFC5627_n19058 (.Y(n24781),
	.A(FE_OFN16326_n19058));
   INVx1_ASAP7_75t_L FE_OFC5626_n19058 (.Y(FE_OFN16326_n19058),
	.A(n19058));
   INVxp33_ASAP7_75t_L FE_OFC5625_n17728 (.Y(n17698),
	.A(n17728));
   BUFx2_ASAP7_75t_L FE_OFC5624_n21899 (.Y(FE_OCPN28358_n21899),
	.A(n21899));
   INVxp67_ASAP7_75t_L FE_OFC5623_n25764 (.Y(n25763),
	.A(n25764));
   INVx3_ASAP7_75t_SL FE_OFC5621_n16774 (.Y(FE_OCPN27631_n16774),
	.A(FE_OCPN27632_n16774));
   INVxp67_ASAP7_75t_L FE_OFC5618_FE_OCPN5180_n18174 (.Y(n24691),
	.A(n18174));
   BUFx2_ASAP7_75t_SL FE_OFC5617_n26842 (.Y(FE_OCPN27940_n26842),
	.A(n26842));
   INVxp67_ASAP7_75t_L FE_OFC5616_n20421 (.Y(n18504),
	.A(n20421));
   INVx1_ASAP7_75t_R FE_OFC5613_FE_OFN16412_w3_26 (.Y(n24470),
	.A(FE_OFN16412_w3_26));
   INVxp67_ASAP7_75t_L FE_OFC5611_n25241 (.Y(FE_OFN28528_n25241),
	.A(n26625));
   INVx1_ASAP7_75t_SL FE_OFC5609_n25241 (.Y(n26625),
	.A(n25241));
   INVxp67_ASAP7_75t_L FE_OFC5601_n19188 (.Y(FE_OFN114_n22512),
	.A(n19188));
   INVxp33_ASAP7_75t_R FE_OFC5598_FE_OCPN28163_FE_OFN99_sa20_5 (.Y(FE_OFN27045_n),
	.A(FE_OCPN28163_FE_OFN99_sa20_5));
   BUFx2_ASAP7_75t_SL FE_OFC5594_n23031 (.Y(FE_OCPN5015_n23031),
	.A(n23031));
   INVx2_ASAP7_75t_SL FE_OFC5593_n26252 (.Y(FE_OFN16311_n26252),
	.A(n26255));
   INVx2_ASAP7_75t_SL FE_OFC5592_n26252 (.Y(n26255),
	.A(n26252));
   INVxp67_ASAP7_75t_R FE_OFC5591_n17261 (.Y(FE_OFN28522_n17261),
	.A(FE_OFN28958_n17261));
   INVxp67_ASAP7_75t_L FE_OFC5589_n24564 (.Y(n19183),
	.A(n24564));
   INVxp67_ASAP7_75t_R FE_OFC5588_n23455 (.Y(n23456),
	.A(FE_OCPN27628_n23455));
   BUFx2_ASAP7_75t_L FE_OFC5587_n23455 (.Y(FE_OCPN27628_n23455),
	.A(n23455));
   INVx1_ASAP7_75t_R FE_OFC5586_n23094 (.Y(n22424),
	.A(n23094));
   INVx1_ASAP7_75t_SL FE_OFC5585_n22353 (.Y(FE_OFN27163_n20304),
	.A(n22353));
   INVx1_ASAP7_75t_R FE_OFC5584_n26007 (.Y(FE_OFN28521_n26007),
	.A(FE_RN_78_0));
   INVxp67_ASAP7_75t_L FE_OFC5583_n26007 (.Y(FE_RN_78_0),
	.A(n26007));
   INVx1_ASAP7_75t_R FE_OFC5582_n22753 (.Y(FE_OFN28520_n22753),
	.A(FE_OCPN27252_n22753));
   INVx1_ASAP7_75t_L FE_OFC5578_n22753 (.Y(FE_OCPN27252_n22753),
	.A(n22753));
   INVxp33_ASAP7_75t_L FE_OFC5573_n22062 (.Y(FE_OFN28515_n22062),
	.A(FE_OFN28924_n25912));
   INVxp67_ASAP7_75t_R FE_OFC5571_FE_OCPN27478_n25011 (.Y(n25010),
	.A(FE_OCPN27478_n25011));
   INVx1_ASAP7_75t_SL FE_OFC5569_n25946 (.Y(FE_OFN16322_n25946),
	.A(n25947));
   INVx2_ASAP7_75t_SL FE_OFC5568_n25946 (.Y(n25947),
	.A(n25946));
   INVxp67_ASAP7_75t_SRAM FE_OFC5565_n19335 (.Y(n18981),
	.A(n19335));
   INVxp33_ASAP7_75t_L FE_OFC5564_n21975 (.Y(n21978),
	.A(n21975));
   INVxp67_ASAP7_75t_L FE_OFC5563_n26155 (.Y(FE_OFN27165_n),
	.A(FE_OFN26542_n26155));
   INVx1_ASAP7_75t_L FE_OFC5562_n26155 (.Y(FE_OFN26542_n26155),
	.A(n23511));
   BUFx3_ASAP7_75t_SL FE_OFC5560_n26336 (.Y(FE_OCPN27991_n26336),
	.A(n26336));
   INVx1_ASAP7_75t_L FE_OFC5557_n20795 (.Y(n20799),
	.A(n20795));
   INVxp67_ASAP7_75t_L FE_OFC5556_n19950 (.Y(n24852),
	.A(n19950));
   INVxp67_ASAP7_75t_L FE_OFC5555_n20470 (.Y(FE_OFN28513_n20470),
	.A(n20481));
   INVx2_ASAP7_75t_SL FE_OFC5554_n20470 (.Y(n20481),
	.A(n20470));
   BUFx2_ASAP7_75t_L FE_OFC5553_n16760 (.Y(FE_OCPN27616_n16760),
	.A(n16760));
   INVxp33_ASAP7_75t_L FE_OFC5551_FE_OCPN27529_sa21_4 (.Y(FE_OFN16267_sa21_4),
	.A(FE_OFN25989_sa21_4));
   INVxp33_ASAP7_75t_L FE_OFC5549_n24157 (.Y(n24159),
	.A(n24157));
   INVxp33_ASAP7_75t_R FE_OFC5548_n15610 (.Y(n14881),
	.A(n15610));
   INVx2_ASAP7_75t_SL FE_OFC5547_n27020 (.Y(FE_OFN28512_n27020),
	.A(n27023));
   INVx2_ASAP7_75t_SL FE_OFC5545_n27020 (.Y(n27023),
	.A(n27020));
   BUFx2_ASAP7_75t_L FE_OFC5543_sa23_5 (.Y(FE_OCPN27482_sa23_5),
	.A(FE_OFN27078_sa23_5));
   INVxp67_ASAP7_75t_R FE_OFC5538_n24855 (.Y(FE_OFN26166_n24855),
	.A(n24855));
   INVxp33_ASAP7_75t_L FE_OFC5537_n25088 (.Y(FE_OFN28511_n25088),
	.A(n24579));
   INVxp67_ASAP7_75t_L FE_OFC5536_n25088 (.Y(n24579),
	.A(n25088));
   INVxp67_ASAP7_75t_L FE_OFC5535_n21074 (.Y(FE_RN_233_0),
	.A(n21074));
   INVxp67_ASAP7_75t_L FE_OFC5534_n21215 (.Y(FE_OFN28510_n21215),
	.A(n21218));
   INVx1_ASAP7_75t_L FE_OFC5533_n21215 (.Y(n21218),
	.A(n21215));
   INVxp67_ASAP7_75t_L FE_OFC5531_n19953 (.Y(n17681),
	.A(n19953));
   INVxp33_ASAP7_75t_L FE_OFC5523_n15661 (.Y(n15662),
	.A(n15661));
   INVxp67_ASAP7_75t_SL FE_OFC5522_n14602 (.Y(n14601),
	.A(n14602));
   INVxp33_ASAP7_75t_L FE_OFC5521_n22194 (.Y(n22204),
	.A(n22194));
   INVx1_ASAP7_75t_SL FE_OFC5520_n24628 (.Y(n24629),
	.A(FE_OFN117_n24628));
   INVx2_ASAP7_75t_SL FE_OFC5519_n24628 (.Y(FE_OFN117_n24628),
	.A(n24628));
   INVxp67_ASAP7_75t_L FE_OFC5518_n26996 (.Y(FE_OFN28506_n26996),
	.A(FE_RN_213_0));
   INVxp67_ASAP7_75t_L FE_OFC5517_n26996 (.Y(FE_RN_213_0),
	.A(n26996));
   INVx1_ASAP7_75t_R FE_OFC5515_n19584 (.Y(n19585),
	.A(n19584));
   BUFx2_ASAP7_75t_SL FE_OFC5514_n16422 (.Y(FE_OCPN27555_n16422),
	.A(n16422));
   INVxp67_ASAP7_75t_L FE_OFC5513_n23488 (.Y(n23492),
	.A(n23488));
   INVx1_ASAP7_75t_SL FE_OFC5512_n25144 (.Y(n25145),
	.A(n25144));
   BUFx2_ASAP7_75t_L FE_OFC5511_n22779 (.Y(FE_OCPN28309_n22779),
	.A(n22779));
   INVxp33_ASAP7_75t_L FE_OFC5510_n18130 (.Y(n18131),
	.A(n18130));
   INVx1_ASAP7_75t_R FE_OFC5509_n23296 (.Y(FE_OFN28505_n23296),
	.A(n21099));
   INVx1_ASAP7_75t_L FE_OFC5508_n23296 (.Y(n21099),
	.A(n23296));
   INVxp67_ASAP7_75t_R FE_OFC5507_n21944 (.Y(n20863),
	.A(n21944));
   INVxp33_ASAP7_75t_L FE_OFC5506_n22039 (.Y(n22040),
	.A(n22039));
   INVx1_ASAP7_75t_L FE_OFC5505_n21349 (.Y(n17496),
	.A(n21349));
   INVx1_ASAP7_75t_SL FE_OFC5504_n26825 (.Y(n26824),
	.A(n26825));
   INVxp33_ASAP7_75t_R FE_OFC5501_n15929 (.Y(n15931),
	.A(n15929));
   INVxp67_ASAP7_75t_L FE_OFC5500_n21904 (.Y(n21907),
	.A(n21904));
   INVxp67_ASAP7_75t_R FE_OFC5499_n19754 (.Y(FE_OFN57_n19754),
	.A(n23121));
   INVx1_ASAP7_75t_SL FE_OFC5498_n19754 (.Y(n23121),
	.A(n19754));
   INVxp67_ASAP7_75t_L FE_OFC5497_n24085 (.Y(FE_RN_187_0),
	.A(n24085));
   INVxp33_ASAP7_75t_R FE_OFC5496_n15809 (.Y(n15042),
	.A(n15809));
   BUFx2_ASAP7_75t_SL FE_OFC5494_n25956 (.Y(FE_OFN16249_n25956),
	.A(n25956));
   INVxp33_ASAP7_75t_L FE_OFC5491_n25526 (.Y(n25527),
	.A(n25526));
   INVx1_ASAP7_75t_SL FE_OFC5490_n15915 (.Y(n15903),
	.A(n15915));
   INVxp33_ASAP7_75t_R FE_OFC5488_FE_OFN26008_n16010 (.Y(FE_OFN26564_n),
	.A(n14919));
   INVxp67_ASAP7_75t_L FE_OFC5487_n14716 (.Y(n14717),
	.A(n14716));
   INVxp33_ASAP7_75t_L FE_OFC5486_n25539 (.Y(n25540),
	.A(n25539));
   INVxp33_ASAP7_75t_R FE_OFC5485_n26596 (.Y(FE_OFN28503_n26596),
	.A(n20828));
   INVx1_ASAP7_75t_SL FE_OFC5484_n26596 (.Y(n20828),
	.A(n26596));
   BUFx2_ASAP7_75t_R FE_OFC5482_n22721 (.Y(FE_OFN25907_sa12_2),
	.A(n22721));
   INVxp33_ASAP7_75t_SL FE_OFC5480_n15055 (.Y(n15056),
	.A(FE_OFN16235_n15055));
   INVxp67_ASAP7_75t_SL FE_OFC5478_FE_OFN16405_n16117 (.Y(FE_OFN16403_n16117),
	.A(FE_OFN16405_n16117));
   INVxp33_ASAP7_75t_R FE_OFC5477_n25865 (.Y(FE_OFN28502_n25865),
	.A(n25996));
   INVxp67_ASAP7_75t_L FE_OFC5475_n15010 (.Y(n15865),
	.A(n15010));
   INVxp33_ASAP7_75t_L FE_OFC5474_n18273 (.Y(n16993),
	.A(n18273));
   INVxp33_ASAP7_75t_L FE_OFC5472_n24241 (.Y(FE_OFN16398_n24241),
	.A(n24241));
   INVxp67_ASAP7_75t_L FE_OFC5470_n19480 (.Y(n18882),
	.A(n19480));
   INVxp33_ASAP7_75t_R FE_OFC5468_FE_OFN26020_n14010 (.Y(FE_OFN16240_n14011),
	.A(FE_OFN28501_FE_OFN26020_n14010));
   BUFx2_ASAP7_75t_SL FE_OFC5467_n18561 (.Y(FE_OCPN27891_n18561),
	.A(n18561));
   INVx1_ASAP7_75t_L FE_OFC5466_n17163 (.Y(n17166),
	.A(n17163));
   INVxp67_ASAP7_75t_L FE_OFC5465_n20813 (.Y(n19505),
	.A(n20813));
   INVxp67_ASAP7_75t_L FE_OFC5464_FE_OCPN5081_n19874 (.Y(n23654),
	.A(n19874));
   INVxp67_ASAP7_75t_L FE_OFC5463_n27011 (.Y(n22417),
	.A(n27011));
   INVxp33_ASAP7_75t_R FE_OFC5462_FE_OCPN5078_n25823 (.Y(FE_OFN28500_FE_OCPN5078_n25823),
	.A(FE_OFN16334_n25823));
   INVxp67_ASAP7_75t_R FE_OFC5461_FE_OCPN5078_n25823 (.Y(FE_OFN16334_n25823),
	.A(n25823));
   INVxp67_ASAP7_75t_L FE_OFC5460_sa00_6 (.Y(FE_OFN28499_sa00_6),
	.A(n17305));
   INVxp67_ASAP7_75t_R FE_OFC5457_sa00_6 (.Y(n17305),
	.A(sa00_6_));
   BUFx2_ASAP7_75t_SL FE_OFC5456_n27143 (.Y(FE_OCPN27235_n27143),
	.A(n27143));
   INVxp33_ASAP7_75t_L FE_OFC5455_n22922 (.Y(n26159),
	.A(n22922));
   INVx1_ASAP7_75t_R FE_OFC5453_n15201 (.Y(FE_OFN28496_n15201),
	.A(n15201));
   INVxp33_ASAP7_75t_L FE_OFC5451_n24584 (.Y(FE_OFN28495_n24584),
	.A(n24601));
   INVxp67_ASAP7_75t_R FE_OFC5449_n24584 (.Y(n24601),
	.A(n24584));
   INVx2_ASAP7_75t_SL FE_OFC5448_n25976 (.Y(FE_OFN16263_n25976),
	.A(n25974));
   BUFx2_ASAP7_75t_SL FE_OFC5447_n25976 (.Y(n25974),
	.A(n25976));
   INVx1_ASAP7_75t_SL FE_OFC5446_n20899 (.Y(n20931),
	.A(n20899));
   BUFx2_ASAP7_75t_SL FE_OFC5441_n23426 (.Y(FE_OCPN27611_n23426),
	.A(n23426));
   HB1xp67_ASAP7_75t_SL FE_OFC5440_n15512 (.Y(FE_OCPN28278_n15512),
	.A(n15512));
   INVxp33_ASAP7_75t_L FE_OFC5439_n24489 (.Y(n16433),
	.A(n24489));
   INVxp33_ASAP7_75t_R FE_OFC5437_n25634 (.Y(n25636),
	.A(n25634));
   BUFx2_ASAP7_75t_SL FE_OFC5436_n16977 (.Y(FE_OCPN27761_n16977),
	.A(n16977));
   INVxp67_ASAP7_75t_L FE_OFC5434_n25738 (.Y(n25742),
	.A(n25738));
   INVxp33_ASAP7_75t_L FE_OFC5433_n16604 (.Y(n16603),
	.A(n16604));
   INVxp67_ASAP7_75t_L FE_OFC5432_n19885 (.Y(n16753),
	.A(n19885));
   HB1xp67_ASAP7_75t_L FE_OFC5431_n23974 (.Y(FE_OFN16421_n23974),
	.A(n23974));
   INVx1_ASAP7_75t_L FE_OFC5430_n23974 (.Y(FE_OFN50_w3_18),
	.A(n23974));
   INVx1_ASAP7_75t_R FE_OFC5429_n18114 (.Y(n18116),
	.A(n18114));
   INVx1_ASAP7_75t_L FE_OFC5428_n26790 (.Y(FE_OCPN27435_n26790),
	.A(n26787));
   BUFx2_ASAP7_75t_SL FE_OFC5427_n26790 (.Y(n26787),
	.A(n26790));
   INVxp33_ASAP7_75t_R FE_OFC5423_n26739 (.Y(FE_OFN171_n26739),
	.A(n26739));
   INVx1_ASAP7_75t_L FE_OFC5422_n24326 (.Y(n16914),
	.A(n24326));
   INVxp33_ASAP7_75t_L FE_OFC5421_n22657 (.Y(n22659),
	.A(n22657));
   BUFx3_ASAP7_75t_L FE_OFC5420_n18016 (.Y(FE_OCPN27617_n18016),
	.A(n18016));
   INVxp33_ASAP7_75t_L FE_OFC5419_n25903 (.Y(n21203),
	.A(n25903));
   INVx4_ASAP7_75t_SL FE_OFC5417_sa31_0 (.Y(FE_OFN28492_sa31_0),
	.A(FE_OFN26095_n16293));
   INVx5_ASAP7_75t_SL FE_OFC5416_sa31_0 (.Y(FE_OFN26095_n16293),
	.A(FE_OFN27116_n16293));
   INVx2_ASAP7_75t_SL FE_OFC5415_sa31_0 (.Y(FE_OFN27116_n16293),
	.A(sa31_0_));
   INVxp67_ASAP7_75t_L FE_OFC5414_n21974 (.Y(n20846),
	.A(n21974));
   BUFx2_ASAP7_75t_SL FE_OFC5410_sa13_3 (.Y(FE_OFN28491_sa13_3),
	.A(FE_OFN28979_n));
   INVx1_ASAP7_75t_L FE_OFC5407_ld_r (.Y(FE_OFN28490_ld_r),
	.A(FE_OFN28485_ld_r));
   INVx3_ASAP7_75t_L FE_OFC5406_ld_r (.Y(FE_OFN28489_ld_r),
	.A(FE_OFN28485_ld_r));
   INVx2_ASAP7_75t_R FE_OFC5404_ld_r (.Y(FE_OFN28487_ld_r),
	.A(FE_OFN17_FE_DBTN0_ld_r));
   INVx1_ASAP7_75t_L FE_OFC5403_ld_r (.Y(FE_OFN28486_ld_r),
	.A(FE_OFN17_FE_DBTN0_ld_r));
   INVxp67_ASAP7_75t_L FE_OFC5402_ld_r (.Y(FE_OFN28485_ld_r),
	.A(FE_OFN15_FE_DBTN0_ld_r));
   BUFx2_ASAP7_75t_R FE_OFC5401_ld_r (.Y(FE_OFN28484_ld_r),
	.A(FE_OFN15_FE_DBTN0_ld_r));
   BUFx2_ASAP7_75t_R FE_OFC5400_ld_r (.Y(FE_OFN28483_ld_r),
	.A(FE_OFN15_FE_DBTN0_ld_r));
   HB1xp67_ASAP7_75t_SL FE_OFC5399_ld_r (.Y(FE_OFN28482_ld_r),
	.A(FE_OFN16214_ld_r));
   INVxp67_ASAP7_75t_R FE_OFC5398_ld_r (.Y(FE_OFN17_FE_DBTN0_ld_r),
	.A(FE_OFN14_FE_DBTN0_ld_r));
   BUFx2_ASAP7_75t_SRAM FE_OFC5397_ld_r (.Y(FE_OFN16_FE_DBTN0_ld_r),
	.A(FE_OFN14_FE_DBTN0_ld_r));
   INVx2_ASAP7_75t_SL FE_OFC5396_ld_r (.Y(FE_OFN15_FE_DBTN0_ld_r),
	.A(FE_OFN13_FE_DBTN0_ld_r));
   INVx2_ASAP7_75t_L FE_OFC5395_ld_r (.Y(FE_OFN16214_ld_r),
	.A(FE_OFN3_ld_r));
   INVx2_ASAP7_75t_R FE_OFC5394_ld_r (.Y(FE_OFN16213_ld_r),
	.A(FE_OFN3_ld_r));
   BUFx2_ASAP7_75t_L FE_OFC5393_ld_r (.Y(FE_OFN14_FE_DBTN0_ld_r),
	.A(FE_DBTN0_ld_r));
   INVx1_ASAP7_75t_L FE_OFC5392_ld_r (.Y(FE_OFN13_FE_DBTN0_ld_r),
	.A(FE_DBTN0_ld_r));
   INVxp33_ASAP7_75t_L FE_OFC5391_ld_r (.Y(FE_OFN3_ld_r),
	.A(FE_OFN12_FE_DBTN0_ld_r));
   INVx1_ASAP7_75t_L FE_OFC5390_ld_r (.Y(FE_DBTN0_ld_r),
	.A(FE_OFN1_ld_r));
   BUFx2_ASAP7_75t_L FE_OFC5389_ld_r (.Y(FE_OFN12_FE_DBTN0_ld_r),
	.A(FE_OFN1_ld_r));
   BUFx2_ASAP7_75t_L FE_OFC5388_ld_r (.Y(FE_OFN1_ld_r),
	.A(ld_r));
   INVxp33_ASAP7_75t_L FE_OFC5384_n15298 (.Y(FE_OFN28481_n15298),
	.A(n15300));
   INVxp67_ASAP7_75t_L FE_OFC5383_n15298 (.Y(n15300),
	.A(n15298));
   INVx2_ASAP7_75t_SL FE_OFC5379_sa32_3 (.Y(FE_OCPN5129_sa32_3),
	.A(sa32_3_));
   HB1xp67_ASAP7_75t_SL FE_OFC5378_n24719 (.Y(FE_OCPN27361_n24719),
	.A(n24719));
   INVx1_ASAP7_75t_L FE_OFC5377_sa30_7 (.Y(FE_OFN28480_sa30_7),
	.A(n19060));
   INVx1_ASAP7_75t_L FE_OFC5376_sa30_7 (.Y(n19060),
	.A(sa30_7_));
   INVxp33_ASAP7_75t_L FE_OFC5375_n26659 (.Y(n26671),
	.A(FE_OCPN27796_n26659));
   INVx2_ASAP7_75t_SL FE_OFC5370_sa13_2 (.Y(FE_OFN16298_sa13_2),
	.A(sa13_2_));
   INVxp33_ASAP7_75t_R FE_OFC5369_n25672 (.Y(FE_OFN16189_n25672),
	.A(FE_OFN16353_n25672));
   BUFx2_ASAP7_75t_L FE_OFC5368_n25672 (.Y(FE_OFN16353_n25672),
	.A(n25672));
   INVx1_ASAP7_75t_SL FE_OFC5367_sa12_3 (.Y(FE_OCPN27368_sa12_3),
	.A(FE_OCPN29485_sa12_3));
   INVx1_ASAP7_75t_L FE_OFC5365_sa12_3 (.Y(FE_OCPN27429_sa12_3),
	.A(FE_OCPN28135_sa12_3));
   INVx2_ASAP7_75t_L FE_OFC5362_n23307 (.Y(FE_OFN26141_n23307),
	.A(n20753));
   INVx2_ASAP7_75t_R FE_OFC5361_n23307 (.Y(FE_RN_0_0),
	.A(n20753));
   INVx2_ASAP7_75t_SL FE_OFC5360_n23307 (.Y(n20753),
	.A(n23307));
   INVxp33_ASAP7_75t_R FE_OFC5359_n16904 (.Y(n16903),
	.A(n16904));
   INVx2_ASAP7_75t_R FE_OFC5357_n15779 (.Y(FE_OFN25928_n15779),
	.A(n15779));
   BUFx3_ASAP7_75t_SL FE_OFC5356_n15779 (.Y(n15835),
	.A(n15779));
   INVxp67_ASAP7_75t_R FE_OFC5355_n15273 (.Y(n14251),
	.A(n15273));
   INVxp33_ASAP7_75t_R FE_OFC5354_n26684 (.Y(n26690),
	.A(FE_OFN16255_n26684));
   INVxp33_ASAP7_75t_L FE_OFC5353_n26684 (.Y(FE_OFN16255_n26684),
	.A(n26684));
   INVxp33_ASAP7_75t_R FE_OFC5350_n17180 (.Y(n17181),
	.A(n17180));
   INVxp33_ASAP7_75t_R FE_OFC5349_n26806 (.Y(FE_OFN16395_n26801),
	.A(n26806));
   BUFx2_ASAP7_75t_L FE_OFC5348_n18333 (.Y(FE_OCPN27792_n18333),
	.A(n18333));
   INVx3_ASAP7_75t_SL FE_OFC5347_n15380 (.Y(n15956),
	.A(n15380));
   INVxp33_ASAP7_75t_L FE_OFC5346_n18438 (.Y(FE_RN_192_0),
	.A(n18438));
   INVxp67_ASAP7_75t_L FE_OFC5345_n13708 (.Y(n13710),
	.A(n13708));
   INVx1_ASAP7_75t_L FE_OFC5344_FE_OCPN27225_n25357 (.Y(FE_OCPN27226_n25357),
	.A(n20355));
   INVx1_ASAP7_75t_R FE_OFC5343_n26802 (.Y(n26803),
	.A(n26802));
   INVxp33_ASAP7_75t_L FE_OFC5342_n19704 (.Y(FE_OFN16402_n19704),
	.A(n19704));
   INVx2_ASAP7_75t_SL FE_OFC5341_n19170 (.Y(FE_OFN26554_n19170),
	.A(n19170));
   INVxp67_ASAP7_75t_L FE_OFC5340_n25888 (.Y(n25889),
	.A(n25888));
   INVxp33_ASAP7_75t_L FE_OFC5339_FE_OCPN5056_n26535 (.Y(n21496),
	.A(FE_OCPN5056_n26535));
   INVx1_ASAP7_75t_R FE_OFC5338_n23853 (.Y(FE_OFN28477_n23853),
	.A(n20623));
   INVxp33_ASAP7_75t_R FE_OFC5336_FE_OCPN27522_n25921 (.Y(n21264),
	.A(FE_OCPN27522_n25921));
   INVxp33_ASAP7_75t_L FE_OFC5335_n22038 (.Y(n22042),
	.A(n22038));
   INVxp67_ASAP7_75t_L FE_OFC5334_sa21_7 (.Y(FE_OFN167_sa21_7),
	.A(sa21_7_));
   INVxp33_ASAP7_75t_R FE_OFC5332_n24529 (.Y(FE_OFN164_n24529),
	.A(n24529));
   INVxp67_ASAP7_75t_L FE_OFC5331_n22728 (.Y(n22731),
	.A(n22728));
   INVxp67_ASAP7_75t_L FE_OFC5330_n22925 (.Y(FE_OFN26127_n22925),
	.A(n19325));
   INVx1_ASAP7_75t_R FE_OFC5329_n22925 (.Y(n19325),
	.A(n22925));
   INVxp33_ASAP7_75t_L FE_OFC5325_n15093 (.Y(n15094),
	.A(n15093));
   INVx1_ASAP7_75t_R FE_OFC5324_n23573 (.Y(FE_OFN28475_n23573),
	.A(n20544));
   INVxp67_ASAP7_75t_L FE_OFC5323_n23573 (.Y(n20544),
	.A(n23573));
   INVx3_ASAP7_75t_SL FE_OFC5322_sa01_5 (.Y(FE_OCPN28217_sa01_5),
	.A(FE_OCPN27403_sa01_5));
   INVx1_ASAP7_75t_SL FE_OFC5320_sa01_5 (.Y(FE_OCPN27403_sa01_5),
	.A(sa01_5_));
   INVxp33_ASAP7_75t_R FE_OFC5319_FE_OCPN5038_n26735 (.Y(FE_OFN28474_FE_OCPN5038_n26735),
	.A(n26736));
   INVxp67_ASAP7_75t_R FE_OFC5318_FE_OCPN5038_n26735 (.Y(n26736),
	.A(FE_OCPN5038_n26735));
   INVx1_ASAP7_75t_L FE_OFC5317_w3_31 (.Y(n26355),
	.A(FE_OCPN28096_w3_31));
   BUFx4f_ASAP7_75t_SL FE_OFC5316_w3_31 (.Y(FE_OCPN28096_w3_31),
	.A(w3_31_));
   INVx1_ASAP7_75t_SL FE_OFC5315_sa00_0 (.Y(FE_OFN42_sa00_0),
	.A(FE_OCPN27818_n17267));
   BUFx6f_ASAP7_75t_SL FE_OFC5314_sa00_0 (.Y(FE_OCPN27818_n17267),
	.A(sa00_0_));
   INVxp33_ASAP7_75t_R FE_OFC5313_n25701 (.Y(n20286),
	.A(n25701));
   INVxp67_ASAP7_75t_R FE_OFC5311_n22438 (.Y(FE_OFN27064_n22438),
	.A(n22438));
   INVxp33_ASAP7_75t_R FE_OFC5310_n19440 (.Y(n19441),
	.A(n19440));
   INVxp33_ASAP7_75t_R FE_OFC5309_n17053 (.Y(n17054),
	.A(n17053));
   BUFx3_ASAP7_75t_SL FE_OFC5306_n19098 (.Y(FE_OCPN27951_n19098),
	.A(n19098));
   INVxp33_ASAP7_75t_R FE_OFC5305_n18964 (.Y(n18965),
	.A(n18964));
   INVxp67_ASAP7_75t_R FE_OFC5304_sa22_7 (.Y(n22300),
	.A(sa22_7_));
   INVxp67_ASAP7_75t_L FE_OFC5303_n16620 (.Y(n16621),
	.A(n16620));
   INVxp67_ASAP7_75t_L FE_OFC5302_n15808 (.Y(FE_OFN16269_n15808),
	.A(n15808));
   HB1xp67_ASAP7_75t_SL FE_OFC5301_n15808 (.Y(FE_OCPN28398_n15808),
	.A(n15808));
   INVxp67_ASAP7_75t_R FE_OFC5300_n15154 (.Y(n14540),
	.A(n15154));
   INVx1_ASAP7_75t_R FE_OFC5299_n20242 (.Y(FE_OFN25890_n23497),
	.A(n20242));
   INVxp33_ASAP7_75t_R FE_OFC5298_n24208 (.Y(FE_OFN26566_n24208),
	.A(n24208));
   INVx3_ASAP7_75t_SL FE_OFC5293_w3_11 (.Y(FE_OCPN28408_FE_OFN16433_w3_11),
	.A(FE_OFN27115_n));
   INVxp33_ASAP7_75t_R FE_OFC5291_FE_OCPN5053_n25832 (.Y(FE_OFN16324_n25832),
	.A(FE_OCPN5053_n25832));
   INVxp33_ASAP7_75t_L FE_OFC5290_n13511 (.Y(n13280),
	.A(n13511));
   INVxp33_ASAP7_75t_L FE_OFC5289_n26536 (.Y(FE_OFN16275_n26536),
	.A(n26541));
   INVxp33_ASAP7_75t_L FE_OFC5288_n26536 (.Y(n26541),
	.A(n26536));
   INVxp33_ASAP7_75t_L FE_OFC5287_n14630 (.Y(n14133),
	.A(n14630));
   INVx2_ASAP7_75t_L FE_OFC5286_n18750 (.Y(n19836),
	.A(FE_OCPN27843_n18750));
   INVxp33_ASAP7_75t_R FE_OFC5284_n16411 (.Y(n16412),
	.A(n16411));
   INVxp33_ASAP7_75t_R FE_OFC5283_FE_OFN128_sa13_7 (.Y(FE_OFN127_sa13_7),
	.A(FE_OFN128_sa13_7));
   INVx1_ASAP7_75t_SL FE_OFC5282_FE_OFN27206_w3_30 (.Y(FE_OFN27209_w3_30),
	.A(FE_OFN27206_w3_30));
   INVxp33_ASAP7_75t_R FE_OFC5281_n18237 (.Y(n18236),
	.A(n18237));
   INVxp33_ASAP7_75t_R FE_OFC5280_n13870 (.Y(n15473),
	.A(FE_OFN29192_n13870));
   INVxp33_ASAP7_75t_SRAM FE_OFC5279_FE_OCPN5105_n25099 (.Y(n19029),
	.A(FE_OCPN5105_n25099));
   BUFx2_ASAP7_75t_SL FE_OFC5278_n18970 (.Y(FE_OCPN27986_n18970),
	.A(n18970));
   INVxp67_ASAP7_75t_R FE_OFC5277_n24668 (.Y(n26823),
	.A(n24668));
   INVx2_ASAP7_75t_SL FE_OFC5275_FE_OFN6_w3_22 (.Y(FE_OFN26091_n24663),
	.A(n24663));
   INVxp33_ASAP7_75t_R FE_OFC5273_n15888 (.Y(n13757),
	.A(n15888));
   INVxp33_ASAP7_75t_R FE_OFC5272_n14913 (.Y(n14723),
	.A(n14913));
   INVxp33_ASAP7_75t_R FE_OFC5271_n20609 (.Y(n20608),
	.A(n20609));
   INVxp33_ASAP7_75t_R FE_OFC5270_FE_OCPN5131_n25916 (.Y(n22118),
	.A(FE_OCPN5131_n25916));
   INVx1_ASAP7_75t_L FE_OFC5265_FE_OCPN27261_sa02_0 (.Y(FE_OCPN27330_n),
	.A(FE_OCPN27261_sa02_0));
   INVxp33_ASAP7_75t_L FE_OFC5262_n25472 (.Y(n25471),
	.A(n25472));
   INVx1_ASAP7_75t_R FE_OFC5261_n13726 (.Y(n15074),
	.A(n13726));
   INVxp67_ASAP7_75t_L FE_OFC5258_FE_OFN16135_sa22_4 (.Y(n21803),
	.A(FE_PSN8315_FE_OFN16135_sa22_4));
   INVxp67_ASAP7_75t_R FE_OFC5257_n22344 (.Y(n20291),
	.A(n22344));
   INVxp67_ASAP7_75t_SL FE_OFC5256_FE_OFN25959_n23011 (.Y(FE_OFN26585_n23011),
	.A(FE_OFN25959_n23011));
   INVx1_ASAP7_75t_SL FE_OFC5255_FE_OFN25959_n23011 (.Y(FE_OFN26587_n23011),
	.A(FE_OFN25959_n23011));
   INVxp33_ASAP7_75t_SRAM FE_OFC5254_n19355 (.Y(n19354),
	.A(n19355));
   INVx2_ASAP7_75t_SL FE_OFC5253_FE_OCPN28006_n17454 (.Y(n19171),
	.A(FE_OCPN28006_n17454));
   INVxp33_ASAP7_75t_R FE_OFC5251_n13613 (.Y(n13379),
	.A(n13613));
   INVxp33_ASAP7_75t_L FE_OFC5250_n16528 (.Y(n16527),
	.A(n16528));
   INVxp67_ASAP7_75t_R FE_OFC5249_n17732 (.Y(FE_OFN25997_n),
	.A(n17732));
   INVx3_ASAP7_75t_SL FE_OFC5242_n26293 (.Y(n20854),
	.A(n26293));
   BUFx2_ASAP7_75t_SL FE_OFC5241_n22034 (.Y(FE_OCPN28086_n22034),
	.A(n22034));
   INVxp33_ASAP7_75t_SL FE_OFC5240_n25437 (.Y(n23972),
	.A(FE_OCPN27282_n25437));
   BUFx3_ASAP7_75t_SL FE_OFC5239_n25437 (.Y(FE_OCPN27282_n25437),
	.A(n25437));
   INVx1_ASAP7_75t_L FE_OFC5233_n25034 (.Y(FE_OFN25946_sa32_6),
	.A(n25034));
   INVx3_ASAP7_75t_SL FE_OFC5232_n19275 (.Y(n22083),
	.A(FE_OCPN27771_n19275));
   INVx3_ASAP7_75t_SL FE_OFC5231_n19275 (.Y(FE_OCPN27771_n19275),
	.A(n19275));
   INVxp67_ASAP7_75t_R FE_OFC5228_n25711 (.Y(n25712),
	.A(n25711));
   INVx2_ASAP7_75t_R FE_OFC5227_n14971 (.Y(n16026),
	.A(n14971));
   INVxp33_ASAP7_75t_L FE_OFC5226_n22043 (.Y(n19336),
	.A(n22043));
   BUFx6f_ASAP7_75t_SL FE_OFC5225_n17986 (.Y(FE_OCPN27675_n17986),
	.A(n17986));
   BUFx3_ASAP7_75t_SL FE_OFC5224_n16976 (.Y(FE_OCPN27836_n16976),
	.A(n16976));
   INVx5_ASAP7_75t_SL FE_OFC5223_FE_OFN8_w3_14 (.Y(FE_OFN26642_w3_14),
	.A(FE_OFN26636_w3_14));
   INVx2_ASAP7_75t_L FE_OFC5222_FE_OFN8_w3_14 (.Y(FE_OFN26641_w3_14),
	.A(FE_OFN26636_w3_14));
   INVxp67_ASAP7_75t_L FE_OFC5221_FE_OFN8_w3_14 (.Y(FE_OFN26640_w3_14),
	.A(FE_OCPN29535_FE_OFN8_w3_14));
   INVx2_ASAP7_75t_L FE_OFC5220_FE_OFN8_w3_14 (.Y(FE_OFN26639_w3_14),
	.A(FE_OCPN29536_FE_OFN8_w3_14));
   INVxp33_ASAP7_75t_R FE_OFC5219_FE_OFN8_w3_14 (.Y(FE_OFN26638_w3_14),
	.A(FE_OCPN29535_FE_OFN8_w3_14));
   INVxp33_ASAP7_75t_R FE_OFC5218_FE_OFN8_w3_14 (.Y(FE_OFN26637_w3_14),
	.A(FE_OFN16417_n));
   INVx2_ASAP7_75t_SL FE_OFC5217_FE_OFN8_w3_14 (.Y(FE_OFN26636_w3_14),
	.A(FE_OFN16417_n));
   INVx1_ASAP7_75t_L FE_OFC5215_FE_OFN8_w3_14 (.Y(FE_OFN26633_w3_14),
	.A(FE_OFN26635_w3_14));
   INVxp33_ASAP7_75t_L FE_OFC5213_n27008 (.Y(FE_OFN16341_n27008),
	.A(n27008));
   INVxp33_ASAP7_75t_R FE_OFC5210_n17489 (.Y(FE_RN_8_0),
	.A(n17489));
   INVx1_ASAP7_75t_SL FE_OFC5209_n21677 (.Y(n20624),
	.A(n21677));
   INVx1_ASAP7_75t_L FE_OFC5208_n24590 (.Y(FE_OFN165_sa12_7),
	.A(n24590));
   INVx1_ASAP7_75t_SL FE_OFC5206_n16331 (.Y(FE_OFN26550_n16331),
	.A(n16331));
   INVx2_ASAP7_75t_R FE_OFC5204_ld (.Y(FE_OFN28472_ld),
	.A(FE_OFN28466_ld));
   INVx1_ASAP7_75t_L FE_OFC5203_ld (.Y(FE_OFN28471_ld),
	.A(FE_OFN28466_ld));
   INVx2_ASAP7_75t_R FE_OFC5202_ld (.Y(FE_OFN28470_ld),
	.A(FE_OFN28465_ld));
   INVx1_ASAP7_75t_R FE_OFC5201_ld (.Y(FE_OFN28469_ld),
	.A(FE_OFN28465_ld));
   HB1xp67_ASAP7_75t_R FE_OFC5200_ld (.Y(FE_OFN28468_ld),
	.A(FE_OFN28461_ld));
   HB1xp67_ASAP7_75t_R FE_OFC5199_ld (.Y(FE_OFN28467_ld),
	.A(FE_OFN28461_ld));
   INVxp33_ASAP7_75t_L FE_OFC5198_ld (.Y(FE_OFN28466_ld),
	.A(FE_OFN28460_ld));
   INVxp33_ASAP7_75t_L FE_OFC5197_ld (.Y(FE_OFN28465_ld),
	.A(FE_OFN26139_n16125));
   HB1xp67_ASAP7_75t_R FE_OFC5196_ld (.Y(FE_OFN28464_ld),
	.A(FE_OFN27_n16125));
   HB1xp67_ASAP7_75t_R FE_OFC5195_ld (.Y(FE_OFN28463_ld),
	.A(FE_OFN25_n16125));
   BUFx2_ASAP7_75t_R FE_OFC5194_ld (.Y(FE_OFN28462_ld),
	.A(FE_OFN25_n16125));
   INVxp67_ASAP7_75t_L FE_OFC5193_ld (.Y(FE_OFN28461_ld),
	.A(FE_OFN26137_n16125));
   INVx1_ASAP7_75t_L FE_OFC5192_ld (.Y(FE_OFN28460_ld),
	.A(FE_OFN26137_n16125));
   INVx1_ASAP7_75t_R FE_OFC5191_ld (.Y(FE_OFN28459_ld),
	.A(FE_OFN24_n16125));
   INVx1_ASAP7_75t_R FE_OFC5190_ld (.Y(FE_OFN28458_ld),
	.A(FE_OFN24_n16125));
   INVx2_ASAP7_75t_SRAM FE_OFC5189_ld (.Y(FE_OFN28457_ld),
	.A(FE_OFN23_n16125));
   INVx1_ASAP7_75t_R FE_OFC5188_ld (.Y(FE_OFN26139_n16125),
	.A(FE_OFN23_n16125));
   INVx2_ASAP7_75t_SRAM FE_OFC5186_ld (.Y(FE_OFN27_n16125),
	.A(FE_OFN23_n16125));
   INVx2_ASAP7_75t_R FE_OFC5185_ld (.Y(FE_OFN26_n16125),
	.A(FE_OFN23_n16125));
   INVx2_ASAP7_75t_R FE_OFC5184_ld (.Y(FE_OFN25_n16125),
	.A(FE_OFN23_n16125));
   INVxp33_ASAP7_75t_L FE_OFC5183_ld (.Y(FE_OFN26137_n16125),
	.A(FE_OFN20_n16125));
   INVxp33_ASAP7_75t_L FE_OFC5182_ld (.Y(FE_OFN24_n16125),
	.A(FE_OFN19_n16125));
   INVx1_ASAP7_75t_R FE_OFC5181_ld (.Y(FE_OFN23_n16125),
	.A(FE_OFN19_n16125));
   INVx2_ASAP7_75t_R FE_OFC5180_ld (.Y(FE_OFN21_n16125),
	.A(FE_OFN18_n16125));
   INVxp33_ASAP7_75t_SRAM FE_OFC5179_ld (.Y(FE_OFN20_n16125),
	.A(ld));
   INVx1_ASAP7_75t_SRAM FE_OFC5178_ld (.Y(FE_OFN19_n16125),
	.A(ld));
   INVxp33_ASAP7_75t_SRAM FE_OFC5177_ld (.Y(FE_OFN18_n16125),
	.A(ld));
   BUFx2_ASAP7_75t_SRAM FE_OFC5176_ld (.Y(n16125),
	.A(ld));
   HB1xp67_ASAP7_75t_SRAM FE_OFC5175_ld (.Y(FE_OFN0_ld),
	.A(ld));
   INVx1_ASAP7_75t_SL FE_OFC5173_n18871 (.Y(FE_OCPN27975_n18871),
	.A(n18871));
   INVx2_ASAP7_75t_SL FE_OFC5169_FE_OCPN27557_sa20_4 (.Y(n20636),
	.A(FE_OCPN27558_sa20_4));
   INVx3_ASAP7_75t_SL FE_OFC5168_FE_OCPN27557_sa20_4 (.Y(FE_OCPN27558_sa20_4),
	.A(FE_OFN16229_sa20_4));
   INVxp67_ASAP7_75t_SL FE_OFC5165_n21643 (.Y(n21225),
	.A(n21643));
   INVx1_ASAP7_75t_L FE_OFC5164_n21643 (.Y(FE_OCPN27531_n21643),
	.A(n21643));
   INVx1_ASAP7_75t_L FE_OFC5162_n18506 (.Y(n24127),
	.A(n18506));
   INVxp33_ASAP7_75t_L FE_OFC5161_n20593 (.Y(n19526),
	.A(n20593));
   INVx1_ASAP7_75t_SL FE_OFC5158_n13348 (.Y(FE_OFN28455_n13348),
	.A(n14535));
   INVxp67_ASAP7_75t_L FE_OFC5156_n13348 (.Y(FE_OFN28453_n13348),
	.A(FE_OFN28454_n13348));
   INVxp67_ASAP7_75t_R FE_OFC5152_FE_OFN16159_w3_24 (.Y(FE_OFN25881_w3_24),
	.A(FE_OFN25880_w3_24));
   INVxp67_ASAP7_75t_L FE_OFC5151_FE_OFN16159_w3_24 (.Y(FE_OFN25880_w3_24),
	.A(FE_OFN16159_w3_24));
   INVxp33_ASAP7_75t_R FE_OFC5150_n23467 (.Y(FE_RN_38_0),
	.A(n23467));
   BUFx2_ASAP7_75t_SL FE_OFC5149_n17170 (.Y(FE_OCPN28137_n17170),
	.A(n17170));
   INVx1_ASAP7_75t_R FE_OFC5148_n17170 (.Y(n17002),
	.A(n17170));
   INVx1_ASAP7_75t_L FE_OFC5147_n16789 (.Y(FE_OCPN27454_n16789),
	.A(n19884));
   INVx2_ASAP7_75t_SL FE_OFC5146_n16789 (.Y(n19884),
	.A(n16789));
   INVx2_ASAP7_75t_L FE_OFC5145_n22224 (.Y(n24367),
	.A(FE_OFN26158_n22224));
   BUFx3_ASAP7_75t_SL FE_OFC5144_n22224 (.Y(FE_OFN26158_n22224),
	.A(n22224));
   INVxp67_ASAP7_75t_L FE_OFC5143_FE_OFN16131_sa12_1 (.Y(FE_OCPN27804_sa12_1),
	.A(FE_OFN26589_sa12_1));
   INVxp67_ASAP7_75t_R FE_OFC5142_FE_OFN16131_sa12_1 (.Y(FE_OFN26589_sa12_1),
	.A(FE_OFN28764_n17928));
   BUFx3_ASAP7_75t_SL FE_OFC5139_n23600 (.Y(FE_OCPN5137_n23600),
	.A(n23600));
   INVx2_ASAP7_75t_L FE_OFC5138_n19005 (.Y(FE_OCPN27881_FE_OFN27126_sa23_3),
	.A(FE_OFN27127_sa23_3));
   INVx2_ASAP7_75t_L FE_OFC5131_n16438 (.Y(FE_OFN27062_n16438),
	.A(FE_OCPN27568_sa33_3));
   INVx5_ASAP7_75t_SL FE_OFC5130_n16438 (.Y(FE_OCPN27568_sa33_3),
	.A(n16438));
   INVx2_ASAP7_75t_SL FE_OFC5129_n16438 (.Y(FE_OFN25938_sa33_3),
	.A(n16438));
   INVx1_ASAP7_75t_SL FE_OFC5126_w3_29 (.Y(FE_OFN27131_w3_29),
	.A(w3_29_));
   INVxp67_ASAP7_75t_L FE_OFC5118_n15506 (.Y(n15735),
	.A(FE_OFN72_n15506));
   INVx1_ASAP7_75t_L FE_OFC5117_n15506 (.Y(FE_OFN72_n15506),
	.A(n15506));
   INVx1_ASAP7_75t_L FE_OFC5116_n13671 (.Y(FE_OFN26059_n),
	.A(FE_OFN16451_n));
   INVx1_ASAP7_75t_SL FE_OFC5115_n13671 (.Y(FE_OFN27085_n),
	.A(n15224));
   INVx1_ASAP7_75t_L FE_OFC5114_n13671 (.Y(FE_OFN16451_n),
	.A(n15224));
   BUFx2_ASAP7_75t_SL FE_OFC5113_n13671 (.Y(n15224),
	.A(n13671));
   INVx1_ASAP7_75t_SL FE_OFC5112_n16271 (.Y(n16272),
	.A(n16271));
   INVx2_ASAP7_75t_L FE_OFC5111_n27179 (.Y(FE_OFN104_n27179),
	.A(n27177));
   BUFx3_ASAP7_75t_SL FE_OFC5110_n27179 (.Y(n27177),
	.A(n27179));
   BUFx2_ASAP7_75t_SL FE_OFC5108_n25483 (.Y(FE_OCPN27467_n25483),
	.A(n25483));
   INVx1_ASAP7_75t_L FE_OFC5107_n16050 (.Y(FE_OFN16360_n16051),
	.A(n16050));
   INVxp67_ASAP7_75t_R FE_OFC5106_FE_OFN27133_n21725 (.Y(n18867),
	.A(FE_OFN27133_n21725));
   INVxp67_ASAP7_75t_L FE_OFC5104_n20369 (.Y(FE_OFN26575_n20369),
	.A(n20369));
   HB1xp67_ASAP7_75t_L FE_OFC5103_n26335 (.Y(FE_OCPN28110_n),
	.A(n26335));
   INVxp33_ASAP7_75t_L FE_OFC5102_w3_7 (.Y(FE_OFN25979_n),
	.A(FE_OCPN29501_FE_OFN28662_w3_7));
   INVxp67_ASAP7_75t_L FE_OFC5100_n18759 (.Y(n17273),
	.A(n18759));
   INVx2_ASAP7_75t_SL FE_OFC5098_sa22_5 (.Y(n18164),
	.A(sa22_5_));
   INVxp67_ASAP7_75t_L FE_OFC5095_n23302 (.Y(FE_OFN26528_n23302),
	.A(FE_OCPN29305_n23302));
   INVx1_ASAP7_75t_SL FE_OFC5093_n22995 (.Y(n22952),
	.A(FE_OFN27056_n22995));
   BUFx3_ASAP7_75t_SL FE_OFC5092_n22995 (.Y(FE_OFN27056_n22995),
	.A(n22995));
   INVxp33_ASAP7_75t_R FE_OFC5091_n25020 (.Y(n25021),
	.A(n25020));
   INVx1_ASAP7_75t_SL FE_OFC5087_n25407 (.Y(FE_OCPN27519_n25407),
	.A(n25407));
   INVxp33_ASAP7_75t_L FE_OFC5086_sa02_5 (.Y(FE_OCPN27579_FE_OFN16138_sa02_5),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5));
   INVx2_ASAP7_75t_L FE_OFC5081_sa33_1 (.Y(n16423),
	.A(FE_OFN28727_sa33_1));
   INVx2_ASAP7_75t_SL FE_OFC5080_FE_OCPN27978_w3_3 (.Y(FE_OFN25887_w3_3),
	.A(FE_OFN26591_w3_3));
   INVx2_ASAP7_75t_SL FE_OFC5079_FE_OCPN27978_w3_3 (.Y(FE_OFN26591_w3_3),
	.A(FE_OFN25886_w3_3));
   INVx3_ASAP7_75t_SL FE_OFC5078_FE_OCPN27978_w3_3 (.Y(n25140),
	.A(FE_OCPN27978_w3_3));
   INVx3_ASAP7_75t_SL FE_OFC5075_sa13_5 (.Y(n16981),
	.A(sa13_5_));
   INVx1_ASAP7_75t_R FE_OFC5059_sa01_0 (.Y(FE_OCPN27810_n),
	.A(FE_OCPN27423_sa01_0));
   BUFx6f_ASAP7_75t_SL FE_OFC5058_sa01_0 (.Y(FE_OCPN27423_sa01_0),
	.A(sa01_0_));
   INVx2_ASAP7_75t_L FE_OFC5057_sa01_1 (.Y(FE_OFN125_sa01_1),
	.A(sa01_1_));
   BUFx2_ASAP7_75t_SL FE_OFC5056_sa33_5 (.Y(FE_OFN26055_n),
	.A(FE_OFN28679_sa33_5));
   INVx2_ASAP7_75t_R FE_OFC5054_FE_OFN21730_sa03_3 (.Y(FE_OFN27125_n21057),
	.A(FE_OFN21730_sa03_3));
   INVx2_ASAP7_75t_L FE_OFC5051_FE_OFN16452_sa30_1 (.Y(n18379),
	.A(FE_OFN16247_sa30_1));
   INVxp67_ASAP7_75t_L FE_OFC5049_sa33_4 (.Y(FE_OCPN27546_sa33_4),
	.A(FE_OCPN27544_sa33_4));
   INVx2_ASAP7_75t_SL FE_OFC5043_sa32_2 (.Y(FE_OFN16128_sa32_2),
	.A(sa32_2_));
   INVx8_ASAP7_75t_SL FE_OFC5038_w3_19 (.Y(FE_OFN26053_n25415),
	.A(FE_OFN26539_w3_19));
   INVx5_ASAP7_75t_SL FE_OFC5034_w3_19 (.Y(FE_OFN26539_w3_19),
	.A(FE_OCPN28093_FE_OFN26534_w3_19));
   INVx2_ASAP7_75t_SL FE_OFC5031_w3_19 (.Y(FE_OCPN28093_FE_OFN26534_w3_19),
	.A(FE_OFN27096_n));
   INVxp33_ASAP7_75t_R FE_OFC5027_sa31_5 (.Y(FE_OFN16315_sa31_5),
	.A(FE_OFN28669_sa31_5));
   INVx1_ASAP7_75t_SL FE_OFC5026_sa31_5 (.Y(FE_OFN26107_sa31_5),
	.A(FE_OFN28669_sa31_5));
   INVxp33_ASAP7_75t_R FE_OFC5025_FE_OCPN27740_sa02_4 (.Y(FE_OCPN28158_n),
	.A(n17760));
   INVx3_ASAP7_75t_SL FE_OFC5023_sa13_0 (.Y(n16982),
	.A(FE_OFN26600_sa13_0));
   INVx2_ASAP7_75t_SL FE_OFC5022_sa13_0 (.Y(FE_OFN26600_sa13_0),
	.A(sa13_0_));
   AOI31xp33_ASAP7_75t_SL FE_RC_750_0 (.Y(n25066),
	.A1(n20400),
	.A2(FE_OFN28558_n23073),
	.A3(n26457),
	.B(n27015));
   AOI31xp33_ASAP7_75t_SL FE_RC_749_0 (.Y(n25564),
	.A1(n25561),
	.A2(n25887),
	.A3(n25562),
	.B(n27095));
   AOI21xp5_ASAP7_75t_SL FE_RC_747_0 (.Y(n15444),
	.A1(FE_OFN26642_w3_14),
	.A2(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(n15927));
   AOI21xp5_ASAP7_75t_L FE_RC_746_0 (.Y(n18058),
	.A1(n25038),
	.A2(n26819),
	.B(n23941));
   AOI31xp67_ASAP7_75t_SL FE_RC_744_0 (.Y(n21078),
	.A1(FE_RN_233_0),
	.A2(n21076),
	.A3(n21077),
	.B(n25420));
   AOI31xp33_ASAP7_75t_L FE_RC_742_0 (.Y(n22476),
	.A1(FE_RN_232_0),
	.A2(n22455),
	.A3(n22456),
	.B(n27004));
   AOI31xp33_ASAP7_75t_L FE_RC_741_0 (.Y(n23115),
	.A1(n23096),
	.A2(n23095),
	.A3(n23097),
	.B(n27004));
   AOI31xp33_ASAP7_75t_L FE_RC_740_0 (.Y(n20534),
	.A1(n20532),
	.A2(n20531),
	.A3(n20533),
	.B(n26959));
   AOI31xp33_ASAP7_75t_L FE_RC_739_0 (.Y(n18852),
	.A1(n18850),
	.A2(n18849),
	.A3(n18851),
	.B(n17584));
   AOI31xp33_ASAP7_75t_SL FE_RC_738_0 (.Y(n19690),
	.A1(n19688),
	.A2(n19687),
	.A3(n19689),
	.B(n24978));
   AOI31xp33_ASAP7_75t_SL FE_RC_736_0 (.Y(n22967),
	.A1(FE_OFN27127_sa23_3),
	.A2(FE_OCPN27482_sa23_5),
	.A3(FE_OCPN29480_n20913),
	.B(n19006));
   AOI21xp33_ASAP7_75t_SL FE_RC_735_0 (.Y(n17255),
	.A1(n19609),
	.A2(FE_OCPN29346_n12998),
	.B(n19605));
   AOI21xp5_ASAP7_75t_SL FE_RC_734_0 (.Y(n20415),
	.A1(n26454),
	.A2(n17321),
	.B(n22582));
   AOI21xp5_ASAP7_75t_SL FE_RC_733_0 (.Y(n20075),
	.A1(n20868),
	.A2(n16299),
	.B(n21963));
   AOI21xp5_ASAP7_75t_SL FE_RC_732_0 (.Y(n19423),
	.A1(FE_OFN16162_n25869),
	.A2(FE_OFN28801_n16978),
	.B(n20491));
   AOI31xp33_ASAP7_75t_SL FE_RC_731_0 (.Y(n15430),
	.A1(n13844),
	.A2(FE_OFN28848_n14912),
	.A3(FE_OFN28884_n),
	.B(n14927));
   AOI21xp5_ASAP7_75t_SL FE_RC_730_0 (.Y(n18639),
	.A1(n21154),
	.A2(FE_OCPN28389_n21479),
	.B(n19836));
   AOI21xp33_ASAP7_75t_R FE_RC_729_0 (.Y(n19879),
	.A1(FE_OFN28778_FE_OCPN28352_n16748),
	.A2(FE_OFN16447_n16749),
	.B(n23925));
   AOI21xp33_ASAP7_75t_L FE_RC_728_0 (.Y(n19043),
	.A1(FE_OFN28818_n17602),
	.A2(n17606),
	.B(n22641));
   AOI21xp5_ASAP7_75t_L FE_RC_727_0 (.Y(n15507),
	.A1(n15694),
	.A2(FE_OCPN27928_FE_OFN4_w3_22),
	.B(n13868));
   XOR2xp5_ASAP7_75t_SL FE_RC_726_0 (.Y(n26783),
	.A(n26780),
	.B(FE_RN_35_0));
   XOR2x1_ASAP7_75t_SL FE_RC_725_0 (.Y(n25812),
	.A(FE_OCPN27321_n26380),
	.B(FE_RN_44_0));
   XOR2xp5_ASAP7_75t_SL FE_RC_724_0 (.Y(n25664),
	.A(FE_OCPN27430_n26334),
	.B(FE_RN_58_0));
   XNOR2xp5_ASAP7_75t_SL FE_RC_722_0 (.Y(FE_RN_35_0),
	.A(n26779),
	.B(n26778));
   XNOR2x1_ASAP7_75t_SL FE_RC_721_0 (.Y(FE_RN_44_0),
	.A(n25810),
	.B(n25809));
   XNOR2xp5_ASAP7_75t_SL FE_RC_720_0 (.Y(FE_RN_58_0),
	.A(n25660),
	.B(n25661));
   INVxp33_ASAP7_75t_L FE_RC_719_0 (.Y(FE_RN_231_0),
	.A(n27091));
   AOI21x1_ASAP7_75t_SL FE_RC_717_0 (.Y(n24511),
	.A1(n24113),
	.A2(n27117),
	.B(n24114));
   AOI31xp67_ASAP7_75t_L FE_RC_716_0 (.Y(n20536),
	.A1(n20504),
	.A2(FE_OCPN5062_n20505),
	.A3(n24166),
	.B(n27095));
   AOI21xp5_ASAP7_75t_SL FE_RC_715_0 (.Y(n23565),
	.A1(n23563),
	.A2(n26770),
	.B(n23564));
   AOI21x1_ASAP7_75t_SL FE_RC_714_0 (.Y(n25805),
	.A1(n26226),
	.A2(FE_OFN16170_n26637),
	.B(n26222));
   AOI31xp33_ASAP7_75t_L FE_RC_713_0 (.Y(n21696),
	.A1(n21694),
	.A2(n23776),
	.A3(n21695),
	.B(n25641));
   AOI31xp33_ASAP7_75t_SL FE_RC_712_0 (.Y(n21335),
	.A1(n21333),
	.A2(n21332),
	.A3(n21334),
	.B(n23467));
   AOI31xp67_ASAP7_75t_L FE_RC_711_0 (.Y(n22324),
	.A1(n22323),
	.A2(n22322),
	.A3(n24699),
	.B(n23345));
   AOI31xp33_ASAP7_75t_SL FE_RC_710_0 (.Y(n15258),
	.A1(n15257),
	.A2(n15255),
	.A3(n15254),
	.B(n15256));
   AOI31xp33_ASAP7_75t_L FE_RC_709_0 (.Y(n22788),
	.A1(n22787),
	.A2(n22786),
	.A3(n25395),
	.B(n24377));
   AOI31xp33_ASAP7_75t_L FE_RC_708_0 (.Y(n21760),
	.A1(n21749),
	.A2(n21748),
	.A3(n21750),
	.B(n23945));
   AOI31xp33_ASAP7_75t_SL FE_RC_707_0 (.Y(n23890),
	.A1(n23868),
	.A2(n23867),
	.A3(n25628),
	.B(n25641));
   AOI31xp33_ASAP7_75t_L FE_RC_706_0 (.Y(n23198),
	.A1(n23196),
	.A2(n23195),
	.A3(FE_PSN8301_n23197),
	.B(n23345));
   AOI31xp67_ASAP7_75t_SL FE_RC_705_0 (.Y(n22325),
	.A1(n22315),
	.A2(n22314),
	.A3(n22316),
	.B(n26889));
   AOI31xp33_ASAP7_75t_SL FE_RC_704_0 (.Y(n22607),
	.A1(n22605),
	.A2(n22604),
	.A3(n22606),
	.B(n26464));
   AOI31xp33_ASAP7_75t_L FE_RC_703_0 (.Y(n20945),
	.A1(n20944),
	.A2(n20943),
	.A3(n26151),
	.B(n26710));
   AOI31xp67_ASAP7_75t_SL FE_RC_702_0 (.Y(n25158),
	.A1(n23232),
	.A2(n23231),
	.A3(n23233),
	.B(n24377));
   AOI31xp67_ASAP7_75t_SL FE_RC_700_0 (.Y(n23906),
	.A1(n21522),
	.A2(FE_OCPN7644_n21523),
	.A3(n21521),
	.B(n25420));
   AOI31xp33_ASAP7_75t_SL FE_RC_699_0 (.Y(n24399),
	.A1(n20397),
	.A2(n22474),
	.A3(n18728),
	.B(n27004));
   AOI31xp33_ASAP7_75t_SL FE_RC_696_0 (.Y(n26031),
	.A1(n22154),
	.A2(n22153),
	.A3(n22155),
	.B(n26687));
   AOI31xp33_ASAP7_75t_SL FE_RC_694_0 (.Y(n23904),
	.A1(FE_RN_230_0),
	.A2(n21516),
	.A3(n21517),
	.B(n23467));
   AOI31xp67_ASAP7_75t_L FE_RC_693_0 (.Y(n24226),
	.A1(n17368),
	.A2(n17367),
	.A3(FE_OCPN29330_n26459),
	.B(n26464));
   AOI31xp33_ASAP7_75t_SL FE_RC_692_0 (.Y(n19566),
	.A1(n20543),
	.A2(n19564),
	.A3(n19565),
	.B(n24377));
   AOI31xp33_ASAP7_75t_SL FE_RC_690_0 (.Y(n14079),
	.A1(n14059),
	.A2(n14058),
	.A3(n14060),
	.B(n13901));
   AOI31xp33_ASAP7_75t_SL FE_RC_688_0 (.Y(n22959),
	.A1(n22958),
	.A2(n22957),
	.A3(n26553),
	.B(n27027));
   AOI31xp33_ASAP7_75t_SL FE_RC_687_0 (.Y(n18907),
	.A1(n18906),
	.A2(n18905),
	.A3(n21277),
	.B(n23945));
   AOI31xp33_ASAP7_75t_SL FE_RC_686_0 (.Y(n22052),
	.A1(n22050),
	.A2(n22049),
	.A3(n22051),
	.B(n26571));
   AOI31xp67_ASAP7_75t_SL FE_RC_685_0 (.Y(n26003),
	.A1(n18945),
	.A2(n25887),
	.A3(n18944),
	.B(n27102));
   AOI31xp33_ASAP7_75t_SL FE_RC_683_0 (.Y(n22263),
	.A1(n22249),
	.A2(n24587),
	.A3(n22246),
	.B(n26607));
   AOI31xp33_ASAP7_75t_SL FE_RC_682_0 (.Y(n22113),
	.A1(n22111),
	.A2(n22110),
	.A3(n22112),
	.B(n27140));
   AOI31xp33_ASAP7_75t_L FE_RC_681_0 (.Y(n21260),
	.A1(n21259),
	.A2(n21258),
	.A3(n23832),
	.B(n25641));
   AOI31xp33_ASAP7_75t_SL FE_RC_680_0 (.Y(n21430),
	.A1(n22487),
	.A2(n21428),
	.A3(n21429),
	.B(n17463));
   AOI31xp33_ASAP7_75t_SL FE_RC_679_0 (.Y(n18292),
	.A1(n18281),
	.A2(n18280),
	.A3(n18282),
	.B(n26959));
   AOI31xp33_ASAP7_75t_SL FE_RC_678_0 (.Y(n23347),
	.A1(n23344),
	.A2(n23343),
	.A3(n23346),
	.B(n23345));
   AOI31xp33_ASAP7_75t_L FE_RC_677_0 (.Y(n19080),
	.A1(n19071),
	.A2(n19070),
	.A3(n22631),
	.B(n26926));
   AOI31xp67_ASAP7_75t_SL FE_RC_675_0 (.Y(n25610),
	.A1(n24488),
	.A2(n24487),
	.A3(n24489),
	.B(n26542));
   AOI31xp33_ASAP7_75t_SL FE_RC_674_0 (.Y(n20122),
	.A1(n20115),
	.A2(n20114),
	.A3(n20116),
	.B(n17584));
   AOI31xp33_ASAP7_75t_SL FE_RC_673_0 (.Y(n25819),
	.A1(n18092),
	.A2(n21935),
	.A3(n21924),
	.B(n26315));
   AOI31xp33_ASAP7_75t_L FE_RC_672_0 (.Y(n24003),
	.A1(n24001),
	.A2(n24000),
	.A3(n24002),
	.B(n24978));
   AOI31xp67_ASAP7_75t_SL FE_RC_671_0 (.Y(n14811),
	.A1(n13867),
	.A2(FE_OFN27096_n),
	.A3(n15729),
	.B(n14810));
   AOI31xp33_ASAP7_75t_SL FE_RC_670_0 (.Y(n19855),
	.A1(n19854),
	.A2(n19852),
	.A3(n19853),
	.B(n26777));
   AOI31xp33_ASAP7_75t_L FE_RC_669_0 (.Y(n23911),
	.A1(n21531),
	.A2(n21529),
	.A3(n21530),
	.B(n23945));
   AOI31xp33_ASAP7_75t_SL FE_RC_668_0 (.Y(n21914),
	.A1(n21913),
	.A2(n21911),
	.A3(n21912),
	.B(n25139));
   AOI21xp5_ASAP7_75t_SL FE_RC_667_0 (.Y(n18485),
	.A1(FE_PSN8308_n22624),
	.A2(n18463),
	.B(n18363));
   AOI31xp33_ASAP7_75t_L FE_RC_666_0 (.Y(n17518),
	.A1(n17480),
	.A2(n17479),
	.A3(n17481),
	.B(n17463));
   AOI31xp33_ASAP7_75t_SL FE_RC_665_0 (.Y(n23520),
	.A1(n23518),
	.A2(n23517),
	.A3(n23519),
	.B(n27027));
   AOI31xp67_ASAP7_75t_SL FE_RC_664_0 (.Y(n19543),
	.A1(FE_OCPN8265_n24362),
	.A2(FE_OCPN27804_sa12_1),
	.A3(FE_OCPN28386_n17899),
	.B(n17962));
   AOI21xp33_ASAP7_75t_SL FE_RC_663_0 (.Y(n23872),
	.A1(n23855),
	.A2(FE_OFN29251_n18536),
	.B(n23764));
   AOI21xp5_ASAP7_75t_SL FE_RC_662_0 (.Y(n16679),
	.A1(FE_OFN28998_n16923),
	.A2(n16479),
	.B(n16466));
   AOI21xp5_ASAP7_75t_SL FE_RC_661_0 (.Y(n20497),
	.A1(FE_OFN16396_n25869),
	.A2(FE_OCPN27859_n25868),
	.B(n19374));
   AOI31xp33_ASAP7_75t_SL FE_RC_660_0 (.Y(n15345),
	.A1(n12994),
	.A2(FE_OCPN27928_FE_OFN4_w3_22),
	.A3(n15536),
	.B(n15344));
   AOI31xp33_ASAP7_75t_SL FE_RC_659_0 (.Y(n16791),
	.A1(FE_OFN62_sa21_3),
	.A2(FE_OCPN27289_sa21_5),
	.A3(FE_OFN25993_n16767),
	.B(n16809));
   AOI31xp33_ASAP7_75t_SL FE_RC_658_0 (.Y(n14887),
	.A1(n15046),
	.A2(n14850),
	.A3(n15585),
	.B(n15881));
   AOI31xp33_ASAP7_75t_L FE_RC_657_0 (.Y(n13621),
	.A1(n13592),
	.A2(n13591),
	.A3(n13593),
	.B(n14585));
   AOI31xp33_ASAP7_75t_L FE_RC_656_0 (.Y(n22294),
	.A1(FE_OCPN27722_n23336),
	.A2(FE_OCPN27673_n18163),
	.A3(FE_OCPN27750_n22293),
	.B(n22292));
   AOI31xp33_ASAP7_75t_SL FE_RC_655_0 (.Y(n20397),
	.A1(FE_OCPN27988_n26454),
	.A2(FE_OFN16141_sa01_3),
	.A3(FE_OCPN27871_n17317),
	.B(n21544));
   AOI21xp5_ASAP7_75t_L FE_RC_654_0 (.Y(n21291),
	.A1(FE_OFN28589_n21048),
	.A2(FE_OCPN27617_n18016),
	.B(n23413));
   AOI21xp5_ASAP7_75t_L FE_RC_653_0 (.Y(n23598),
	.A1(n23208),
	.A2(FE_OCPN27429_sa12_3),
	.B(n22255));
   AOI21xp5_ASAP7_75t_L FE_RC_652_0 (.Y(n17482),
	.A1(FE_OCPN27562_n17447),
	.A2(n19206),
	.B(n19229));
   AOI31xp33_ASAP7_75t_L FE_RC_651_0 (.Y(n22012),
	.A1(FE_OCPN27727_n22964),
	.A2(FE_OCPN27627_sa23_1),
	.A3(n18971),
	.B(n22008));
   AOI31xp33_ASAP7_75t_SL FE_RC_650_0 (.Y(n15646),
	.A1(n15590),
	.A2(n15593),
	.A3(n15594),
	.B(FE_OFN28682_n15888));
   AOI21xp33_ASAP7_75t_L FE_RC_649_0 (.Y(n18595),
	.A1(FE_OFN29140_n18527),
	.A2(FE_OFN27083_n),
	.B(FE_OFN26150_n21253));
   AOI21xp5_ASAP7_75t_L FE_RC_648_0 (.Y(n23414),
	.A1(FE_OCPN28214_n21500),
	.A2(FE_OCPN27617_n18016),
	.B(n17989));
   AOI21xp5_ASAP7_75t_SL FE_RC_647_0 (.Y(n26451),
	.A1(n23059),
	.A2(FE_OCPN27988_n26454),
	.B(n23062));
   AOI21xp5_ASAP7_75t_SL FE_RC_646_0 (.Y(n21002),
	.A1(n20982),
	.A2(FE_OFN28812_FE_OCPN27261_sa02_0),
	.B(n22060));
   AOI31xp33_ASAP7_75t_SL FE_RC_645_0 (.Y(n13278),
	.A1(n13643),
	.A2(n15224),
	.A3(FE_OFN28496_n15201),
	.B(n13276));
   AOI31xp67_ASAP7_75t_SL FE_RC_644_0 (.Y(n18825),
	.A1(FE_OCPN28245_n),
	.A2(FE_OFN69_sa32_4),
	.A3(n19938),
	.B(n17689));
   AOI31xp33_ASAP7_75t_SL FE_RC_643_0 (.Y(n19873),
	.A1(FE_OFN29023_n16750),
	.A2(FE_OFN29066_FE_OCPN27328_sa21_2),
	.A3(FE_OCPN29418_n),
	.B(n20005));
   AOI31xp67_ASAP7_75t_L FE_RC_642_0 (.Y(n19096),
	.A1(FE_OFN28835_n),
	.A2(FE_OCPN29370_FE_OFN28744),
	.A3(FE_OCPN27819_n17245),
	.B(n21163));
   AOI31xp33_ASAP7_75t_SL FE_RC_641_0 (.Y(n16525),
	.A1(FE_OFN26060_sa31_4),
	.A2(n20868),
	.A3(FE_OCPN29483_FE_OFN26014_sa31_3),
	.B(n21964));
   AOI21xp5_ASAP7_75t_L FE_RC_640_0 (.Y(n17146),
	.A1(n25869),
	.A2(n25868),
	.B(n17082));
   AOI21xp33_ASAP7_75t_L FE_RC_639_0 (.Y(n22134),
	.A1(FE_OFN25901_n22133),
	.A2(n21625),
	.B(n21604));
   AOI21xp5_ASAP7_75t_L FE_RC_638_0 (.Y(n16341),
	.A1(FE_OCPN27516_n26292),
	.A2(n21989),
	.B(n16306));
   AOI21xp5_ASAP7_75t_SL FE_RC_637_0 (.Y(n22689),
	.A1(FE_OFN28778_FE_OCPN28352_n16748),
	.A2(FE_OCPN28298_n),
	.B(n20325));
   AOI21xp5_ASAP7_75t_L FE_RC_636_0 (.Y(n18472),
	.A1(n17602),
	.A2(n25108),
	.B(n22614));
   AOI21xp5_ASAP7_75t_L FE_RC_635_0 (.Y(n18861),
	.A1(FE_OCPN8247_n21317),
	.A2(FE_OFN29158_n18860),
	.B(n23455));
   AOI21xp5_ASAP7_75t_SL FE_RC_634_0 (.Y(n19386),
	.A1(FE_OFN28801_n16978),
	.A2(n19376),
	.B(n18919));
   AOI21x1_ASAP7_75t_SL FE_RC_633_0 (.Y(n20258),
	.A1(n19019),
	.A2(FE_OFN29003_n23491),
	.B(n23472));
   AOI31xp33_ASAP7_75t_L FE_RC_632_0 (.Y(n20051),
	.A1(FE_OCPN27444_n20064),
	.A2(FE_OFN29016_n16512),
	.A3(n16493),
	.B(n25319));
   AOI31xp33_ASAP7_75t_SL FE_RC_631_0 (.Y(n18871),
	.A1(n21500),
	.A2(n18016),
	.A3(FE_OCPN5195_FE_OFN25874_sa03_2),
	.B(n21027));
   AOI31xp33_ASAP7_75t_SL FE_RC_630_0 (.Y(n20272),
	.A1(n18971),
	.A2(FE_OCPN27627_sa23_1),
	.A3(n19313),
	.B(n25711));
   AOI31xp33_ASAP7_75t_SL FE_RC_629_0 (.Y(n15782),
	.A1(FE_OFN26058_w3_1),
	.A2(FE_OFN28829_n),
	.A3(n25140),
	.B(n15019));
   AOI31xp33_ASAP7_75t_L FE_RC_628_0 (.Y(n15946),
	.A1(FE_OFN28659_n15934),
	.A2(FE_OFN27115_n),
	.A3(FE_OCPN29534_FE_OFN8_w3_14),
	.B(n14115));
   AOI21xp5_ASAP7_75t_SL FE_RC_627_0 (.Y(n20847),
	.A1(FE_OCPN27516_n26292),
	.A2(n16299),
	.B(n20033));
   AOI21xp5_ASAP7_75t_L FE_RC_626_0 (.Y(n24473),
	.A1(FE_OCPN28021_n21445),
	.A2(FE_OCPN27819_n17245),
	.B(n21444));
   AOI21xp5_ASAP7_75t_L FE_RC_625_0 (.Y(n23551),
	.A1(n16418),
	.A2(FE_OFN28998_n16923),
	.B(n23537));
   AOI21xp5_ASAP7_75t_SL FE_RC_624_0 (.Y(n21644),
	.A1(n18583),
	.A2(FE_OFN28988_n18597),
	.B(n23775));
   AOI21x1_ASAP7_75t_SL FE_RC_623_0 (.Y(n19164),
	.A1(n22505),
	.A2(n17446),
	.B(n21358));
   AOI21xp5_ASAP7_75t_L FE_RC_622_0 (.Y(n22346),
	.A1(FE_OFN28778_FE_OCPN28352_n16748),
	.A2(FE_OFN29023_n16750),
	.B(n17872));
   AOI31xp33_ASAP7_75t_SL FE_RC_621_0 (.Y(n20249),
	.A1(FE_OCPN27986_n18970),
	.A2(FE_OFN29001_n23491),
	.A3(FE_OCPN27916_n),
	.B(n20265));
   AOI31xp33_ASAP7_75t_SL FE_RC_620_0 (.Y(n20449),
	.A1(n21591),
	.A2(n17603),
	.A3(FE_OFN26597_n),
	.B(n19037));
   AOI21xp5_ASAP7_75t_L FE_RC_619_0 (.Y(n19603),
	.A1(n17254),
	.A2(FE_OFN28835_n),
	.B(n17258));
   AOI21xp5_ASAP7_75t_SL FE_RC_618_0 (.Y(n15585),
	.A1(FE_OFN25912_n15848),
	.A2(n13741),
	.B(n13776));
   AOI21xp5_ASAP7_75t_SL FE_RC_617_0 (.Y(n15347),
	.A1(FE_OFN26539_w3_19),
	.A2(FE_OFN26045_n25377),
	.B(FE_OFN26091_n24663));
   AOI21x1_ASAP7_75t_SL FE_RC_616_0 (.Y(n22758),
	.A1(FE_OFN28739_n17898),
	.A2(n25741),
	.B(n20556));
   AOI31xp33_ASAP7_75t_SL FE_RC_615_0 (.Y(n14566),
	.A1(FE_OCPN27659_w3_25),
	.A2(n25675),
	.A3(FE_OFN27206_w3_30),
	.B(FE_OFN27061_n15239));
   AOI21xp5_ASAP7_75t_SL FE_RC_614_0 (.Y(n15386),
	.A1(FE_OFN27115_n),
	.A2(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(n15414));
   AOI21x1_ASAP7_75t_L FE_RC_613_0 (.Y(n15338),
	.A1(FE_OFN28706_n),
	.A2(FE_OFN26539_w3_19),
	.B(FE_OFN5_w3_22));
   AOI21x1_ASAP7_75t_L FE_RC_612_0 (.Y(n15146),
	.A1(FE_OCPN29350_w3_25),
	.A2(n25675),
	.B(FE_OFN27209_w3_30));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5199_n21457 (.Y(FE_OCPN5199_n21457),
	.A(n21457));
   HB1xp67_ASAP7_75t_R FE_OCPC5198_n25566 (.Y(FE_OCPN5198_n25566),
	.A(n25566));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5178_n25039 (.Y(FE_OCPN5178_n25039),
	.A(FE_OCPN8263_n25039));
   BUFx2_ASAP7_75t_SL FE_OCPC5172_n26281 (.Y(FE_OCPN5172_n26281),
	.A(n26281));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5166_n27203 (.Y(FE_OCPN5166_n27203),
	.A(FE_OCPN29445_n27203));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5158_n24742 (.Y(FE_OCPN5158_n24742),
	.A(n24742));
   HB1xp67_ASAP7_75t_R FE_OCPC5156_n23958 (.Y(FE_OCPN5156_n23958),
	.A(n23958));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5147_n18548 (.Y(FE_OCPN5147_n18548),
	.A(n18548));
   HB1xp67_ASAP7_75t_SL FE_OCPC5146_n26207 (.Y(FE_OCPN5146_n26207),
	.A(n26207));
   HB1xp67_ASAP7_75t_L FE_OCPC5140_n21049 (.Y(FE_OCPN5140_n21049),
	.A(n21049));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5139_n24167 (.Y(FE_OCPN5139_n24167),
	.A(n24167));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5133_n26620 (.Y(FE_OCPN5133_n26620),
	.A(n26620));
   HB1xp67_ASAP7_75t_R FE_OCPC5132_n23890 (.Y(FE_OCPN5132_n23890),
	.A(n23890));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5131_n25916 (.Y(FE_OCPN5131_n25916),
	.A(n25916));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5116_n25443 (.Y(FE_OCPN5116_n25443),
	.A(n25443));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5115_n25574 (.Y(FE_OCPN5115_n25574),
	.A(n25574));
   HB1xp67_ASAP7_75t_L FE_OCPC5110_n23721 (.Y(FE_OCPN5110_n23721),
	.A(n23721));
   HB1xp67_ASAP7_75t_R FE_OCPC5109_n26551 (.Y(FE_OCPN5109_n26551),
	.A(n26551));
   HB1xp67_ASAP7_75t_R FE_OCPC5107_n24418 (.Y(FE_OCPN5107_n24418),
	.A(n24418));
   HB1xp67_ASAP7_75t_L FE_OCPC5106_n25999 (.Y(FE_OCPN5106_n25999),
	.A(n25999));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5105_n25099 (.Y(FE_OCPN5105_n25099),
	.A(n25099));
   HB1xp67_ASAP7_75t_L FE_OCPC5099_n24677 (.Y(FE_OCPN5099_n24677),
	.A(n24677));
   HB1xp67_ASAP7_75t_SL FE_OCPC5088_n27079 (.Y(FE_OCPN5088_n27079),
	.A(FE_OCPN27391_n27079));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5086_n26050 (.Y(FE_OCPN5086_n26050),
	.A(n26050));
   HB1xp67_ASAP7_75t_R FE_OCPC5082_n22663 (.Y(FE_OCPN5082_n22663),
	.A(n22663));
   HB1xp67_ASAP7_75t_SL FE_OCPC5080_n25758 (.Y(FE_OCPN5080_n25758),
	.A(n25758));
   BUFx2_ASAP7_75t_L FE_OCPC5079_n20287 (.Y(FE_OCPN5079_n20287),
	.A(n20287));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5077_n25855 (.Y(FE_OCPN5077_n25855),
	.A(n25855));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5076_n24192 (.Y(FE_OCPN5076_n24192),
	.A(n24192));
   HB1xp67_ASAP7_75t_R FE_OCPC5073_n24996 (.Y(FE_OCPN5073_n24996),
	.A(n24996));
   HB1xp67_ASAP7_75t_SL FE_OCPC5068_n25984 (.Y(FE_OCPN5068_n25984),
	.A(n25984));
   BUFx3_ASAP7_75t_SL FE_OCPC5019_n26728 (.Y(FE_OCPN27787_n26728),
	.A(n26728));
   INVxp67_ASAP7_75t_L FE_OCPC5018_sa23_1 (.Y(FE_OCPN27956_n),
	.A(FE_OCPN27627_sa23_1));
   BUFx6f_ASAP7_75t_SL FE_OCPC5017_sa23_1 (.Y(FE_OCPN27627_sa23_1),
	.A(sa23_1_));
   HB1xp67_ASAP7_75t_R FE_OCPC5062_n20505 (.Y(FE_OCPN5062_n20505),
	.A(n20505));
   HB1xp67_ASAP7_75t_R FE_OCPC5056_n26535 (.Y(FE_OCPN5056_n26535),
	.A(n26535));
   HB1xp67_ASAP7_75t_L FE_OCPC5053_n25832 (.Y(FE_OCPN5053_n25832),
	.A(n25832));
   HB1xp67_ASAP7_75t_R FE_OCPC5051_n25883 (.Y(FE_OCPN5051_n25883),
	.A(n25883));
   HB1xp67_ASAP7_75t_SL FE_OCPC5043_n26230 (.Y(FE_OCPN5043_n26230),
	.A(n26230));
   HB1xp67_ASAP7_75t_R FE_OCPC5041_n26726 (.Y(FE_OCPN5041_n26726),
	.A(n26726));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5038_n26735 (.Y(FE_OCPN5038_n26735),
	.A(n26735));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC5020_n27079 (.Y(FE_OCPN5020_n27079),
	.A(n27079));
   OAI21x1_ASAP7_75t_SL FE_RC_611_0 (.Y(n15915),
	.A1(n25648),
	.A2(n15902),
	.B(n15901));
   OR3x1_ASAP7_75t_SL FE_RC_609_0 (.Y(FE_RN_229_0),
	.A(n22775),
	.B(n22774),
	.C(n23573));
   INVx3_ASAP7_75t_L FE_RC_605_0 (.Y(n25741),
	.A(FE_RN_228_0));
   OR3x1_ASAP7_75t_SL FE_RC_604_0 (.Y(FE_RN_228_0),
	.A(FE_OFN25908_sa12_2),
	.B(FE_OCPN29499_FE_OFN16131_sa12_1),
	.C(FE_OFN29225_sa12_0));
   AOI31xp33_ASAP7_75t_L FE_RC_603_0 (.Y(n23549),
	.A1(n17416),
	.A2(FE_OFN28771_n),
	.A3(FE_OCPN29487_FE_OFN28694_sa33_4),
	.B(n16871));
   INVxp33_ASAP7_75t_R FE_RC_601_0 (.Y(FE_RN_226_0),
	.A(FE_OFN21_n16125));
   NAND2xp33_ASAP7_75t_SRAM FE_RC_600_0 (.Y(FE_RN_227_0),
	.A(n21957),
	.B(FE_RN_226_0));
   OAI21x1_ASAP7_75t_SL FE_RC_599_0 (.Y(n16081),
	.A1(FE_OFN21_n16125),
	.A2(n16082),
	.B(FE_RN_227_0));
   OR3x1_ASAP7_75t_L FE_RC_598_0 (.Y(FE_RN_224_0),
	.A(n22045),
	.B(FE_OFN29151_n22988),
	.C(n22989));
   NOR3xp33_ASAP7_75t_SL FE_RC_597_0 (.Y(n22994),
	.A(FE_RN_224_0),
	.B(n19340),
	.C(n19339));
   AOI31xp33_ASAP7_75t_SL FE_RC_596_0 (.Y(n21808),
	.A1(n21806),
	.A2(n21807),
	.A3(n21805),
	.B(n26889));
   NOR3xp33_ASAP7_75t_SL FE_RC_594_0 (.Y(n20694),
	.A(n23885),
	.B(n26900),
	.C(n20692));
   NAND3xp33_ASAP7_75t_SL FE_RC_593_0 (.Y(n16855),
	.A(n16417),
	.B(n17416),
	.C(FE_OFN28771_n));
   OAI21xp5_ASAP7_75t_SL FE_RC_592_0 (.Y(n646),
	.A1(FE_OCPN29428_FE_OFN27131_w3_29),
	.A2(FE_OFN16253_n16189),
	.B(n16188));
   BUFx4f_ASAP7_75t_SL FE_OCPC5012_n23392 (.Y(FE_OCPN28447_n23392),
	.A(n23392));
   AND2x2_ASAP7_75t_SRAM FE_RC_591_0 (.Y(FE_RN_223_0),
	.A(n26621),
	.B(n26620));
   NAND2xp5_ASAP7_75t_SL FE_RC_590_0 (.Y(n26618),
	.A(FE_RN_223_0),
	.B(n26619));
   AOI31xp33_ASAP7_75t_SL FE_RC_588_0 (.Y(n16824),
	.A1(n17830),
	.A2(n16823),
	.A3(n16822),
	.B(n25585));
   NOR3xp33_ASAP7_75t_L FE_RC_586_0 (.Y(n24597),
	.A(n24598),
	.B(FE_OCPN27723_n),
	.C(n25484));
   BUFx2_ASAP7_75t_SL FE_OCPC5009_n428 (.Y(FE_OCPN28444_n428),
	.A(n428));
   BUFx3_ASAP7_75t_SL FE_OCPC5007_n27056 (.Y(FE_OCPN28442_n27056),
	.A(n27056));
   OAI21x1_ASAP7_75t_SL FE_RC_583_0 (.Y(n27110),
	.A1(n25568),
	.A2(FE_RN_137_0),
	.B(n25567));
   NOR3xp33_ASAP7_75t_SL FE_RC_579_0 (.Y(n15749),
	.A(n15283),
	.B(n13870),
	.C(FE_OFN28_w3_23));
   NOR3xp33_ASAP7_75t_SL FE_RC_578_0 (.Y(n17918),
	.A(n22734),
	.B(n23590),
	.C(n22730));
   AOI31xp33_ASAP7_75t_SL FE_RC_577_0 (.Y(n23846),
	.A1(n25628),
	.A2(n23845),
	.A3(n25630),
	.B(n26517));
   OAI21xp5_ASAP7_75t_SL FE_RC_576_0 (.Y(n25784),
	.A1(n25780),
	.A2(FE_RN_219_0),
	.B(n25779));
   HB1xp67_ASAP7_75t_R FE_OCPC5003_n27080 (.Y(FE_OCPN28438_n27080),
	.A(n27080));
   AOI31xp33_ASAP7_75t_SL FE_RC_575_0 (.Y(n23465),
	.A1(n23453),
	.A2(n23454),
	.A3(n23452),
	.B(n23945));
   OAI21x1_ASAP7_75t_SL FE_RC_573_0 (.Y(n26944),
	.A1(FE_RN_121_0),
	.A2(n25538),
	.B(n25537));
   NAND3x1_ASAP7_75t_L FE_RC_572_0 (.Y(n25277),
	.A(n17778),
	.B(n22890),
	.C(n22554));
   NOR3xp33_ASAP7_75t_L FE_RC_571_0 (.Y(n16378),
	.A(n27070),
	.B(n20078),
	.C(n16496));
   AOI31xp33_ASAP7_75t_SL FE_RC_570_0 (.Y(n25291),
	.A1(n19437),
	.A2(n19438),
	.A3(n19436),
	.B(n26959));
   OR3x1_ASAP7_75t_SL FE_RC_567_0 (.Y(FE_RN_222_0),
	.A(FE_OFN28712_n),
	.B(FE_OFN28_w3_23),
	.C(FE_OFN28683_w3_21));
   BUFx4f_ASAP7_75t_SL FE_OCPC4999_n17546 (.Y(FE_OCPN28434_n17546),
	.A(n17546));
   HB1xp67_ASAP7_75t_L FE_OCPC4996_n21734 (.Y(FE_OCPN28431_n21734),
	.A(n21734));
   HB1xp67_ASAP7_75t_L FE_OCPC4992_n25064 (.Y(FE_OCPN28427_n25064),
	.A(n25064));
   BUFx2_ASAP7_75t_L FE_OCPC4988_n18836 (.Y(FE_OCPN28423_n18836),
	.A(n18836));
   AND2x2_ASAP7_75t_L FE_RC_564_0 (.Y(FE_RN_220_0),
	.A(n26407),
	.B(n25510));
   OAI21xp5_ASAP7_75t_SL FE_RC_563_0 (.Y(n26654),
	.A1(FE_RN_220_0),
	.A2(n25195),
	.B(n25194));
   HB1xp67_ASAP7_75t_R FE_OCPC4983_n19586 (.Y(FE_OCPN28418_n19586),
	.A(n19586));
   AND2x2_ASAP7_75t_SL FE_RC_562_0 (.Y(FE_RN_219_0),
	.A(FE_OCPN27787_n26728),
	.B(FE_OFN28489_ld_r));
   HB1xp67_ASAP7_75t_R FE_OCPC4698_n25497 (.Y(FE_OCPN4698_n25497),
	.A(n25497));
   HB1xp67_ASAP7_75t_L FE_OCPC4685_n15658 (.Y(FE_OCPN4685_n15658),
	.A(n15658));
   HB1xp67_ASAP7_75t_R FE_OCPC4680_n21317 (.Y(FE_OCPN4680_n21317),
	.A(n21317));
   BUFx2_ASAP7_75t_L FE_OCPC4951_n17899 (.Y(FE_OCPN28386_n17899),
	.A(n17899));
   HB1xp67_ASAP7_75t_R FE_OCPC4948_n24808 (.Y(FE_OCPN28383_n24808),
	.A(n26683));
   BUFx2_ASAP7_75t_L FE_OCPC4946_n26660 (.Y(FE_OCPN28381_n26660),
	.A(n26660));
   BUFx2_ASAP7_75t_SL FE_OCPC4945_n22433 (.Y(FE_OCPN28380_n22433),
	.A(n22433));
   BUFx2_ASAP7_75t_L FE_OCPC4943_n22632 (.Y(FE_OCPN28378_n22632),
	.A(n22632));
   AND2x2_ASAP7_75t_SRAM FE_RC_560_0 (.Y(FE_RN_218_0),
	.A(FE_OCPN29586_n26857),
	.B(n25044));
   OAI21x1_ASAP7_75t_SL FE_RC_559_0 (.Y(n25423),
	.A1(FE_RN_218_0),
	.A2(n23935),
	.B(n23934));
   HB1xp67_ASAP7_75t_SL FE_OCPC4931_n25329 (.Y(FE_OCPN28366_n25329),
	.A(n25329));
   BUFx3_ASAP7_75t_L FE_OCPC4928_n22979 (.Y(FE_OCPN28363_n22979),
	.A(n22979));
   HB1xp67_ASAP7_75t_L FE_OCPC4922_n22882 (.Y(FE_OCPN28357_n22882),
	.A(n22882));
   BUFx3_ASAP7_75t_SL FE_OCPC4920_n26909 (.Y(FE_OCPN28355_n26909),
	.A(n26910));
   HB1xp67_ASAP7_75t_L FE_OCPC4919_n16677 (.Y(FE_OCPN28354_n16677),
	.A(n16677));
   BUFx3_ASAP7_75t_SL FE_OCPC4918_n18534 (.Y(FE_OCPN28353_n18534),
	.A(n18534));
   OA21x2_ASAP7_75t_SRAM FE_RC_558_0 (.Y(FE_RN_217_0),
	.A1(w2_4_),
	.A2(text_in_r_36_),
	.B(n26209));
   NOR2x1p5_ASAP7_75t_SL FE_RC_557_0 (.Y(n500),
	.A(FE_RN_217_0),
	.B(n26208));
   HB1xp67_ASAP7_75t_SL FE_OCPC4911_n24051 (.Y(FE_OCPN28346_n24051),
	.A(n24051));
   HB1xp67_ASAP7_75t_R FE_OCPC4893_n25953 (.Y(FE_OCPN28328_n25953),
	.A(n25953));
   AO21x1_ASAP7_75t_SL FE_RC_556_0 (.Y(FE_RN_216_0),
	.A1(n27117),
	.A2(n26531),
	.B(FE_OCPN29389_n26528));
   NAND2xp5_ASAP7_75t_SL FE_RC_555_0 (.Y(n24304),
	.A(FE_RN_216_0),
	.B(n25252));
   BUFx2_ASAP7_75t_L FE_OCPC4887_n18141 (.Y(FE_OCPN28322_n18141),
	.A(n18141));
   BUFx4_ASAP7_75t_SL FE_OCPC4886_n21341 (.Y(FE_OCPN28321_n21341),
	.A(n21341));
   HB1xp67_ASAP7_75t_R FE_OCPC4885_n25954 (.Y(FE_OCPN28320_n25954),
	.A(n25954));
   HB1xp67_ASAP7_75t_R FE_OCPC4881_n26980 (.Y(FE_OCPN28316_n26980),
	.A(n26980));
   INVx3_ASAP7_75t_SL FE_OCPC4879_n20842 (.Y(FE_OCPN28314_n20842),
	.A(FE_OCPN28312_n20842));
   INVx1_ASAP7_75t_SL FE_OCPC4877_n20842 (.Y(FE_OCPN28312_n20842),
	.A(n20842));
   BUFx3_ASAP7_75t_SL FE_OCPC4872_n26491 (.Y(FE_OCPN28307_n26491),
	.A(n26491));
   HB1xp67_ASAP7_75t_SL FE_OCPC4870_n26451 (.Y(FE_OCPN28305_n26451),
	.A(n26451));
   BUFx2_ASAP7_75t_SL FE_OCPC4868_n20961 (.Y(FE_OCPN28303_n20961),
	.A(n20961));
   NAND2xp5_ASAP7_75t_L FE_RC_554_0 (.Y(n26180),
	.A(FE_RN_210_0),
	.B(n20486));
   NAND2xp5_ASAP7_75t_SL FE_RC_552_0 (.Y(FE_RN_205_0),
	.A(FE_RN_210_0),
	.B(FE_RN_206_0));
   NAND2x1_ASAP7_75t_SL FE_RC_550_0 (.Y(FE_RN_206_0),
	.A(n26183),
	.B(FE_OFN16163_n26584));
   INVxp67_ASAP7_75t_L FE_RC_549_0 (.Y(FE_RN_207_0),
	.A(FE_RN_206_0));
   INVxp33_ASAP7_75t_R FE_RC_548_0 (.Y(FE_RN_208_0),
	.A(n20487));
   INVxp33_ASAP7_75t_R FE_RC_547_0 (.Y(FE_RN_209_0),
	.A(n26926));
   NAND2xp5_ASAP7_75t_L FE_RC_546_0 (.Y(FE_RN_210_0),
	.A(FE_RN_208_0),
	.B(FE_RN_209_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_545_0 (.Y(FE_RN_211_0),
	.A(FE_RN_210_0),
	.B(n20486));
   NOR2x1_ASAP7_75t_SL FE_RC_544_0 (.Y(FE_RN_212_0),
	.A(FE_RN_207_0),
	.B(FE_RN_211_0));
   INVxp33_ASAP7_75t_R FE_RC_542_0 (.Y(FE_RN_214_0),
	.A(FE_OFN16169_n26567));
   NOR2xp33_ASAP7_75t_R FE_RC_541_0 (.Y(FE_RN_215_0),
	.A(FE_RN_213_0),
	.B(FE_RN_214_0));
   OAI21xp5_ASAP7_75t_SL FE_RC_540_0 (.Y(n25449),
	.A1(FE_OFN28512_n27020),
	.A2(FE_RN_215_0),
	.B(FE_RN_212_0));
   INVxp33_ASAP7_75t_L FE_RC_539_0 (.Y(FE_RN_195_0),
	.A(n20203));
   NOR2xp33_ASAP7_75t_L FE_RC_538_0 (.Y(n20992),
	.A(FE_RN_195_0),
	.B(FE_RN_202_0));
   INVxp67_ASAP7_75t_L FE_RC_537_0 (.Y(FE_RN_196_0),
	.A(n20990));
   INVxp67_ASAP7_75t_SL FE_RC_536_0 (.Y(FE_RN_197_0),
	.A(n20206));
   NAND2xp5_ASAP7_75t_R FE_RC_535_0 (.Y(FE_RN_198_0),
	.A(n20204),
	.B(FE_RN_197_0));
   NOR2xp33_ASAP7_75t_SL FE_RC_533_0 (.Y(FE_RN_200_0),
	.A(FE_RN_198_0),
	.B(FE_OFN28924_n25912));
   NAND2xp5_ASAP7_75t_SL FE_RC_531_0 (.Y(FE_RN_202_0),
	.A(FE_RN_200_0),
	.B(FE_RN_201_0));
   NOR2xp67_ASAP7_75t_SL FE_RC_530_0 (.Y(FE_RN_203_0),
	.A(FE_RN_196_0),
	.B(FE_RN_202_0));
   AOI31xp33_ASAP7_75t_SL FE_RC_529_0 (.Y(n21006),
	.A1(FE_RN_203_0),
	.A2(n20991),
	.A3(n20203),
	.B(n27140));
   INVxp67_ASAP7_75t_R FE_RC_526_0 (.Y(FE_RN_193_0),
	.A(n18439));
   NOR4xp25_ASAP7_75t_L FE_RC_525_0 (.Y(FE_RN_194_0),
	.A(FE_RN_193_0),
	.B(FE_RN_192_0),
	.C(FE_RN_191_0),
	.D(FE_OCPN29577_n24298));
   OAI21xp5_ASAP7_75t_SL FE_RC_524_0 (.Y(n26766),
	.A1(FE_RN_194_0),
	.A2(n24331),
	.B(n18448));
   INVxp33_ASAP7_75t_L FE_RC_522_0 (.Y(FE_RN_188_0),
	.A(n19137));
   NAND4xp25_ASAP7_75t_SL FE_RC_520_0 (.Y(FE_RN_190_0),
	.A(n19133),
	.B(n19131),
	.C(n19132),
	.D(n18653));
   OR3x1_ASAP7_75t_SL FE_RC_519_0 (.Y(n21180),
	.A(FE_RN_190_0),
	.B(FE_RN_188_0),
	.C(FE_RN_187_0));
   INVxp33_ASAP7_75t_R FE_RC_518_0 (.Y(FE_RN_179_0),
	.A(n26857));
   INVxp67_ASAP7_75t_SL FE_RC_517_0 (.Y(FE_RN_180_0),
	.A(n23050));
   INVxp33_ASAP7_75t_R FE_RC_516_0 (.Y(FE_RN_181_0),
	.A(n23051));
   AOI21xp5_ASAP7_75t_SL FE_RC_515_0 (.Y(FE_RN_182_0),
	.A1(FE_RN_181_0),
	.A2(FE_RN_180_0),
	.B(FE_RN_179_0));
   INVxp33_ASAP7_75t_R FE_RC_514_0 (.Y(FE_RN_183_0),
	.A(n25139));
   INVxp33_ASAP7_75t_L FE_RC_513_0 (.Y(FE_RN_184_0),
	.A(n23046));
   AOI21xp33_ASAP7_75t_L FE_RC_512_0 (.Y(FE_RN_185_0),
	.A1(n23041),
	.A2(n23042),
	.B(FE_RN_184_0));
   NAND2xp5_ASAP7_75t_R FE_RC_511_0 (.Y(FE_RN_186_0),
	.A(n23048),
	.B(FE_RN_185_0));
   AOI21x1_ASAP7_75t_SL FE_RC_510_0 (.Y(n26335),
	.A1(FE_RN_186_0),
	.A2(FE_RN_183_0),
	.B(FE_RN_182_0));
   NAND2x1_ASAP7_75t_SL FE_RC_509_0 (.Y(FE_OCPN27772_n24234),
	.A(FE_RN_175_0),
	.B(n20948));
   INVxp67_ASAP7_75t_SL FE_RC_508_0 (.Y(FE_RN_170_0),
	.A(n20948));
   NOR2xp33_ASAP7_75t_L FE_RC_506_0 (.Y(n24602),
	.A(FE_RN_170_0),
	.B(FE_RN_171_0));
   INVxp33_ASAP7_75t_R FE_RC_504_0 (.Y(FE_RN_173_0),
	.A(n27027));
   NAND2xp33_ASAP7_75t_L FE_RC_503_0 (.Y(FE_RN_174_0),
	.A(n20949),
	.B(n22957));
   NAND2xp5_ASAP7_75t_R FE_RC_502_0 (.Y(FE_RN_175_0),
	.A(FE_RN_173_0),
	.B(FE_RN_174_0));
   AOI21xp33_ASAP7_75t_R FE_RC_500_0 (.Y(FE_RN_177_0),
	.A1(n24038),
	.A2(n24037),
	.B(FE_RN_171_0));
   NAND2xp33_ASAP7_75t_SL FE_RC_499_0 (.Y(FE_RN_178_0),
	.A(n24033),
	.B(FE_RN_177_0));
   OAI21xp5_ASAP7_75t_SL FE_RC_498_0 (.Y(n25488),
	.A1(FE_RN_178_0),
	.A2(FE_RN_170_0),
	.B(n24035));
   NOR2x1p5_ASAP7_75t_SL FE_RC_497_0 (.Y(n18526),
	.A(n18551),
	.B(FE_OFN28536_sa20_2));
   NOR2xp33_ASAP7_75t_SL FE_RC_496_0 (.Y(FE_RN_164_0),
	.A(FE_OFN28536_sa20_2),
	.B(n18551));
   NAND3xp33_ASAP7_75t_L FE_RC_495_0 (.Y(FE_OCPN27591_n23742),
	.A(FE_RN_164_0),
	.B(n21195),
	.C(FE_OFN29150_sa20_5));
   INVxp67_ASAP7_75t_R FE_RC_493_0 (.Y(FE_RN_166_0),
	.A(n18551));
   NAND4xp25_ASAP7_75t_SRAM FE_RC_492_0 (.Y(FE_OCPN28246_n),
	.A(FE_RN_166_0),
	.B(n18533),
	.C(n21195),
	.D(FE_OFN29150_sa20_5));
   NAND4xp25_ASAP7_75t_L FE_RC_489_0 (.Y(FE_RN_169_0),
	.A(FE_OFN29150_sa20_5),
	.B(n21195),
	.C(n18533),
	.D(FE_RN_166_0));
   NAND2x1_ASAP7_75t_SL FE_RC_488_0 (.Y(n23879),
	.A(n23710),
	.B(FE_RN_169_0));
   NOR2xp33_ASAP7_75t_L FE_RC_486_0 (.Y(FE_RN_159_0),
	.A(n22407),
	.B(n22406));
   INVxp33_ASAP7_75t_L FE_RC_485_0 (.Y(FE_RN_160_0),
	.A(n22405));
   NOR2xp33_ASAP7_75t_R FE_RC_484_0 (.Y(FE_RN_161_0),
	.A(FE_RN_159_0),
	.B(FE_RN_160_0));
   AOI31xp33_ASAP7_75t_SL FE_RC_483_0 (.Y(FE_RN_162_0),
	.A1(n22403),
	.A2(n22402),
	.A3(n22401),
	.B(n23899));
   AOI21xp5_ASAP7_75t_L FE_RC_482_0 (.Y(FE_RN_163_0),
	.A1(n22409),
	.A2(n22410),
	.B(n26346));
   OR3x2_ASAP7_75t_SL FE_RC_481_0 (.Y(n25667),
	.A(FE_RN_163_0),
	.B(FE_RN_162_0),
	.C(FE_RN_161_0));
   AO21x1_ASAP7_75t_L FE_RC_480_0 (.Y(FE_RN_154_0),
	.A1(n21143),
	.A2(n23165),
	.B(n26889));
   OAI21xp5_ASAP7_75t_SL FE_RC_479_0 (.Y(FE_RN_155_0),
	.A1(n21140),
	.A2(n21141),
	.B(n26878));
   NAND2xp33_ASAP7_75t_L FE_RC_478_0 (.Y(FE_RN_156_0),
	.A(n22868),
	.B(n21137));
   INVxp67_ASAP7_75t_L FE_RC_477_0 (.Y(FE_RN_157_0),
	.A(n21138));
   NOR2xp33_ASAP7_75t_SL FE_RC_476_0 (.Y(FE_RN_158_0),
	.A(FE_RN_156_0),
	.B(FE_RN_157_0));
   OAI21xp33_ASAP7_75t_SRAM FE_RC_474_0 (.Y(FE_RN_149_0),
	.A1(text_in_r_65_),
	.A2(w1_1_),
	.B(n27036));
   NOR2xp33_ASAP7_75t_R FE_RC_473_0 (.Y(FE_RN_150_0),
	.A(FE_OCPN27519_n25407),
	.B(FE_OFN12_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL FE_RC_471_0 (.Y(FE_RN_152_0),
	.A(FE_RN_150_0),
	.B(FE_RN_151_0));
   NOR2xp33_ASAP7_75t_SL FE_RC_470_0 (.Y(FE_RN_153_0),
	.A(n27033),
	.B(n27031));
   OA21x2_ASAP7_75t_SL FE_RC_469_0 (.Y(n469),
	.A1(FE_RN_153_0),
	.A2(FE_RN_152_0),
	.B(FE_RN_149_0));
   NAND2xp5_ASAP7_75t_L FE_RC_466_0 (.Y(FE_RN_147_0),
	.A(n16379),
	.B(n16380));
   NAND2xp5_ASAP7_75t_SL FE_RC_465_0 (.Y(FE_RN_148_0),
	.A(n16382),
	.B(FE_RN_147_0));
   AOI31xp33_ASAP7_75t_SL FE_RC_464_0 (.Y(n24192),
	.A1(FE_RN_148_0),
	.A2(n26296),
	.A3(n26045),
	.B(n27075));
   AND4x1_ASAP7_75t_L FE_RC_463_0 (.Y(FE_RN_146_0),
	.A(n22621),
	.B(n21609),
	.C(n21613),
	.D(n21611));
   AOI31xp33_ASAP7_75t_SL FE_RC_462_0 (.Y(n25116),
	.A1(FE_RN_146_0),
	.A2(n24030),
	.A3(n21615),
	.B(n24800));
   AND2x2_ASAP7_75t_L FE_RC_461_0 (.Y(FE_RN_145_0),
	.A(FE_OFN16176_n27207),
	.B(n26196));
   OAI21x1_ASAP7_75t_SL FE_RC_460_0 (.Y(n26649),
	.A1(FE_RN_145_0),
	.A2(n26195),
	.B(n26194));
   AOI31xp33_ASAP7_75t_SL FE_RC_459_0 (.Y(FE_RN_142_0),
	.A1(FE_OFN27148_sa32_3),
	.A2(FE_OCPN29459_n),
	.A3(n17529),
	.B(n24869));
   INVxp67_ASAP7_75t_L FE_RC_458_0 (.Y(FE_RN_143_0),
	.A(n24868));
   NAND4xp25_ASAP7_75t_SL FE_RC_457_0 (.Y(FE_RN_144_0),
	.A(FE_RN_143_0),
	.B(n24866),
	.C(n24867),
	.D(FE_RN_142_0));
   NOR2x1_ASAP7_75t_SL FE_RC_456_0 (.Y(n17678),
	.A(FE_RN_144_0),
	.B(n24864));
   BUFx2_ASAP7_75t_SL FE_OCPC4854_n20235 (.Y(FE_OCPN28289_n20235),
	.A(n20235));
   HB1xp67_ASAP7_75t_SL FE_OCPC4844_n26675 (.Y(FE_OCPN28279_n),
	.A(n26675));
   AND2x2_ASAP7_75t_R FE_RC_455_0 (.Y(FE_RN_141_0),
	.A(n26249),
	.B(n26248));
   OAI21x1_ASAP7_75t_SL FE_RC_454_0 (.Y(n26713),
	.A1(FE_RN_141_0),
	.A2(n25766),
	.B(n25765));
   OR2x2_ASAP7_75t_R FE_RC_453_0 (.Y(FE_RN_140_0),
	.A(n20551),
	.B(FE_OFN28520_n22753));
   NOR2x1_ASAP7_75t_L FE_RC_452_0 (.Y(n24046),
	.A(FE_RN_140_0),
	.B(n20810));
   AND2x2_ASAP7_75t_L FE_RC_451_0 (.Y(FE_RN_139_0),
	.A(n26770),
	.B(n26769));
   OAI21xp5_ASAP7_75t_SL FE_RC_450_0 (.Y(n26779),
	.A1(FE_RN_139_0),
	.A2(n26768),
	.B(n26767));
   XOR2xp5_ASAP7_75t_SL FE_RC_449_0 (.Y(FE_RN_138_0),
	.A(n26838),
	.B(FE_OCPN27497_n25431));
   XNOR2xp5_ASAP7_75t_SL FE_RC_448_0 (.Y(n25436),
	.A(FE_RN_138_0),
	.B(n25430));
   AND2x2_ASAP7_75t_L FE_RC_447_0 (.Y(FE_RN_137_0),
	.A(n27183),
	.B(n27182));
   AND2x2_ASAP7_75t_SRAM FE_RC_445_0 (.Y(FE_RN_136_0),
	.A(n26282),
	.B(FE_OCPN5172_n26281));
   OAI21xp5_ASAP7_75t_SL FE_RC_444_0 (.Y(n26176),
	.A1(FE_RN_136_0),
	.A2(n26174),
	.B(n26173));
   AND2x2_ASAP7_75t_SRAM FE_RC_443_0 (.Y(FE_RN_135_0),
	.A(n26819),
	.B(FE_OCPN8227_n25950));
   OAI21x1_ASAP7_75t_SL FE_RC_442_0 (.Y(n25952),
	.A1(FE_RN_135_0),
	.A2(n25949),
	.B(n25948));
   OA21x2_ASAP7_75t_SRAM FE_RC_441_0 (.Y(FE_RN_134_0),
	.A1(w2_17_),
	.A2(text_in_r_49_),
	.B(n27149));
   NOR2x1_ASAP7_75t_SL FE_RC_440_0 (.Y(n434),
	.A(FE_RN_134_0),
	.B(n27148));
   XNOR2xp5_ASAP7_75t_SL FE_RC_439_0 (.Y(FE_RN_133_0),
	.A(n26260),
	.B(n26259));
   XOR2xp5_ASAP7_75t_SL FE_RC_438_0 (.Y(n26263),
	.A(FE_RN_133_0),
	.B(n26261));
   AND2x2_ASAP7_75t_L FE_RC_437_0 (.Y(FE_RN_132_0),
	.A(FE_OFN16148_n25466),
	.B(FE_OFN29051_n25465));
   OAI21x1_ASAP7_75t_SL FE_RC_436_0 (.Y(n26349),
	.A1(FE_RN_132_0),
	.A2(n24906),
	.B(n24905));
   OR2x2_ASAP7_75t_SL FE_RC_435_0 (.Y(FE_RN_131_0),
	.A(n18023),
	.B(n18024));
   NOR2x1p5_ASAP7_75t_SL FE_RC_434_0 (.Y(n21531),
	.A(FE_RN_131_0),
	.B(n23460));
   AND2x2_ASAP7_75t_L FE_RC_433_0 (.Y(FE_RN_130_0),
	.A(n14817),
	.B(n14816));
   OAI21xp5_ASAP7_75t_SL FE_RC_432_0 (.Y(n14819),
	.A1(FE_RN_130_0),
	.A2(n13901),
	.B(n14815));
   OR2x2_ASAP7_75t_L FE_RC_431_0 (.Y(FE_RN_129_0),
	.A(n17463),
	.B(n24556));
   AND2x2_ASAP7_75t_SL FE_RC_429_0 (.Y(FE_RN_128_0),
	.A(n26322),
	.B(n26323));
   NOR2x1p5_ASAP7_75t_SL FE_RC_428_0 (.Y(n26495),
	.A(FE_RN_128_0),
	.B(n26319));
   XOR2x2_ASAP7_75t_SL FE_RC_427_0 (.Y(FE_RN_127_0),
	.A(n26519),
	.B(n26518));
   XNOR2xp5_ASAP7_75t_SL FE_RC_426_0 (.Y(n26522),
	.A(FE_RN_127_0),
	.B(n26520));
   OR2x2_ASAP7_75t_SRAM FE_RC_425_0 (.Y(FE_RN_126_0),
	.A(n26926),
	.B(n26995));
   OR2x2_ASAP7_75t_SL FE_RC_423_0 (.Y(FE_RN_125_0),
	.A(n24457),
	.B(n24456));
   AOI21x1_ASAP7_75t_SL FE_RC_422_0 (.Y(FE_OCPN27306_n334),
	.A1(FE_RN_125_0),
	.A2(FE_OFN16432_w3_16),
	.B(n24455));
   AO21x1_ASAP7_75t_SL FE_RC_421_0 (.Y(FE_RN_124_0),
	.A1(n26934),
	.A2(n26933),
	.B(n26932));
   NAND2xp5_ASAP7_75t_SL FE_RC_420_0 (.Y(n430),
	.A(FE_RN_124_0),
	.B(n26931));
   BUFx2_ASAP7_75t_L FE_OCPC4833_n19911 (.Y(FE_OCPN28268_n19911),
	.A(n19911));
   BUFx3_ASAP7_75t_SL FE_OCPC4831_n20920 (.Y(FE_OCPN28266_n20920),
	.A(n20920));
   AND2x2_ASAP7_75t_L FE_RC_419_0 (.Y(FE_RN_123_0),
	.A(n18043),
	.B(n21750));
   AOI21xp5_ASAP7_75t_SL FE_RC_418_0 (.Y(n23941),
	.A1(n18044),
	.A2(FE_RN_123_0),
	.B(n23467));
   AND2x2_ASAP7_75t_SRAM FE_RC_417_0 (.Y(FE_RN_122_0),
	.A(n27183),
	.B(n27182));
   OAI21xp5_ASAP7_75t_SL FE_RC_416_0 (.Y(n27185),
	.A1(FE_RN_122_0),
	.A2(n27181),
	.B(n27180));
   HB1xp67_ASAP7_75t_L FE_OCPC4822_n23689 (.Y(FE_OCPN28257_n23689),
	.A(n23689));
   AND2x2_ASAP7_75t_L FE_RC_415_0 (.Y(FE_RN_121_0),
	.A(n26915),
	.B(n26914));
   BUFx2_ASAP7_75t_L FE_OCPC4815_n19573 (.Y(FE_OCPN28250_n19573),
	.A(n19573));
   HB1xp67_ASAP7_75t_L FE_OCPC4813_n17971 (.Y(FE_OCPN28248_n17971),
	.A(n17971));
   BUFx2_ASAP7_75t_SL FE_OCPC4806_n22142 (.Y(FE_OCPN28241_n22142),
	.A(n22142));
   NOR2xp33_ASAP7_75t_SL FE_RC_413_0 (.Y(FE_RN_120_0),
	.A(FE_OFN1_ld_r),
	.B(n26654));
   INVxp67_ASAP7_75t_SL FE_RC_412_0 (.Y(FE_RN_119_0),
	.A(FE_RN_120_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_411_0 (.Y(n26652),
	.A(FE_RN_119_0),
	.B(n26653));
   BUFx2_ASAP7_75t_L FE_OCPC4797_n17949 (.Y(FE_OCPN28232_n17949),
	.A(n17949));
   AND2x2_ASAP7_75t_L FE_RC_410_0 (.Y(FE_RN_118_0),
	.A(n27117),
	.B(n26531));
   BUFx2_ASAP7_75t_SL FE_OCPC4794_n17529 (.Y(FE_OCPN28229_n17529),
	.A(n17529));
   AND2x2_ASAP7_75t_SRAM FE_RC_408_0 (.Y(FE_RN_117_0),
	.A(FE_OCPN29587_n26857),
	.B(FE_OFN29242_n26856));
   OAI21xp5_ASAP7_75t_L FE_RC_407_0 (.Y(n26859),
	.A1(FE_RN_117_0),
	.A2(n26855),
	.B(n26854));
   BUFx2_ASAP7_75t_L FE_OCPC4779_n21500 (.Y(FE_OCPN28214_n21500),
	.A(n21500));
   BUFx3_ASAP7_75t_SL FE_OCPC4769_n20526 (.Y(FE_OCPN28204_n20526),
	.A(n20526));
   BUFx6f_ASAP7_75t_SL FE_OCPC4767_n16991 (.Y(FE_OCPN28202_n16991),
	.A(n16991));
   AND2x2_ASAP7_75t_SRAM FE_RC_406_0 (.Y(FE_RN_116_0),
	.A(n18940),
	.B(n18272));
   NAND2x1p5_ASAP7_75t_L FE_RC_405_0 (.Y(n25282),
	.A(FE_RN_116_0),
	.B(n18271));
   AND2x2_ASAP7_75t_SRAM FE_RC_404_0 (.Y(FE_RN_115_0),
	.A(n27117),
	.B(n26531));
   OAI21xp5_ASAP7_75t_SL FE_RC_403_0 (.Y(n26533),
	.A1(FE_RN_115_0),
	.A2(n26530),
	.B(n26529));
   OR2x2_ASAP7_75t_SRAM FE_RC_402_0 (.Y(FE_RN_114_0),
	.A(w2_1_),
	.B(text_in_r_33_));
   AND2x2_ASAP7_75t_SRAM FE_RC_400_0 (.Y(FE_RN_113_0),
	.A(FE_OFN28565_n26845),
	.B(FE_OFN28489_ld_r));
   OAI21x1_ASAP7_75t_SL FE_RC_399_0 (.Y(n26849),
	.A1(FE_RN_113_0),
	.A2(n26844),
	.B(n26843));
   AND2x2_ASAP7_75t_SRAM FE_RC_398_0 (.Y(FE_RN_112_0),
	.A(n26139),
	.B(n26138));
   OAI21x1_ASAP7_75t_SL FE_RC_397_0 (.Y(n26472),
	.A1(FE_RN_112_0),
	.A2(n24427),
	.B(n24426));
   AND2x2_ASAP7_75t_R FE_RC_396_0 (.Y(FE_RN_111_0),
	.A(n27183),
	.B(n24178));
   OAI21xp5_ASAP7_75t_SL FE_RC_395_0 (.Y(n26420),
	.A1(FE_RN_111_0),
	.A2(n24177),
	.B(n24176));
   AND2x2_ASAP7_75t_L FE_RC_394_0 (.Y(FE_RN_110_0),
	.A(n26915),
	.B(n26753));
   XNOR2xp5_ASAP7_75t_SL FE_RC_392_0 (.Y(FE_RN_109_0),
	.A(n24846),
	.B(n24845));
   XOR2x2_ASAP7_75t_SL FE_RC_391_0 (.Y(n24849),
	.A(FE_RN_109_0),
	.B(FE_OCPN27446_n24847));
   AND2x2_ASAP7_75t_R FE_RC_390_0 (.Y(FE_RN_108_0),
	.A(n22690),
	.B(n17869));
   NAND2xp5_ASAP7_75t_SL FE_RC_389_0 (.Y(n22704),
	.A(FE_RN_108_0),
	.B(n17868));
   HB1xp67_ASAP7_75t_L FE_OCPC4761_n22547 (.Y(FE_OCPN28196_n22547),
	.A(n22547));
   HB1xp67_ASAP7_75t_SL FE_OCPC4754_n20491 (.Y(FE_OCPN28189_n20491),
	.A(n20491));
   HB1xp67_ASAP7_75t_R FE_OCPC4752_n16806 (.Y(FE_OCPN28187_n16806),
	.A(n16806));
   BUFx2_ASAP7_75t_SL FE_OCPC4751_n16123 (.Y(FE_OCPN28186_n16123),
	.A(n16123));
   BUFx2_ASAP7_75t_SL FE_OCPC4740_n21818 (.Y(FE_OCPN28175_n21818),
	.A(n21818));
   HB1xp67_ASAP7_75t_R FE_OCPC4738_n27153 (.Y(FE_OCPN28173_n27153),
	.A(n27153));
   AND2x2_ASAP7_75t_SRAM FE_RC_388_0 (.Y(FE_RN_107_0),
	.A(n25367),
	.B(n25366));
   BUFx2_ASAP7_75t_SL FE_OCPC4728_FE_OFN99_sa20_5 (.Y(FE_OCPN28163_FE_OFN99_sa20_5),
	.A(FE_OCPN27633_sa20_5));
   HB1xp67_ASAP7_75t_SL FE_OCPC4721_n26304 (.Y(FE_OCPN28156_n26304),
	.A(n26304));
   HB1xp67_ASAP7_75t_L FE_OCPC4715_n27152 (.Y(FE_OCPN28150_n27152),
	.A(n27152));
   HB1xp67_ASAP7_75t_SL FE_OCPC4714_n17121 (.Y(FE_OCPN28149_n17121),
	.A(n17121));
   HB1xp67_ASAP7_75t_SL FE_OCPC4705_FE_OFN133_n24306 (.Y(FE_OCPN28140_FE_OFN133_n24306),
	.A(FE_OFN133_n24306));
   BUFx2_ASAP7_75t_SL FE_OCPC4703_n26654 (.Y(FE_OCPN28138_n26654),
	.A(n26654));
   AO21x1_ASAP7_75t_R FE_RC_386_0 (.Y(FE_RN_106_0),
	.A1(n25307),
	.A2(n17821),
	.B(n26976));
   NAND2x1p5_ASAP7_75t_SL FE_RC_385_0 (.Y(n27212),
	.A(FE_RN_106_0),
	.B(n17820));
   AND2x2_ASAP7_75t_R FE_RC_384_0 (.Y(FE_RN_105_0),
	.A(n26942),
	.B(n26941));
   OAI21x1_ASAP7_75t_SL FE_RC_383_0 (.Y(n27143),
	.A1(FE_RN_105_0),
	.A2(n26940),
	.B(n26939));
   OR2x2_ASAP7_75t_SRAM FE_RC_382_0 (.Y(FE_RN_104_0),
	.A(n17506),
	.B(n26739));
   AOI21x1_ASAP7_75t_SL FE_RC_381_0 (.Y(n26741),
	.A1(FE_RN_104_0),
	.A2(n26738),
	.B(n26737));
   AND2x2_ASAP7_75t_SRAM FE_RC_380_0 (.Y(FE_RN_103_0),
	.A(n26770),
	.B(n26769));
   OAI21x1_ASAP7_75t_SL FE_RC_379_0 (.Y(n26393),
	.A1(FE_RN_103_0),
	.A2(n26391),
	.B(n26390));
   AND2x2_ASAP7_75t_SRAM FE_RC_378_0 (.Y(FE_RN_102_0),
	.A(n26819),
	.B(FE_OCPN8227_n25950));
   OAI21x1_ASAP7_75t_SL FE_RC_377_0 (.Y(n25778),
	.A1(FE_RN_102_0),
	.A2(n24879),
	.B(n24878));
   OA21x2_ASAP7_75t_R FE_RC_376_0 (.Y(FE_RN_101_0),
	.A1(n25331),
	.A2(n25330),
	.B(n26323));
   NOR2x1p5_ASAP7_75t_SL FE_RC_375_0 (.Y(n26749),
	.A(FE_RN_101_0),
	.B(n25921));
   OA21x2_ASAP7_75t_L FE_RC_374_0 (.Y(FE_RN_100_0),
	.A1(n18346),
	.A2(n18345),
	.B(n22405));
   NOR2x1_ASAP7_75t_SL FE_RC_373_0 (.Y(n25146),
	.A(FE_RN_100_0),
	.B(n25020));
   AND2x2_ASAP7_75t_SL FE_RC_372_0 (.Y(FE_RN_99_0),
	.A(n27133),
	.B(n27132));
   OAI21x1_ASAP7_75t_SL FE_RC_371_0 (.Y(n482),
	.A1(FE_RN_99_0),
	.A2(n27131),
	.B(n27130));
   AND2x2_ASAP7_75t_L FE_RC_370_0 (.Y(FE_RN_98_0),
	.A(FE_OFN16177_n27207),
	.B(n26057));
   OAI21x1_ASAP7_75t_SL FE_RC_369_0 (.Y(n27178),
	.A1(FE_RN_98_0),
	.A2(n25344),
	.B(n25343));
   AO21x1_ASAP7_75t_SL FE_RC_368_0 (.Y(FE_RN_97_0),
	.A1(n25731),
	.A2(n25730),
	.B(n25729));
   NAND2x1p5_ASAP7_75t_SL FE_RC_367_0 (.Y(n453),
	.A(FE_RN_97_0),
	.B(n25728));
   AND2x2_ASAP7_75t_R FE_RC_366_0 (.Y(FE_RN_96_0),
	.A(n26282),
	.B(n26250));
   OAI21xp5_ASAP7_75t_SL FE_RC_365_0 (.Y(n25754),
	.A1(FE_RN_96_0),
	.A2(n25753),
	.B(n25752));
   AND2x2_ASAP7_75t_SRAM FE_RC_364_0 (.Y(FE_RN_95_0),
	.A(FE_OFN16329_n27151),
	.B(FE_OFN28483_ld_r));
   OAI21xp5_ASAP7_75t_SL FE_RC_363_0 (.Y(n26647),
	.A1(FE_RN_95_0),
	.A2(n26643),
	.B(n26642));
   AO21x1_ASAP7_75t_R FE_RC_362_0 (.Y(FE_RN_94_0),
	.A1(n24571),
	.A2(n24570),
	.B(n17463));
   NAND2x1_ASAP7_75t_SL FE_RC_361_0 (.Y(n26268),
	.A(FE_RN_94_0),
	.B(n24569));
   XOR2xp5_ASAP7_75t_SL FE_RC_360_0 (.Y(FE_RN_93_0),
	.A(n26891),
	.B(n26890));
   XNOR2x1_ASAP7_75t_SL FE_RC_359_0 (.Y(n26894),
	.A(FE_RN_93_0),
	.B(FE_OCPN28122_n27157));
   AND2x2_ASAP7_75t_SL FE_RC_358_0 (.Y(FE_RN_92_0),
	.A(n25901),
	.B(n18595));
   NAND2xp5_ASAP7_75t_SL FE_RC_357_0 (.Y(n18596),
	.A(FE_RN_92_0),
	.B(n18594));
   AO21x1_ASAP7_75t_L FE_RC_356_0 (.Y(FE_RN_91_0),
	.A1(FE_OCPN29425_n24172),
	.A2(n24171),
	.B(n27102));
   NAND2x1_ASAP7_75t_SL FE_RC_355_0 (.Y(n26236),
	.A(FE_RN_91_0),
	.B(n24170));
   OA21x2_ASAP7_75t_SRAM FE_RC_354_0 (.Y(FE_RN_90_0),
	.A1(w0_4_),
	.A2(text_in_r_100_),
	.B(n25814));
   NOR2x2_ASAP7_75t_SL FE_RC_353_0 (.Y(n497),
	.A(FE_RN_90_0),
	.B(n25813));
   OR2x2_ASAP7_75t_L FE_RC_352_0 (.Y(FE_RN_89_0),
	.A(FE_OFN28561_n25419),
	.B(n25420));
   NAND2x1_ASAP7_75t_SL FE_RC_351_0 (.Y(n25657),
	.A(FE_RN_89_0),
	.B(FE_OCPN27682_n25414));
   AO21x1_ASAP7_75t_SL FE_RC_350_0 (.Y(FE_RN_88_0),
	.A1(n19904),
	.A2(n19903),
	.B(n25585));
   NAND2x1_ASAP7_75t_SL FE_RC_349_0 (.Y(n25379),
	.A(FE_RN_88_0),
	.B(n19902));
   OA21x2_ASAP7_75t_SRAM FE_RC_348_0 (.Y(FE_RN_87_0),
	.A1(w0_1_),
	.A2(text_in_r_97_),
	.B(n25272));
   NOR2x1p5_ASAP7_75t_SL FE_RC_347_0 (.Y(n431),
	.A(FE_RN_87_0),
	.B(n25271));
   AND2x2_ASAP7_75t_SRAM FE_RC_346_0 (.Y(FE_RN_86_0),
	.A(n26942),
	.B(n26201));
   AND2x2_ASAP7_75t_R FE_RC_344_0 (.Y(FE_RN_85_0),
	.A(n26249),
	.B(n25736));
   OAI21x1_ASAP7_75t_SL FE_RC_343_0 (.Y(n25688),
	.A1(FE_RN_85_0),
	.A2(n24385),
	.B(n24384));
   XOR2xp5_ASAP7_75t_SL FE_RC_342_0 (.Y(FE_RN_84_0),
	.A(n26727),
	.B(n26726));
   XNOR2xp5_ASAP7_75t_SL FE_RC_341_0 (.Y(n26731),
	.A(FE_RN_84_0),
	.B(n26728));
   XNOR2xp5_ASAP7_75t_SL FE_RC_340_0 (.Y(FE_RN_83_0),
	.A(n26326),
	.B(n26325));
   XOR2xp5_ASAP7_75t_SL FE_RC_339_0 (.Y(n26329),
	.A(FE_RN_83_0),
	.B(n26324));
   OR2x2_ASAP7_75t_SL FE_RC_338_0 (.Y(FE_RN_82_0),
	.A(n26119),
	.B(n26118));
   AOI21x1_ASAP7_75t_SL FE_RC_337_0 (.Y(FE_OCPN27530_n362),
	.A1(FE_RN_82_0),
	.A2(w0_0_),
	.B(n26117));
   AND2x2_ASAP7_75t_SRAM FE_RC_336_0 (.Y(FE_RN_81_0),
	.A(FE_OCPN28328_n25953),
	.B(FE_OCPN28320_n25954));
   NAND2xp5_ASAP7_75t_SL FE_RC_335_0 (.Y(n25951),
	.A(FE_RN_81_0),
	.B(n25952));
   XOR2xp5_ASAP7_75t_SL FE_RC_334_0 (.Y(FE_RN_80_0),
	.A(n25388),
	.B(n25387));
   XNOR2x1_ASAP7_75t_SL FE_RC_333_0 (.Y(n25392),
	.A(FE_RN_80_0),
	.B(FE_OCPN27292_n25389));
   INVxp33_ASAP7_75t_R FE_RC_332_0 (.Y(FE_RN_77_0),
	.A(n27168));
   NAND2xp33_ASAP7_75t_R FE_RC_330_0 (.Y(FE_RN_79_0),
	.A(FE_RN_77_0),
	.B(FE_RN_78_0));
   OAI221xp5_ASAP7_75t_SL FE_RC_329_0 (.Y(n20891),
	.A1(n20890),
	.A2(n27168),
	.B1(n26404),
	.B2(n27168),
	.C(FE_RN_79_0));
   HB1xp67_ASAP7_75t_SL FE_OCPC4688_n27047 (.Y(FE_OCPN28123_n27047),
	.A(n24306));
   AND2x2_ASAP7_75t_SRAM FE_RC_327_0 (.Y(FE_RN_76_0),
	.A(n26651),
	.B(FE_OCPN29471_n24175));
   NAND2xp5_ASAP7_75t_SL FE_RC_326_0 (.Y(n25511),
	.A(FE_RN_76_0),
	.B(n25512));
   NOR3x2_ASAP7_75t_SL FE_RC_325_0 (.Y(n18919),
	.A(FE_OCPN29544_n20527),
	.B(FE_OCPN29369_n16982),
	.C(FE_OFN29243_n17065));
   INVx1_ASAP7_75t_SL FE_OCPC4685_n16975 (.Y(FE_OCPN28120_n16975),
	.A(n16975));
   NAND2xp5_ASAP7_75t_SL FE_RC_323_0 (.Y(FE_RN_73_0),
	.A(n25150),
	.B(n25151));
   OAI21xp5_ASAP7_75t_SL FE_RC_322_0 (.Y(FE_RN_74_0),
	.A1(n25150),
	.A2(n25151),
	.B(FE_RN_73_0));
   OAI21xp5_ASAP7_75t_SL FE_RC_319_0 (.Y(n26319),
	.A1(n25641),
	.A2(n18611),
	.B(n18610));
   AOI31xp33_ASAP7_75t_SL FE_RC_318_0 (.Y(n25229),
	.A1(n17026),
	.A2(n17025),
	.A3(n19372),
	.B(n27095));
   OAI21xp5_ASAP7_75t_SL FE_RC_316_0 (.Y(n25452),
	.A1(n23622),
	.A2(n24377),
	.B(n24387));
   NAND3x2_ASAP7_75t_SL FE_RC_315_0 (.Y(n18263),
	.A(FE_OFN29234_n16996),
	.B(FE_OCPN29351_FE_OFN26116_sa13_1),
	.C(FE_OCPN27902_n20514));
   AND2x2_ASAP7_75t_L FE_RC_314_0 (.Y(FE_RN_71_0),
	.A(n25575),
	.B(n24749));
   NOR2x2_ASAP7_75t_SL FE_RC_313_0 (.Y(n25133),
	.A(FE_RN_71_0),
	.B(FE_OCPN29262_n24750));
   INVx1_ASAP7_75t_SL FE_RC_310_0 (.Y(FE_RN_66_0),
	.A(FE_RN_69_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_309_0 (.Y(FE_RN_67_0),
	.A(FE_OCPN28355_n26909),
	.B(FE_RN_66_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_308_0 (.Y(FE_RN_68_0),
	.A(n25938),
	.B(n25939));
   OAI21xp33_ASAP7_75t_SL FE_RC_307_0 (.Y(FE_RN_69_0),
	.A1(n25938),
	.A2(n25939),
	.B(FE_RN_68_0));
   OAI21xp5_ASAP7_75t_SL FE_RC_305_0 (.Y(n25942),
	.A1(FE_RN_66_0),
	.A2(FE_OCPN28355_n26909),
	.B(FE_RN_67_0));
   HB1xp67_ASAP7_75t_L FE_OCPC4680_n25293 (.Y(FE_OCPN28115_n25293),
	.A(n25293));
   NAND2xp5_ASAP7_75t_SL FE_RC_301_0 (.Y(FE_RN_64_0),
	.A(n20499),
	.B(n20498));
   NOR2xp33_ASAP7_75t_SL FE_RC_299_0 (.Y(FE_RN_65_0),
	.A(FE_RN_63_0),
	.B(FE_RN_64_0));
   BUFx3_ASAP7_75t_SL FE_OCPC4677_n26664 (.Y(FE_OCPN28112_n26664),
	.A(n26664));
   INVxp33_ASAP7_75t_L FE_OCPC4676_n19091 (.Y(FE_OCPN28111_n19091),
	.A(n18743));
   INVx2_ASAP7_75t_SL FE_OCPC4675_n19091 (.Y(n18743),
	.A(n19091));
   BUFx2_ASAP7_75t_SL FE_OCPC4670_n23504 (.Y(FE_OCPN28107_n23504),
	.A(n23504));
   HB1xp67_ASAP7_75t_R FE_OCPC4662_n25470 (.Y(FE_OCPN28100_n25470),
	.A(n25470));
   BUFx2_ASAP7_75t_SL FE_OCPC4650_n25431 (.Y(FE_OCPN27497_n25431),
	.A(n25431));
   INVxp67_ASAP7_75t_L FE_OCPC4649_n24904 (.Y(n24902),
	.A(n24904));
   INVx1_ASAP7_75t_L FE_OCPC4648_n23913 (.Y(FE_OCPN28089_n23913),
	.A(n23913));
   INVxp33_ASAP7_75t_SRAM FE_OCPC4640_n26574 (.Y(FE_OCPN28083_n26574),
	.A(n26575));
   BUFx3_ASAP7_75t_SL FE_OCPC4637_n21860 (.Y(FE_OCPN28082_n21860),
	.A(n21860));
   HB1xp67_ASAP7_75t_L FE_OCPC4631_n24296 (.Y(FE_OCPN28078_n24296),
	.A(n24296));
   HB1xp67_ASAP7_75t_SL FE_OCPC4630_n25488 (.Y(FE_OCPN28077_n),
	.A(n25488));
   HB1xp67_ASAP7_75t_L FE_OCPC4629_FE_OFN9_w3_6 (.Y(FE_OCPN28076_FE_OFN9_w3_6),
	.A(FE_OFN28699_w3_6));
   BUFx3_ASAP7_75t_SL FE_OCPC4628_n16048 (.Y(FE_OCPN28075_n16048),
	.A(n16048));
   HB1xp67_ASAP7_75t_L FE_OCPC4623_w3_3 (.Y(FE_OCPN28072_w3_3),
	.A(w3_3_));
   BUFx3_ASAP7_75t_SL FE_OCPC4622_n25092 (.Y(FE_OCPN28071_n25092),
	.A(n25092));
   NOR2xp33_ASAP7_75t_L FE_RC_298_0 (.Y(FE_RN_61_0),
	.A(FE_OFN27096_n),
	.B(FE_OFN27214_w3_17));
   INVx1_ASAP7_75t_SL FE_RC_297_0 (.Y(FE_RN_62_0),
	.A(n15514));
   OR2x2_ASAP7_75t_SL FE_RC_296_0 (.Y(n13874),
	.A(FE_RN_62_0),
	.B(FE_RN_61_0));
   OR3x1_ASAP7_75t_SL FE_RC_295_0 (.Y(n13869),
	.A(FE_OFN16426_w3_20),
	.B(FE_OFN28683_w3_21),
	.C(FE_OFN28_w3_23));
   OAI21xp5_ASAP7_75t_L FE_RC_294_0 (.Y(n24915),
	.A1(FE_OCPN8244_n25778),
	.A2(n24916),
	.B(FE_OFN28490_ld_r));
   OAI21xp33_ASAP7_75t_SL FE_RC_292_0 (.Y(n654),
	.A1(FE_OCPN29571_n26355),
	.A2(FE_OFN25904_n16143),
	.B(n16142));
   OR3x1_ASAP7_75t_L FE_RC_290_0 (.Y(FE_RN_60_0),
	.A(n16351),
	.B(n20043),
	.C(n18088));
   BUFx3_ASAP7_75t_SL FE_OCPC4616_n15774 (.Y(FE_OCPN28065_n15774),
	.A(n15774));
   NOR3xp33_ASAP7_75t_L FE_RC_289_0 (.Y(n26035),
	.A(FE_OCPN27373_n26172),
	.B(n26037),
	.C(n26036));
   HB1xp67_ASAP7_75t_R FE_OCPC4612_n20076 (.Y(FE_OCPN28061_n20076),
	.A(n20076));
   OAI21xp5_ASAP7_75t_L FE_RC_282_0 (.Y(n26097),
	.A1(FE_OCPN28140_FE_OFN133_n24306),
	.A2(FE_OCPN5045_n26098),
	.B(FE_OFN28483_ld_r));
   INVx4_ASAP7_75t_SL FE_OCPC4598_n17301 (.Y(n19097),
	.A(n17301));
   INVx1_ASAP7_75t_L FE_OCPC4597_n17750 (.Y(n17752),
	.A(n17750));
   BUFx2_ASAP7_75t_L FE_OCPC4572_n19766 (.Y(FE_OCPN28040_n19766),
	.A(n19766));
   BUFx2_ASAP7_75t_L FE_OCPC4569_n22855 (.Y(FE_OCPN28037_n22855),
	.A(n22855));
   HB1xp67_ASAP7_75t_R FE_OCPC4555_n25770 (.Y(FE_OCPN28023_n25770),
	.A(n25770));
   BUFx4f_ASAP7_75t_SL FE_OCPC4551_n21445 (.Y(FE_OCPN28021_n21445),
	.A(n21445));
   BUFx2_ASAP7_75t_SL FE_OCPC4547_n18548 (.Y(FE_OCPN28017_n18548),
	.A(n18548));
   HB1xp67_ASAP7_75t_SL FE_OCPC4546_n21124 (.Y(FE_OCPN28016_n21124),
	.A(n21124));
   BUFx3_ASAP7_75t_L FE_OCPC4538_n16290 (.Y(FE_OCPN28008_n16290),
	.A(n16290));
   BUFx4f_ASAP7_75t_SL FE_OCPC4536_n17454 (.Y(FE_OCPN28006_n17454),
	.A(n17454));
   OR3x1_ASAP7_75t_SL FE_RC_280_0 (.Y(FE_RN_54_0),
	.A(n18651),
	.B(FE_OCPN29291_n17282),
	.C(FE_OCPN29411_n));
   BUFx2_ASAP7_75t_L FE_OCPC4530_n22450 (.Y(FE_OCPN28000_n22450),
	.A(n22450));
   OAI21xp5_ASAP7_75t_SL FE_RC_279_0 (.Y(n25348),
	.A1(FE_OCPN7629_FE_OFN105_n27178),
	.A2(n25349),
	.B(FE_OFN16215_ld_r));
   BUFx4f_ASAP7_75t_SL FE_OCPC4528_n18019 (.Y(FE_OCPN27998_n18019),
	.A(n18019));
   HB1xp67_ASAP7_75t_SL FE_OCPC4520_FE_OFN16132_sa03_5 (.Y(FE_OCPN27990_FE_OFN16132_sa03_5),
	.A(FE_OFN28689_sa03_5));
   BUFx2_ASAP7_75t_L FE_OCPC4515_n24831 (.Y(FE_OCPN27985_n24831),
	.A(n24831));
   OR3x1_ASAP7_75t_SL FE_RC_277_0 (.Y(FE_RN_53_0),
	.A(n16343),
	.B(n16342),
	.C(n21982));
   HB1xp67_ASAP7_75t_SL FE_OCPC4509_FE_OFN16147_sa22_1 (.Y(FE_OCPN27979_FE_OFN16147_sa22_1),
	.A(FE_OCPN29269_sa22_1));
   BUFx5_ASAP7_75t_SL FE_OCPC4508_w3_3 (.Y(FE_OCPN27978_w3_3),
	.A(w3_3_));
   BUFx3_ASAP7_75t_SL FE_OCPC4501_n21627 (.Y(FE_OCPN27971_n21627),
	.A(n21627));
   BUFx2_ASAP7_75t_SL FE_OCPC4493_n18473 (.Y(FE_OCPN27966_n18473),
	.A(n18473));
   NAND3xp33_ASAP7_75t_SL FE_RC_276_0 (.Y(n25050),
	.A(n25053),
	.B(n25052),
	.C(n25051));
   INVxp33_ASAP7_75t_R FE_OCPC4481_sa23_1 (.Y(n23510),
	.A(FE_OCPN27627_sa23_1));
   INVx1_ASAP7_75t_SL FE_OCPC4477_n22945 (.Y(FE_OFN25883_n22945),
	.A(n22945));
   HB1xp67_ASAP7_75t_SL FE_OCPC4471_FE_OFN26173_n21511 (.Y(FE_OCPN27948_FE_OFN26173_n21511),
	.A(FE_OFN29182_n21708));
   AND2x2_ASAP7_75t_L FE_RC_275_0 (.Y(FE_RN_52_0),
	.A(n25591),
	.B(n25592));
   NAND2xp5_ASAP7_75t_SL FE_RC_274_0 (.Y(n25590),
	.A(FE_RN_52_0),
	.B(n26852));
   HB1xp67_ASAP7_75t_SL FE_OCPC4452_FE_OFN4_w3_22 (.Y(FE_OCPN27929_FE_OFN4_w3_22),
	.A(FE_OFN4_w3_22));
   HB1xp67_ASAP7_75t_SL FE_OCPC4451_FE_OFN4_w3_22 (.Y(FE_OCPN27928_FE_OFN4_w3_22),
	.A(FE_OFN4_w3_22));
   BUFx3_ASAP7_75t_SL FE_OCPC4441_n20155 (.Y(FE_OCPN27919_n20155),
	.A(n20155));
   HB1xp67_ASAP7_75t_R FE_OCPC4438_sa23_2 (.Y(FE_OCPN27916_n),
	.A(FE_OFN29191_sa23_2));
   BUFx2_ASAP7_75t_L FE_OCPC4422_n19223 (.Y(FE_OCPN27903_n19223),
	.A(n19223));
   BUFx2_ASAP7_75t_SL FE_OCPC4415_n18583 (.Y(FE_OCPN27896_n18583),
	.A(n18583));
   BUFx3_ASAP7_75t_SL FE_OCPC4407_sa12_2 (.Y(FE_OCPN27888_sa12_2),
	.A(sa12_2_));
   BUFx2_ASAP7_75t_SL FE_OCPC4406_n17331 (.Y(FE_OCPN27887_n17331),
	.A(n17331));
   BUFx2_ASAP7_75t_SL FE_OCPC4401_n26717 (.Y(FE_OCPN27884_n26717),
	.A(n26717));
   BUFx4f_ASAP7_75t_SL FE_OCPC4399_n18829 (.Y(FE_OCPN27882_n18829),
	.A(n18829));
   BUFx2_ASAP7_75t_L FE_OCPC4387_n17317 (.Y(FE_OCPN27871_n17317),
	.A(n17317));
   BUFx3_ASAP7_75t_SL FE_OCPC4341_n25169 (.Y(FE_OCPN27825_n25169),
	.A(n25169));
   BUFx2_ASAP7_75t_L FE_OCPC4335_n17245 (.Y(FE_OCPN27819_n17245),
	.A(n17245));
   INVxp67_ASAP7_75t_L FE_OCPC4333_n23960 (.Y(n23959),
	.A(n23960));
   HB1xp67_ASAP7_75t_SL FE_OCPC4308_n23375 (.Y(FE_OCPN27807_n23375),
	.A(n23375));
   INVxp67_ASAP7_75t_SL FE_OCPC4306_n25497 (.Y(FE_OCPN27806_n25497),
	.A(n25497));
   INVx2_ASAP7_75t_SL FE_OCPC4300_sa12_1 (.Y(FE_OFN16131_sa12_1),
	.A(sa12_1_));
   INVxp33_ASAP7_75t_R FE_RC_273_0 (.Y(FE_RN_46_0),
	.A(n26607));
   INVxp67_ASAP7_75t_L FE_RC_272_0 (.Y(FE_RN_47_0),
	.A(n23616));
   NAND2xp5_ASAP7_75t_L FE_RC_271_0 (.Y(FE_RN_48_0),
	.A(FE_RN_46_0),
	.B(FE_RN_47_0));
   INVxp33_ASAP7_75t_R FE_RC_270_0 (.Y(FE_RN_49_0),
	.A(n26607));
   INVxp33_ASAP7_75t_L FE_RC_269_0 (.Y(FE_RN_50_0),
	.A(n23617));
   NAND2xp33_ASAP7_75t_L FE_RC_268_0 (.Y(FE_RN_51_0),
	.A(FE_RN_49_0),
	.B(FE_RN_50_0));
   OAI211xp5_ASAP7_75t_SL FE_RC_267_0 (.Y(n23619),
	.A1(n26607),
	.A2(n23618),
	.B(FE_RN_51_0),
	.C(FE_RN_48_0));
   INVx2_ASAP7_75t_SL FE_OCPC4274_sa00_3 (.Y(FE_OCPN27337_n19149),
	.A(sa00_3_));
   HB1xp67_ASAP7_75t_L FE_OCPC4269_n16490 (.Y(FE_OCPN27786_n16490),
	.A(n16490));
   HB1xp67_ASAP7_75t_L FE_OCPC4263_n16873 (.Y(FE_OCPN27782_n16873),
	.A(n16873));
   HB1xp67_ASAP7_75t_L FE_OCPC4261_n20083 (.Y(FE_OCPN27780_n20083),
	.A(n20083));
   HB1xp67_ASAP7_75t_L FE_OCPC4251_n22070 (.Y(FE_OCPN27773_n22070),
	.A(n22070));
   INVx5_ASAP7_75t_SL FE_OCPC4249_sa02_0 (.Y(FE_OCPN27261_sa02_0),
	.A(FE_OCPN27276_sa02_0));
   HB1xp67_ASAP7_75t_SL FE_OCPC4236_FE_OFN16265_n26527 (.Y(FE_OCPN27765_FE_OFN16265_n26527),
	.A(FE_OFN16265_n26527));
   BUFx2_ASAP7_75t_L FE_OCPC4235_n22152 (.Y(FE_OCPN27764_n22152),
	.A(n22152));
   BUFx3_ASAP7_75t_SL FE_OCPC4228_n21819 (.Y(FE_OCPN27757_n21819),
	.A(n21819));
   HB1xp67_ASAP7_75t_L FE_OCPC4214_n22009 (.Y(FE_OCPN27743_n22009),
	.A(n22009));
   BUFx3_ASAP7_75t_SL FE_OCPC4201_n17996 (.Y(FE_OCPN27733_n17996),
	.A(n17996));
   BUFx4f_ASAP7_75t_SL FE_OCPC4197_n17464 (.Y(FE_OCPN27730_n17464),
	.A(n17464));
   BUFx2_ASAP7_75t_L FE_OCPC4196_n24362 (.Y(FE_OCPN27729_n24362),
	.A(n24362));
   BUFx2_ASAP7_75t_L FE_OCPC4194_n22964 (.Y(FE_OCPN27727_n22964),
	.A(n22964));
   HB1xp67_ASAP7_75t_L FE_OCPC4190_n25485 (.Y(FE_OCPN27723_n),
	.A(n25485));
   BUFx2_ASAP7_75t_L FE_OCPC4189_n23336 (.Y(FE_OCPN27722_n23336),
	.A(n23336));
   BUFx2_ASAP7_75t_SL FE_OCPC4188_n23336 (.Y(FE_OCPN27721_n23336),
	.A(n23336));
   BUFx2_ASAP7_75t_SL FE_OCPC4170_n19847 (.Y(FE_OCPN27703_n19847),
	.A(n19847));
   BUFx2_ASAP7_75t_SL FE_OCPC4160_n16309 (.Y(FE_OCPN27697_n16309),
	.A(n16309));
   BUFx2_ASAP7_75t_SL FE_OCPC4153_n16757 (.Y(FE_OCPN27690_n16757),
	.A(n16757));
   HB1xp67_ASAP7_75t_L FE_OCPC4152_n20172 (.Y(FE_OCPN27689_n20172),
	.A(n20172));
   INVxp33_ASAP7_75t_L FE_OCPC4147_n17139 (.Y(FE_OCPN27684_n17139),
	.A(n17004));
   INVx1_ASAP7_75t_SL FE_OCPC4146_n17139 (.Y(n17004),
	.A(n17139));
   BUFx2_ASAP7_75t_L FE_OCPC4135_n18163 (.Y(FE_OCPN27673_n18163),
	.A(FE_OFN28688_sa22_2));
   NOR3xp33_ASAP7_75t_L FE_RC_266_0 (.Y(n24994),
	.A(n24992),
	.B(n24991),
	.C(n24993));
   HB1xp67_ASAP7_75t_L FE_OCPC4127_w3_25 (.Y(FE_OCPN27665_w3_25),
	.A(FE_OCPN27655_w3_25));
   BUFx3_ASAP7_75t_SL FE_OCPC4121_w3_25 (.Y(FE_OCPN27659_w3_25),
	.A(FE_OCPN27655_w3_25));
   BUFx5_ASAP7_75t_SL FE_OCPC4118_w3_25 (.Y(FE_OCPN27656_w3_25),
	.A(w3_25_));
   INVx3_ASAP7_75t_L FE_OCPC4117_w3_25 (.Y(FE_OCPN27655_w3_25),
	.A(w3_25_));
   BUFx3_ASAP7_75t_SL FE_OCPC4106_n17236 (.Y(FE_OCPN27649_n17236),
	.A(n17236));
   INVxp33_ASAP7_75t_L FE_RC_258_0 (.Y(FE_RN_39_0),
	.A(n19483));
   NAND2xp33_ASAP7_75t_L FE_RC_257_0 (.Y(FE_RN_40_0),
	.A(FE_RN_38_0),
	.B(FE_RN_39_0));
   BUFx2_ASAP7_75t_SL FE_OCPC4089_n26223 (.Y(n26222),
	.A(n26223));
   BUFx3_ASAP7_75t_SL FE_OCPC4088_n21725 (.Y(FE_OFN27133_n21725),
	.A(n21725));
   INVxp67_ASAP7_75t_L FE_OCPC4084_n26851 (.Y(FE_OCPN27295_n26851),
	.A(n26851));
   BUFx3_ASAP7_75t_SL FE_OCPC4083_n26851 (.Y(n26852),
	.A(n26851));
   INVx1_ASAP7_75t_SL FE_OCPC4079_n26428 (.Y(n26427),
	.A(n26428));
   HB1xp67_ASAP7_75t_L FE_OCPC4063_n25589 (.Y(FE_OCPN27629_n25589),
	.A(n25589));
   BUFx3_ASAP7_75t_SL FE_OCPC4040_n23869 (.Y(FE_OCPN27606_n23869),
	.A(n23869));
   BUFx2_ASAP7_75t_L FE_OCPC4027_n16908 (.Y(FE_OCPN27593_n16908),
	.A(n16908));
   AND2x2_ASAP7_75t_R FE_RC_255_0 (.Y(FE_RN_37_0),
	.A(n26412),
	.B(FE_OCPN29443_n25507));
   NAND2xp5_ASAP7_75t_L FE_RC_254_0 (.Y(n26410),
	.A(FE_RN_37_0),
	.B(FE_OCPN7589_n26420));
   BUFx3_ASAP7_75t_SL FE_OCPC4018_n19824 (.Y(FE_OCPN27588_n19824),
	.A(n19824));
   BUFx3_ASAP7_75t_SL FE_OCPC4015_sa02_1 (.Y(FE_OCPN27585_sa02_1),
	.A(sa02_1_));
   INVx1_ASAP7_75t_SL FE_OCPC4014_sa02_1 (.Y(FE_OCPN27572_sa02_1),
	.A(sa02_1_));
   HB1xp67_ASAP7_75t_L FE_OCPC4012_n22497 (.Y(FE_OCPN27584_n22497),
	.A(n22497));
   INVxp67_ASAP7_75t_L FE_OCPC4010_n25935 (.Y(FE_OFN27142_n25934),
	.A(n25935));
   BUFx3_ASAP7_75t_SL FE_OCPC4004_n26389 (.Y(FE_OCPN27310_n26389),
	.A(n26389));
   OAI22xp33_ASAP7_75t_L FE_RC_253_0 (.Y(n22379),
	.A1(FE_OCPN28229_n17529),
	.A2(n20107),
	.B1(n22392),
	.B2(n20107));
   BUFx2_ASAP7_75t_L FE_OCPC3996_FE_OFN16132_sa03_5 (.Y(FE_OCPN27483_FE_OFN16132_sa03_5),
	.A(FE_OFN28689_sa03_5));
   INVxp67_ASAP7_75t_SL FE_OCPC3994_n27151 (.Y(FE_OFN16331_n27151),
	.A(n27151));
   HB1xp67_ASAP7_75t_SL FE_OCPC3993_n27151 (.Y(FE_OFN16329_n27151),
	.A(n27151));
   NAND3x1_ASAP7_75t_SL FE_RC_252_0 (.Y(n16421),
	.A(FE_OFN28694_sa33_4),
	.B(FE_OCPN27568_sa33_3),
	.C(FE_OFN28679_sa33_5));
   BUFx3_ASAP7_75t_SL FE_OCPC3987_n16913 (.Y(FE_OCPN27460_n16913),
	.A(n16913));
   HB1xp67_ASAP7_75t_L FE_OCPC3985_n20196 (.Y(FE_OCPN27574_n20196),
	.A(FE_OCPN27573_n20196));
   BUFx3_ASAP7_75t_SL FE_OCPC3984_n20196 (.Y(FE_OCPN27573_n20196),
	.A(n20196));
   INVx3_ASAP7_75t_L FE_OCPC3972_n17791 (.Y(FE_OCPN27570_n17791),
	.A(n17791));
   INVx3_ASAP7_75t_SL FE_OCPC3961_sa33_3 (.Y(n16438),
	.A(sa33_3_));
   HB1xp67_ASAP7_75t_SRAM FE_OCPC3948_n25755 (.Y(FE_OCPN27560_n25755),
	.A(FE_OCPN27322_n25755));
   OAI21xp5_ASAP7_75t_SL FE_RC_245_0 (.Y(n25650),
	.A1(n25651),
	.A2(n25652),
	.B(FE_OFN16215_ld_r));
   BUFx2_ASAP7_75t_SL FE_OCPC3940_n17843 (.Y(FE_OCPN27556_n17843),
	.A(n17843));
   NAND2xp5_ASAP7_75t_SL FE_RC_243_0 (.Y(FE_RN_27_0),
	.A(n27142),
	.B(FE_RN_26_0));
   OAI21xp5_ASAP7_75t_SL FE_RC_238_0 (.Y(n27146),
	.A1(FE_RN_26_0),
	.A2(n27142),
	.B(FE_RN_27_0));
   INVx1_ASAP7_75t_SL FE_OCPC3907_n25383 (.Y(n25384),
	.A(n25383));
   BUFx6f_ASAP7_75t_SL FE_OCPC3895_sa00_5 (.Y(FE_OCPN27227_sa00_5),
	.A(sa00_5_));
   INVx1_ASAP7_75t_SL FE_OCPC3894_sa00_5 (.Y(FE_OCPN27224_sa00_5),
	.A(sa00_5_));
   NAND2xp33_ASAP7_75t_SL FE_RC_236_0 (.Y(FE_RN_23_0),
	.A(FE_OCPN27678_n26227),
	.B(n26128));
   OAI21xp33_ASAP7_75t_SL FE_RC_235_0 (.Y(FE_RN_24_0),
	.A1(FE_OCPN27678_n26227),
	.A2(n26128),
	.B(FE_RN_23_0));
   INVx2_ASAP7_75t_SL FE_OCPC3889_sa21_4 (.Y(FE_OCPN27388_FE_OFN25990_sa21_4),
	.A(sa21_4_));
   INVx2_ASAP7_75t_SL FE_OCPC3883_sa02_0 (.Y(FE_OCPN27276_sa02_0),
	.A(sa02_0_));
   INVxp67_ASAP7_75t_SL FE_OCPC3878_n25362 (.Y(n25360),
	.A(n25362));
   HB1xp67_ASAP7_75t_R FE_OCPC3876_n25921 (.Y(FE_OCPN27522_n25921),
	.A(n25921));
   HB1xp67_ASAP7_75t_L FE_OCPC3875_n18163 (.Y(FE_OCPN27521_n18163),
	.A(FE_OFN28688_sa22_2));
   BUFx4f_ASAP7_75t_SL FE_OCPC3872_n17251 (.Y(FE_OCPN27518_n17251),
	.A(n17251));
   BUFx6f_ASAP7_75t_SL FE_OCPC3866_sa11_2 (.Y(FE_OCPN27512_sa11_2),
	.A(sa11_2_));
   BUFx3_ASAP7_75t_SL FE_OCPC3861_n25695 (.Y(FE_OCPN27507_n25695),
	.A(n25695));
   BUFx2_ASAP7_75t_SL FE_OCPC3859_n24684 (.Y(FE_OCPN27505_n24684),
	.A(n24684));
   BUFx3_ASAP7_75t_SL FE_OCPC3850_n21820 (.Y(FE_OCPN27496_n21820),
	.A(n21820));
   BUFx3_ASAP7_75t_SL FE_OCPC3848_n26479 (.Y(FE_OCPN27494_n26479),
	.A(n26479));
   BUFx2_ASAP7_75t_SL FE_OCPC3844_n18798 (.Y(FE_OCPN27490_n18798),
	.A(n18798));
   AND2x2_ASAP7_75t_SRAM FE_RC_232_0 (.Y(FE_RN_21_0),
	.A(n20333),
	.B(n19884));
   NAND2x1_ASAP7_75t_SL FE_RC_231_0 (.Y(n25578),
	.A(FE_RN_21_0),
	.B(n19883));
   HB1xp67_ASAP7_75t_SL FE_OCPC3832_n25011 (.Y(FE_OCPN27478_n25011),
	.A(n25011));
   HB1xp67_ASAP7_75t_L FE_OCPC3830_n26852 (.Y(FE_OCPN27476_n26852),
	.A(FE_OCPN27295_n26851));
   HB1xp67_ASAP7_75t_L FE_OCPC3812_n24891 (.Y(FE_OCPN27458_n24891),
	.A(n24891));
   HB1xp67_ASAP7_75t_R FE_OCPC3805_n26236 (.Y(FE_OCPN27451_n26236),
	.A(n26236));
   BUFx3_ASAP7_75t_SL FE_OCPC3799_n26837 (.Y(FE_OCPN27445_n26837),
	.A(n26837));
   HB1xp67_ASAP7_75t_SL FE_OCPC3796_n27202 (.Y(FE_OCPN27442_n27202),
	.A(n27202));
   BUFx2_ASAP7_75t_L FE_OCPC3795_n25688 (.Y(FE_OCPN27441_n25688),
	.A(n25688));
   BUFx2_ASAP7_75t_L FE_OCPC3778_n22560 (.Y(FE_OCPN27424_n22560),
	.A(n22560));
   BUFx2_ASAP7_75t_SL FE_OCPC3775_n25768 (.Y(FE_OCPN27421_n25768),
	.A(n25768));
   BUFx2_ASAP7_75t_SL FE_OCPC3774_n18794 (.Y(FE_OCPN27420_n18794),
	.A(n18794));
   BUFx3_ASAP7_75t_SL FE_OCPC3753_n22598 (.Y(FE_OCPN27399_n22598),
	.A(n22598));
   BUFx3_ASAP7_75t_SL FE_OCPC3745_n27079 (.Y(FE_OCPN27391_n27079),
	.A(n27079));
   BUFx3_ASAP7_75t_SL FE_OCPC3738_n22888 (.Y(FE_OCPN27384_n22888),
	.A(n22888));
   BUFx3_ASAP7_75t_SL FE_OCPC3728_n26394 (.Y(FE_OCPN27374_n26394),
	.A(n26394));
   BUFx2_ASAP7_75t_SL FE_OCPC3720_n26326 (.Y(FE_OCPN27366_n26326),
	.A(n26326));
   BUFx2_ASAP7_75t_SL FE_OCPC3717_n26649 (.Y(FE_OCPN27363_n26649),
	.A(n26649));
   BUFx2_ASAP7_75t_SL FE_OCPC3716_n25679 (.Y(FE_OCPN27362_n25679),
	.A(n25679));
   HB1xp67_ASAP7_75t_SL FE_OCPC3713_n26726 (.Y(FE_OCPN27359_n26726),
	.A(n26726));
   BUFx2_ASAP7_75t_SL FE_OCPC3687_n25250 (.Y(FE_OCPN27333_n25250),
	.A(n25250));
   BUFx3_ASAP7_75t_SL FE_OCPC3674_n410 (.Y(FE_OCPN27320_n410),
	.A(n410));
   BUFx2_ASAP7_75t_L FE_OCPC3670_n25849 (.Y(FE_OCPN27316_n25849),
	.A(n25849));
   BUFx2_ASAP7_75t_SL FE_OCPC3643_sa21_5 (.Y(FE_OCPN27289_sa21_5),
	.A(n16783));
   BUFx3_ASAP7_75t_SL FE_OCPC3638_n26633 (.Y(FE_OCPN27284_n26633),
	.A(n26633));
   BUFx2_ASAP7_75t_SL FE_OCPC3637_n26867 (.Y(FE_OCPN27283_n26867),
	.A(n26867));
   BUFx2_ASAP7_75t_SL FE_OCPC3628_n26394 (.Y(FE_OCPN27274_n26394),
	.A(FE_OCPN27374_n26394));
   BUFx2_ASAP7_75t_SL FE_OCPC3621_n18794 (.Y(FE_OCPN27267_n18794),
	.A(n18794));
   BUFx2_ASAP7_75t_SL FE_OCPC3607_n17923 (.Y(FE_OCPN27253_n17923),
	.A(n17923));
   BUFx3_ASAP7_75t_SL FE_OCPC3600_n22663 (.Y(FE_OCPN27246_n22663),
	.A(n22663));
   BUFx3_ASAP7_75t_SL FE_OCPC3588_n26837 (.Y(FE_OCPN27234_n26837),
	.A(FE_OCPN27445_n26837));
   INVx1_ASAP7_75t_SL FE_RC_230_0 (.Y(FE_RN_16_0),
	.A(FE_RN_19_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_229_0 (.Y(FE_RN_17_0),
	.A(FE_OCPN7657_n26213),
	.B(FE_RN_16_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_228_0 (.Y(FE_RN_18_0),
	.A(n26214),
	.B(n26215));
   OAI21xp33_ASAP7_75t_SL FE_RC_227_0 (.Y(FE_RN_19_0),
	.A1(n26214),
	.A2(n26215),
	.B(FE_RN_18_0));
   OAI21xp5_ASAP7_75t_SL FE_RC_225_0 (.Y(n26217),
	.A1(FE_RN_16_0),
	.A2(FE_OCPN7657_n26213),
	.B(FE_RN_17_0));
   NAND2xp33_ASAP7_75t_L FE_RC_222_0 (.Y(FE_RN_15_0),
	.A(FE_OFN16315_sa31_5),
	.B(FE_OFN28933_n16321));
   NOR2x1_ASAP7_75t_L FE_RC_221_0 (.Y(n18072),
	.A(FE_RN_15_0),
	.B(n21981));
   INVxp33_ASAP7_75t_L FE_RC_220_0 (.Y(FE_RN_10_0),
	.A(n18837));
   NOR2xp33_ASAP7_75t_L FE_RC_219_0 (.Y(FE_RN_11_0),
	.A(FE_OFN27148_sa32_3),
	.B(n19721));
   INVx1_ASAP7_75t_SL FE_RC_218_0 (.Y(n18846),
	.A(FE_RN_12_0));
   NAND2xp5_ASAP7_75t_SL FE_RC_217_0 (.Y(FE_RN_12_0),
	.A(FE_RN_10_0),
	.B(FE_RN_11_0));
   NOR2xp33_ASAP7_75t_L FE_RC_216_0 (.Y(FE_RN_7_0),
	.A(n21844),
	.B(n21819));
   INVx2_ASAP7_75t_L FE_RC_214_0 (.Y(n21406),
	.A(FE_RN_9_0));
   NAND2xp5_ASAP7_75t_L FE_RC_213_0 (.Y(FE_RN_9_0),
	.A(FE_RN_7_0),
	.B(FE_RN_8_0));
   NOR2x1_ASAP7_75t_SL FE_RC_211_0 (.Y(FE_RN_6_0),
	.A(FE_OFN29249_n),
	.B(FE_OCPN29260_sa00_5));
   AND2x4_ASAP7_75t_SL FE_RC_210_0 (.Y(n17245),
	.A(n17248),
	.B(FE_RN_6_0));
   AOI21xp5_ASAP7_75t_SL FE_RC_209_0 (.Y(n15370),
	.A1(n25931),
	.A2(n15371),
	.B(n16125));
   AOI21xp33_ASAP7_75t_SL FE_RC_208_0 (.Y(n16174),
	.A1(n26512),
	.A2(n16175),
	.B(ld));
   AOI21xp33_ASAP7_75t_SL FE_RC_206_0 (.Y(n595),
	.A1(key_40_),
	.A2(ld),
	.B(n16272));
   AOI21xp5_ASAP7_75t_SL FE_RC_205_0 (.Y(n16090),
	.A1(n25247),
	.A2(n16091),
	.B(FE_OFN21_n16125));
   AOI21x1_ASAP7_75t_SL FE_RC_204_0 (.Y(n15909),
	.A1(n26310),
	.A2(n15910),
	.B(ld));
   AOI31xp33_ASAP7_75t_SL FE_RC_203_0 (.Y(n23669),
	.A1(n23667),
	.A2(n23666),
	.A3(n23668),
	.B(n25585));
   AOI21xp5_ASAP7_75t_SL FE_RC_202_0 (.Y(n19081),
	.A1(n19079),
	.A2(FE_OFN16163_n26584),
	.B(n19080));
   AOI31xp33_ASAP7_75t_L FE_RC_200_0 (.Y(n21336),
	.A1(n21316),
	.A2(n21315),
	.A3(FE_OCPN7644_n21523),
	.B(n23945));
   AOI21xp5_ASAP7_75t_L FE_RC_198_0 (.Y(n571),
	.A1(key_44_),
	.A2(ld),
	.B(n16202));
   AOI21xp5_ASAP7_75t_SL FE_RC_197_0 (.Y(n583),
	.A1(key_42_),
	.A2(ld),
	.B(n16223));
   AOI21xp5_ASAP7_75t_SL FE_RC_196_0 (.Y(n16133),
	.A1(n25841),
	.A2(n16134),
	.B(ld));
   AOI21xp5_ASAP7_75t_SL FE_RC_195_0 (.Y(n16178),
	.A1(n26018),
	.A2(n16179),
	.B(n16125));
   AOI21x1_ASAP7_75t_SL FE_RC_194_0 (.Y(n16102),
	.A1(n26656),
	.A2(n16103),
	.B(FE_OFN0_ld));
   AOI21xp5_ASAP7_75t_SL FE_RC_193_0 (.Y(n16193),
	.A1(n26416),
	.A2(n16194),
	.B(FE_OFN21_n16125));
   AOI21x1_ASAP7_75t_SL FE_RC_192_0 (.Y(n26574),
	.A1(FE_OCPN29352_n25173),
	.A2(n26282),
	.B(n25174));
   AOI21xp5_ASAP7_75t_SL FE_RC_191_0 (.Y(n23466),
	.A1(n23464),
	.A2(n26819),
	.B(n23465));
   AOI31xp33_ASAP7_75t_L FE_RC_190_0 (.Y(n19746),
	.A1(n19744),
	.A2(n19743),
	.A3(n19745),
	.B(n26346));
   AOI21xp33_ASAP7_75t_L FE_RC_189_0 (.Y(n23114),
	.A1(n23112),
	.A2(FE_OCPN8226_n23113),
	.B(n26464));
   AOI21xp5_ASAP7_75t_SL FE_RC_188_0 (.Y(n22571),
	.A1(n22569),
	.A2(n27216),
	.B(n22570));
   AOI21xp5_ASAP7_75t_SL FE_RC_187_0 (.Y(n24569),
	.A1(n19236),
	.A2(n26082),
	.B(n19237));
   AOI21xp5_ASAP7_75t_SL FE_RC_186_0 (.Y(n25040),
	.A1(n17231),
	.A2(n24974),
	.B(n17232));
   AOI21xp33_ASAP7_75t_SL FE_RC_184_0 (.Y(n17597),
	.A1(n17596),
	.A2(n18813),
	.B(n17584));
   AOI21xp5_ASAP7_75t_SL FE_RC_183_0 (.Y(n14403),
	.A1(n14400),
	.A2(n15757),
	.B(n14401));
   AOI31xp33_ASAP7_75t_SL FE_RC_181_0 (.Y(n20280),
	.A1(n20279),
	.A2(n20278),
	.A3(n24218),
	.B(n26710));
   AOI31xp33_ASAP7_75t_SRAM FE_RC_180_0 (.Y(n20475),
	.A1(n20452),
	.A2(n20478),
	.A3(n20476),
	.B(n26926));
   AOI31xp33_ASAP7_75t_SL FE_RC_179_0 (.Y(n19497),
	.A1(n19477),
	.A2(n19476),
	.A3(n21026),
	.B(n23945));
   AOI31xp33_ASAP7_75t_L FE_RC_178_0 (.Y(n22360),
	.A1(n22347),
	.A2(n22346),
	.A3(n22348),
	.B(n24263));
   AOI31xp33_ASAP7_75t_SL FE_RC_177_0 (.Y(n20696),
	.A1(n20694),
	.A2(n20693),
	.A3(n20695),
	.B(n25641));
   AOI31xp33_ASAP7_75t_R FE_RC_175_0 (.Y(n15053),
	.A1(n15040),
	.A2(n15030),
	.A3(n15031),
	.B(n15881));
   AOI31xp33_ASAP7_75t_L FE_RC_174_0 (.Y(n13948),
	.A1(n15922),
	.A2(FE_OFN29063_n25433),
	.A3(FE_OCPN29521_n24755),
	.B(n13939));
   AOI31xp33_ASAP7_75t_L FE_RC_173_0 (.Y(n14727),
	.A1(n15973),
	.A2(n15922),
	.A3(FE_OCPN29521_n24755),
	.B(n14726));
   AOI21xp5_ASAP7_75t_L FE_RC_172_0 (.Y(n15726),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(FE_OFN25915_n15514),
	.B(n15713));
   AOI31xp67_ASAP7_75t_L FE_RC_171_0 (.Y(n15589),
	.A1(FE_OFN28829_n),
	.A2(FE_OFN26057_w3_1),
	.A3(FE_OFN29209_FE_OCPN27978_w3_3),
	.B(n14410));
   AOI31xp67_ASAP7_75t_SL FE_RC_170_0 (.Y(n14215),
	.A1(FE_OFN26532_n13766),
	.A2(n15835),
	.A3(FE_OFN28747_n),
	.B(n14211));
   AOI21xp5_ASAP7_75t_SL FE_RC_169_0 (.Y(n26065),
	.A1(FE_OCPN27562_n17447),
	.A2(FE_OFN29061_n22505),
	.B(n17507));
   AOI21xp5_ASAP7_75t_SL FE_RC_168_0 (.Y(n15162),
	.A1(FE_OCPN27655_w3_25),
	.A2(FE_OFN27208_w3_30),
	.B(n14504));
   AOI21xp5_ASAP7_75t_SL FE_RC_167_0 (.Y(n22516),
	.A1(FE_OCPN27229_sa11_2),
	.A2(n21834),
	.B(n24565));
   AOI21x1_ASAP7_75t_SL FE_RC_165_0 (.Y(n26488),
	.A1(text_in_r_112_),
	.A2(FE_OFN2_ld_r),
	.B(n26483));
   AOI21xp5_ASAP7_75t_SL FE_RC_164_0 (.Y(n26450),
	.A1(text_in_r_95_),
	.A2(FE_OFN16213_ld_r),
	.B(n26444));
   AOI21xp5_ASAP7_75t_SL FE_RC_162_0 (.Y(n16183),
	.A1(n16184),
	.A2(w2_6_),
	.B(FE_OFN21_n16125));
   AOI21xp5_ASAP7_75t_SL FE_RC_161_0 (.Y(n25413),
	.A1(text_in_r_79_),
	.A2(FE_OFN16214_ld_r),
	.B(n25408));
   AOI21xp5_ASAP7_75t_SL FE_RC_160_0 (.Y(n26063),
	.A1(text_in_r_63_),
	.A2(FE_OFN1_ld_r),
	.B(n26058));
   AOI21xp5_ASAP7_75t_L FE_RC_157_0 (.Y(n559),
	.A1(key_46_),
	.A2(FE_OFN21_n16125),
	.B(n16095));
   AOI21xp5_ASAP7_75t_SL FE_RC_156_0 (.Y(n26357),
	.A1(text_in_r_31_),
	.A2(FE_OFN28482_ld_r),
	.B(n26352));
   BUFx4f_ASAP7_75t_SL FE_RC_155_0 (.Y(FE_OFN16246_n16113),
	.A(n16113));
   AOI21xp5_ASAP7_75t_SL FE_RC_154_0 (.Y(n25731),
	.A1(text_in_r_80_),
	.A2(FE_OFN16214_ld_r),
	.B(n25726));
   AOI21x1_ASAP7_75t_SL FE_RC_153_0 (.Y(n16242),
	.A1(n27219),
	.A2(n16243),
	.B(ld));
   AOI21xp5_ASAP7_75t_L FE_RC_152_0 (.Y(n607),
	.A1(key_45_),
	.A2(ld),
	.B(FE_OCPN29452_n16240));
   AOI21x1_ASAP7_75t_SL FE_RC_151_0 (.Y(n24315),
	.A1(FE_OCPN7622_n24526),
	.A2(n27127),
	.B(FE_OCPN27402_n24523));
   AOI21xp5_ASAP7_75t_SL FE_RC_150_0 (.Y(n15366),
	.A1(n24200),
	.A2(n15367),
	.B(ld));
   AOI21x1_ASAP7_75t_SL FE_RC_149_0 (.Y(n16144),
	.A1(n27135),
	.A2(n16145),
	.B(FE_OFN0_ld));
   AOI21x1_ASAP7_75t_SL FE_RC_148_0 (.Y(n24537),
	.A1(n24309),
	.A2(n26770),
	.B(n24310));
   AOI21xp5_ASAP7_75t_SL FE_RC_147_0 (.Y(n16267),
	.A1(n27173),
	.A2(n16268),
	.B(FE_OFN21_n16125));
   AOI21x1_ASAP7_75t_SL FE_RC_146_0 (.Y(n24827),
	.A1(n26818),
	.A2(n26819),
	.B(n26815));
   AOI21xp33_ASAP7_75t_SL FE_RC_145_0 (.Y(n16068),
	.A1(n27195),
	.A2(n16069),
	.B(ld));
   AOI21x1_ASAP7_75t_L FE_RC_144_0 (.Y(n26253),
	.A1(n26250),
	.A2(n26282),
	.B(n26251));
   AOI21xp5_ASAP7_75t_SL FE_RC_143_0 (.Y(n25168),
	.A1(n25164),
	.A2(n25682),
	.B(n25165));
   AOI21x1_ASAP7_75t_SL FE_RC_141_0 (.Y(n26508),
	.A1(n25860),
	.A2(n27216),
	.B(n25861));
   OR2x2_ASAP7_75t_SL FE_RC_139_0 (.Y(n25748),
	.A(n17982),
	.B(n17981));
   AOI21xp5_ASAP7_75t_L FE_RC_138_0 (.Y(n21997),
	.A1(n21995),
	.A2(n26407),
	.B(n21996));
   INVxp33_ASAP7_75t_L FE_RC_135_0 (.Y(FE_RN_4_0),
	.A(n22205));
   AOI31xp33_ASAP7_75t_SL FE_RC_133_0 (.Y(n23564),
	.A1(n23547),
	.A2(n23546),
	.A3(FE_OFN28648_n23549),
	.B(n23548));
   AOI21x1_ASAP7_75t_L FE_RC_132_0 (.Y(n26937),
	.A1(n27206),
	.A2(FE_OFN16177_n27207),
	.B(FE_OCPN29445_n27203));
   AOI21xp5_ASAP7_75t_L FE_RC_131_0 (.Y(n22713),
	.A1(n22711),
	.A2(n25575),
	.B(n22712));
   AOI21x1_ASAP7_75t_SL FE_RC_130_0 (.Y(n24816),
	.A1(n25455),
	.A2(n26139),
	.B(n25452));
   AOI21x1_ASAP7_75t_SL FE_RC_129_0 (.Y(n25144),
	.A1(n25038),
	.A2(n26819),
	.B(n25039));
   AOI21x1_ASAP7_75t_SL FE_RC_128_0 (.Y(n21007),
	.A1(n21005),
	.A2(n27183),
	.B(n21006));
   AOI21x1_ASAP7_75t_SL FE_RC_127_0 (.Y(n25827),
	.A1(n25824),
	.A2(n26407),
	.B(n25825));
   AOI21x1_ASAP7_75t_SL FE_RC_126_0 (.Y(n26704),
	.A1(n25680),
	.A2(n25682),
	.B(n25681));
   AOI21x1_ASAP7_75t_SL FE_RC_125_0 (.Y(n24382),
	.A1(n26583),
	.A2(FE_OFN16163_n26584),
	.B(FE_OFN29029_n26579));
   AOI31xp67_ASAP7_75t_SL FE_RC_123_0 (.Y(n21080),
	.A1(n21056),
	.A2(n23438),
	.A3(n21332),
	.B(n23467));
   AOI31xp33_ASAP7_75t_SL FE_RC_121_0 (.Y(n18660),
	.A1(FE_RN_3_0),
	.A2(n18658),
	.A3(n18744),
	.B(n26777));
   AOI31xp33_ASAP7_75t_SL FE_RC_120_0 (.Y(n25557),
	.A1(n17085),
	.A2(n17084),
	.A3(n19370),
	.B(n27102));
   AOI21xp5_ASAP7_75t_SL FE_RC_119_0 (.Y(n15762),
	.A1(n15736),
	.A2(n13867),
	.B(n15737));
   AOI31xp33_ASAP7_75t_SL FE_RC_118_0 (.Y(n24622),
	.A1(n18423),
	.A2(n18422),
	.A3(n18424),
	.B(n26542));
   AOI31xp33_ASAP7_75t_SL FE_RC_116_0 (.Y(n22712),
	.A1(n22702),
	.A2(n22701),
	.A3(n22703),
	.B(n25585));
   AOI31xp33_ASAP7_75t_L FE_RC_115_0 (.Y(n20121),
	.A1(n20120),
	.A2(n26347),
	.A3(n22395),
	.B(n23899));
   AOI21xp5_ASAP7_75t_SL FE_RC_113_0 (.Y(n18398),
	.A1(n18396),
	.A2(n26584),
	.B(n18397));
   AOI21xp5_ASAP7_75t_SL FE_RC_112_0 (.Y(n14320),
	.A1(n14318),
	.A2(n13867),
	.B(n14319));
   AOI31xp33_ASAP7_75t_L FE_RC_110_0 (.Y(n27019),
	.A1(FE_OFN28576_n27003),
	.A2(n27002),
	.A3(n27005),
	.B(n27004));
   AOI31xp67_ASAP7_75t_SL FE_RC_109_0 (.Y(n22961),
	.A1(n22941),
	.A2(n22940),
	.A3(n22942),
	.B(n26710));
   AOI31xp33_ASAP7_75t_SL FE_RC_108_0 (.Y(n25574),
	.A1(n19900),
	.A2(n19899),
	.A3(n19901),
	.B(n24263));
   AOI31xp33_ASAP7_75t_SL FE_RC_107_0 (.Y(n25215),
	.A1(n19283),
	.A2(n22559),
	.A3(n22077),
	.B(n27140));
   AOI31xp33_ASAP7_75t_SL FE_RC_104_0 (.Y(n22517),
	.A1(n22515),
	.A2(n22514),
	.A3(FE_OCPN29416_n22516),
	.B(n17463));
   AOI31xp33_ASAP7_75t_SL FE_RC_103_0 (.Y(n24740),
	.A1(n23154),
	.A2(n23153),
	.A3(n23155),
	.B(n24978));
   AOI31xp33_ASAP7_75t_SL FE_RC_102_0 (.Y(n20351),
	.A1(n20350),
	.A2(n20349),
	.A3(n24281),
	.B(n25585));
   AOI31xp33_ASAP7_75t_L FE_RC_100_0 (.Y(n24337),
	.A1(n16899),
	.A2(n16898),
	.A3(n18138),
	.B(n26542));
   AOI31xp33_ASAP7_75t_SL FE_RC_98_0 (.Y(n22477),
	.A1(n22446),
	.A2(n22445),
	.A3(n27017),
	.B(n26464));
   AOI21xp5_ASAP7_75t_SL FE_RC_97_0 (.Y(n20825),
	.A1(n20823),
	.A2(n20824),
	.B(n24377));
   AOI21xp5_ASAP7_75t_L FE_RC_96_0 (.Y(n22361),
	.A1(n22359),
	.A2(n25575),
	.B(n22360));
   AOI21xp5_ASAP7_75t_SL FE_RC_95_0 (.Y(n13929),
	.A1(n13927),
	.A2(n15757),
	.B(n13928));
   AOI21xp5_ASAP7_75t_L FE_RC_94_0 (.Y(n21759),
	.A1(n21757),
	.A2(n21758),
	.B(n23467));
   AOI31xp33_ASAP7_75t_L FE_RC_93_0 (.Y(n21996),
	.A1(n21985),
	.A2(n21984),
	.A3(n21986),
	.B(n27168));
   AOI31xp33_ASAP7_75t_SL FE_RC_92_0 (.Y(n18608),
	.A1(n18607),
	.A2(n21258),
	.A3(n21238),
	.B(n26517));
   AOI31xp33_ASAP7_75t_SL FE_RC_91_0 (.Y(n19958),
	.A1(n19957),
	.A2(n19956),
	.A3(n24852),
	.B(n17584));
   AOI31xp33_ASAP7_75t_SL FE_RC_90_0 (.Y(n19616),
	.A1(n19614),
	.A2(n19613),
	.A3(n19615),
	.B(n21493));
   AOI31xp33_ASAP7_75t_SL FE_RC_89_0 (.Y(n19027),
	.A1(n19026),
	.A2(n26549),
	.A3(n19010),
	.B(n26710));
   AOI31xp33_ASAP7_75t_SL FE_RC_86_0 (.Y(n21337),
	.A1(n21289),
	.A2(n21721),
	.A3(n24834),
	.B(n25420));
   AOI31xp67_ASAP7_75t_SL FE_RC_85_0 (.Y(n21079),
	.A1(n21064),
	.A2(n21063),
	.A3(n21065),
	.B(n23945));
   AOI21xp5_ASAP7_75t_SL FE_RC_84_0 (.Y(n14732),
	.A1(n15983),
	.A2(n14731),
	.B(n14730));
   AOI21xp5_ASAP7_75t_L FE_RC_83_0 (.Y(n22264),
	.A1(n22262),
	.A2(n25682),
	.B(n22263));
   AOI31xp33_ASAP7_75t_SL FE_RC_82_0 (.Y(n17733),
	.A1(n19697),
	.A2(n17710),
	.A3(n22378),
	.B(n23899));
   AOI31xp33_ASAP7_75t_SL FE_RC_81_0 (.Y(n17889),
	.A1(n17888),
	.A2(n17887),
	.A3(n22348),
	.B(n24263));
   AOI31xp33_ASAP7_75t_SL FE_RC_80_0 (.Y(n21863),
	.A1(n21862),
	.A2(n24571),
	.A3(n21857),
	.B(n26078));
   AOI31xp33_ASAP7_75t_SL FE_RC_78_0 (.Y(n21761),
	.A1(n21737),
	.A2(n21736),
	.A3(n24245),
	.B(n25420));
   AOI31xp33_ASAP7_75t_SL FE_RC_76_0 (.Y(n24796),
	.A1(n24794),
	.A2(n24793),
	.A3(n24795),
	.B(n26687));
   INVxp67_ASAP7_75t_SL FE_RC_73_0 (.Y(FE_RN_1_0),
	.A(n23770));
   AOI31xp33_ASAP7_75t_SL FE_RC_72_0 (.Y(n23785),
	.A1(FE_RN_1_0),
	.A2(n23771),
	.A3(n23872),
	.B(n25641));
   AOI31xp33_ASAP7_75t_SL FE_RC_71_0 (.Y(n15708),
	.A1(n15706),
	.A2(n12994),
	.A3(n15757),
	.B(n15707));
   AOI21xp5_ASAP7_75t_L FE_RC_70_0 (.Y(n13542),
	.A1(n13525),
	.A2(n13526),
	.B(n15238));
   AOI21xp5_ASAP7_75t_SL FE_RC_69_0 (.Y(n18801),
	.A1(n19712),
	.A2(FE_OFN69_sa32_4),
	.B(n18797));
   AOI21xp5_ASAP7_75t_SL FE_RC_68_0 (.Y(n18851),
	.A1(FE_OCPN28434_n17546),
	.A2(n18298),
	.B(n18323));
   AOI21xp5_ASAP7_75t_SL FE_RC_67_0 (.Y(n15707),
	.A1(n15703),
	.A2(n15705),
	.B(n15704));
   AOI31xp33_ASAP7_75t_SL FE_RC_66_0 (.Y(n16666),
	.A1(n16665),
	.A2(n23140),
	.A3(n23992),
	.B(n25139));
   AOI31xp33_ASAP7_75t_L FE_RC_65_0 (.Y(n18291),
	.A1(n18290),
	.A2(n20497),
	.A3(n25562),
	.B(n27095));
   AOI31xp33_ASAP7_75t_SL FE_RC_64_0 (.Y(n20179),
	.A1(n22065),
	.A2(n20177),
	.A3(n20178),
	.B(n27140));
   AOI31xp33_ASAP7_75t_SL FE_RC_63_0 (.Y(n15883),
	.A1(n15880),
	.A2(n15879),
	.A3(n15882),
	.B(n15881));
   AOI31xp33_ASAP7_75t_SL FE_RC_62_0 (.Y(n13363),
	.A1(n13357),
	.A2(n13356),
	.A3(n13358),
	.B(n15259));
   AOI31xp33_ASAP7_75t_SL FE_RC_60_0 (.Y(n14730),
	.A1(n14728),
	.A2(n14727),
	.A3(n14729),
	.B(n15969));
   AND2x2_ASAP7_75t_SL FE_RC_59_0 (.Y(n17530),
	.A(n19700),
	.B(n17713));
   AOI21xp5_ASAP7_75t_L FE_RC_58_0 (.Y(n15348),
	.A1(n15347),
	.A2(n15729),
	.B(n15346));
   AOI21xp5_ASAP7_75t_SL FE_RC_57_0 (.Y(n23341),
	.A1(FE_OCPN27721_n23336),
	.A2(FE_OFN25952_n22312),
	.B(n21121));
   AOI31xp33_ASAP7_75t_SL FE_RC_56_0 (.Y(n15137),
	.A1(n15090),
	.A2(n15089),
	.A3(n15091),
	.B(n15881));
   AOI31xp33_ASAP7_75t_SL FE_RC_55_0 (.Y(n14461),
	.A1(n14459),
	.A2(n14833),
	.A3(n14460),
	.B(n15888));
   AOI31xp33_ASAP7_75t_SL FE_RC_54_0 (.Y(n14956),
	.A1(n14953),
	.A2(n14952),
	.A3(n14954),
	.B(n16023));
   AOI31xp33_ASAP7_75t_SL FE_RC_53_0 (.Y(n13992),
	.A1(n13990),
	.A2(n13989),
	.A3(n13991),
	.B(n15969));
   AOI31xp33_ASAP7_75t_SL FE_RC_52_0 (.Y(n15437),
	.A1(n15431),
	.A2(n15430),
	.A3(n15432),
	.B(n16026));
   AOI31xp33_ASAP7_75t_SL FE_RC_51_0 (.Y(n25762),
	.A1(n17670),
	.A2(n17669),
	.A3(n24581),
	.B(n26926));
   AOI31xp33_ASAP7_75t_SL FE_RC_49_0 (.Y(n13467),
	.A1(n13445),
	.A2(n13444),
	.A3(n13446),
	.B(n13689));
   OR3x1_ASAP7_75t_L FE_RC_48_0 (.Y(n18434),
	.A(n16469),
	.B(n16852),
	.C(n16720));
   AOI21xp5_ASAP7_75t_SL FE_RC_47_0 (.Y(n23284),
	.A1(n21815),
	.A2(n19171),
	.B(n17500));
   AOI21xp5_ASAP7_75t_SL FE_RC_46_0 (.Y(n13693),
	.A1(n13688),
	.A2(n13690),
	.B(n13689));
   AOI31xp33_ASAP7_75t_L FE_RC_45_0 (.Y(n13928),
	.A1(n13913),
	.A2(n13912),
	.A3(n13914),
	.B(n15704));
   AOI31xp33_ASAP7_75t_L FE_RC_43_0 (.Y(n23310),
	.A1(FE_RN_0_0),
	.A2(FE_OFN26133_sa22_3),
	.A3(FE_PSN8315_FE_OFN16135_sa22_4),
	.B(n23309));
   AOI31xp33_ASAP7_75t_SL FE_RC_42_0 (.Y(n26945),
	.A1(n16352),
	.A2(n26296),
	.A3(n26294),
	.B(n26315));
   AOI31xp33_ASAP7_75t_L FE_RC_41_0 (.Y(n13789),
	.A1(n13787),
	.A2(n13786),
	.A3(n13788),
	.B(n15881));
   OR3x1_ASAP7_75t_R FE_RC_40_0 (.Y(n23145),
	.A(n23139),
	.B(n23138),
	.C(n23137));
   AOI21xp5_ASAP7_75t_SL FE_RC_39_0 (.Y(n23882),
	.A1(FE_OFN29081_n18526),
	.A2(FE_OFN29140_n18527),
	.B(n20624));
   AOI21xp33_ASAP7_75t_L FE_RC_38_0 (.Y(n14447),
	.A1(FE_OFN25900_w3_4),
	.A2(n14976),
	.B(n14446));
   AOI31xp33_ASAP7_75t_SL FE_RC_37_0 (.Y(n20791),
	.A1(FE_OFN26125_n22742),
	.A2(FE_OFN25907_sa12_2),
	.A3(FE_OCPN27804_sa12_1),
	.B(n22739));
   AOI31xp33_ASAP7_75t_SL FE_RC_36_0 (.Y(n14646),
	.A1(n14639),
	.A2(n14638),
	.A3(n14640),
	.B(n15969));
   AOI21xp33_ASAP7_75t_SRAM FE_RC_35_0 (.Y(n18824),
	.A1(n17525),
	.A2(n18799),
	.B(n18798));
   AOI21xp5_ASAP7_75t_L FE_RC_34_0 (.Y(n18302),
	.A1(FE_OCPN28229_n17529),
	.A2(FE_OCPN28434_n17546),
	.B(n24855));
   AOI31xp33_ASAP7_75t_SL FE_RC_33_0 (.Y(n21090),
	.A1(n18162),
	.A2(n18176),
	.A3(FE_OCPN27979_FE_OFN16147_sa22_1),
	.B(n22857));
   AOI31xp33_ASAP7_75t_SL FE_RC_32_0 (.Y(n20935),
	.A1(n18970),
	.A2(FE_OCPN27482_sa23_5),
	.A3(n20933),
	.B(n20932));
   AOI31xp33_ASAP7_75t_SL FE_RC_31_0 (.Y(n15218),
	.A1(n13596),
	.A2(FE_OFN26567_n),
	.A3(FE_OCPN27665_w3_25),
	.B(n13655));
   AOI31xp33_ASAP7_75t_L FE_RC_30_0 (.Y(n15321),
	.A1(n15528),
	.A2(FE_OFN26091_n24663),
	.A3(n15536),
	.B(n15320));
   AOI31xp33_ASAP7_75t_SL FE_RC_29_0 (.Y(n14947),
	.A1(FE_OFN28659_n15934),
	.A2(FE_OFN29125_n),
	.A3(FE_OCPN29535_FE_OFN8_w3_14),
	.B(n14946));
   OR2x2_ASAP7_75t_SL FE_RC_28_0 (.Y(n19552),
	.A(n20554),
	.B(n17970));
   AOI21xp5_ASAP7_75t_L FE_RC_27_0 (.Y(n19875),
	.A1(FE_OFN28529_n16774),
	.A2(FE_OFN28778_FE_OCPN28352_n16748),
	.B(n19874));
   AOI21xp5_ASAP7_75t_L FE_RC_26_0 (.Y(n17964),
	.A1(n23587),
	.A2(n24364),
	.B(n22750));
   AOI21xp33_ASAP7_75t_R FE_RC_25_0 (.Y(n25284),
	.A1(n19376),
	.A2(FE_OFN29234_n16996),
	.B(n17067));
   AOI21xp33_ASAP7_75t_SL FE_RC_24_0 (.Y(n15222),
	.A1(FE_OFN27211_w3_30),
	.A2(FE_OCPN27656_w3_25),
	.B(n14514));
   AOI21x1_ASAP7_75t_SL FE_RC_23_0 (.Y(n15492),
	.A1(FE_OFN26053_n25415),
	.A2(FE_OFN28551_FE_OFN26114_n),
	.B(n13869));
   AOI31xp33_ASAP7_75t_SRAM FE_RC_22_0 (.Y(n14444),
	.A1(n14442),
	.A2(n15835),
	.A3(n13771),
	.B(n14443));
   AOI31xp67_ASAP7_75t_L FE_RC_21_0 (.Y(n20469),
	.A1(n22125),
	.A2(FE_OCPN28378_n22632),
	.A3(n18463),
	.B(n22168));
   AOI31xp67_ASAP7_75t_SL FE_RC_20_0 (.Y(n22110),
	.A1(FE_OCPN29469_n17747),
	.A2(FE_OCPN27634_n20169),
	.A3(FE_OFN26159_n22080),
	.B(n20152));
   AOI21xp5_ASAP7_75t_L FE_RC_19_0 (.Y(n15487),
	.A1(FE_OFN26053_n25415),
	.A2(FE_OFN26045_n25377),
	.B(FE_OFN26091_n24663));
   AOI21xp33_ASAP7_75t_L FE_RC_18_0 (.Y(n20454),
	.A1(FE_OFN28610_n22125),
	.A2(n25108),
	.B(n18362));
   AOI21xp5_ASAP7_75t_SL FE_RC_17_0 (.Y(n15609),
	.A1(n15817),
	.A2(FE_OFN28671_FE_OCPN28076),
	.B(n15808));
   AOI21xp5_ASAP7_75t_SL FE_RC_16_0 (.Y(n15586),
	.A1(n15842),
	.A2(n13739),
	.B(n15858));
   AOI31xp33_ASAP7_75t_SL FE_RC_15_0 (.Y(n21183),
	.A1(FE_OFN28835_n),
	.A2(n17254),
	.A3(FE_OCPN27908_FE_OFN16156_sa00_2),
	.B(n18656));
   AOI31xp33_ASAP7_75t_SL FE_RC_14_0 (.Y(n20924),
	.A1(FE_OCPN27986_n18970),
	.A2(FE_OFN28580_n23491),
	.A3(FE_OCPN29374_FE_OFN29191_sa23_2),
	.B(n20903));
   AOI31xp67_ASAP7_75t_L FE_RC_13_0 (.Y(n15216),
	.A1(FE_OCPN27655_w3_25),
	.A2(FE_OFN26049_w3_27),
	.A3(FE_OFN27212_w3_30),
	.B(n13636));
   AOI31xp33_ASAP7_75t_R FE_RC_12_0 (.Y(n20499),
	.A1(n16975),
	.A2(n16980),
	.A3(FE_OFN28979_n),
	.B(n18921));
   AOI31xp33_ASAP7_75t_SL FE_RC_11_0 (.Y(n19176),
	.A1(n19171),
	.A2(FE_OCPN28321_n21341),
	.A3(FE_OFN94_sa11_5),
	.B(n22497));
   AOI31xp33_ASAP7_75t_SL FE_RC_10_0 (.Y(n21667),
	.A1(n18529),
	.A2(n18583),
	.A3(FE_OFN29131_FE_OCPN27371_sa20_2),
	.B(n18603));
   AOI21xp5_ASAP7_75t_SL FE_RC_8_0 (.Y(n18214),
	.A1(FE_OFN26141_n23307),
	.A2(n23336),
	.B(n20726));
   AOI21x1_ASAP7_75t_L FE_RC_7_0 (.Y(n22507),
	.A1(FE_OCPN29435_n17445),
	.A2(FE_OCPN5021_n17446),
	.B(n21822));
   AOI31xp33_ASAP7_75t_L FE_RC_6_0 (.Y(n23800),
	.A1(n21195),
	.A2(n20617),
	.A3(FE_OCPN28163_FE_OFN99_sa20_5),
	.B(n21648));
   AOI31xp33_ASAP7_75t_R FE_RC_5_0 (.Y(n13503),
	.A1(n13596),
	.A2(FE_OFN16437_n),
	.A3(n15145),
	.B(n15189));
   AOI21x1_ASAP7_75t_SL FE_RC_4_0 (.Y(n13766),
	.A1(FE_OCPN27978_w3_3),
	.A2(FE_OFN26057_w3_1),
	.B(n15862));
   AOI21xp33_ASAP7_75t_L FE_RC_3_0 (.Y(n15189),
	.A1(FE_OCPN27655_w3_25),
	.A2(FE_OCPN8232_FE_OFN27206_w3_30),
	.B(n14535));
   INVx4_ASAP7_75t_SL FE_OFC3557_n16100 (.Y(n16099),
	.A(FE_OFN26541_n16100));
   INVx2_ASAP7_75t_SL FE_OFC3556_n16100 (.Y(FE_OFN26541_n16100),
	.A(n16100));
   INVx1_ASAP7_75t_SL FE_OFC3549_n15770 (.Y(n15771),
	.A(FE_OFN25891_n15770));
   INVx2_ASAP7_75t_SL FE_OFC3548_n15770 (.Y(FE_OFN25891_n15770),
	.A(n15770));
   INVx1_ASAP7_75t_L FE_OFC3547_n16189 (.Y(FE_OFN26630_n16190),
	.A(n16189));
   INVx1_ASAP7_75t_SL FE_OFC3545_n16247 (.Y(n16244),
	.A(n16247));
   INVx4_ASAP7_75t_SL FE_OFC3525_w3_17 (.Y(FE_OFN27214_w3_17),
	.A(FE_OFN26041_w3_17));
   INVx1_ASAP7_75t_R FE_OFC3523_w3_17 (.Y(n25377),
	.A(FE_OFN28674_n));
   INVx3_ASAP7_75t_SL FE_OFC3522_w3_17 (.Y(FE_OFN26041_w3_17),
	.A(w3_17_));
   INVx1_ASAP7_75t_SL FE_OFC3508_n16052 (.Y(FE_OFN16262_n16052),
	.A(n16053));
   INVx2_ASAP7_75t_SL FE_OFC3507_n16052 (.Y(n16053),
	.A(n16052));
   HB1xp67_ASAP7_75t_SL FE_OFC3506_w3_30 (.Y(FE_OFN27212_w3_30),
	.A(FE_OFN27208_w3_30));
   INVx3_ASAP7_75t_SL FE_OFC3505_w3_30 (.Y(FE_OFN27211_w3_30),
	.A(FE_OFN27207_w3_30));
   INVx3_ASAP7_75t_SL FE_OFC3504_w3_30 (.Y(FE_OFN27210_w3_30),
	.A(FE_OFN27207_w3_30));
   INVx1_ASAP7_75t_L FE_OFC3502_w3_30 (.Y(FE_OFN27208_w3_30),
	.A(FE_OFN26076_w3_30));
   BUFx5_ASAP7_75t_SL FE_OFC3501_w3_30 (.Y(FE_OFN27207_w3_30),
	.A(n24688));
   INVx2_ASAP7_75t_SL FE_OFC3500_w3_30 (.Y(FE_OFN27206_w3_30),
	.A(n24688));
   INVxp67_ASAP7_75t_SL FE_OFC3497_w3_30 (.Y(FE_OFN26076_w3_30),
	.A(n24688));
   INVx2_ASAP7_75t_SL FE_OFC3496_w3_30 (.Y(n24688),
	.A(w3_30_));
   INVx2_ASAP7_75t_L FE_OFC3492_w3_27 (.Y(FE_OFN26051_w3_27),
	.A(n25675));
   BUFx4f_ASAP7_75t_SL FE_OFC3491_w3_27 (.Y(FE_OFN26049_w3_27),
	.A(n25675));
   INVx1_ASAP7_75t_L FE_OFC3490_w3_27 (.Y(FE_OFN26048_w3_27),
	.A(n25675));
   BUFx6f_ASAP7_75t_SL FE_OFC3489_w3_27 (.Y(n25675),
	.A(w3_27_));
   BUFx5_ASAP7_75t_SL FE_OFC3488_n16749 (.Y(FE_OFN16447_n16749),
	.A(n16749));
   BUFx2_ASAP7_75t_SL FE_OFC3486_w3_20 (.Y(FE_OFN16426_w3_20),
	.A(w3_20_));
   INVx2_ASAP7_75t_SL FE_OFC3485_w3_20 (.Y(FE_OFN25909_w3_20),
	.A(w3_20_));
   BUFx6f_ASAP7_75t_SL FE_OFC3481_w3_22 (.Y(FE_OFN4_w3_22),
	.A(w3_22_));
   INVx3_ASAP7_75t_L FE_OFC3452_n16447 (.Y(FE_OFN26545_n16447),
	.A(n16946));
   BUFx3_ASAP7_75t_SL FE_OFC3451_n16447 (.Y(n16946),
	.A(n16447));
   BUFx2_ASAP7_75t_L FE_OFC3435_n23315 (.Y(FE_OFN27173_n),
	.A(n23315));
   INVxp33_ASAP7_75t_L FE_OFC3434_n23315 (.Y(FE_OFN16450_n23315),
	.A(n23315));
   INVxp67_ASAP7_75t_R FE_OFC3433_n20209 (.Y(FE_OFN41_n20971),
	.A(n20209));
   INVxp33_ASAP7_75t_R FE_OFC3431_n17441 (.Y(FE_OFN27172_n17441),
	.A(n24310));
   INVx1_ASAP7_75t_SL FE_OFC3420_n24006 (.Y(n24007),
	.A(n24006));
   INVx2_ASAP7_75t_SL FE_OFC3419_n26683 (.Y(FE_OFN27169_n26683),
	.A(n26683));
   INVx1_ASAP7_75t_L FE_OFC3416_n16334 (.Y(n16361),
	.A(n16334));
   INVx2_ASAP7_75t_SL FE_OFC3411_n17995 (.Y(n18034),
	.A(n17995));
   INVx2_ASAP7_75t_L FE_OFC3406_n18710 (.Y(n17386),
	.A(FE_OCPN29406_n18710));
   INVxp67_ASAP7_75t_L FE_OFC3400_n22136 (.Y(FE_OFN26037_n22144),
	.A(n22136));
   INVx2_ASAP7_75t_SL FE_OFC3397_n15714 (.Y(FE_OFN25915_n15514),
	.A(n15714));
   INVx2_ASAP7_75t_SL FE_OFC3391_n20304 (.Y(n22353),
	.A(n20304));
   INVx3_ASAP7_75t_SL FE_OFC3380_n23928 (.Y(FE_OFN27157_n23928),
	.A(n23633));
   HB1xp67_ASAP7_75t_L FE_OFC3374_w3_6 (.Y(FE_OFN27156_n),
	.A(FE_OFN28695_n));
   BUFx3_ASAP7_75t_SL FE_OFC3373_w3_6 (.Y(FE_OFN26531_n),
	.A(FE_OFN28699_w3_6));
   INVx2_ASAP7_75t_SL FE_OFC3357_n17315 (.Y(FE_OFN25950_sa01_2),
	.A(FE_OFN28672_sa01_2));
   INVxp33_ASAP7_75t_R FE_OFC3354_n16837 (.Y(n16691),
	.A(n16837));
   INVx1_ASAP7_75t_L FE_OFC3348_n22175 (.Y(n22189),
	.A(n22175));
   INVxp67_ASAP7_75t_R FE_OFC3347_n18789 (.Y(n18790),
	.A(n18789));
   INVx2_ASAP7_75t_SL FE_OFC3330_n25934 (.Y(n25935),
	.A(n25934));
   INVxp67_ASAP7_75t_L FE_OFC3322_n24012 (.Y(n24995),
	.A(n24012));
   INVxp67_ASAP7_75t_L FE_OFC3319_n15385 (.Y(n14939),
	.A(n15385));
   INVxp67_ASAP7_75t_R FE_OFC3317_n15992 (.Y(FE_OFN27136_n15992),
	.A(n15992));
   INVx2_ASAP7_75t_SL FE_OFC3316_n15992 (.Y(FE_OFN27135_n15992),
	.A(n15992));
   INVx1_ASAP7_75t_R FE_OFC3297_n19552 (.Y(FE_OFN26023_n20807),
	.A(n19552));
   BUFx3_ASAP7_75t_SL FE_OFC3294_n25869 (.Y(FE_OFN16162_n25869),
	.A(n25869));
   BUFx2_ASAP7_75t_SL FE_OFC3293_n13876 (.Y(FE_OFN16210_n13876),
	.A(n13876));
   INVx1_ASAP7_75t_SL FE_OFC3270_n23101 (.Y(FE_OFN16208_n23101),
	.A(n23107));
   BUFx3_ASAP7_75t_SL FE_OFC3269_n23101 (.Y(n23107),
	.A(n23101));
   BUFx12f_ASAP7_75t_SL FE_OFC3266_n21057 (.Y(FE_OFN21730_sa03_3),
	.A(sa03_3_));
   INVxp33_ASAP7_75t_R FE_OFC3258_n14663 (.Y(FE_OFN16274_n14664),
	.A(FE_OFN16273_n14664));
   INVx2_ASAP7_75t_L FE_OFC3253_n26971 (.Y(FE_OFN108_n26971),
	.A(FE_OCPN27624_n26971));
   BUFx2_ASAP7_75t_SL FE_OFC3241_w3_1 (.Y(FE_OFN27124_w3_1),
	.A(n24831));
   INVx2_ASAP7_75t_SL FE_OFC3240_w3_1 (.Y(FE_OFN26058_w3_1),
	.A(n24831));
   BUFx2_ASAP7_75t_L FE_OFC3239_w3_1 (.Y(FE_OFN26057_w3_1),
	.A(n24831));
   BUFx6f_ASAP7_75t_SL FE_OFC3238_w3_1 (.Y(n24831),
	.A(w3_1_));
   BUFx2_ASAP7_75t_SL FE_OFC3215_sa22_3 (.Y(n23308),
	.A(sa22_3_));
   BUFx3_ASAP7_75t_SL FE_OFC3214_sa22_3 (.Y(FE_OFN26136_sa22_3),
	.A(sa22_3_));
   INVx1_ASAP7_75t_SL FE_OFC3213_sa22_3 (.Y(FE_OFN26133_sa22_3),
	.A(sa22_3_));
   INVx2_ASAP7_75t_SL FE_OFC3209_n17329 (.Y(FE_OFN25878_n17329),
	.A(n17329));
   INVxp67_ASAP7_75t_R FE_OFC3202_n15197 (.Y(FE_OFN16201_n15197),
	.A(n15197));
   HB1xp67_ASAP7_75t_R FE_OFC3190_n (.Y(FE_OFN27111_n),
	.A(FE_OFN16459_n));
   INVxp67_ASAP7_75t_R FE_OFC3169_n24956 (.Y(n24960),
	.A(n24956));
   INVxp33_ASAP7_75t_L FE_OFC3165_n17265 (.Y(n17266),
	.A(n17265));
   INVx1_ASAP7_75t_L FE_OFC3160_n20305 (.Y(n20307),
	.A(n20305));
   INVxp67_ASAP7_75t_L FE_OFC3159_n22660 (.Y(n17847),
	.A(n22660));
   INVxp67_ASAP7_75t_L FE_OFC3158_n23558 (.Y(FE_OFN27090_n23558),
	.A(FE_OFN27089_n23558));
   INVx1_ASAP7_75t_R FE_OFC3154_n22808 (.Y(FE_OFN16304_n22808),
	.A(n23182));
   INVx1_ASAP7_75t_SL FE_OFC3153_n22808 (.Y(n23182),
	.A(n22808));
   INVx1_ASAP7_75t_SRAM FE_OFC3152_n23754 (.Y(FE_OFN27088_n23754),
	.A(n23754));
   INVxp67_ASAP7_75t_L FE_OFC3143_n23774 (.Y(FE_OFN27083_n),
	.A(n20670));
   BUFx2_ASAP7_75t_SL FE_OFC3141_n25377 (.Y(FE_OFN27082_n25377),
	.A(FE_OFN28706_n));
   INVxp33_ASAP7_75t_R FE_OFC3128_n23409 (.Y(FE_OFN27075_n23409),
	.A(n25606));
   BUFx2_ASAP7_75t_L FE_OFC3126_n13868 (.Y(FE_OFN27074_n13868),
	.A(n13868));
   INVx1_ASAP7_75t_SL FE_OFC3125_n13868 (.Y(FE_OFN25981_n13868),
	.A(n13868));
   INVx2_ASAP7_75t_L FE_OFC3116_n20866 (.Y(FE_OFN26570_n20866),
	.A(FE_OFN26569_n20866));
   INVx4_ASAP7_75t_SL FE_OFC3106_n13869 (.Y(FE_OFN27066_n13869),
	.A(n15480));
   BUFx3_ASAP7_75t_SL FE_OFC3105_n13869 (.Y(n15480),
	.A(n13869));
   INVx2_ASAP7_75t_SL FE_OFC3103_n17059 (.Y(n25545),
	.A(n17059));
   INVxp67_ASAP7_75t_L FE_OFC3102_n17203 (.Y(n17205),
	.A(n17203));
   INVx1_ASAP7_75t_SL FE_OFC3079_n13662 (.Y(FE_OFN27057_n13662),
	.A(n13662));
   INVx2_ASAP7_75t_L FE_OFC3071_n15034 (.Y(FE_OFN26532_n13766),
	.A(n15034));
   INVxp67_ASAP7_75t_L FE_OFC3065_n13648 (.Y(n13500),
	.A(n13648));
   INVx1_ASAP7_75t_L FE_OFC3053_n22765 (.Y(n22767),
	.A(n22765));
   INVxp33_ASAP7_75t_R FE_OFC3052_n20170 (.Y(FE_OFN152_n20170),
	.A(n20170));
   INVx1_ASAP7_75t_L FE_OFC3051_n24340 (.Y(n24341),
	.A(n24340));
   INVxp33_ASAP7_75t_L FE_OFC3048_n16469 (.Y(n16470),
	.A(n16469));
   INVxp67_ASAP7_75t_L FE_OFC3047_n17833 (.Y(n20323),
	.A(n17833));
   BUFx2_ASAP7_75t_SL FE_OFC3034_n15236 (.Y(n13596),
	.A(n15236));
   INVx1_ASAP7_75t_SL FE_OFC3030_n15862 (.Y(n13736),
	.A(n15862));
   INVx1_ASAP7_75t_SL FE_OFC3029_n13534 (.Y(n13386),
	.A(n13534));
   INVxp67_ASAP7_75t_L FE_OFC3018_n24378 (.Y(FE_OFN26140_n23585),
	.A(n24378));
   INVx2_ASAP7_75t_L FE_OFC3014_n19573 (.Y(FE_OFN16216_n19573),
	.A(FE_OCPN28250_n19573));
   INVx2_ASAP7_75t_L FE_OFC3012_n27164 (.Y(FE_OFN26650_n27164),
	.A(n27163));
   BUFx3_ASAP7_75t_SL FE_OFC3011_n27164 (.Y(n27163),
	.A(n27164));
   INVxp67_ASAP7_75t_R FE_OFC2997_n18263 (.Y(n18264),
	.A(n18263));
   INVxp67_ASAP7_75t_R FE_OFC2996_w3_15 (.Y(FE_OFN26129_w3_15),
	.A(FE_OCPN29427_w3_15));
   INVxp33_ASAP7_75t_R FE_OFC2993_n15665 (.Y(n13882),
	.A(n15665));
   INVxp67_ASAP7_75t_R FE_OFC2990_n25905 (.Y(FE_OFN16301_n25905),
	.A(FE_OCPN28366_n25329));
   INVx1_ASAP7_75t_SL FE_OFC2989_n25905 (.Y(n25329),
	.A(n25905));
   INVx1_ASAP7_75t_L FE_OFC2987_n16159 (.Y(FE_OFN26646_n16159),
	.A(FE_OFN16251_n16162));
   INVx2_ASAP7_75t_SL FE_OFC2986_n16159 (.Y(FE_OFN16251_n16162),
	.A(n16159));
   HB1xp67_ASAP7_75t_SL FE_OFC2984_w3_6 (.Y(FE_OFN26645_n),
	.A(FE_OFN28699_w3_6));
   INVx2_ASAP7_75t_L FE_OFC2975_n15200 (.Y(FE_OFN16193_n15200),
	.A(n15200));
   INVxp33_ASAP7_75t_R FE_OFC2964_w3_14 (.Y(FE_OFN26634_w3_14),
	.A(FE_OFN26637_w3_14));
   INVx2_ASAP7_75t_SL FE_OFC2956_w3_14 (.Y(FE_OFN8_w3_14),
	.A(w3_14_));
   INVx2_ASAP7_75t_SL FE_OFC2947_w3_9 (.Y(FE_OFN16184_w3_9),
	.A(FE_OFN16182_w3_9));
   INVx2_ASAP7_75t_SL FE_OFC2941_n26088 (.Y(FE_OFN25973_n26087),
	.A(n26088));
   BUFx3_ASAP7_75t_SL FE_OFC2927_n16575 (.Y(n23980),
	.A(n16575));
   INVx1_ASAP7_75t_SL FE_OFC2926_n16575 (.Y(FE_OFN25956_n16575),
	.A(n16575));
   INVxp67_ASAP7_75t_R FE_OFC2920_n25782 (.Y(FE_OFN26163_w3_13),
	.A(FE_OFN26162_w3_13));
   INVx1_ASAP7_75t_L FE_OFC2919_n25782 (.Y(FE_OFN26162_w3_13),
	.A(n25782));
   INVx2_ASAP7_75t_L FE_OFC2902_n26478 (.Y(n26742),
	.A(FE_OCPN29274_n26478));
   INVx2_ASAP7_75t_SL FE_OFC2899_n24537 (.Y(FE_OFN26546_n24537),
	.A(n24537));
   INVx1_ASAP7_75t_SL FE_OFC2898_n26491 (.Y(FE_OFN25911_n26491),
	.A(FE_OCPN28307_n26491));
   BUFx3_ASAP7_75t_SL FE_OFC2895_n23837 (.Y(n23677),
	.A(n23837));
   INVxp33_ASAP7_75t_R FE_OFC2890_n24644 (.Y(FE_OFN26553_n24644),
	.A(n17560));
   BUFx5_ASAP7_75t_SL FE_OFC2889_n24644 (.Y(n17560),
	.A(n24644));
   INVx1_ASAP7_75t_SL FE_OFC2877_n21253 (.Y(FE_OFN26150_n21253),
	.A(n18570));
   INVx2_ASAP7_75t_SL FE_OFC2869_sa31_4 (.Y(FE_OFN26629_sa31_4),
	.A(FE_OFN26595_sa31_4));
   INVx1_ASAP7_75t_SL FE_OFC2865_sa31_4 (.Y(FE_OFN26060_sa31_4),
	.A(FE_OFN26595_sa31_4));
   BUFx3_ASAP7_75t_L FE_OFC2839_n16010 (.Y(FE_OFN26007_n16010),
	.A(n16010));
   INVxp67_ASAP7_75t_L FE_OFC2838_n16010 (.Y(n14919),
	.A(n16010));
   INVx2_ASAP7_75t_SL FE_OFC2823_n26527 (.Y(FE_OFN25927_n26527),
	.A(FE_OFN16265_n26527));
   BUFx3_ASAP7_75t_SL FE_OFC2821_n26527 (.Y(FE_OFN16265_n26527),
	.A(n26527));
   HB1xp67_ASAP7_75t_R FE_OFC2798_w3_20 (.Y(FE_OFN26614_n),
	.A(FE_OFN16426_w3_20));
   INVx2_ASAP7_75t_SL FE_OFC2764_n23011 (.Y(FE_OFN25959_n23011),
	.A(sa10_5_));
   INVx1_ASAP7_75t_L FE_OFC2763_n13602 (.Y(n13605),
	.A(n13602));
   INVx1_ASAP7_75t_L FE_OFC2758_n24458 (.Y(n23149),
	.A(n24458));
   INVxp33_ASAP7_75t_R FE_OFC2744_n23913 (.Y(FE_OFN26578_n23913),
	.A(FE_OCPN28089_n23913));
   INVx1_ASAP7_75t_R FE_OFC2737_n21224 (.Y(n21240),
	.A(n21224));
   INVx1_ASAP7_75t_L FE_OFC2723_n19405 (.Y(FE_OFN26572_n19405),
	.A(n19405));
   INVx1_ASAP7_75t_SL FE_OFC2717_n20866 (.Y(FE_OFN26569_n20866),
	.A(n20866));
   INVx2_ASAP7_75t_SL FE_OFC2708_n13646 (.Y(FE_OFN25966_n13646),
	.A(n15203));
   INVx2_ASAP7_75t_SL FE_OFC2707_n13646 (.Y(n15203),
	.A(n13646));
   HB1xp67_ASAP7_75t_SL FE_OFC2705_n15195 (.Y(FE_OFN26567_n),
	.A(FE_OFN25875_n15227));
   INVx1_ASAP7_75t_SL FE_OFC2704_n15195 (.Y(FE_OFN16225_n15195),
	.A(FE_OFN25875_n15227));
   INVx2_ASAP7_75t_L FE_OFC2703_n15195 (.Y(FE_OFN25875_n15227),
	.A(n15195));
   INVxp67_ASAP7_75t_R FE_OFC2696_n19229 (.Y(n19231),
	.A(n19229));
   INVxp33_ASAP7_75t_R FE_OFC2685_n26754 (.Y(FE_OFN26559_n26754),
	.A(FE_OCPN29356_n27110));
   INVxp33_ASAP7_75t_L FE_OFC2678_n20546 (.Y(n20547),
	.A(n20546));
   INVx1_ASAP7_75t_SL FE_OFC2665_n14545 (.Y(FE_OFN26552_n14545),
	.A(n13556));
   INVx2_ASAP7_75t_SL FE_OFC2664_n14545 (.Y(n13556),
	.A(n14545));
   INVxp67_ASAP7_75t_L FE_OFC2659_n20666 (.Y(n20669),
	.A(n20666));
   INVxp67_ASAP7_75t_SL FE_OFC2658_n24174 (.Y(n24173),
	.A(n24174));
   INVxp33_ASAP7_75t_L FE_OFC2619_n17964 (.Y(n17936),
	.A(n17964));
   BUFx3_ASAP7_75t_SL FE_OFC2614_n13766 (.Y(n15034),
	.A(n13766));
   INVx4_ASAP7_75t_SL FE_OFC2600_n21511 (.Y(n21708),
	.A(n21511));
   INVxp33_ASAP7_75t_R FE_OFC2584_w3_13 (.Y(FE_OFN26164_w3_13),
	.A(FE_OFN26163_w3_13));
   INVx2_ASAP7_75t_SL FE_OFC2581_w3_13 (.Y(n25782),
	.A(w3_13_));
   INVx1_ASAP7_75t_R FE_OFC2571_n23812 (.Y(n23815),
	.A(n23812));
   INVxp67_ASAP7_75t_SL FE_OFC2565_sa12_2 (.Y(FE_OFN25906_sa12_2),
	.A(sa12_2_));
   BUFx3_ASAP7_75t_SL FE_OFC2564_sa12_2 (.Y(FE_OFN25908_sa12_2),
	.A(FE_OCPN27888_sa12_2));
   BUFx6f_ASAP7_75t_SL FE_OFC2530_n18774 (.Y(n19817),
	.A(n18774));
   INVx1_ASAP7_75t_L FE_OFC2522_n14924 (.Y(n15921),
	.A(n14924));
   INVx1_ASAP7_75t_SL FE_OFC2513_n23585 (.Y(n24378),
	.A(n23585));
   INVx1_ASAP7_75t_L FE_OFC2487_n17802 (.Y(FE_OFN26033_n20197),
	.A(n17802));
   BUFx2_ASAP7_75t_L FE_OFC2483_n22742 (.Y(FE_OFN26125_n22742),
	.A(n22742));
   INVx3_ASAP7_75t_SL FE_OFC2482_n22742 (.Y(n23217),
	.A(n22742));
   INVxp33_ASAP7_75t_L FE_OFC2472_n20440 (.Y(n20441),
	.A(n20440));
   INVxp67_ASAP7_75t_R FE_OFC2471_n20985 (.Y(n20986),
	.A(n20985));
   INVxp67_ASAP7_75t_L FE_OFC2455_n25787 (.Y(n21360),
	.A(n25787));
   INVx2_ASAP7_75t_SL FE_OFC2445_n26087 (.Y(n26088),
	.A(n26087));
   INVxp33_ASAP7_75t_L FE_OFC2444_n15275 (.Y(n15277),
	.A(n15275));
   INVx1_ASAP7_75t_L FE_OFC2436_n26502 (.Y(n27147),
	.A(FE_OCPN29397_n26502));
   INVx2_ASAP7_75t_L FE_OFC2424_n13876 (.Y(n15683),
	.A(n13876));
   BUFx4f_ASAP7_75t_SL FE_OFC2422_n22133 (.Y(FE_OFN25901_n22133),
	.A(n22133));
   INVxp33_ASAP7_75t_R FE_OFC2407_sa13_1 (.Y(FE_OFN16445_sa13_1),
	.A(FE_OFN26061_n));
   INVx1_ASAP7_75t_SL FE_OFC2402_n27123 (.Y(FE_OFN25963_n27123),
	.A(n27123));
   INVxp33_ASAP7_75t_L FE_OFC2401_n26316 (.Y(FE_OFN26019_n26319),
	.A(n26319));
   INVx1_ASAP7_75t_SL FE_OFC2380_n26788 (.Y(n26789),
	.A(n26788));
   BUFx2_ASAP7_75t_SL FE_OFC2379_n26788 (.Y(FE_OFN16283_n26788),
	.A(n26788));
   INVx1_ASAP7_75t_SL FE_OFC2358_n13288 (.Y(n15182),
	.A(n13288));
   INVxp67_ASAP7_75t_L FE_OFC2354_n15848 (.Y(FE_OFN26110_n15848),
	.A(FE_OFN25912_n15848));
   INVx2_ASAP7_75t_SL FE_OFC2353_n15848 (.Y(FE_OFN25912_n15848),
	.A(n15639));
   BUFx2_ASAP7_75t_SL FE_OFC2352_n15848 (.Y(n15639),
	.A(n15848));
   INVxp33_ASAP7_75t_L FE_OFC2349_w3_1 (.Y(FE_OFN16423_n24831),
	.A(FE_OFN26058_w3_1));
   INVx1_ASAP7_75t_L FE_OFC2344_n18213 (.Y(FE_OFN26009_n18213),
	.A(n18213));
   INVx2_ASAP7_75t_SL FE_OFC2324_n15257 (.Y(n15155),
	.A(n15257));
   BUFx3_ASAP7_75t_SL FE_OFC2322_n13659 (.Y(n14593),
	.A(n13659));
   INVx1_ASAP7_75t_SL FE_OFC2310_w3_9 (.Y(FE_OFN16182_w3_9),
	.A(w3_9_));
   INVxp67_ASAP7_75t_L FE_OFC2304_w3_20 (.Y(FE_OFN26072_n26720),
	.A(FE_OFN25909_w3_20));
   INVx1_ASAP7_75t_SL FE_OFC2295_n24803 (.Y(FE_OFN16297_n24803),
	.A(n24803));
   INVx1_ASAP7_75t_SL FE_OFC2288_n26602 (.Y(n26601),
	.A(FE_OCPN29335_n));
   INVxp67_ASAP7_75t_L FE_OFC2287_n26602 (.Y(FE_OFN16227_n26602),
	.A(FE_OCPN27419_n26602));
   HB1xp67_ASAP7_75t_SL FE_OFC2255_w3_4 (.Y(FE_OFN26073_n),
	.A(FE_OFN25900_w3_4));
   BUFx3_ASAP7_75t_SL FE_OFC2236_sa01_3 (.Y(FE_OFN26054_sa01_3),
	.A(sa01_3_));
   INVxp33_ASAP7_75t_L FE_OFC2218_n19464 (.Y(n19473),
	.A(n19464));
   INVxp67_ASAP7_75t_SL FE_OFC2217_n24887 (.Y(FE_OFN26038_n24887),
	.A(n24887));
   INVx1_ASAP7_75t_L FE_OFC2213_n22144 (.Y(n22136),
	.A(n22144));
   INVx1_ASAP7_75t_L FE_OFC2204_n20197 (.Y(n17802),
	.A(n20197));
   INVx1_ASAP7_75t_SL FE_OFC2203_n20230 (.Y(FE_OFN26032_n20230),
	.A(n20230));
   INVxp33_ASAP7_75t_L FE_OFC2200_n18472 (.Y(n17604),
	.A(n18472));
   INVxp67_ASAP7_75t_SL FE_OFC2193_n26903 (.Y(n26901),
	.A(n26903));
   INVxp67_ASAP7_75t_L FE_OFC2192_n24206 (.Y(n24207),
	.A(n24206));
   INVxp33_ASAP7_75t_R FE_OFC2189_n25368 (.Y(FE_OFN26030_n25368),
	.A(n25369));
   INVxp67_ASAP7_75t_L FE_OFC2187_n25368 (.Y(n25369),
	.A(n25368));
   INVxp67_ASAP7_75t_SL FE_OFC2183_n24034 (.Y(n24033),
	.A(n24034));
   INVx4_ASAP7_75t_SL FE_OFC2182_n23306 (.Y(n18162),
	.A(FE_OCPN29478_n23306));
   INVxp67_ASAP7_75t_SL FE_OFC2178_n17971 (.Y(n17972),
	.A(FE_OCPN28248_n17971));
   INVxp67_ASAP7_75t_L FE_OFC2177_n20646 (.Y(n18538),
	.A(n20646));
   INVx1_ASAP7_75t_SL FE_OFC2163_n16253 (.Y(FE_OFN26021_n16253),
	.A(n16253));
   INVxp33_ASAP7_75t_R FE_OFC2161_n18418 (.Y(n24484),
	.A(FE_OFN16218_n18418));
   INVx1_ASAP7_75t_SL FE_OFC2160_n18418 (.Y(FE_OFN16218_n18418),
	.A(n18418));
   INVxp33_ASAP7_75t_L FE_OFC2157_n25582 (.Y(n25583),
	.A(n25582));
   INVxp33_ASAP7_75t_SRAM FE_OFC2152_n16237 (.Y(n16139),
	.A(n16237));
   INVxp33_ASAP7_75t_L FE_OFC2151_n24268 (.Y(FE_OFN168_n24268),
	.A(n24268));
   INVx1_ASAP7_75t_SL FE_OFC2136_n27208 (.Y(FE_OFN26012_n27208),
	.A(n27208));
   INVxp67_ASAP7_75t_R FE_OFC2135_n27208 (.Y(n25311),
	.A(n27208));
   INVx1_ASAP7_75t_L FE_OFC2133_n20971 (.Y(n20209),
	.A(n20971));
   INVx1_ASAP7_75t_SL FE_OFC2131_n24953 (.Y(n21881),
	.A(n24953));
   INVxp33_ASAP7_75t_R FE_OFC2126_n24733 (.Y(n23122),
	.A(n24733));
   INVxp67_ASAP7_75t_L FE_OFC2119_n25612 (.Y(n25611),
	.A(n25612));
   INVx1_ASAP7_75t_SL FE_OFC2118_n25001 (.Y(n24999),
	.A(n25001));
   INVxp67_ASAP7_75t_R FE_OFC2114_n15992 (.Y(FE_OFN26003_n15992),
	.A(FE_OFN27136_n15992));
   INVxp67_ASAP7_75t_L FE_OFC2108_n19067 (.Y(n17665),
	.A(n19067));
   INVxp67_ASAP7_75t_R FE_OFC2095_n22122 (.Y(n22126),
	.A(n22122));
   INVxp67_ASAP7_75t_SL FE_OFC2094_n24743 (.Y(n24744),
	.A(n24743));
   INVx1_ASAP7_75t_L FE_OFC2092_sa32_7 (.Y(n17732),
	.A(FE_OFN136_sa32_7));
   INVxp67_ASAP7_75t_L FE_OFC2091_n26006 (.Y(FE_OFN25996_n26006),
	.A(n24180));
   INVx2_ASAP7_75t_SL FE_OFC2090_n26006 (.Y(n24180),
	.A(n26006));
   INVxp33_ASAP7_75t_L FE_OFC2078_n17815 (.Y(FE_OFN68_sa02_6),
	.A(n17815));
   INVxp33_ASAP7_75t_R FE_OFC2068_n23322 (.Y(FE_OFN16407_n23322),
	.A(FE_OFN25987_n23322));
   INVx1_ASAP7_75t_SL FE_OFC2058_n24816 (.Y(n24817),
	.A(n24816));
   INVxp67_ASAP7_75t_L FE_OFC2043_n18302 (.Y(n18303),
	.A(n18302));
   INVxp33_ASAP7_75t_R FE_OFC2037_n23023 (.Y(FE_OFN16377_n23998),
	.A(n23998));
   INVx1_ASAP7_75t_SL FE_OFC2035_n20056 (.Y(FE_OFN25972_n20056),
	.A(n20056));
   INVxp33_ASAP7_75t_SRAM FE_OFC2033_n14472 (.Y(FE_OFN25971_n14472),
	.A(n13723));
   INVxp33_ASAP7_75t_L FE_OFC2031_sa31_6 (.Y(FE_OFN25970_n),
	.A(n16377));
   INVxp67_ASAP7_75t_R FE_OFC2030_sa31_6 (.Y(n16377),
	.A(FE_OFN134_sa31_6));
   INVx1_ASAP7_75t_L FE_OFC2023_n22668 (.Y(FE_OFN25968_n22668),
	.A(n22675));
   INVx1_ASAP7_75t_SL FE_OFC2022_n22668 (.Y(n22675),
	.A(n22668));
   INVxp33_ASAP7_75t_R FE_OFC2021_n17109 (.Y(n17110),
	.A(n17109));
   INVx2_ASAP7_75t_L FE_OFC2008_w3_8 (.Y(FE_OFN25961_w3_8),
	.A(w3_8_));
   INVx2_ASAP7_75t_SL FE_OFC2005_n16434 (.Y(n16923),
	.A(n16434));
   BUFx8_ASAP7_75t_SL FE_OFC2002_n23011 (.Y(FE_OFN130_sa10_5),
	.A(sa10_5_));
   INVxp67_ASAP7_75t_L FE_OFC1999_n21412 (.Y(n21368),
	.A(n21412));
   INVx1_ASAP7_75t_SL FE_OFC1992_n25122 (.Y(FE_OFN25955_n25122),
	.A(n25123));
   INVx2_ASAP7_75t_SL FE_OFC1991_n25122 (.Y(n25123),
	.A(n25122));
   INVx1_ASAP7_75t_SL FE_OFC1983_n21351 (.Y(n21352),
	.A(n21351));
   INVx1_ASAP7_75t_L FE_OFC1965_sa32_6 (.Y(n25034),
	.A(sa32_6_));
   INVxp67_ASAP7_75t_L FE_OFC1964_n23270 (.Y(n23257),
	.A(n23270));
   INVxp33_ASAP7_75t_R FE_OFC1959_n22768 (.Y(n22737),
	.A(n22768));
   INVx1_ASAP7_75t_R FE_OFC1957_n22857 (.Y(n23311),
	.A(n22857));
   INVxp67_ASAP7_75t_R FE_OFC1955_n24621 (.Y(FE_OFN25940_n24621),
	.A(n18434));
   INVx1_ASAP7_75t_SL FE_OFC1939_n18859 (.Y(n18880),
	.A(n18859));
   INVxp33_ASAP7_75t_R FE_OFC1937_w3_26 (.Y(FE_OFN25934_n),
	.A(n24470));
   INVxp67_ASAP7_75t_L FE_OFC1904_n21788 (.Y(n21790),
	.A(n21788));
   INVxp33_ASAP7_75t_L FE_OFC1899_n21308 (.Y(n21311),
	.A(n21308));
   BUFx6f_ASAP7_75t_SL FE_OFC1893_sa11_3 (.Y(n19170),
	.A(sa11_3_));
   INVx1_ASAP7_75t_L FE_OFC1892_n15995 (.Y(FE_OFN25920_n15995),
	.A(n15374));
   INVx1_ASAP7_75t_SL FE_OFC1890_n15995 (.Y(n15374),
	.A(n15995));
   INVx1_ASAP7_75t_SL FE_OFC1875_n20527 (.Y(FE_OFN16319_n20527),
	.A(FE_OCPN29544_n20527));
   BUFx2_ASAP7_75t_SL FE_OFC1872_n15514 (.Y(n15714),
	.A(n15514));
   INVx1_ASAP7_75t_R FE_OFC1858_n23693 (.Y(n23803),
	.A(n23693));
   INVx1_ASAP7_75t_L FE_OFC1840_n17691 (.Y(FE_OFN16231_n17691),
	.A(n17691));
   INVxp67_ASAP7_75t_L FE_OFC1839_n22290 (.Y(n22291),
	.A(n22290));
   BUFx2_ASAP7_75t_SL FE_OFC1829_w3_4 (.Y(FE_OFN25900_w3_4),
	.A(FE_OFN25896_w3_4));
   INVxp67_ASAP7_75t_R FE_OFC1828_w3_4 (.Y(FE_OFN25899_w3_4),
	.A(FE_OFN25896_w3_4));
   INVx1_ASAP7_75t_L FE_OFC1826_w3_4 (.Y(FE_OFN25897_w3_4),
	.A(FE_OFN25896_w3_4));
   INVx2_ASAP7_75t_SL FE_OFC1825_w3_4 (.Y(FE_OFN25896_w3_4),
	.A(w3_4_));
   INVx2_ASAP7_75t_L FE_OFC1822_n13662 (.Y(FE_OFN25895_n13662),
	.A(FE_OFN27057_n13662));
   INVx1_ASAP7_75t_SRAM FE_OFC1817_n23413 (.Y(n21045),
	.A(n23413));
   INVx1_ASAP7_75t_L FE_OFC1813_n15214 (.Y(FE_OFN16145_n15214),
	.A(n15233));
   INVx2_ASAP7_75t_L FE_OFC1812_n15214 (.Y(FE_OFN16437_n),
	.A(FE_OFN25893_n15214));
   INVx1_ASAP7_75t_SL FE_OFC1805_n23497 (.Y(n20242),
	.A(n23497));
   INVx1_ASAP7_75t_SL FE_OFC1770_n15501 (.Y(n14778),
	.A(n15501));
   INVx1_ASAP7_75t_SL FE_OFC1769_n14044 (.Y(n13917),
	.A(n14044));
   INVx1_ASAP7_75t_L FE_OFC1767_n16262 (.Y(FE_OFN25882_n16262),
	.A(FE_OFN16370_n16261));
   INVx2_ASAP7_75t_SL FE_OFC1766_n16262 (.Y(FE_OFN16370_n16261),
	.A(n16262));
   INVxp33_ASAP7_75t_R FE_OFC1762_n23055 (.Y(n23054),
	.A(n23055));
   INVx3_ASAP7_75t_SL FE_OFC1752_n15343 (.Y(n12994),
	.A(n15343));
   INVx2_ASAP7_75t_L FE_OFC1751_n14573 (.Y(n15145),
	.A(n14573));
   INVxp33_ASAP7_75t_R FE_OFC1745_w3_24 (.Y(n26798),
	.A(FE_OFN25881_w3_24));
   INVx1_ASAP7_75t_R FE_OFC1744_w3_24 (.Y(FE_OFN16159_w3_24),
	.A(w3_24_));
   INVxp67_ASAP7_75t_L FE_OFC1715_n15422 (.Y(n15975),
	.A(FE_OFN28758_n15422));
   INVx3_ASAP7_75t_SL FE_OFC1709_n22855 (.Y(n23315),
	.A(n22855));
   INVxp33_ASAP7_75t_R FE_OFC1683_w3_9 (.Y(FE_OFN16448_n),
	.A(FE_OFN16459_n));
   INVxp67_ASAP7_75t_R FE_OFC1675_n13655 (.Y(FE_OFN16236_n13655),
	.A(n13655));
   INVx1_ASAP7_75t_SRAM FE_OFC1664_sa13_6 (.Y(n19359),
	.A(FE_OFN16389_n19359));
   INVxp67_ASAP7_75t_R FE_OFC1663_sa13_6 (.Y(FE_OFN16389_n19359),
	.A(sa13_6_));
   INVxp67_ASAP7_75t_R FE_OFC1620_w3_21 (.Y(FE_OFN16441_w3_21),
	.A(n25961));
   INVxp67_ASAP7_75t_R FE_OFC1611_w3_16 (.Y(FE_OFN16432_w3_16),
	.A(FE_OFN16431_w3_16));
   INVxp67_ASAP7_75t_R FE_OFC1610_w3_16 (.Y(FE_OFN16431_w3_16),
	.A(FE_OFN28701_w3_16));
   HB1xp67_ASAP7_75t_L FE_OFC1592_n26687 (.Y(FE_OFN16413_n26687),
	.A(n26687));
   BUFx2_ASAP7_75t_R FE_OFC1591_w3_26 (.Y(FE_OFN16412_w3_26),
	.A(w3_26_));
   HB1xp67_ASAP7_75t_L FE_OFC1590_n15884 (.Y(FE_OFN16411_n15884),
	.A(n15884));
   INVxp33_ASAP7_75t_R FE_OFC1583_n18030 (.Y(FE_OFN156_sa03_6),
	.A(sa03_6_));
   INVx1_ASAP7_75t_L FE_OFC1581_n24705 (.Y(n26875),
	.A(n24705));
   HB1xp67_ASAP7_75t_SL FE_OFC1563_n25869 (.Y(FE_OFN16396_n25869),
	.A(FE_OFN16162_n25869));
   INVxp33_ASAP7_75t_L FE_OFC1558_n26801 (.Y(n26806),
	.A(n26801));
   INVxp33_ASAP7_75t_R FE_OFC1553_n23904 (.Y(n23907),
	.A(n23904));
   INVx1_ASAP7_75t_SL FE_OFC1550_n22490 (.Y(n21377),
	.A(n22490));
   INVx3_ASAP7_75t_SL FE_OFC1537_sa32_1 (.Y(n17526),
	.A(sa32_1_));
   INVxp67_ASAP7_75t_SL FE_OFC1536_n21158 (.Y(n21160),
	.A(n21158));
   INVx1_ASAP7_75t_SL FE_OFC1532_n20584 (.Y(FE_OFN16380_n20584),
	.A(n20584));
   INVxp33_ASAP7_75t_L FE_OFC1528_n23030 (.Y(FE_OFN16378_n23030),
	.A(n16612));
   INVx1_ASAP7_75t_L FE_OFC1527_n23030 (.Y(n16612),
	.A(n23030));
   INVxp33_ASAP7_75t_SRAM FE_OFC1526_n16258 (.Y(n16164),
	.A(n16258));
   INVxp33_ASAP7_75t_R FE_OFC1512_n22565 (.Y(n22566),
	.A(n22565));
   INVx1_ASAP7_75t_SL FE_OFC1510_n16261 (.Y(n16262),
	.A(n16261));
   INVxp67_ASAP7_75t_R FE_OFC1503_n17129 (.Y(n17036),
	.A(n17129));
   INVx2_ASAP7_75t_SL FE_OFC1502_n25922 (.Y(n25923),
	.A(n25922));
   INVxp33_ASAP7_75t_L FE_OFC1500_n21973 (.Y(FE_OFN16367_n21973),
	.A(n20865));
   INVxp67_ASAP7_75t_R FE_OFC1477_n19485 (.Y(n21753),
	.A(n19485));
   INVxp33_ASAP7_75t_L FE_OFC1451_n19960 (.Y(FE_OFN16349_n19960),
	.A(n17530));
   INVxp67_ASAP7_75t_L FE_OFC1447_n15949 (.Y(n15950),
	.A(n15949));
   INVxp33_ASAP7_75t_L FE_OFC1435_n16106 (.Y(n15907),
	.A(n16106));
   INVxp67_ASAP7_75t_L FE_OFC1429_n13329 (.Y(n13330),
	.A(n13329));
   INVxp67_ASAP7_75t_R FE_OFC1427_n16563 (.Y(FE_OFN59_sa10_7),
	.A(n16563));
   INVx1_ASAP7_75t_SL FE_OFC1371_n22115 (.Y(n20974),
	.A(n22115));
   INVx1_ASAP7_75t_SL FE_OFC1368_n21650 (.Y(n20680),
	.A(n21650));
   INVxp33_ASAP7_75t_R FE_OFC1366_w3_0 (.Y(FE_OFN16313_w3_0),
	.A(n25596));
   INVx1_ASAP7_75t_L FE_OFC1365_w3_0 (.Y(n25596),
	.A(w3_0_));
   INVxp67_ASAP7_75t_R FE_OFC1364_n22943 (.Y(n22944),
	.A(n22943));
   INVxp33_ASAP7_75t_L FE_OFC1349_n16186 (.Y(n16120),
	.A(n16186));
   INVx2_ASAP7_75t_SL FE_OFC1346_n16150 (.Y(n16152),
	.A(n16150));
   INVxp67_ASAP7_75t_L FE_OFC1343_n15798 (.Y(n15076),
	.A(n15798));
   INVx1_ASAP7_75t_R FE_OFC1342_n15984 (.Y(FE_OFN16305_n15984),
	.A(n14615));
   INVx1_ASAP7_75t_L FE_OFC1341_n15984 (.Y(n14615),
	.A(n15984));
   INVxp33_ASAP7_75t_L FE_OFC1340_n19161 (.Y(FE_OFN150_sa11_7),
	.A(n19161));
   INVxp67_ASAP7_75t_R FE_OFC1334_n19101 (.Y(n18616),
	.A(n19101));
   INVx1_ASAP7_75t_L FE_OFC1327_n14826 (.Y(FE_OFN56_n14826),
	.A(n14826));
   INVxp67_ASAP7_75t_L FE_OFC1311_n25175 (.Y(FE_OFN16292_n25175),
	.A(n25748));
   BUFx6f_ASAP7_75t_SL FE_OFC1306_n23774 (.Y(n20670),
	.A(n23774));
   INVxp33_ASAP7_75t_L FE_OFC1303_n24205 (.Y(n24208),
	.A(n24205));
   INVxp67_ASAP7_75t_SL FE_OFC1297_n15652 (.Y(n15653),
	.A(n15652));
   INVxp33_ASAP7_75t_R FE_OFC1295_n18707 (.Y(n18708),
	.A(n18707));
   INVxp67_ASAP7_75t_L FE_OFC1280_n14099 (.Y(n13986),
	.A(n14099));
   INVxp33_ASAP7_75t_L FE_OFC1273_n15492 (.Y(n14755),
	.A(n15492));
   INVxp33_ASAP7_75t_R FE_OFC1272_n26011 (.Y(FE_OFN16281_n26011),
	.A(n26012));
   INVx1_ASAP7_75t_SL FE_OFC1271_n26011 (.Y(n26012),
	.A(n26011));
   INVxp67_ASAP7_75t_L FE_OFC1267_n24483 (.Y(n24486),
	.A(n24483));
   INVxp33_ASAP7_75t_L FE_OFC1263_w3_5 (.Y(FE_OFN16278_w3_5),
	.A(FE_OFN16276_w3_5));
   INVx1_ASAP7_75t_R FE_OFC1261_w3_5 (.Y(FE_OFN16276_w3_5),
	.A(FE_OFN29052_w3_5));
   INVxp67_ASAP7_75t_R FE_OFC1250_sa33_6 (.Y(FE_OFN174_sa33_6),
	.A(sa33_6_));
   INVxp67_ASAP7_75t_L FE_OFC1247_n26814 (.Y(FE_OFN16271_n26814),
	.A(n26815));
   INVx3_ASAP7_75t_SL FE_OFC1245_n26814 (.Y(n26815),
	.A(n26814));
   INVxp33_ASAP7_75t_R FE_OFC1240_sa13_3 (.Y(n17091),
	.A(FE_OFN16268_sa13_3));
   INVxp33_ASAP7_75t_R FE_OFC1236_n24419 (.Y(n24045),
	.A(n24419));
   INVxp33_ASAP7_75t_R FE_OFC1235_n23929 (.Y(n23930),
	.A(n23929));
   INVxp67_ASAP7_75t_L FE_OFC1234_n16208 (.Y(n16200),
	.A(n16208));
   INVxp33_ASAP7_75t_L FE_OFC1200_n15789 (.Y(n15793),
	.A(n15789));
   INVx1_ASAP7_75t_SL FE_OFC1198_n16162 (.Y(n16159),
	.A(n16162));
   INVxp67_ASAP7_75t_R FE_OFC1185_n13665 (.Y(n15159),
	.A(n13665));
   INVx1_ASAP7_75t_R FE_OFC1169_n17020 (.Y(FE_OFN128_sa13_7),
	.A(n17020));
   INVx1_ASAP7_75t_SL FE_OFC1166_n14171 (.Y(n14174),
	.A(n14171));
   INVxp67_ASAP7_75t_L FE_OFC1165_n16870 (.Y(n24335),
	.A(n16870));
   INVxp67_ASAP7_75t_R FE_OFC1164_n13290 (.Y(n13291),
	.A(n13290));
   INVx2_ASAP7_75t_SL FE_OFC1162_n16048 (.Y(n16047),
	.A(FE_OCPN28075_n16048));
   INVxp33_ASAP7_75t_R FE_OFC1159_n23299 (.Y(n23305),
	.A(n23299));
   INVx1_ASAP7_75t_L FE_OFC1157_n14005 (.Y(FE_OFN16239_n14005),
	.A(n14004));
   BUFx2_ASAP7_75t_SL FE_OFC1156_n14005 (.Y(n14004),
	.A(n14005));
   INVxp33_ASAP7_75t_L FE_OFC1148_sa30_6 (.Y(n17629),
	.A(sa30_6_));
   INVxp67_ASAP7_75t_R FE_OFC1139_n24474 (.Y(n21446),
	.A(n24474));
   INVxp67_ASAP7_75t_L FE_OFC1138_n14775 (.Y(n14776),
	.A(n14775));
   INVxp67_ASAP7_75t_SL FE_OFC1121_n22720 (.Y(n23224),
	.A(n22720));
   INVx1_ASAP7_75t_L FE_OFC1115_n21234 (.Y(n23691),
	.A(n21234));
   INVxp67_ASAP7_75t_SL FE_OFC1113_n16097 (.Y(n16096),
	.A(FE_OCPN29581_n16097));
   INVxp67_ASAP7_75t_R FE_OFC1109_n16857 (.Y(n16860),
	.A(FE_OFN79_n16857));
   INVx1_ASAP7_75t_SL FE_OFC1108_n16857 (.Y(FE_OFN79_n16857),
	.A(n16857));
   INVxp33_ASAP7_75t_R FE_OFC1107_n25881 (.Y(n18917),
	.A(n25881));
   INVxp33_ASAP7_75t_L FE_OFC1105_sa23_7 (.Y(FE_OFN162_sa23_7),
	.A(sa23_7_));
   HB1xp67_ASAP7_75t_SL FE_OFC1087_ld_r (.Y(FE_OFN16215_ld_r),
	.A(FE_DBTN0_ld_r));
   INVx1_ASAP7_75t_SL FE_OFC1078_n25805 (.Y(n25806),
	.A(n25805));
   INVxp67_ASAP7_75t_SL FE_OFC1068_n14178 (.Y(n14179),
	.A(n14178));
   INVxp33_ASAP7_75t_R FE_OFC1067_n19394 (.Y(n19393),
	.A(n19394));
   INVxp33_ASAP7_75t_R FE_OFC1060_n15407 (.Y(n15408),
	.A(n15407));
   INVxp67_ASAP7_75t_L FE_OFC1059_n13532 (.Y(n13535),
	.A(n13532));
   INVxp33_ASAP7_75t_L FE_OFC1057_n23992 (.Y(FE_OFN169_n23992),
	.A(n23992));
   INVxp33_ASAP7_75t_L FE_OFC1054_n23483 (.Y(n23485),
	.A(n23483));
   INVxp67_ASAP7_75t_L FE_OFC1047_n20915 (.Y(n19339),
	.A(n20915));
   INVxp33_ASAP7_75t_R FE_OFC1046_n14485 (.Y(n13554),
	.A(n14485));
   INVxp33_ASAP7_75t_L FE_OFC1045_n20219 (.Y(n20218),
	.A(n20219));
   INVxp33_ASAP7_75t_R FE_OFC1043_n15780 (.Y(n15783),
	.A(n15780));
   INVxp33_ASAP7_75t_L FE_OFC1042_n18517 (.Y(n18516),
	.A(n18517));
   INVxp67_ASAP7_75t_R FE_OFC1039_n13904 (.Y(n13881),
	.A(n13904));
   INVxp67_ASAP7_75t_R FE_OFC1036_n19447 (.Y(n18004),
	.A(n19447));
   INVxp33_ASAP7_75t_R FE_OFC1033_n20070 (.Y(n20071),
	.A(n20070));
   INVxp33_ASAP7_75t_L FE_OFC1029_n19434 (.Y(n18952),
	.A(n19434));
   INVxp33_ASAP7_75t_L FE_OFC1026_n25793 (.Y(n21401),
	.A(n25793));
   INVxp33_ASAP7_75t_L FE_OFC1025_n15296 (.Y(n15297),
	.A(n15296));
   INVxp33_ASAP7_75t_R FE_OFC1019_n16158 (.Y(n16066),
	.A(n16158));
   INVx1_ASAP7_75t_L FE_OFC1015_n23487 (.Y(n20911),
	.A(n23487));
   INVxp67_ASAP7_75t_R FE_OFC1006_n15870 (.Y(n15875),
	.A(n15870));
   INVxp67_ASAP7_75t_L FE_OFC1005_n22134 (.Y(n17623),
	.A(n22134));
   INVxp67_ASAP7_75t_L FE_OFC1001_n15402 (.Y(n13816),
	.A(n15402));
   INVxp33_ASAP7_75t_L FE_OFC1000_n24473 (.Y(n24475),
	.A(n24473));
   INVxp67_ASAP7_75t_R FE_OFC984_n16023 (.Y(n14183),
	.A(n16023));
   INVxp67_ASAP7_75t_R FE_OFC981_sa32_7 (.Y(FE_OFN136_sa32_7),
	.A(sa32_7_));
   INVxp33_ASAP7_75t_L FE_OFC969_n23246 (.Y(n22480),
	.A(n23246));
   INVxp67_ASAP7_75t_R FE_OFC961_sa31_6 (.Y(FE_OFN16197_sa31_6),
	.A(FE_OFN25970_n));
   INVxp33_ASAP7_75t_R FE_OFC959_sa31_6 (.Y(FE_OFN134_sa31_6),
	.A(sa31_6_));
   INVx2_ASAP7_75t_SL FE_OFC947_n13771 (.Y(FE_OFN16195_n13771),
	.A(n13771));
   INVx2_ASAP7_75t_SL FE_OFC946_n13771 (.Y(n13729),
	.A(n13771));
   BUFx2_ASAP7_75t_SL FE_OFC929_n15180 (.Y(n15200),
	.A(n15180));
   BUFx2_ASAP7_75t_R FE_OFC911_n26542 (.Y(FE_OFN16180_n26542),
	.A(n26542));
   INVxp67_ASAP7_75t_R FE_OFC910_w3_19 (.Y(FE_OFN16179_w3_19),
	.A(FE_OFN16178_w3_19));
   INVxp33_ASAP7_75t_L FE_OFC909_w3_19 (.Y(FE_OFN16178_w3_19),
	.A(FE_OFN27096_n));
   HB1xp67_ASAP7_75t_R FE_OFC908_n27207 (.Y(FE_OFN16177_n27207),
	.A(n27207));
   BUFx2_ASAP7_75t_SRAM FE_OFC907_n27207 (.Y(FE_OFN16176_n27207),
	.A(n27207));
   BUFx2_ASAP7_75t_SRAM FE_OFC901_n26637 (.Y(FE_OFN16170_n26637),
	.A(n26637));
   BUFx2_ASAP7_75t_SRAM FE_OFC900_n26567 (.Y(FE_OFN16169_n26567),
	.A(n26567));
   HB1xp67_ASAP7_75t_R FE_OFC895_n25081 (.Y(FE_OFN16164_n25081),
	.A(n25081));
   BUFx2_ASAP7_75t_R FE_OFC894_n26584 (.Y(FE_OFN16163_n26584),
	.A(n26584));
   BUFx2_ASAP7_75t_R FE_OFC889_n26959 (.Y(FE_OFN16158_n26959),
	.A(n26959));
   HB1xp67_ASAP7_75t_L FE_OFC879_n25466 (.Y(FE_OFN16148_n25466),
	.A(n25466));
   INVx4_ASAP7_75t_SL FE_OFC872_sa01_3 (.Y(FE_OFN16141_sa01_3),
	.A(FE_OFN26132_sa01_3));
   BUFx6f_ASAP7_75t_SL FE_OFC866_sa22_4 (.Y(FE_OFN16135_sa22_4),
	.A(sa22_4_));
   INVxp67_ASAP7_75t_R FE_OFC854_sa12_6 (.Y(FE_OFN175_sa12_6),
	.A(n17915));
   INVxp67_ASAP7_75t_L FE_OFC853_sa12_6 (.Y(n17915),
	.A(sa12_6_));
   INVxp33_ASAP7_75t_R FE_OFC851_sa33_6 (.Y(FE_OFN173_sa33_6),
	.A(FE_OFN174_sa33_6));
   INVxp33_ASAP7_75t_R FE_OFC837_sa12_7 (.Y(FE_OFN166_sa12_7),
	.A(FE_OFN165_sa12_7));
   INVxp67_ASAP7_75t_R FE_OFC835_sa12_7 (.Y(n24590),
	.A(sa12_7_));
   INVxp67_ASAP7_75t_R FE_OFC832_sa00_7 (.Y(FE_OFN163_sa00_7),
	.A(sa00_7_));
   INVxp33_ASAP7_75t_L FE_OFC821_n21965 (.Y(n21967),
	.A(n21965));
   INVxp33_ASAP7_75t_R FE_OFC815_n26898 (.Y(n23848),
	.A(FE_OCPN7621_n26898));
   INVxp67_ASAP7_75t_R FE_OFC808_sa11_7 (.Y(n19161),
	.A(sa11_7_));
   INVxp33_ASAP7_75t_L FE_OFC795_n23942 (.Y(n18002),
	.A(n23942));
   INVxp33_ASAP7_75t_R FE_OFC794_w3_2 (.Y(FE_OFN140_w3_2),
	.A(n23937));
   INVxp67_ASAP7_75t_R FE_OFC792_w3_2 (.Y(n23937),
	.A(w3_2_));
   INVxp33_ASAP7_75t_R FE_OFC791_n25231 (.Y(n16995),
	.A(n25231));
   HB1xp67_ASAP7_75t_L FE_OFC784_n26172 (.Y(n26171),
	.A(FE_OCPN27373_n26172));
   INVx3_ASAP7_75t_SL FE_OFC781_n24306 (.Y(FE_OFN133_n24306),
	.A(n24306));
   INVxp67_ASAP7_75t_SRAM FE_OFC777_sa10_6 (.Y(FE_OFN131_sa10_6),
	.A(sa10_6_));
   INVxp67_ASAP7_75t_R FE_OFC769_sa13_7 (.Y(n17020),
	.A(sa13_7_));
   INVxp33_ASAP7_75t_R FE_OFC748_n26594 (.Y(n26595),
	.A(n26594));
   INVxp67_ASAP7_75t_L FE_OFC744_n26120 (.Y(n24612),
	.A(n26120));
   INVxp33_ASAP7_75t_L FE_OFC739_n27187 (.Y(FE_OFN116_n27187),
	.A(FE_OFN115_n27187));
   INVx1_ASAP7_75t_L FE_OFC734_n27072 (.Y(n25338),
	.A(n27072));
   INVx1_ASAP7_75t_R FE_OFC731_n22512 (.Y(n19188),
	.A(n22512));
   INVxp67_ASAP7_75t_SL FE_OFC730_n21162 (.Y(n21186),
	.A(n21162));
   INVxp67_ASAP7_75t_R FE_OFC729_n23432 (.Y(n23435),
	.A(n23432));
   INVxp67_ASAP7_75t_SL FE_OFC722_n22536 (.Y(n20145),
	.A(n22536));
   INVxp67_ASAP7_75t_R FE_OFC718_n20932 (.Y(n19317),
	.A(n20932));
   INVxp33_ASAP7_75t_L FE_OFC714_n22745 (.Y(FE_OFN107_n22745),
	.A(n22745));
   INVx2_ASAP7_75t_SL FE_OFC710_n24511 (.Y(n24510),
	.A(n24511));
   INVxp67_ASAP7_75t_L FE_OFC709_n27031 (.Y(n24603),
	.A(n27031));
   INVxp33_ASAP7_75t_R FE_OFC708_n19828 (.Y(n19829),
	.A(n19828));
   INVxp33_ASAP7_75t_R FE_OFC704_n25563 (.Y(n19392),
	.A(n25563));
   INVxp33_ASAP7_75t_L FE_OFC696_n25279 (.Y(n19415),
	.A(n25279));
   INVxp33_ASAP7_75t_R FE_OFC689_w3_12 (.Y(FE_OFN102_w3_12),
	.A(FE_OCPN29520_n24755));
   BUFx6f_ASAP7_75t_L FE_OFC687_w3_12 (.Y(n24755),
	.A(w3_12_));
   INVx1_ASAP7_75t_SL FE_OFC681_n21049 (.Y(n21052),
	.A(n21049));
   INVxp33_ASAP7_75t_L FE_OFC679_n22435 (.Y(n20410),
	.A(n22435));
   INVxp33_ASAP7_75t_L FE_OFC673_n25223 (.Y(n25224),
	.A(n25223));
   INVxp67_ASAP7_75t_L FE_OFC671_n24381 (.Y(n23576),
	.A(n24381));
   INVxp67_ASAP7_75t_R FE_OFC657_sa33_7 (.Y(FE_OFN90_sa33_7),
	.A(n16468));
   INVxp67_ASAP7_75t_R FE_OFC654_sa33_7 (.Y(n16468),
	.A(sa33_7_));
   INVx2_ASAP7_75t_SL FE_OFC648_n24449 (.Y(n24450),
	.A(n24449));
   INVxp67_ASAP7_75t_SL FE_OFC647_n16203 (.Y(n16198),
	.A(n16203));
   INVxp33_ASAP7_75t_L FE_OFC642_n19618 (.Y(n19621),
	.A(n19618));
   INVxp33_ASAP7_75t_L FE_OFC630_n24000 (.Y(n23022),
	.A(n24000));
   INVx2_ASAP7_75t_SL FE_OFC609_n21942 (.Y(n20039),
	.A(n21942));
   INVxp33_ASAP7_75t_R FE_OFC608_n24759 (.Y(n18510),
	.A(n24759));
   INVxp33_ASAP7_75t_L FE_OFC603_n24344 (.Y(n24346),
	.A(n24344));
   INVx1_ASAP7_75t_L FE_OFC599_n26704 (.Y(n26705),
	.A(n26704));
   INVxp33_ASAP7_75t_L FE_OFC597_n25199 (.Y(n17040),
	.A(FE_OCPN8234_n25199));
   INVx1_ASAP7_75t_SL FE_OFC595_n15138 (.Y(n15139),
	.A(n15138));
   INVxp33_ASAP7_75t_R FE_OFC591_w2_20 (.Y(FE_OFN70_w2_20),
	.A(w2_20_));
   INVxp67_ASAP7_75t_L FE_OFC589_n19598 (.Y(n19600),
	.A(n19598));
   INVx1_ASAP7_75t_SL FE_OFC581_n16148 (.Y(n16149),
	.A(n16148));
   INVx1_ASAP7_75t_L FE_OFC580_n22349 (.Y(n16795),
	.A(n22349));
   INVxp67_ASAP7_75t_R FE_OFC572_w1_25 (.Y(FE_OFN66_w1_25),
	.A(w1_25_));
   INVxp33_ASAP7_75t_L FE_OFC569_n23882 (.Y(n23883),
	.A(n23882));
   INVxp33_ASAP7_75t_R FE_OFC562_w0_31 (.Y(FE_OFN64_w0_31),
	.A(n26811));
   INVxp33_ASAP7_75t_L FE_OFC561_w0_31 (.Y(n26811),
	.A(w0_31_));
   INVxp67_ASAP7_75t_R FE_OFC559_n23443 (.Y(n23444),
	.A(n23443));
   INVx1_ASAP7_75t_SL FE_OFC557_n16156 (.Y(n16153),
	.A(n16156));
   INVxp67_ASAP7_75t_L FE_OFC554_n20268 (.Y(n20269),
	.A(n20268));
   INVx1_ASAP7_75t_SL FE_OFC548_sa21_3 (.Y(FE_OFN62_sa21_3),
	.A(FE_OFN28678_sa21_3));
   INVxp33_ASAP7_75t_L FE_OFC541_n19603 (.Y(n19604),
	.A(n19603));
   INVx1_ASAP7_75t_SL FE_OFC530_n26467 (.Y(n26466),
	.A(n26467));
   INVxp33_ASAP7_75t_SRAM FE_OFC527_n16131 (.Y(n16056),
	.A(n16131));
   INVxp33_ASAP7_75t_L FE_OFC526_n25635 (.Y(n23795),
	.A(n25635));
   INVxp33_ASAP7_75t_SRAM FE_OFC525_n15904 (.Y(n14408),
	.A(n15904));
   INVx1_ASAP7_75t_SL FE_OFC523_n27007 (.Y(FE_OFN60_n27007),
	.A(n27007));
   BUFx2_ASAP7_75t_L FE_OFC522_n27007 (.Y(n22597),
	.A(n27007));
   INVxp33_ASAP7_75t_L FE_OFC518_sa10_7 (.Y(n16563),
	.A(sa10_7_));
   INVxp67_ASAP7_75t_L FE_OFC517_n23203 (.Y(n20735),
	.A(n23203));
   INVxp33_ASAP7_75t_L FE_OFC513_n25022 (.Y(n25023),
	.A(n25022));
   INVxp67_ASAP7_75t_SL FE_OFC512_n24671 (.Y(n19805),
	.A(n24671));
   INVxp67_ASAP7_75t_L FE_OFC509_n22928 (.Y(n22931),
	.A(n22928));
   INVx3_ASAP7_75t_SL FE_OFC508_n26837 (.Y(n26838),
	.A(FE_OCPN27445_n26837));
   INVxp67_ASAP7_75t_L FE_OFC507_n19481 (.Y(n18013),
	.A(n19481));
   INVxp33_ASAP7_75t_R FE_OFC503_w1_4 (.Y(FE_OFN58_w1_4),
	.A(n26243));
   INVxp67_ASAP7_75t_R FE_OFC502_w1_4 (.Y(n26243),
	.A(w1_4_));
   INVx1_ASAP7_75t_SL FE_OFC501_n22355 (.Y(n20340),
	.A(n22355));
   INVx1_ASAP7_75t_R FE_OFC499_n22825 (.Y(n22829),
	.A(n22825));
   INVx1_ASAP7_75t_SL FE_OFC494_n24336 (.Y(n24338),
	.A(n24336));
   INVxp33_ASAP7_75t_L FE_OFC488_sa01_7 (.Y(n17392),
	.A(sa01_7_));
   INVxp67_ASAP7_75t_SL FE_OFC485_n22547 (.Y(n22549),
	.A(n22547));
   INVxp33_ASAP7_75t_L FE_OFC476_n21121 (.Y(n21113),
	.A(n21121));
   INVx1_ASAP7_75t_L FE_OFC475_n16406 (.Y(n16362),
	.A(n16406));
   INVx1_ASAP7_75t_L FE_OFC461_sa22_2 (.Y(FE_OFN54_sa22_2),
	.A(FE_OFN28688_sa22_2));
   INVxp67_ASAP7_75t_L FE_OFC457_n26553 (.Y(n23486),
	.A(n26553));
   INVxp33_ASAP7_75t_R FE_OFC451_w0_8 (.Y(FE_OFN53_w0_8),
	.A(n26744));
   INVxp33_ASAP7_75t_L FE_OFC450_w0_8 (.Y(n26744),
	.A(w0_8_));
   INVxp67_ASAP7_75t_L FE_OFC449_n19848 (.Y(n19849),
	.A(n19848));
   INVxp33_ASAP7_75t_R FE_OFC441_w3_18 (.Y(FE_OFN51_w3_18),
	.A(FE_OFN16421_n23974));
   INVx1_ASAP7_75t_L FE_OFC439_w3_18 (.Y(n23974),
	.A(w3_18_));
   INVxp33_ASAP7_75t_L FE_OFC437_n16216 (.Y(n16136),
	.A(n16216));
   INVxp33_ASAP7_75t_R FE_OFC433_w0_23 (.Y(FE_OFN49_w0_23),
	.A(n27064));
   INVxp67_ASAP7_75t_R FE_OFC432_w0_23 (.Y(n27064),
	.A(w0_23_));
   INVxp33_ASAP7_75t_L FE_OFC431_w0_30 (.Y(n26645),
	.A(w0_30_));
   INVxp67_ASAP7_75t_L FE_OFC430_n13695 (.Y(n15254),
	.A(n13695));
   INVxp33_ASAP7_75t_R FE_OFC429_w0_2 (.Y(FE_OFN48_w0_2),
	.A(n24531));
   INVxp67_ASAP7_75t_R FE_OFC428_w0_2 (.Y(n24531),
	.A(w0_2_));
   INVxp67_ASAP7_75t_R FE_OFC426_n19824 (.Y(n19826),
	.A(n19824));
   INVxp33_ASAP7_75t_R FE_OFC425_n24298 (.Y(n16681),
	.A(FE_OCPN29577_n24298));
   INVxp33_ASAP7_75t_L FE_OFC424_sa31_7 (.Y(n16344),
	.A(sa31_7_));
   INVxp33_ASAP7_75t_R FE_OFC419_w1_2 (.Y(FE_OFN47_w1_2),
	.A(n26185));
   INVxp67_ASAP7_75t_L FE_OFC418_w1_2 (.Y(n26185),
	.A(w1_2_));
   INVx1_ASAP7_75t_SL FE_OFC417_n21488 (.Y(n24094),
	.A(n21488));
   INVx1_ASAP7_75t_SL FE_OFC416_n16182 (.Y(n16184),
	.A(n16182));
   INVxp33_ASAP7_75t_R FE_OFC415_w0_12 (.Y(FE_OFN46_w0_12),
	.A(n26130));
   INVxp67_ASAP7_75t_R FE_OFC414_w0_12 (.Y(n26130),
	.A(w0_12_));
   INVx1_ASAP7_75t_L FE_OFC413_n25827 (.Y(n25826),
	.A(n25827));
   INVxp67_ASAP7_75t_R FE_OFC412_sa23_6 (.Y(FE_OFN45_sa23_6),
	.A(n26562));
   INVxp67_ASAP7_75t_L FE_OFC411_sa23_6 (.Y(n26562),
	.A(sa23_6_));
   INVxp33_ASAP7_75t_L FE_OFC406_n25601 (.Y(n24477),
	.A(n25601));
   INVx1_ASAP7_75t_L FE_OFC401_n26311 (.Y(n26946),
	.A(n26311));
   INVx2_ASAP7_75t_SL FE_OFC399_n26633 (.Y(n26631),
	.A(FE_OCPN27284_n26633));
   INVxp67_ASAP7_75t_SL FE_OFC398_n14967 (.Y(n14966),
	.A(n14967));
   INVxp33_ASAP7_75t_L FE_OFC393_w0_29 (.Y(n26385),
	.A(w0_29_));
   INVxp33_ASAP7_75t_L FE_OFC391_w0_26 (.Y(n26396),
	.A(w0_26_));
   INVxp33_ASAP7_75t_L FE_OFC389_w0_24 (.Y(n26436),
	.A(w0_24_));
   INVx1_ASAP7_75t_SL FE_OFC388_n24809 (.Y(n24807),
	.A(n24809));
   INVx1_ASAP7_75t_SL FE_OFC386_n20507 (.Y(n17134),
	.A(n20507));
   INVxp33_ASAP7_75t_R FE_OFC383_n21195 (.Y(n18574),
	.A(n21195));
   INVxp67_ASAP7_75t_R FE_OFC381_w1_3 (.Y(n26578),
	.A(w1_3_));
   INVxp33_ASAP7_75t_R FE_OFC380_w0_9 (.Y(FE_OFN44_w0_9),
	.A(n24320));
   INVxp67_ASAP7_75t_R FE_OFC379_w0_9 (.Y(n24320),
	.A(w0_9_));
   INVxp33_ASAP7_75t_L FE_OFC376_w0_10 (.Y(FE_OFN43_w0_10),
	.A(n24641));
   INVxp67_ASAP7_75t_R FE_OFC375_w0_10 (.Y(n24641),
	.A(w0_10_));
   INVx1_ASAP7_75t_R FE_OFC367_n16114 (.Y(n16115),
	.A(FE_OCPN29550_n16114));
   INVxp67_ASAP7_75t_SL FE_OFC352_n26253 (.Y(n26254),
	.A(n26253));
   INVx1_ASAP7_75t_SL FE_OFC351_n22456 (.Y(n24393),
	.A(n22456));
   INVx1_ASAP7_75t_SL FE_OFC348_n25133 (.Y(n25134),
	.A(n25133));
   INVxp33_ASAP7_75t_L FE_OFC345_sa20_6 (.Y(n24154),
	.A(sa20_6_));
   INVxp67_ASAP7_75t_SL FE_OFC336_n14819 (.Y(n14818),
	.A(n14819));
   INVxp67_ASAP7_75t_R FE_OFC333_w1_1 (.Y(n26991),
	.A(w1_1_));
   INVxp67_ASAP7_75t_R FE_OFC329_w0_14 (.Y(n24495),
	.A(w0_14_));
   INVxp33_ASAP7_75t_L FE_OFC328_n15872 (.Y(n15873),
	.A(n15872));
   INVxp33_ASAP7_75t_R FE_OFC327_n15658 (.Y(n15659),
	.A(n15658));
   INVxp33_ASAP7_75t_L FE_OFC324_w2_9 (.Y(n25346),
	.A(w2_9_));
   INVxp67_ASAP7_75t_R FE_OFC322_w1_22 (.Y(n24073),
	.A(w1_22_));
   INVxp67_ASAP7_75t_SL FE_OFC312_n13795 (.Y(n13794),
	.A(n13795));
   INVxp33_ASAP7_75t_L FE_OFC311_n19910 (.Y(n18834),
	.A(n19910));
   INVxp67_ASAP7_75t_L FE_OFC308_n26937 (.Y(n26935),
	.A(n26937));
   INVx1_ASAP7_75t_L FE_OFC304_n19404 (.Y(n25290),
	.A(n19404));
   INVxp67_ASAP7_75t_R FE_OFC302_w1_21 (.Y(n24435),
	.A(w1_21_));
   INVxp67_ASAP7_75t_L FE_OFC301_n16094 (.Y(n16095),
	.A(n16094));
   INVxp67_ASAP7_75t_L FE_OFC300_n22670 (.Y(n22671),
	.A(n22670));
   INVxp33_ASAP7_75t_L FE_OFC299_w0_4 (.Y(n25802),
	.A(w0_4_));
   INVx1_ASAP7_75t_L FE_OFC295_n16720 (.Y(n18128),
	.A(n16720));
   INVx1_ASAP7_75t_SL FE_OFC293_n24891 (.Y(n17830),
	.A(n24891));
   INVxp33_ASAP7_75t_L FE_OFC283_w0_15 (.Y(n26272),
	.A(w0_15_));
   INVxp67_ASAP7_75t_SL FE_OFC281_n25193 (.Y(n25192),
	.A(n25193));
   INVxp33_ASAP7_75t_R FE_OFC278_n15040 (.Y(n15041),
	.A(n15040));
   INVxp67_ASAP7_75t_SRAM FE_OFC276_w0_3 (.Y(n26772),
	.A(w0_3_));
   INVxp67_ASAP7_75t_R FE_OFC275_w2_27 (.Y(n25570),
	.A(w2_27_));
   INVx1_ASAP7_75t_L FE_OFC272_n19551 (.Y(n17931),
	.A(n19551));
   INVxp67_ASAP7_75t_L FE_OFC265_w2_11 (.Y(n26963),
	.A(w2_11_));
   INVx1_ASAP7_75t_SL FE_OFC262_n27012 (.Y(n17337),
	.A(n27012));
   INVxp67_ASAP7_75t_SL FE_OFC260_n16037 (.Y(n16038),
	.A(n16037));
   INVxp67_ASAP7_75t_SL FE_OFC259_n26349 (.Y(n24907),
	.A(n26349));
   INVxp33_ASAP7_75t_L FE_OFC257_w0_1 (.Y(n25265),
	.A(w0_1_));
   INVxp33_ASAP7_75t_L FE_OFC256_w0_7 (.Y(n26544),
	.A(w0_7_));
   INVxp33_ASAP7_75t_R FE_OFC253_w1_28 (.Y(n26142),
	.A(w1_28_));
   INVxp67_ASAP7_75t_R FE_OFC252_w1_17 (.Y(n26210),
	.A(w1_17_));
   INVxp33_ASAP7_75t_R FE_OFC246_n25220 (.Y(n17050),
	.A(n25220));
   INVxp33_ASAP7_75t_L FE_OFC244_w0_25 (.Y(n24575),
	.A(w0_25_));
   INVxp67_ASAP7_75t_R FE_OFC243_w1_5 (.Y(n24149),
	.A(w1_5_));
   INVxp67_ASAP7_75t_R FE_OFC239_w2_3 (.Y(n26310),
	.A(w2_3_));
   INVx2_ASAP7_75t_L FE_OFC236_n16080 (.Y(n16082),
	.A(n16080));
   INVxp67_ASAP7_75t_R FE_OFC235_w0_19 (.Y(FE_OFN40_w0_19),
	.A(n26221));
   INVxp67_ASAP7_75t_L FE_OFC234_w0_19 (.Y(n26221),
	.A(w0_19_));
   INVx1_ASAP7_75t_L FE_OFC232_n21619 (.Y(n22626),
	.A(n21619));
   INVxp67_ASAP7_75t_R FE_OFC231_w2_5 (.Y(n24200),
	.A(w2_5_));
   INVxp33_ASAP7_75t_R FE_OFC229_w0_21 (.Y(FE_OFN39_w0_21),
	.A(n24358));
   INVxp67_ASAP7_75t_R FE_OFC228_w0_21 (.Y(n24358),
	.A(w0_21_));
   INVxp67_ASAP7_75t_R FE_OFC222_w1_23 (.Y(n24608),
	.A(w1_23_));
   INVxp67_ASAP7_75t_R FE_OFC221_w0_13 (.Y(n27160),
	.A(w0_13_));
   INVx1_ASAP7_75t_L FE_OFC218_n27058 (.Y(n27057),
	.A(n27058));
   INVxp67_ASAP7_75t_SL FE_OFC216_n13406 (.Y(n13405),
	.A(n13406));
   INVxp67_ASAP7_75t_L FE_OFC215_n16110 (.Y(n16104),
	.A(n16110));
   INVxp33_ASAP7_75t_L FE_OFC213_w0_17 (.Y(FE_OFN38_w0_17),
	.A(n25975));
   INVxp67_ASAP7_75t_L FE_OFC212_w0_17 (.Y(n25975),
	.A(w0_17_));
   INVxp67_ASAP7_75t_R FE_OFC211_w0_28 (.Y(n26375),
	.A(w0_28_));
   INVx1_ASAP7_75t_SL FE_OFC209_n15627 (.Y(n15817),
	.A(n15627));
   INVxp33_ASAP7_75t_R FE_OFC205_w3_23 (.Y(n26831),
	.A(FE_OCPN29502_w3_23));
   INVx1_ASAP7_75t_SL FE_OFC201_n17939 (.Y(n17941),
	.A(n17939));
   INVx1_ASAP7_75t_SL FE_OFC200_n23376 (.Y(n23377),
	.A(n23376));
   INVxp67_ASAP7_75t_R FE_OFC195_w1_11 (.Y(n25690),
	.A(w1_11_));
   INVxp67_ASAP7_75t_L FE_OFC194_n15453 (.Y(n15411),
	.A(n15453));
   INVxp33_ASAP7_75t_L FE_OFC193_n20814 (.Y(n22743),
	.A(n20814));
   INVxp67_ASAP7_75t_R FE_OFC188_w1_13 (.Y(n25774),
	.A(w1_13_));
   INVxp67_ASAP7_75t_R FE_OFC186_w2_1 (.Y(n25931),
	.A(w2_1_));
   INVxp33_ASAP7_75t_R FE_OFC185_w1_19 (.Y(n25732),
	.A(w1_19_));
   INVxp67_ASAP7_75t_SL FE_OFC184_n13544 (.Y(n13545),
	.A(n13544));
   INVx2_ASAP7_75t_SL FE_OFC183_n18161 (.Y(n21770),
	.A(n18161));
   INVxp67_ASAP7_75t_SL FE_OFC182_n15892 (.Y(n15891),
	.A(n15892));
   INVxp67_ASAP7_75t_R FE_OFC181_w0_5 (.Y(n27129),
	.A(w0_5_));
   INVxp67_ASAP7_75t_SL FE_OFC179_n14467 (.Y(n14466),
	.A(n14467));
   INVx1_ASAP7_75t_L FE_OFC176_n25077 (.Y(n25076),
	.A(n25077));
   INVxp67_ASAP7_75t_R FE_OFC175_w1_12 (.Y(n25128),
	.A(w1_12_));
   INVxp67_ASAP7_75t_R FE_OFC174_w0_6 (.Y(n24506),
	.A(w0_6_));
   INVx1_ASAP7_75t_SL FE_OFC173_n19791 (.Y(n19649),
	.A(n19791));
   INVxp67_ASAP7_75t_R FE_OFC171_w1_9 (.Y(n24821),
	.A(w1_9_));
   INVxp67_ASAP7_75t_R FE_OFC170_w1_18 (.Y(n24412),
	.A(w1_18_));
   INVxp67_ASAP7_75t_R FE_OFC169_w2_17 (.Y(n27135),
	.A(w2_17_));
   INVxp67_ASAP7_75t_SL FE_OFC166_n14084 (.Y(n14083),
	.A(n14084));
   INVxp67_ASAP7_75t_L FE_OFC163_n15491 (.Y(n14383),
	.A(n15491));
   INVx1_ASAP7_75t_L FE_OFC161_n23581 (.Y(n22735),
	.A(n23581));
   INVx1_ASAP7_75t_SL FE_OFC159_n24382 (.Y(n24383),
	.A(n24382));
   INVx2_ASAP7_75t_L FE_OFC155_n26721 (.Y(n26722),
	.A(n26721));
   INVxp67_ASAP7_75t_R FE_OFC151_w0_18 (.Y(n24118),
	.A(w0_18_));
   INVxp67_ASAP7_75t_L FE_OFC149_w2_12 (.Y(n26018),
	.A(w2_12_));
   INVxp67_ASAP7_75t_R FE_OFC148_u0_r0_rcnt_0 (.Y(n16286),
	.A(u0_r0_rcnt_0_));
   INVx1_ASAP7_75t_R FE_OFC147_n25834 (.Y(n25833),
	.A(n25834));
   INVxp67_ASAP7_75t_L FE_OFC146_w2_4 (.Y(n26202),
	.A(w2_4_));
   INVxp67_ASAP7_75t_L FE_OFC144_w2_2 (.Y(n25648),
	.A(w2_2_));
   INVxp67_ASAP7_75t_R FE_OFC143_w0_22 (.Y(n25616),
	.A(w0_22_));
   INVxp67_ASAP7_75t_R FE_OFC142_n23206 (.Y(n23209),
	.A(n23206));
   INVxp67_ASAP7_75t_L FE_OFC138_n15188 (.Y(n13310),
	.A(n15188));
   INVx1_ASAP7_75t_R FE_OFC137_n19478 (.Y(n18895),
	.A(n19478));
   INVxp67_ASAP7_75t_R FE_OFC133_w0_27 (.Y(n24721),
	.A(w0_27_));
   INVxp67_ASAP7_75t_R FE_OFC132_w0_11 (.Y(n26095),
	.A(w0_11_));
   INVxp33_ASAP7_75t_R FE_OFC128_w3_22 (.Y(FE_OFN34_w3_22),
	.A(FE_OFN7_w3_22));
   INVxp33_ASAP7_75t_L FE_OFC125_w3_22 (.Y(FE_OFN7_w3_22),
	.A(FE_OCPN7623_FE_OFN4_w3_22));
   INVxp67_ASAP7_75t_R FE_OFC120_w1_20 (.Y(n26698),
	.A(w1_20_));
   INVxp67_ASAP7_75t_R FE_OFC118_w0_20 (.Y(n26884),
	.A(w0_20_));
   INVxp67_ASAP7_75t_R FE_OFC108_w0_16 (.Y(n26486),
	.A(w0_16_));
   INVxp67_ASAP7_75t_L FE_OFC105_n15560 (.Y(n15559),
	.A(n15560));
   INVxp33_ASAP7_75t_R FE_OFC103_n25901 (.Y(n21202),
	.A(n25901));
   INVxp67_ASAP7_75t_SL FE_OFC102_n14323 (.Y(n14324),
	.A(n14323));
   INVx2_ASAP7_75t_L FE_OFC99_n16991 (.Y(n17060),
	.A(FE_OCPN28202_n16991));
   INVx2_ASAP7_75t_SL FE_OFC98_n23036 (.Y(n24959),
	.A(n23036));
   INVxp67_ASAP7_75t_R FE_OFC96_n20344 (.Y(n20346),
	.A(n20344));
   INVx1_ASAP7_75t_SL FE_OFC94_n15466 (.Y(n15465),
	.A(n15466));
   INVxp67_ASAP7_75t_SL FE_OFC91_n13630 (.Y(n13629),
	.A(n13630));
   INVxp67_ASAP7_75t_L FE_OFC89_n23335 (.Y(n23187),
	.A(n23335));
   INVx1_ASAP7_75t_L FE_OFC88_n15187 (.Y(n14572),
	.A(n15187));
   INVx1_ASAP7_75t_SL FE_OFC79_n16507 (.Y(n16289),
	.A(n16507));
   INVxp67_ASAP7_75t_R FE_OFC78_n18988 (.Y(n18974),
	.A(n18988));
   INVx2_ASAP7_75t_L FE_OFC60_n22888 (.Y(n17780),
	.A(FE_OCPN27384_n22888));
   INVx2_ASAP7_75t_L FE_OFC53_n15774 (.Y(n15773),
	.A(FE_OCPN28065_n15774));
   INVx1_ASAP7_75t_SL FE_OFC52_n22957 (.Y(n18998),
	.A(n22957));
   INVx1_ASAP7_75t_SL FE_OFC50_n27056 (.Y(n25251),
	.A(n27056));
   INVx1_ASAP7_75t_SL FE_OFC49_n26749 (.Y(n26747),
	.A(n26749));
   INVx1_ASAP7_75t_L FE_OFC34_n15856 (.Y(n14855),
	.A(n15856));
   INVxp67_ASAP7_75t_SL FE_OFC33_n15061 (.Y(n13751),
	.A(n15061));
   BUFx2_ASAP7_75t_R FE_OFC22_n16125 (.Y(FE_OFN22_n16125),
	.A(FE_OFN19_n16125));
   BUFx2_ASAP7_75t_L FE_OFC2_ld_r (.Y(FE_OFN2_ld_r),
	.A(FE_OFN13_FE_DBTN0_ld_r));
   DFFHQNx1_ASAP7_75t_SRAM dcnt_reg_3_ (.QN(dcnt_3_),
	.CLK(CTS_39),
	.D(n928));
   DFFHQNx1_ASAP7_75t_SRAM dcnt_reg_2_ (.QN(dcnt_2_),
	.CLK(CTS_39),
	.D(n926));
   DFFHQNx1_ASAP7_75t_SRAM dcnt_reg_1_ (.QN(dcnt_1_),
	.CLK(CTS_39),
	.D(n924));
   DFFHQNx1_ASAP7_75t_SRAM done_reg (.QN(done),
	.CLK(CTS_39),
	.D(n923));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_127_ (.QN(text_in_r_127_),
	.CLK(CTS_39),
	.D(n921));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_126_ (.QN(text_in_r_126_),
	.CLK(CTS_39),
	.D(n919));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_125_ (.QN(text_in_r_125_),
	.CLK(CTS_39),
	.D(n917));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_124_ (.QN(text_in_r_124_),
	.CLK(CTS_39),
	.D(n915));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_123_ (.QN(text_in_r_123_),
	.CLK(CTS_39),
	.D(n913));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_122_ (.QN(text_in_r_122_),
	.CLK(CTS_39),
	.D(n911));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_121_ (.QN(text_in_r_121_),
	.CLK(CTS_39),
	.D(n909));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_120_ (.QN(text_in_r_120_),
	.CLK(CTS_39),
	.D(n907));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_119_ (.QN(text_in_r_119_),
	.CLK(CTS_38),
	.D(n905));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_118_ (.QN(text_in_r_118_),
	.CLK(CTS_38),
	.D(n903));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_117_ (.QN(text_in_r_117_),
	.CLK(CTS_38),
	.D(n901));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_116_ (.QN(text_in_r_116_),
	.CLK(CTS_38),
	.D(n899));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_115_ (.QN(text_in_r_115_),
	.CLK(CTS_38),
	.D(n897));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_114_ (.QN(text_in_r_114_),
	.CLK(CTS_38),
	.D(n895));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_113_ (.QN(text_in_r_113_),
	.CLK(CTS_37),
	.D(n893));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_112_ (.QN(text_in_r_112_),
	.CLK(CTS_38),
	.D(n891));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_111_ (.QN(text_in_r_111_),
	.CLK(CTS_38),
	.D(n889));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_110_ (.QN(text_in_r_110_),
	.CLK(CTS_38),
	.D(n887));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_109_ (.QN(text_in_r_109_),
	.CLK(CTS_39),
	.D(n885));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_108_ (.QN(text_in_r_108_),
	.CLK(CTS_38),
	.D(n883));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_107_ (.QN(text_in_r_107_),
	.CLK(CTS_39),
	.D(n881));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_106_ (.QN(text_in_r_106_),
	.CLK(CTS_33),
	.D(n879));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_105_ (.QN(text_in_r_105_),
	.CLK(CTS_38),
	.D(n877));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_104_ (.QN(text_in_r_104_),
	.CLK(CTS_39),
	.D(n875));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_103_ (.QN(text_in_r_103_),
	.CLK(CTS_38),
	.D(n873));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_102_ (.QN(text_in_r_102_),
	.CLK(CTS_38),
	.D(n871));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_101_ (.QN(text_in_r_101_),
	.CLK(CTS_38),
	.D(n869));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_100_ (.QN(text_in_r_100_),
	.CLK(CTS_38),
	.D(n867));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_99_ (.QN(text_in_r_99_),
	.CLK(CTS_38),
	.D(n865));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_98_ (.QN(text_in_r_98_),
	.CLK(CTS_38),
	.D(n863));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_97_ (.QN(text_in_r_97_),
	.CLK(CTS_38),
	.D(n861));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_96_ (.QN(text_in_r_96_),
	.CLK(CTS_38),
	.D(n859));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_95_ (.QN(text_in_r_95_),
	.CLK(CTS_32),
	.D(n857));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_94_ (.QN(text_in_r_94_),
	.CLK(CTS_32),
	.D(n855));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_93_ (.QN(text_in_r_93_),
	.CLK(CTS_32),
	.D(n853));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_92_ (.QN(text_in_r_92_),
	.CLK(CTS_32),
	.D(n851));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_91_ (.QN(text_in_r_91_),
	.CLK(CTS_32),
	.D(n849));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_90_ (.QN(text_in_r_90_),
	.CLK(CTS_32),
	.D(n847));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_89_ (.QN(text_in_r_89_),
	.CLK(CTS_32),
	.D(n845));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_88_ (.QN(text_in_r_88_),
	.CLK(CTS_32),
	.D(n843));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_87_ (.QN(text_in_r_87_),
	.CLK(CTS_31),
	.D(n841));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_86_ (.QN(text_in_r_86_),
	.CLK(CTS_32),
	.D(n839));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_85_ (.QN(text_in_r_85_),
	.CLK(CTS_32),
	.D(n837));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_84_ (.QN(text_in_r_84_),
	.CLK(CTS_36),
	.D(n835));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_83_ (.QN(text_in_r_83_),
	.CLK(CTS_36),
	.D(n833));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_82_ (.QN(text_in_r_82_),
	.CLK(CTS_32),
	.D(n831));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_81_ (.QN(text_in_r_81_),
	.CLK(CTS_31),
	.D(n829));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_80_ (.QN(text_in_r_80_),
	.CLK(CTS_31),
	.D(n827));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_79_ (.QN(text_in_r_79_),
	.CLK(CTS_36),
	.D(n825));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_78_ (.QN(text_in_r_78_),
	.CLK(CTS_36),
	.D(n823));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_77_ (.QN(text_in_r_77_),
	.CLK(CTS_36),
	.D(n821));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_76_ (.QN(text_in_r_76_),
	.CLK(CTS_36),
	.D(n819));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_75_ (.QN(text_in_r_75_),
	.CLK(CTS_32),
	.D(n817));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_74_ (.QN(text_in_r_74_),
	.CLK(CTS_36),
	.D(n815));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_73_ (.QN(text_in_r_73_),
	.CLK(CTS_36),
	.D(n813));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_72_ (.QN(text_in_r_72_),
	.CLK(CTS_36),
	.D(n811));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_71_ (.QN(text_in_r_71_),
	.CLK(CTS_33),
	.D(n809));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_70_ (.QN(text_in_r_70_),
	.CLK(CTS_33),
	.D(n807));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_69_ (.QN(text_in_r_69_),
	.CLK(CTS_32),
	.D(n805));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_68_ (.QN(text_in_r_68_),
	.CLK(CTS_31),
	.D(n803));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_67_ (.QN(text_in_r_67_),
	.CLK(CTS_31),
	.D(n801));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_66_ (.QN(text_in_r_66_),
	.CLK(CTS_31),
	.D(n799));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_65_ (.QN(text_in_r_65_),
	.CLK(CTS_31),
	.D(n797));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_64_ (.QN(text_in_r_64_),
	.CLK(CTS_31),
	.D(n795));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_63_ (.QN(text_in_r_63_),
	.CLK(CTS_34),
	.D(n793));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_62_ (.QN(text_in_r_62_),
	.CLK(CTS_34),
	.D(n791));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_61_ (.QN(text_in_r_61_),
	.CLK(CTS_34),
	.D(n789));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_60_ (.QN(text_in_r_60_),
	.CLK(CTS_33),
	.D(n787));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_59_ (.QN(text_in_r_59_),
	.CLK(CTS_34),
	.D(n785));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_58_ (.QN(text_in_r_58_),
	.CLK(CTS_34),
	.D(n783));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_57_ (.QN(text_in_r_57_),
	.CLK(CTS_34),
	.D(n781));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_56_ (.QN(text_in_r_56_),
	.CLK(CTS_34),
	.D(n779));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_55_ (.QN(text_in_r_55_),
	.CLK(CTS_33),
	.D(n777));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_54_ (.QN(text_in_r_54_),
	.CLK(CTS_33),
	.D(n775));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_53_ (.QN(text_in_r_53_),
	.CLK(CTS_33),
	.D(n773));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_52_ (.QN(text_in_r_52_),
	.CLK(CTS_33),
	.D(n771));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_51_ (.QN(text_in_r_51_),
	.CLK(CTS_33),
	.D(n769));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_50_ (.QN(text_in_r_50_),
	.CLK(CTS_34),
	.D(n767));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_49_ (.QN(text_in_r_49_),
	.CLK(CTS_33),
	.D(n765));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_48_ (.QN(text_in_r_48_),
	.CLK(CTS_33),
	.D(n763));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_47_ (.QN(text_in_r_47_),
	.CLK(CTS_34),
	.D(n761));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_46_ (.QN(text_in_r_46_),
	.CLK(CTS_33),
	.D(n759));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_45_ (.QN(text_in_r_45_),
	.CLK(CTS_34),
	.D(n757));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_44_ (.QN(text_in_r_44_),
	.CLK(CTS_34),
	.D(n755));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_43_ (.QN(text_in_r_43_),
	.CLK(CTS_34),
	.D(n753));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_42_ (.QN(text_in_r_42_),
	.CLK(CTS_34),
	.D(n751));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_41_ (.QN(text_in_r_41_),
	.CLK(CTS_34),
	.D(n749));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_40_ (.QN(text_in_r_40_),
	.CLK(CTS_34),
	.D(n747));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_39_ (.QN(text_in_r_39_),
	.CLK(CTS_33),
	.D(n745));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_38_ (.QN(text_in_r_38_),
	.CLK(CTS_33),
	.D(n743));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_37_ (.QN(text_in_r_37_),
	.CLK(CTS_33),
	.D(n741));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_36_ (.QN(text_in_r_36_),
	.CLK(CTS_33),
	.D(n739));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_35_ (.QN(text_in_r_35_),
	.CLK(CTS_33),
	.D(n737));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_34_ (.QN(text_in_r_34_),
	.CLK(CTS_34),
	.D(n735));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_33_ (.QN(text_in_r_33_),
	.CLK(CTS_33),
	.D(n733));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_32_ (.QN(text_in_r_32_),
	.CLK(CTS_33),
	.D(n731));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_31_ (.QN(text_in_r_31_),
	.CLK(CTS_37),
	.D(n729));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_30_ (.QN(text_in_r_30_),
	.CLK(CTS_37),
	.D(n727));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_29_ (.QN(text_in_r_29_),
	.CLK(CTS_37),
	.D(n725));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_28_ (.QN(text_in_r_28_),
	.CLK(CTS_37),
	.D(n723));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_27_ (.QN(text_in_r_27_),
	.CLK(CTS_37),
	.D(n721));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_26_ (.QN(text_in_r_26_),
	.CLK(CTS_37),
	.D(n719));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_25_ (.QN(text_in_r_25_),
	.CLK(CTS_37),
	.D(n717));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_24_ (.QN(text_in_r_24_),
	.CLK(CTS_37),
	.D(n715));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_23_ (.QN(text_in_r_23_),
	.CLK(CTS_36),
	.D(n713));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_22_ (.QN(text_in_r_22_),
	.CLK(CTS_37),
	.D(n711));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_21_ (.QN(text_in_r_21_),
	.CLK(CTS_36),
	.D(n709));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_20_ (.QN(text_in_r_20_),
	.CLK(CTS_36),
	.D(n707));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_19_ (.QN(text_in_r_19_),
	.CLK(CTS_36),
	.D(n705));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_18_ (.QN(text_in_r_18_),
	.CLK(CTS_36),
	.D(n703));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_17_ (.QN(text_in_r_17_),
	.CLK(CTS_36),
	.D(n701));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_16_ (.QN(text_in_r_16_),
	.CLK(CTS_36),
	.D(n699));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_15_ (.QN(text_in_r_15_),
	.CLK(CTS_36),
	.D(n697));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_14_ (.QN(text_in_r_14_),
	.CLK(CTS_36),
	.D(n695));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_13_ (.QN(text_in_r_13_),
	.CLK(CTS_36),
	.D(n693));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_12_ (.QN(text_in_r_12_),
	.CLK(CTS_36),
	.D(n691));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_11_ (.QN(text_in_r_11_),
	.CLK(CTS_36),
	.D(n689));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_10_ (.QN(text_in_r_10_),
	.CLK(CTS_36),
	.D(n687));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_9_ (.QN(text_in_r_9_),
	.CLK(CTS_36),
	.D(n685));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_8_ (.QN(text_in_r_8_),
	.CLK(CTS_36),
	.D(n683));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_7_ (.QN(text_in_r_7_),
	.CLK(CTS_36),
	.D(n681));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_6_ (.QN(text_in_r_6_),
	.CLK(CTS_37),
	.D(n679));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_5_ (.QN(text_in_r_5_),
	.CLK(CTS_37),
	.D(n677));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_4_ (.QN(text_in_r_4_),
	.CLK(CTS_37),
	.D(n675));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_3_ (.QN(text_in_r_3_),
	.CLK(CTS_37),
	.D(n673));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_2_ (.QN(text_in_r_2_),
	.CLK(CTS_37),
	.D(n671));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_1_ (.QN(text_in_r_1_),
	.CLK(CTS_37),
	.D(n669));
   DFFHQNx1_ASAP7_75t_SRAM text_in_r_reg_0_ (.QN(text_in_r_0_),
	.CLK(CTS_36),
	.D(n667));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_rcnt_reg_0_ (.QN(u0_r0_rcnt_0_),
	.CLK(CTS_39),
	.D(n666));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_rcnt_reg_1_ (.QN(u0_r0_rcnt_1_),
	.CLK(CTS_39),
	.D(n665));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_rcnt_reg_3_ (.QN(u0_r0_rcnt_3_),
	.CLK(CTS_39),
	.D(n663));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_24_ (.QN(u0_rcon_24_),
	.CLK(CTS_39),
	.D(n662));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_25_ (.QN(u0_rcon_25_),
	.CLK(CTS_39),
	.D(n661));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_26_ (.QN(u0_rcon_26_),
	.CLK(CTS_39),
	.D(n660));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_27_ (.QN(u0_rcon_27_),
	.CLK(CTS_39),
	.D(n659));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_28_ (.QN(u0_rcon_28_),
	.CLK(CTS_39),
	.D(n658));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_29_ (.QN(u0_rcon_29_),
	.CLK(CTS_39),
	.D(n657));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_30_ (.QN(u0_rcon_30_),
	.CLK(CTS_39),
	.D(n656));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_out_reg_31_ (.QN(u0_rcon_31_),
	.CLK(CTS_39),
	.D(n655));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__6_ (.QN(w3_6_),
	.CLK(CTS_31),
	.D(n649));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__22_ (.QN(w3_22_),
	.CLK(CTS_33),
	.D(n647));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__14_ (.QN(w3_14_),
	.CLK(CTS_31),
	.D(n644));
   DFFHQNx2_ASAP7_75t_L u0_w_reg_3__8_ (.QN(w3_8_),
	.CLK(CTS_31),
	.D(n632));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__24_ (.QN(w3_24_),
	.CLK(CTS_37),
	.D(n630));
   DFFHQNx2_ASAP7_75t_L u0_w_reg_3__0_ (.QN(w3_0_),
	.CLK(CTS_36),
	.D(n625));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__16_ (.QN(w2_16_),
	.CLK(CTS_33),
	.D(n622));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__16_ (.QN(w1_16_),
	.CLK(CTS_31),
	.D(n621));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__16_ (.QN(w0_16_),
	.CLK(CTS_31),
	.D(n620));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__9_ (.QN(w2_9_),
	.CLK(CTS_31),
	.D(n619));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__9_ (.QN(w1_9_),
	.CLK(CTS_31),
	.D(n618));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__9_ (.QN(w0_9_),
	.CLK(CTS_38),
	.D(n617));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__0_ (.QN(w2_0_),
	.CLK(CTS_33),
	.D(n616));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__0_ (.QN(w1_0_),
	.CLK(CTS_31),
	.D(n615));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__0_ (.QN(w0_0_),
	.CLK(CTS_37),
	.D(n614));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__25_ (.QN(w2_25_),
	.CLK(CTS_33),
	.D(n613));
   DFFHQNx2_ASAP7_75t_L u0_w_reg_1__25_ (.QN(w1_25_),
	.CLK(CTS_34),
	.D(n612));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__25_ (.QN(w0_25_),
	.CLK(CTS_39),
	.D(n611));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_2__17_ (.QN(w2_17_),
	.CLK(CTS_33),
	.D(n610));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__17_ (.QN(w1_17_),
	.CLK(CTS_31),
	.D(n609));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__17_ (.QN(w0_17_),
	.CLK(CTS_31),
	.D(n608));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__13_ (.QN(w2_13_),
	.CLK(CTS_33),
	.D(n607));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__13_ (.QN(w1_13_),
	.CLK(CTS_31),
	.D(n606));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__13_ (.QN(w0_13_),
	.CLK(CTS_38),
	.D(n605));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__3_ (.QN(w2_3_),
	.CLK(CTS_33),
	.D(n604));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__3_ (.QN(w1_3_),
	.CLK(CTS_33),
	.D(n603));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__3_ (.QN(w0_3_),
	.CLK(CTS_38),
	.D(n602));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__24_ (.QN(w2_24_),
	.CLK(CTS_34),
	.D(n601));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__24_ (.QN(w1_24_),
	.CLK(CTS_34),
	.D(n600));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__24_ (.QN(w0_24_),
	.CLK(CTS_39),
	.D(n599));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_2__19_ (.QN(w2_19_),
	.CLK(CTS_33),
	.D(n598));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__19_ (.QN(w1_19_),
	.CLK(CTS_31),
	.D(n597));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__19_ (.QN(w0_19_),
	.CLK(CTS_31),
	.D(n596));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__8_ (.QN(w2_8_),
	.CLK(CTS_34),
	.D(n595));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__8_ (.QN(w1_8_),
	.CLK(CTS_31),
	.D(n594));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__8_ (.QN(w0_8_),
	.CLK(CTS_38),
	.D(n593));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__1_ (.QN(w2_1_),
	.CLK(CTS_33),
	.D(n592));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__1_ (.QN(w1_1_),
	.CLK(CTS_31),
	.D(n591));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__1_ (.QN(w0_1_),
	.CLK(CTS_38),
	.D(n590));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__26_ (.QN(w2_26_),
	.CLK(CTS_33),
	.D(n589));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__26_ (.QN(w1_26_),
	.CLK(CTS_33),
	.D(n588));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__26_ (.QN(w0_26_),
	.CLK(CTS_39),
	.D(n587));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__18_ (.QN(w2_18_),
	.CLK(CTS_34),
	.D(n586));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__18_ (.QN(w1_18_),
	.CLK(CTS_32),
	.D(n585));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__18_ (.QN(w0_18_),
	.CLK(CTS_31),
	.D(n584));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__10_ (.QN(w2_10_),
	.CLK(CTS_34),
	.D(n583));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__10_ (.QN(w1_10_),
	.CLK(CTS_31),
	.D(n582));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__10_ (.QN(w0_10_),
	.CLK(CTS_38),
	.D(n581));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__2_ (.QN(w2_2_),
	.CLK(CTS_33),
	.D(n580));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__2_ (.QN(w1_2_),
	.CLK(CTS_31),
	.D(n579));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__2_ (.QN(w0_2_),
	.CLK(CTS_38),
	.D(n578));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__27_ (.QN(w2_27_),
	.CLK(CTS_33),
	.D(n577));
   DFFHQNx2_ASAP7_75t_SRAM u0_w_reg_1__27_ (.QN(w1_27_),
	.CLK(CTS_34),
	.D(n576));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__27_ (.QN(w0_27_),
	.CLK(CTS_39),
	.D(n575));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_2__20_ (.QN(w2_20_),
	.CLK(CTS_31),
	.D(n574));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__20_ (.QN(w1_20_),
	.CLK(CTS_31),
	.D(n573));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__20_ (.QN(w0_20_),
	.CLK(CTS_31),
	.D(n572));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__12_ (.QN(w2_12_),
	.CLK(CTS_33),
	.D(n571));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__12_ (.QN(w1_12_),
	.CLK(CTS_31),
	.D(n570));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__12_ (.QN(w0_12_),
	.CLK(CTS_38),
	.D(n569));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__4_ (.QN(w2_4_),
	.CLK(CTS_33),
	.D(n568));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__4_ (.QN(w1_4_),
	.CLK(CTS_31),
	.D(n567));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__4_ (.QN(w0_4_),
	.CLK(CTS_37),
	.D(n566));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__28_ (.QN(w2_28_),
	.CLK(CTS_33),
	.D(n565));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__28_ (.QN(w1_28_),
	.CLK(CTS_33),
	.D(n564));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__28_ (.QN(w0_28_),
	.CLK(CTS_39),
	.D(n563));
   DFFHQNx2_ASAP7_75t_R u0_w_reg_2__21_ (.QN(w2_21_),
	.CLK(CTS_33),
	.D(n562));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__21_ (.QN(w1_21_),
	.CLK(CTS_32),
	.D(n561));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__21_ (.QN(w0_21_),
	.CLK(CTS_31),
	.D(n560));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__14_ (.QN(w2_14_),
	.CLK(CTS_33),
	.D(n559));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__14_ (.QN(w1_14_),
	.CLK(CTS_31),
	.D(n558));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__14_ (.QN(w0_14_),
	.CLK(CTS_38),
	.D(n557));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__5_ (.QN(w2_5_),
	.CLK(CTS_33),
	.D(n556));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__5_ (.QN(w1_5_),
	.CLK(CTS_31),
	.D(n555));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__5_ (.QN(w0_5_),
	.CLK(CTS_38),
	.D(n554));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_2__29_ (.QN(w2_29_),
	.CLK(CTS_33),
	.D(n553));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__29_ (.QN(w1_29_),
	.CLK(CTS_33),
	.D(n552));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__29_ (.QN(w0_29_),
	.CLK(CTS_39),
	.D(n551));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__22_ (.QN(w2_22_),
	.CLK(CTS_33),
	.D(n550));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__22_ (.QN(w1_22_),
	.CLK(CTS_32),
	.D(n549));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__22_ (.QN(w0_22_),
	.CLK(CTS_31),
	.D(n548));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__11_ (.QN(w2_11_),
	.CLK(CTS_33),
	.D(n547));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__11_ (.QN(w1_11_),
	.CLK(CTS_31),
	.D(n546));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__11_ (.QN(w0_11_),
	.CLK(CTS_38),
	.D(n545));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__6_ (.QN(w2_6_),
	.CLK(CTS_31),
	.D(n544));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__6_ (.QN(w1_6_),
	.CLK(CTS_33),
	.D(n543));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__6_ (.QN(w0_6_),
	.CLK(CTS_38),
	.D(n542));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_2__30_ (.QN(w2_30_),
	.CLK(CTS_38),
	.D(n541));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__30_ (.QN(w1_30_),
	.CLK(CTS_38),
	.D(n540));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__30_ (.QN(w0_30_),
	.CLK(CTS_39),
	.D(n539));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_2__23_ (.QN(w2_23_),
	.CLK(CTS_33),
	.D(n538));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_1__23_ (.QN(w1_23_),
	.CLK(CTS_31),
	.D(n537));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__23_ (.QN(w0_23_),
	.CLK(CTS_31),
	.D(n536));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__15_ (.QN(w2_15_),
	.CLK(CTS_33),
	.D(n535));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__15_ (.QN(w1_15_),
	.CLK(CTS_31),
	.D(n534));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__15_ (.QN(w0_15_),
	.CLK(CTS_38),
	.D(n533));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_2__7_ (.QN(w2_7_),
	.CLK(CTS_31),
	.D(n532));
   DFFHQNx1_ASAP7_75t_R u0_w_reg_1__7_ (.QN(w1_7_),
	.CLK(CTS_31),
	.D(n531));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__7_ (.QN(w0_7_),
	.CLK(CTS_38),
	.D(n530));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_2__31_ (.QN(w2_31_),
	.CLK(CTS_33),
	.D(n529));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_1__31_ (.QN(w1_31_),
	.CLK(CTS_33),
	.D(n528));
   DFFHQNx1_ASAP7_75t_SRAM u0_w_reg_0__31_ (.QN(w0_31_),
	.CLK(CTS_39),
	.D(n527));
   DFFHQNx1_ASAP7_75t_L sa30_reg_7_ (.QN(sa30_7_),
	.CLK(CTS_38),
	.D(n525));
   DFFHQNx2_ASAP7_75t_L sa31_reg_7_ (.QN(sa31_7_),
	.CLK(CTS_33),
	.D(n524));
   DFFHQNx2_ASAP7_75t_L sa32_reg_7_ (.QN(sa32_7_),
	.CLK(CTS_33),
	.D(n523));
   DFFHQNx1_ASAP7_75t_L sa33_reg_7_ (.QN(sa33_7_),
	.CLK(CTS_36),
	.D(n522));
   DFFHQNx1_ASAP7_75t_L sa30_reg_6_ (.QN(sa30_6_),
	.CLK(CTS_33),
	.D(n521));
   DFFHQNx1_ASAP7_75t_L sa21_reg_7_ (.QN(sa21_7_),
	.CLK(CTS_36),
	.D(n520));
   DFFHQNx1_ASAP7_75t_L sa22_reg_7_ (.QN(sa22_7_),
	.CLK(CTS_33),
	.D(n516));
   DFFHQNx1_ASAP7_75t_L sa31_reg_6_ (.QN(sa31_6_),
	.CLK(CTS_33),
	.D(n511));
   DFFHQNx1_ASAP7_75t_R sa12_reg_6_ (.QN(sa12_6_),
	.CLK(CTS_33),
	.D(n510));
   DFFHQNx1_ASAP7_75t_L sa22_reg_6_ (.QN(sa22_6_),
	.CLK(CTS_33),
	.D(n507));
   DFFHQNx1_ASAP7_75t_L sa10_reg_7_ (.QN(sa10_7_),
	.CLK(CTS_38),
	.D(n506));
   DFFHQNx1_ASAP7_75t_L sa33_reg_6_ (.QN(sa33_6_),
	.CLK(CTS_37),
	.D(n505));
   DFFHQNx2_ASAP7_75t_L sa32_reg_6_ (.QN(sa32_6_),
	.CLK(CTS_33),
	.D(n503));
   DFFHQNx2_ASAP7_75t_L sa13_reg_6_ (.QN(sa13_6_),
	.CLK(CTS_37),
	.D(n502));
   DFFHQNx1_ASAP7_75t_L sa02_reg_7_ (.QN(sa02_7_),
	.CLK(CTS_34),
	.D(n501));
   DFFHQNx1_ASAP7_75t_L sa21_reg_6_ (.QN(sa21_6_),
	.CLK(CTS_36),
	.D(n496));
   DFFHQNx1_ASAP7_75t_L sa13_reg_7_ (.QN(sa13_7_),
	.CLK(CTS_36),
	.D(n495));
   DFFHQNx2_ASAP7_75t_L sa01_reg_7_ (.QN(sa01_7_),
	.CLK(CTS_32),
	.D(n493));
   DFFHQNx2_ASAP7_75t_L sa01_reg_6_ (.QN(sa01_6_),
	.CLK(CTS_32),
	.D(n490));
   DFFHQNx1_ASAP7_75t_L sa11_reg_6_ (.QN(sa11_6_),
	.CLK(CTS_36),
	.D(n489));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_6_ (.QN(sa20_6_),
	.CLK(CTS_38),
	.D(n488));
   DFFHQNx2_ASAP7_75t_L sa11_reg_7_ (.QN(sa11_7_),
	.CLK(CTS_33),
	.D(n486));
   DFFHQNx2_ASAP7_75t_L sa00_reg_6_ (.QN(sa00_6_),
	.CLK(CTS_39),
	.D(n485));
   DFFHQNx2_ASAP7_75t_L sa02_reg_6_ (.QN(sa02_6_),
	.CLK(CTS_34),
	.D(n473));
   DFFHQNx1_ASAP7_75t_L sa03_reg_7_ (.QN(sa03_7_),
	.CLK(CTS_37),
	.D(n460));
   DFFHQNx2_ASAP7_75t_L sa03_reg_6_ (.QN(sa03_6_),
	.CLK(CTS_37),
	.D(n445));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_34_ (.QN(text_out_34_),
	.CLK(CTS_34),
	.D(n439));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_36_ (.QN(text_out_36_),
	.CLK(CTS_34),
	.D(n438));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_35_ (.QN(text_out_35_),
	.CLK(CTS_34),
	.D(n437));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_32_ (.QN(text_out_32_),
	.CLK(CTS_34),
	.D(n436));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_33_ (.QN(text_out_33_),
	.CLK(CTS_34),
	.D(n435));
   DFFHQNx1_ASAP7_75t_SL sa33_reg_1_ (.QN(sa33_1_),
	.CLK(CTS_38),
	.D(FE_OCPN29565_n432));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_12_ (.QN(text_out_12_),
	.CLK(CTS_36),
	.D(n423));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_9_ (.QN(text_out_9_),
	.CLK(CTS_36),
	.D(n422));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_8_ (.QN(text_out_8_),
	.CLK(CTS_36),
	.D(n421));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_10_ (.QN(text_out_10_),
	.CLK(CTS_36),
	.D(n420));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_11_ (.QN(text_out_11_),
	.CLK(CTS_36),
	.D(n419));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_3_ (.QN(text_out_3_),
	.CLK(CTS_36),
	.D(n415));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_0_ (.QN(text_out_0_),
	.CLK(CTS_36),
	.D(n414));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_1_ (.QN(text_out_1_),
	.CLK(CTS_36),
	.D(n413));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_2_ (.QN(text_out_2_),
	.CLK(CTS_37),
	.D(n412));
   DFFHQNx2_ASAP7_75t_SL sa02_reg_1_ (.QN(sa02_1_),
	.CLK(CTS_34),
	.D(n409));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_80_ (.QN(text_out_80_),
	.CLK(CTS_32),
	.D(n407));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_81_ (.QN(text_out_81_),
	.CLK(CTS_32),
	.D(n406));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_86_ (.QN(text_out_86_),
	.CLK(CTS_32),
	.D(n404));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_84_ (.QN(text_out_84_),
	.CLK(CTS_32),
	.D(n403));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_82_ (.QN(text_out_82_),
	.CLK(CTS_32),
	.D(n402));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_83_ (.QN(text_out_83_),
	.CLK(CTS_32),
	.D(n400));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_91_ (.QN(text_out_91_),
	.CLK(CTS_32),
	.D(n398));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_88_ (.QN(text_out_88_),
	.CLK(CTS_32),
	.D(n397));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_93_ (.QN(text_out_93_),
	.CLK(CTS_32),
	.D(n396));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_89_ (.QN(text_out_89_),
	.CLK(CTS_32),
	.D(n395));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_90_ (.QN(text_out_90_),
	.CLK(CTS_32),
	.D(n394));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_79_ (.QN(text_out_79_),
	.CLK(CTS_32),
	.D(n389));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_73_ (.QN(text_out_73_),
	.CLK(CTS_32),
	.D(n388));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_72_ (.QN(text_out_72_),
	.CLK(CTS_32),
	.D(n387));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_74_ (.QN(text_out_74_),
	.CLK(CTS_36),
	.D(n385));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_75_ (.QN(text_out_75_),
	.CLK(CTS_36),
	.D(n384));
   DFFHQNx1_ASAP7_75t_SL sa33_reg_0_ (.QN(sa33_0_),
	.CLK(CTS_38),
	.D(FE_OCPN29556_n383));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_101_ (.QN(text_out_101_),
	.CLK(CTS_39),
	.D(n382));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_100_ (.QN(text_out_100_),
	.CLK(CTS_38),
	.D(n381));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_99_ (.QN(text_out_99_),
	.CLK(CTS_38),
	.D(n380));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_96_ (.QN(text_out_96_),
	.CLK(CTS_38),
	.D(n379));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_97_ (.QN(text_out_97_),
	.CLK(CTS_38),
	.D(n378));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_98_ (.QN(text_out_98_),
	.CLK(CTS_38),
	.D(n377));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_47_ (.QN(text_out_47_),
	.CLK(CTS_34),
	.D(n374));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_41_ (.QN(text_out_41_),
	.CLK(CTS_34),
	.D(n373));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_45_ (.QN(text_out_45_),
	.CLK(CTS_34),
	.D(n372));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_40_ (.QN(text_out_40_),
	.CLK(CTS_34),
	.D(n371));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_111_ (.QN(text_out_111_),
	.CLK(CTS_39),
	.D(n369));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_107_ (.QN(text_out_107_),
	.CLK(CTS_39),
	.D(n368));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_104_ (.QN(text_out_104_),
	.CLK(CTS_38),
	.D(n367));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_106_ (.QN(text_out_106_),
	.CLK(CTS_38),
	.D(n366));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_109_ (.QN(text_out_109_),
	.CLK(CTS_39),
	.D(n365));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_105_ (.QN(text_out_105_),
	.CLK(CTS_38),
	.D(n364));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_43_ (.QN(text_out_43_),
	.CLK(CTS_34),
	.D(n363));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_67_ (.QN(text_out_67_),
	.CLK(CTS_31),
	.D(n361));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_64_ (.QN(text_out_64_),
	.CLK(CTS_31),
	.D(n360));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_117_ (.QN(text_out_117_),
	.CLK(CTS_38),
	.D(n358));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_116_ (.QN(text_out_116_),
	.CLK(CTS_38),
	.D(n357));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_112_ (.QN(text_out_112_),
	.CLK(CTS_38),
	.D(n356));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_115_ (.QN(text_out_115_),
	.CLK(CTS_38),
	.D(n354));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_113_ (.QN(text_out_113_),
	.CLK(CTS_38),
	.D(n353));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_120_ (.QN(text_out_120_),
	.CLK(CTS_39),
	.D(n351));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_114_ (.QN(text_out_114_),
	.CLK(CTS_38),
	.D(n349));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_65_ (.QN(text_out_65_),
	.CLK(CTS_32),
	.D(n348));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_66_ (.QN(text_out_66_),
	.CLK(CTS_32),
	.D(n347));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_71_ (.QN(text_out_71_),
	.CLK(CTS_31),
	.D(n346));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_121_ (.QN(text_out_121_),
	.CLK(CTS_39),
	.D(n345));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_19_ (.QN(text_out_19_),
	.CLK(CTS_37),
	.D(n343));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_20_ (.QN(text_out_20_),
	.CLK(CTS_37),
	.D(n342));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_16_ (.QN(text_out_16_),
	.CLK(CTS_37),
	.D(n341));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_18_ (.QN(text_out_18_),
	.CLK(CTS_37),
	.D(n339));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_17_ (.QN(text_out_17_),
	.CLK(CTS_37),
	.D(n338));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_25_ (.QN(text_out_25_),
	.CLK(CTS_37),
	.D(n336));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_24_ (.QN(text_out_24_),
	.CLK(CTS_37),
	.D(n335));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_48_ (.QN(text_out_48_),
	.CLK(CTS_34),
	.D(n333));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_49_ (.QN(text_out_49_),
	.CLK(CTS_34),
	.D(n331));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_50_ (.QN(text_out_50_),
	.CLK(CTS_34),
	.D(n330));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_56_ (.QN(text_out_56_),
	.CLK(CTS_34),
	.D(n328));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_57_ (.QN(text_out_57_),
	.CLK(CTS_34),
	.D(n327));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_59_ (.QN(text_out_59_),
	.CLK(CTS_34),
	.D(n326));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_51_ (.QN(text_out_51_),
	.CLK(CTS_33),
	.D(n325));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_122_ (.QN(text_out_122_),
	.CLK(CTS_39),
	.D(n324));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_123_ (.QN(text_out_123_),
	.CLK(CTS_39),
	.D(n323));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_126_ (.QN(text_out_126_),
	.CLK(CTS_39),
	.D(n322));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_125_ (.QN(text_out_125_),
	.CLK(CTS_39),
	.D(n321));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_21_ (.QN(text_out_21_),
	.CLK(CTS_37),
	.D(n320));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_61_ (.QN(text_out_61_),
	.CLK(CTS_34),
	.D(n319));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_26_ (.QN(text_out_26_),
	.CLK(CTS_37),
	.D(n318));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_27_ (.QN(text_out_27_),
	.CLK(CTS_37),
	.D(n317));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_29_ (.QN(text_out_29_),
	.CLK(CTS_37),
	.D(n316));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_7_ (.QN(text_out_7_),
	.CLK(CTS_36),
	.D(n315));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_58_ (.QN(text_out_58_),
	.CLK(CTS_34),
	.D(n314));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_52_ (.QN(text_out_52_),
	.CLK(CTS_33),
	.D(n313));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_4_ (.QN(text_out_4_),
	.CLK(CTS_36),
	.D(n312));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_53_ (.QN(text_out_53_),
	.CLK(CTS_33),
	.D(n311));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_55_ (.QN(text_out_55_),
	.CLK(CTS_33),
	.D(n310));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_68_ (.QN(text_out_68_),
	.CLK(CTS_32),
	.D(n309));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_103_ (.QN(text_out_103_),
	.CLK(CTS_38),
	.D(n308));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_13_ (.QN(text_out_13_),
	.CLK(CTS_36),
	.D(n307));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_37_ (.QN(text_out_37_),
	.CLK(CTS_33),
	.D(n306));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_92_ (.QN(text_out_92_),
	.CLK(CTS_32),
	.D(n305));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_76_ (.QN(text_out_76_),
	.CLK(CTS_32),
	.D(n304));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_28_ (.QN(text_out_28_),
	.CLK(CTS_37),
	.D(n303));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_30_ (.QN(text_out_30_),
	.CLK(CTS_37),
	.D(n302));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_31_ (.QN(text_out_31_),
	.CLK(CTS_37),
	.D(n301));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_23_ (.QN(text_out_23_),
	.CLK(CTS_37),
	.D(n300));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_39_ (.QN(text_out_39_),
	.CLK(CTS_34),
	.D(n299));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_85_ (.QN(text_out_85_),
	.CLK(CTS_32),
	.D(n298));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_42_ (.QN(text_out_42_),
	.CLK(CTS_34),
	.D(n297));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_127_ (.QN(text_out_127_),
	.CLK(CTS_39),
	.D(n296));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_124_ (.QN(text_out_124_),
	.CLK(CTS_39),
	.D(n295));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_94_ (.QN(text_out_94_),
	.CLK(CTS_32),
	.D(n294));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_95_ (.QN(text_out_95_),
	.CLK(CTS_32),
	.D(n293));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_44_ (.QN(text_out_44_),
	.CLK(CTS_34),
	.D(n292));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_22_ (.QN(text_out_22_),
	.CLK(CTS_37),
	.D(n291));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_108_ (.QN(text_out_108_),
	.CLK(CTS_38),
	.D(n290));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_63_ (.QN(text_out_63_),
	.CLK(CTS_34),
	.D(n289));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_60_ (.QN(text_out_60_),
	.CLK(CTS_33),
	.D(n288));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_77_ (.QN(text_out_77_),
	.CLK(CTS_36),
	.D(n287));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_78_ (.QN(text_out_78_),
	.CLK(CTS_32),
	.D(n286));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_5_ (.QN(text_out_5_),
	.CLK(CTS_36),
	.D(n285));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_62_ (.QN(text_out_62_),
	.CLK(CTS_34),
	.D(n284));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_54_ (.QN(text_out_54_),
	.CLK(CTS_34),
	.D(n283));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_6_ (.QN(text_out_6_),
	.CLK(CTS_36),
	.D(n282));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_46_ (.QN(text_out_46_),
	.CLK(CTS_33),
	.D(n281));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_102_ (.QN(text_out_102_),
	.CLK(CTS_38),
	.D(n280));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_14_ (.QN(text_out_14_),
	.CLK(CTS_36),
	.D(n279));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_110_ (.QN(text_out_110_),
	.CLK(CTS_38),
	.D(n278));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_69_ (.QN(text_out_69_),
	.CLK(CTS_32),
	.D(n277));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_118_ (.QN(text_out_118_),
	.CLK(CTS_38),
	.D(n276));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_70_ (.QN(text_out_70_),
	.CLK(CTS_31),
	.D(n275));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_87_ (.QN(text_out_87_),
	.CLK(CTS_32),
	.D(n274));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_38_ (.QN(text_out_38_),
	.CLK(CTS_33),
	.D(n273));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_15_ (.QN(text_out_15_),
	.CLK(CTS_36),
	.D(n272));
   DFFHQNx1_ASAP7_75t_SRAM text_out_reg_119_ (.QN(text_out_119_),
	.CLK(CTS_38),
	.D(n271));
   DFFHQNx1_ASAP7_75t_SRAM dcnt_reg_0_ (.QN(dcnt_0_),
	.CLK(CTS_39),
	.D(n930));
   DFFHQNx1_ASAP7_75t_SRAM u0_r0_rcnt_reg_2_ (.QN(u0_r0_rcnt_2_),
	.CLK(CTS_39),
	.D(n664));
   DFFHQNx2_ASAP7_75t_SL u0_w_reg_3__21_ (.QN(w3_21_),
	.CLK(CTS_39),
	.D(n643));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_3__2_ (.QN(w3_2_),
	.CLK(CTS_36),
	.D(n637));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__10_ (.QN(w3_10_),
	.CLK(CTS_31),
	.D(n636));
   DFFHQNx2_ASAP7_75t_SL u0_w_reg_3__18_ (.QN(w3_18_),
	.CLK(CTS_39),
	.D(n635));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_3__26_ (.QN(w3_26_),
	.CLK(CTS_37),
	.D(n634));
   DFFHQNx1_ASAP7_75t_SL sa13_reg_4_ (.QN(sa13_4_),
	.CLK(CTS_31),
	.D(n517));
   DFFHQNx3_ASAP7_75t_L sa20_reg_7_ (.QN(sa20_7_),
	.CLK(CTS_33),
	.D(n504));
   DFFHQNx1_ASAP7_75t_L sa23_reg_6_ (.QN(sa23_6_),
	.CLK(CTS_36),
	.D(n499));
   DFFHQNx1_ASAP7_75t_SL sa12_reg_3_ (.QN(sa12_3_),
	.CLK(CTS_32),
	.D(FE_OCPN29417_n455));
   DFFHQNx1_ASAP7_75t_SL sa00_reg_4_ (.QN(sa00_4_),
	.CLK(CTS_39),
	.D(n452));
   DFFHQNx2_ASAP7_75t_L sa10_reg_6_ (.QN(sa10_6_),
	.CLK(CTS_38),
	.D(n446));
   DFFHQNx1_ASAP7_75t_SL sa03_reg_4_ (.QN(sa03_4_),
	.CLK(CTS_37),
	.D(n429));
   DFFHQNx1_ASAP7_75t_SL sa13_reg_3_ (.QN(sa13_3_),
	.CLK(CTS_31),
	.D(FE_OCPN29256_n418));
   DFFHQNx1_ASAP7_75t_SL sa01_reg_5_ (.QN(sa01_5_),
	.CLK(CTS_32),
	.D(n454));
   DFFHQNx1_ASAP7_75t_SL sa12_reg_5_ (.QN(sa12_5_),
	.CLK(CTS_32),
	.D(n491));
   DFFHQNx1_ASAP7_75t_SL sa10_reg_0_ (.QN(sa10_0_),
	.CLK(CTS_37),
	.D(n350));
   DFFHQNx1_ASAP7_75t_SL sa21_reg_0_ (.QN(sa21_0_),
	.CLK(CTS_36),
	.D(n430));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_5_ (.QN(sa20_5_),
	.CLK(CTS_33),
	.D(n466));
   DFFHQNx1_ASAP7_75t_L sa32_reg_4_ (.QN(sa32_4_),
	.CLK(CTS_36),
	.D(n500));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_1_ (.QN(sa20_1_),
	.CLK(CTS_33),
	.D(n456));
   DFFHQNx1_ASAP7_75t_SL sa30_reg_1_ (.QN(sa30_1_),
	.CLK(CTS_31),
	.D(n431));
   DFFHQNx1_ASAP7_75t_SL sa01_reg_3_ (.QN(sa01_3_),
	.CLK(CTS_32),
	.D(n399));
   DFFHQNx1_ASAP7_75t_SL sa03_reg_1_ (.QN(sa03_1_),
	.CLK(CTS_37),
	.D(n337));
   DFFHQNx2_ASAP7_75t_L sa12_reg_7_ (.QN(sa12_7_),
	.CLK(CTS_33),
	.D(n487));
   DFFHQNx1_ASAP7_75t_SL sa31_reg_5_ (.QN(sa31_5_),
	.CLK(CTS_34),
	.D(FE_OCPN29355_n492));
   DFFHQNx1_ASAP7_75t_SL sa21_reg_1_ (.QN(sa21_1_),
	.CLK(CTS_36),
	.D(n433));
   DFFHQNx1_ASAP7_75t_SL sa11_reg_0_ (.QN(sa11_0_),
	.CLK(CTS_31),
	.D(n453));
   DFFHQNx1_ASAP7_75t_SL sa21_reg_3_ (.QN(sa21_3_),
	.CLK(CTS_36),
	.D(n463));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_4_ (.QN(sa20_4_),
	.CLK(CTS_33),
	.D(n515));
   DFFHQNx1_ASAP7_75t_SL sa23_reg_3_ (.QN(sa23_3_),
	.CLK(CTS_36),
	.D(n442));
   DFFHQNx2_ASAP7_75t_SL sa11_reg_3_ (.QN(sa11_3_),
	.CLK(CTS_31),
	.D(n359));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__1_ (.QN(w3_1_),
	.CLK(CTS_38),
	.D(n633));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__5_ (.QN(w3_5_),
	.CLK(CTS_31),
	.D(n645));
   DFFHQNx1_ASAP7_75t_SRAM ld_r_reg (.QN(ld_r),
	.CLK(CTS_34),
	.D(FE_OFN28459_ld));
   DFFHQNx1_ASAP7_75t_SL sa31_reg_4_ (.QN(sa31_4_),
	.CLK(CTS_33),
	.D(n508));
   DFFHQNx2_ASAP7_75t_SL sa21_reg_2_ (.QN(sa21_2_),
	.CLK(CTS_36),
	.D(n424));
   DFFHQNx1_ASAP7_75t_SL sa00_reg_0_ (.QN(sa00_0_),
	.CLK(CTS_39),
	.D(n355));
   DFFHQNx2_ASAP7_75t_SL sa30_reg_5_ (.QN(sa30_5_),
	.CLK(CTS_33),
	.D(n482));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__17_ (.QN(w3_17_),
	.CLK(CTS_39),
	.D(n627));
   DFFHQNx1_ASAP7_75t_SL sa01_reg_0_ (.QN(sa01_0_),
	.CLK(CTS_32),
	.D(n509));
   DFFHQNx1_ASAP7_75t_SL sa02_reg_0_ (.QN(sa02_0_),
	.CLK(CTS_34),
	.D(n332));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_3__31_ (.QN(w3_31_),
	.CLK(CTS_37),
	.D(n654));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__28_ (.QN(w3_28_),
	.CLK(CTS_37),
	.D(n642));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__13_ (.QN(w3_13_),
	.CLK(CTS_36),
	.D(n628));
   DFFHQNx1_ASAP7_75t_SL sa11_reg_4_ (.QN(sa11_4_),
	.CLK(CTS_31),
	.D(n498));
   DFFHQNx1_ASAP7_75t_SL sa32_reg_5_ (.QN(sa32_5_),
	.CLK(CTS_31),
	.D(n475));
   DFFHQNx1_ASAP7_75t_SL sa02_reg_5_ (.QN(sa02_5_),
	.CLK(CTS_34),
	.D(n472));
   DFFHQNx1_ASAP7_75t_SL sa32_reg_3_ (.QN(sa32_3_),
	.CLK(CTS_31),
	.D(n471));
   DFFHQNx1_ASAP7_75t_SL sa22_reg_3_ (.QN(sa22_3_),
	.CLK(CTS_34),
	.D(n467));
   DFFHQNx1_ASAP7_75t_SL sa32_reg_2_ (.QN(sa32_2_),
	.CLK(CTS_31),
	.D(n465));
   DFFHQNx1_ASAP7_75t_SL sa33_reg_3_ (.QN(sa33_3_),
	.CLK(CTS_37),
	.D(n459));
   DFFHQNx1_ASAP7_75t_SL sa31_reg_0_ (.QN(sa31_0_),
	.CLK(CTS_34),
	.D(FE_OCPN29364_n448));
   DFFHQNx1_ASAP7_75t_SL sa22_reg_2_ (.QN(sa22_2_),
	.CLK(CTS_34),
	.D(n447));
   DFFHQNx1_ASAP7_75t_SL sa03_reg_5_ (.QN(sa03_5_),
	.CLK(CTS_37),
	.D(n444));
   DFFHQNx1_ASAP7_75t_SL sa01_reg_4_ (.QN(sa01_4_),
	.CLK(CTS_32),
	.D(n441));
   DFFHQNx1_ASAP7_75t_SL sa12_reg_1_ (.QN(sa12_1_),
	.CLK(CTS_32),
	.D(n434));
   DFFHQNx1_ASAP7_75t_SL sa22_reg_0_ (.QN(sa22_0_),
	.CLK(CTS_34),
	.D(n427));
   DFFHQNx1_ASAP7_75t_SL sa32_reg_0_ (.QN(sa32_0_),
	.CLK(CTS_31),
	.D(FE_OCPN29589_n426));
   DFFHQNx2_ASAP7_75t_SL sa32_reg_1_ (.QN(sa32_1_),
	.CLK(CTS_36),
	.D(n416));
   DFFHQNx2_ASAP7_75t_SL sa01_reg_1_ (.QN(sa01_1_),
	.CLK(CTS_32),
	.D(n405));
   DFFHQNx1_ASAP7_75t_SL sa23_reg_0_ (.QN(sa23_0_),
	.CLK(CTS_36),
	.D(n390));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_0_ (.QN(sa20_0_),
	.CLK(CTS_33),
	.D(n375));
   DFFHQNx1_ASAP7_75t_SL sa22_reg_1_ (.QN(sa22_1_),
	.CLK(CTS_34),
	.D(n370));
   DFFHQNx1_ASAP7_75t_SL sa00_reg_1_ (.QN(sa00_1_),
	.CLK(CTS_39),
	.D(n352));
   DFFHQNx1_ASAP7_75t_SL sa13_reg_0_ (.QN(sa13_0_),
	.CLK(CTS_31),
	.D(FE_OCPN27306_n334));
   DFFHQNx1_ASAP7_75t_SL sa10_reg_1_ (.QN(sa10_1_),
	.CLK(CTS_37),
	.D(n344));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__12_ (.QN(w3_12_),
	.CLK(CTS_31),
	.D(n640));
   DFFHQNx1_ASAP7_75t_L u0_w_reg_3__16_ (.QN(w3_16_),
	.CLK(CTS_33),
	.D(n623));
   DFFHQNx2_ASAP7_75t_L sa00_reg_7_ (.QN(sa00_7_),
	.CLK(CTS_39),
	.D(n526));
   DFFHQNx1_ASAP7_75t_SL sa22_reg_5_ (.QN(sa22_5_),
	.CLK(CTS_33),
	.D(n480));
   DFFHQNx1_ASAP7_75t_SL sa21_reg_4_ (.QN(sa21_4_),
	.CLK(CTS_36),
	.D(n518));
   DFFHQNx1_ASAP7_75t_SL sa31_reg_2_ (.QN(sa31_2_),
	.CLK(CTS_33),
	.D(n481));
   DFFHQNx1_ASAP7_75t_SL sa02_reg_4_ (.QN(sa02_4_),
	.CLK(CTS_34),
	.D(n468));
   DFFHQNx1_ASAP7_75t_SL sa33_reg_5_ (.QN(sa33_5_),
	.CLK(CTS_38),
	.D(FE_OCPN29588_n457));
   DFFHQNx1_ASAP7_75t_SL sa33_reg_4_ (.QN(sa33_4_),
	.CLK(CTS_38),
	.D(n462));
   DFFHQNx2_ASAP7_75t_SL u0_w_reg_3__23_ (.QN(w3_23_),
	.CLK(CTS_39),
	.D(n651));
   DFFHQNx1_ASAP7_75t_SL sa02_reg_2_ (.QN(sa02_2_),
	.CLK(CTS_34),
	.D(n329));
   DFFHQNx1_ASAP7_75t_SL sa22_reg_4_ (.QN(sa22_4_),
	.CLK(CTS_34),
	.D(n514));
   DFFHQNx1_ASAP7_75t_SL sa12_reg_0_ (.QN(sa12_0_),
	.CLK(CTS_32),
	.D(FE_OCPN29434_n408));
   DFFHQNx1_ASAP7_75t_SL sa13_reg_2_ (.QN(sa13_2_),
	.CLK(CTS_31),
	.D(FE_OCPN28444_n428));
   DFFHQNx1_ASAP7_75t_L sa01_reg_2_ (.QN(sa01_2_),
	.CLK(CTS_32),
	.D(n401));
   DFFHQNx1_ASAP7_75t_SL sa02_reg_3_ (.QN(sa02_3_),
	.CLK(CTS_34),
	.D(n417));
   DFFHQNx1_ASAP7_75t_SL sa31_reg_3_ (.QN(sa31_3_),
	.CLK(CTS_33),
	.D(n440));
   DFFHQNx1_ASAP7_75t_SL sa10_reg_3_ (.QN(sa10_3_),
	.CLK(CTS_37),
	.D(n461));
   DFFHQNx2_ASAP7_75t_SL sa33_reg_2_ (.QN(sa33_2_),
	.CLK(CTS_37),
	.D(n477));
   DFFHQNx1_ASAP7_75t_SL sa03_reg_2_ (.QN(sa03_2_),
	.CLK(CTS_37),
	.D(n411));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__29_ (.QN(w3_29_),
	.CLK(CTS_37),
	.D(n646));
   DFFHQNx1_ASAP7_75t_L sa23_reg_7_ (.QN(sa23_7_),
	.CLK(CTS_36),
	.D(n512));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__4_ (.QN(w3_4_),
	.CLK(CTS_31),
	.D(n641));
   DFFHQNx1_ASAP7_75t_SL sa12_reg_4_ (.QN(sa12_4_),
	.CLK(CTS_32),
	.D(n494));
   DFFHQNx1_ASAP7_75t_SL sa00_reg_2_ (.QN(sa00_2_),
	.CLK(CTS_39),
	.D(n376));
   DFFHQNx2_ASAP7_75t_SL u0_w_reg_3__25_ (.QN(w3_25_),
	.CLK(CTS_37),
	.D(n626));
   DFFHQNx2_ASAP7_75t_SL sa00_reg_5_ (.QN(sa00_5_),
	.CLK(CTS_39),
	.D(n392));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__27_ (.QN(w3_27_),
	.CLK(CTS_38),
	.D(n638));
   DFFHQNx1_ASAP7_75t_SL sa00_reg_3_ (.QN(sa00_3_),
	.CLK(CTS_39),
	.D(n451));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__30_ (.QN(w3_30_),
	.CLK(CTS_38),
	.D(n650));
   DFFHQNx1_ASAP7_75t_SL sa03_reg_0_ (.QN(sa03_0_),
	.CLK(CTS_37),
	.D(n340));
   DFFHQNx1_ASAP7_75t_SL sa13_reg_5_ (.QN(sa13_5_),
	.CLK(CTS_33),
	.D(FE_OCPN29257_n474));
   DFFHQNx1_ASAP7_75t_SL sa21_reg_5_ (.QN(sa21_5_),
	.CLK(CTS_36),
	.D(n478));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_3_ (.QN(sa20_3_),
	.CLK(CTS_33),
	.D(n450));
   DFFHQNx1_ASAP7_75t_SL sa30_reg_2_ (.QN(sa30_2_),
	.CLK(CTS_33),
	.D(FE_OCPN29394_n479));
   DFFHQNx1_ASAP7_75t_SL sa13_reg_1_ (.QN(sa13_1_),
	.CLK(CTS_31),
	.D(FE_OCPN27320_n410));
   DFFHQNx1_ASAP7_75t_SL sa11_reg_1_ (.QN(sa11_1_),
	.CLK(CTS_31),
	.D(n386));
   DFFHQNx2_ASAP7_75t_SL sa03_reg_3_ (.QN(sa03_3_),
	.CLK(CTS_37),
	.D(n443));
   DFFHQNx1_ASAP7_75t_SL sa23_reg_4_ (.QN(sa23_4_),
	.CLK(CTS_36),
	.D(n519));
   DFFHQNx1_ASAP7_75t_SL sa23_reg_1_ (.QN(sa23_1_),
	.CLK(CTS_36),
	.D(n425));
   DFFHQNx1_ASAP7_75t_SL sa11_reg_5_ (.QN(sa11_5_),
	.CLK(CTS_31),
	.D(FE_OCPN29393_n483));
   DFFHQNx1_ASAP7_75t_SL sa30_reg_4_ (.QN(sa30_4_),
	.CLK(CTS_33),
	.D(n497));
   DFFHQNx2_ASAP7_75t_SL sa30_reg_0_ (.QN(sa30_0_),
	.CLK(CTS_33),
	.D(FE_OCPN27530_n362));
   DFFHQNx1_ASAP7_75t_SL sa23_reg_2_ (.QN(sa23_2_),
	.CLK(CTS_36),
	.D(n470));
   DFFHQNx1_ASAP7_75t_SL sa11_reg_2_ (.QN(sa11_2_),
	.CLK(CTS_31),
	.D(FE_OCPN29552_n393));
   DFFHQNx1_ASAP7_75t_SL sa12_reg_2_ (.QN(sa12_2_),
	.CLK(CTS_32),
	.D(FE_OCPN29590_n449));
   DFFHQNx1_ASAP7_75t_SL sa23_reg_5_ (.QN(sa23_5_),
	.CLK(CTS_36),
	.D(n464));
   DFFHQNx1_ASAP7_75t_SL sa31_reg_1_ (.QN(sa31_1_),
	.CLK(CTS_34),
	.D(n469));
   DFFHQNx1_ASAP7_75t_SL sa10_reg_5_ (.QN(sa10_5_),
	.CLK(CTS_37),
	.D(FE_OCPN29442_n458));
   DFFHQNx1_ASAP7_75t_SL sa20_reg_2_ (.QN(sa20_2_),
	.CLK(CTS_33),
	.D(n476));
   DFFHQNx1_ASAP7_75t_SL sa10_reg_2_ (.QN(sa10_2_),
	.CLK(CTS_37),
	.D(n391));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__15_ (.QN(w3_15_),
	.CLK(CTS_31),
	.D(n652));
   DFFHQNx1_ASAP7_75t_SL sa30_reg_3_ (.QN(sa30_3_),
	.CLK(CTS_31),
	.D(FE_OCPN29574_n484));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__9_ (.QN(w3_9_),
	.CLK(CTS_31),
	.D(n624));
   DFFHQNx1_ASAP7_75t_SL sa10_reg_4_ (.QN(sa10_4_),
	.CLK(CTS_37),
	.D(n513));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__20_ (.QN(w3_20_),
	.CLK(CTS_39),
	.D(n639));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__19_ (.QN(w3_19_),
	.CLK(CTS_39),
	.D(n631));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__11_ (.QN(w3_11_),
	.CLK(CTS_31),
	.D(n648));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__7_ (.QN(w3_7_),
	.CLK(CTS_31),
	.D(n653));
   DFFHQNx1_ASAP7_75t_SL u0_w_reg_3__3_ (.QN(w3_3_),
	.CLK(CTS_38),
	.D(n629));
   NOR2x1_ASAP7_75t_SL U13400 (.Y(n26192),
	.A(n26003),
	.B(n26002));
   NOR2xp33_ASAP7_75t_R U13402 (.Y(n25466),
	.A(sa03_7_),
	.B(FE_OFN156_sa03_6));
   NOR2x1p5_ASAP7_75t_SL U13403 (.Y(n21906),
	.A(FE_OFN29255_n),
	.B(n16629));
   NOR2x1p5_ASAP7_75t_L U13404 (.Y(n26100),
	.A(FE_OCPN27951_n19098),
	.B(FE_OFN29062_n18651));
   NOR2x1_ASAP7_75t_L U13406 (.Y(n24726),
	.A(n23981),
	.B(n16648));
   NAND3x1_ASAP7_75t_SL U13407 (.Y(n15813),
	.A(FE_OCPN8252_FE_OFN28661_w3_7),
	.B(FE_OFN25900_w3_4),
	.C(FE_OFN29052_w3_5));
   NOR2x1p5_ASAP7_75t_L U13408 (.Y(n13844),
	.A(FE_OFN28715_w3_15),
	.B(FE_OCPN29570_n15423));
   NOR2x1_ASAP7_75t_L U13409 (.Y(n13741),
	.A(n24831),
	.B(FE_OCPN28076_FE_OFN9_w3_6));
   NOR2x1_ASAP7_75t_SL U13411 (.Y(n20476),
	.A(n18457),
	.B(n18456));
   NOR2x2_ASAP7_75t_SL U13412 (.Y(n18008),
	.A(FE_OCPN27599_n18875),
	.B(n17996));
   NOR2x1_ASAP7_75t_SL U13413 (.Y(n21715),
	.A(n18875),
	.B(n17993));
   NOR2x1_ASAP7_75t_SL U13415 (.Y(n16750),
	.A(FE_OCPN29293_FE_OFN28678_sa21_3),
	.B(n16806));
   NOR2x1_ASAP7_75t_SL U13416 (.Y(n17757),
	.A(FE_OCPN27261_sa02_0),
	.B(FE_OFN29049_n17756));
   NAND2x2_ASAP7_75t_SL U13417 (.Y(n13771),
	.A(FE_OCPN27985_n24831),
	.B(FE_OFN25887_w3_3));
   NOR2x1_ASAP7_75t_SL U13418 (.Y(n17546),
	.A(FE_OFN27148_sa32_3),
	.B(n18837));
   INVxp67_ASAP7_75t_R U13421 (.Y(n24913),
	.A(FE_OFN26531_n));
   NOR2x1p5_ASAP7_75t_SL U13422 (.Y(n18971),
	.A(FE_OFN29191_sa23_2),
	.B(FE_OFN29189_sa23_0));
   NOR2x1p5_ASAP7_75t_L U13423 (.Y(n18529),
	.A(FE_OCPN29380_sa20_1),
	.B(FE_OCPN28223_FE_OFN27219_n18522));
   NOR2x1_ASAP7_75t_L U13424 (.Y(n18016),
	.A(FE_OCPN27483_FE_OFN16132_sa03_5),
	.B(n18029));
   NOR2x1p5_ASAP7_75t_L U13425 (.Y(n19019),
	.A(FE_OCPN29373_FE_OFN29191_sa23_2),
	.B(n23504));
   NOR2x1_ASAP7_75t_SL U13426 (.Y(n17898),
	.A(FE_OCPN29494_sa12_4),
	.B(n17949));
   NAND2x1p5_ASAP7_75t_L U13427 (.Y(n13805),
	.A(FE_OCPN29427_w3_15),
	.B(n15924));
   NOR2xp67_ASAP7_75t_SL U13428 (.Y(n21734),
	.A(n18875),
	.B(n21725));
   NOR2x1p5_ASAP7_75t_SL U13429 (.Y(n16300),
	.A(FE_OCPN29482_FE_OFN26014_sa31_3),
	.B(FE_OFN28669_sa31_5));
   NOR2x1p5_ASAP7_75t_SL U13430 (.Y(n21553),
	.A(FE_OFN16141_sa01_3),
	.B(FE_OCPN28217_sa01_5));
   NOR2x1p5_ASAP7_75t_SL U13431 (.Y(n18532),
	.A(FE_OCPN27371_sa20_2),
	.B(FE_OCPN28223_FE_OFN27219_n18522));
   NOR2x1p5_ASAP7_75t_SL U13432 (.Y(n22632),
	.A(FE_OCPN29431_sa30_3),
	.B(n17618));
   NOR2x1p5_ASAP7_75t_SL U13433 (.Y(n15922),
	.A(FE_OCPN28402_w3_13),
	.B(FE_OFN27200_n));
   NOR2x2_ASAP7_75t_SL U13434 (.Y(n17453),
	.A(FE_OCPN27229_sa11_2),
	.B(n21818));
   NOR2x2_ASAP7_75t_L U13436 (.Y(n16299),
	.A(FE_OFN28669_sa31_5),
	.B(n16321));
   NOR2x1p5_ASAP7_75t_SL U13437 (.Y(n17602),
	.A(FE_OFN28895_sa30_2),
	.B(n19051));
   NOR2x2_ASAP7_75t_SL U13438 (.Y(n18583),
	.A(FE_OFN28791_n),
	.B(n18571));
   NOR2x1p5_ASAP7_75t_SL U13439 (.Y(n19725),
	.A(FE_OFN27148_sa32_3),
	.B(FE_OCPN27499_FE_OFN16151_sa32_5));
   NOR3xp33_ASAP7_75t_SL U13440 (.Y(n23644),
	.A(FE_OFN25989_sa21_4),
	.B(FE_OFN28678_sa21_3),
	.C(n16783));
   NOR2x1p5_ASAP7_75t_SL U13441 (.Y(n17529),
	.A(FE_OFN28892_n),
	.B(n17566));
   NOR2x1p5_ASAP7_75t_SL U13442 (.Y(n16430),
	.A(FE_OFN25938_sa33_3),
	.B(n16677));
   NOR2x1p5_ASAP7_75t_SL U13443 (.Y(n16760),
	.A(FE_OCPN27327_sa21_2),
	.B(FE_OFN28903_sa21_0));
   NOR2x1p5_ASAP7_75t_SL U13444 (.Y(n22745),
	.A(FE_OFN25908_sa12_2),
	.B(n17971));
   NOR2x1p5_ASAP7_75t_L U13446 (.Y(n12998),
	.A(FE_OCPN27227_sa00_5),
	.B(n17282));
   NOR3xp33_ASAP7_75t_SL U13447 (.Y(n13671),
	.A(FE_OFN28571_w3_28),
	.B(FE_OCPN28096_w3_31),
	.C(FE_OCPN29428_FE_OFN27131_w3_29));
   NOR2x2_ASAP7_75t_L U13448 (.Y(n16975),
	.A(FE_OFN16181_sa13_5),
	.B(FE_OFN27186_sa13_4));
   NOR2x1p5_ASAP7_75t_SL U13449 (.Y(n22543),
	.A(n17760),
	.B(FE_OCPN27566_FE_OFN16138_sa02_5));
   NOR2x1p5_ASAP7_75t_SL U13450 (.Y(n16295),
	.A(FE_OFN100_sa31_1),
	.B(FE_OFN26095_n16293));
   NOR2x1p5_ASAP7_75t_SL U13451 (.Y(n16983),
	.A(FE_OFN28478_sa13_2),
	.B(n17079));
   TIEHIx1_ASAP7_75t_L U13452 (.H(n22528));
   O2A1O1Ixp33_ASAP7_75t_L U13454 (.Y(n13312),
	.A1(n14479),
	.A2(n15203),
	.B(FE_OFN26104_n13659),
	.C(n13637));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13455 (.Y(n14053),
	.A1(FE_OFN27151_n),
	.A2(FE_OFN28706_n),
	.B(n15339),
	.C(FE_OFN16352_n14289));
   O2A1O1Ixp5_ASAP7_75t_SL U13456 (.Y(n14392),
	.A1(FE_OFN27151_n),
	.A2(n15694),
	.B(n15484),
	.C(FE_OFN16210_n13876));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13457 (.Y(n14375),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(FE_OFN25915_n15514),
	.B(FE_PSN8334_n15539),
	.C(FE_OFN16352_n14289));
   O2A1O1Ixp33_ASAP7_75t_L U13458 (.Y(n13610),
	.A1(n14514),
	.A2(FE_OFN27085_n),
	.B(n13609),
	.C(n15238));
   OAI21xp33_ASAP7_75t_SL U13459 (.Y(n15346),
	.A1(n15744),
	.A2(n15480),
	.B(n15345));
   OAI21xp5_ASAP7_75t_SL U13461 (.Y(n15711),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(n15694),
	.B(n15492));
   INVx1_ASAP7_75t_SL U13463 (.Y(n13614),
	.A(n13610));
   OAI22xp5_ASAP7_75t_L U13464 (.Y(n13516),
	.A1(FE_OFN27211_w3_30),
	.A2(n14592),
	.B1(FE_OFN26051_w3_27),
	.B2(n14592));
   NAND2xp33_ASAP7_75t_L U13466 (.Y(n14115),
	.A(n14114),
	.B(n14113));
   OAI21xp33_ASAP7_75t_SL U13467 (.Y(n15350),
	.A1(n15349),
	.A2(n15710),
	.B(n15348));
   NAND2xp5_ASAP7_75t_R U13468 (.Y(n15108),
	.A(n15033),
	.B(FE_OFN25918_n15813));
   NAND2xp5_ASAP7_75t_L U13469 (.Y(n15491),
	.A(n15757),
	.B(n12994));
   NAND2xp5_ASAP7_75t_L U13471 (.Y(n17811),
	.A(n17810),
	.B(n17809));
   NAND2xp5_ASAP7_75t_SL U13473 (.Y(n22290),
	.A(n18205),
	.B(n18204));
   NAND2xp5_ASAP7_75t_SL U13477 (.Y(n14595),
	.A(n14533),
	.B(n14532));
   NAND2xp5_ASAP7_75t_SL U13478 (.Y(n14217),
	.A(n14216),
	.B(n14215));
   OAI22xp33_ASAP7_75t_SL U13479 (.Y(n15829),
	.A1(FE_OFN28671_FE_OCPN28076),
	.A2(n15033),
	.B1(n13771),
	.B2(n15033));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13481 (.Y(n13772),
	.A1(FE_OFN28671_FE_OCPN28076),
	.A2(n15817),
	.B(n13771),
	.C(FE_OFN28691_n13725));
   O2A1O1Ixp33_ASAP7_75t_L U13482 (.Y(n13878),
	.A1(FE_OFN26045_n25377),
	.A2(FE_OFN26091_n24663),
	.B(n15668),
	.C(n15747));
   OAI22xp33_ASAP7_75t_L U13483 (.Y(n15024),
	.A1(n15859),
	.A2(n15021),
	.B1(n15020),
	.B2(n15021));
   O2A1O1Ixp33_ASAP7_75t_L U13484 (.Y(n15594),
	.A1(n24831),
	.A2(n15809),
	.B(n15588),
	.C(n15587));
   NAND2x1_ASAP7_75t_L U13485 (.Y(n14929),
	.A(FE_OFN26642_w3_14),
	.B(FE_OFN28856_n15450));
   O2A1O1Ixp33_ASAP7_75t_SL U13486 (.Y(n13699),
	.A1(n13669),
	.A2(FE_OFN27085_n),
	.B(n13668),
	.C(n15238));
   O2A1O1Ixp33_ASAP7_75t_SL U13487 (.Y(n15019),
	.A1(FE_OFN26058_w3_1),
	.A2(n25140),
	.B(FE_OFN28829_n),
	.C(n15028));
   O2A1O1Ixp5_ASAP7_75t_SL U13488 (.Y(n18284),
	.A1(FE_OFN16319_n20527),
	.A2(FE_OFN28801_n16978),
	.B(FE_OCPN28212_n16980),
	.C(n18283));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13489 (.Y(n19250),
	.A1(FE_OFN28704_FE_OCPN27740_sa02_4),
	.A2(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(FE_OCPN27566_FE_OFN16138_sa02_5),
	.C(FE_OFN28961_n17744));
   INVx1_ASAP7_75t_SL U13490 (.Y(n18207),
	.A(n23309));
   NAND2xp5_ASAP7_75t_SL U13492 (.Y(n19551),
	.A(n22251),
	.B(n19503));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13494 (.Y(n13773),
	.A1(FE_OFN28671_FE_OCPN28076),
	.A2(FE_OFN26532_n13766),
	.B(FE_OFN28831_n15838),
	.C(n13772));
   NAND2xp5_ASAP7_75t_SL U13495 (.Y(n14545),
	.A(n13421),
	.B(n15197));
   OAI21x1_ASAP7_75t_SL U13497 (.Y(n15856),
	.A1(FE_OFN28671_FE_OCPN28076),
	.A2(FE_OFN26532_n13766),
	.B(n14442));
   O2A1O1Ixp5_ASAP7_75t_SL U13499 (.Y(n14672),
	.A1(n15438),
	.A2(FE_OFN109_n15994),
	.B(FE_OFN28544_n13805),
	.C(n14667));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13500 (.Y(n15673),
	.A1(FE_OFN5_w3_22),
	.A2(FE_OFN26053_n25415),
	.B(FE_OFN26045_n25377),
	.C(n13869));
   O2A1O1Ixp33_ASAP7_75t_SL U13502 (.Y(n19175),
	.A1(n17444),
	.A2(n23355),
	.B(n21365),
	.C(n23262));
   NAND2xp5_ASAP7_75t_SL U13503 (.Y(n22645),
	.A(n22615),
	.B(n18370));
   NAND2x1_ASAP7_75t_SL U13504 (.Y(n23701),
	.A(n21664),
	.B(n23871));
   NAND2x1_ASAP7_75t_SL U13507 (.Y(n20318),
	.A(n20002),
	.B(n19889));
   O2A1O1Ixp33_ASAP7_75t_SL U13512 (.Y(n17034),
	.A1(FE_OCPN28137_n17170),
	.A2(FE_OFN26170_n19361),
	.B(FE_OFN16162_n25869),
	.C(n20529));
   NAND2xp5_ASAP7_75t_L U13513 (.Y(n20427),
	.A(n17602),
	.B(n25108));
   OAI21xp5_ASAP7_75t_SL U13516 (.Y(n21241),
	.A1(FE_OCPN28353_n18534),
	.A2(n20670),
	.B(n23750));
   NAND2x1p5_ASAP7_75t_SL U13517 (.Y(n18602),
	.A(FE_OCPN27558_sa20_4),
	.B(FE_OCPN27633_sa20_5));
   O2A1O1Ixp5_ASAP7_75t_SL U13519 (.Y(n22946),
	.A1(FE_OCPN27955_n22945),
	.A2(FE_OFN29026_n20911),
	.B(FE_OFN28580_n23491),
	.C(n22944));
   NAND2xp33_ASAP7_75t_L U13521 (.Y(n22185),
	.A(n24220),
	.B(n22468));
   NAND2xp5_ASAP7_75t_L U13522 (.Y(n19736),
	.A(n19731),
	.B(n19733));
   NAND2xp5_ASAP7_75t_SL U13523 (.Y(n19874),
	.A(n19894),
	.B(n19974));
   NAND2xp5_ASAP7_75t_SL U13525 (.Y(n17291),
	.A(n17290),
	.B(n17289));
   O2A1O1Ixp33_ASAP7_75t_SL U13526 (.Y(n14815),
	.A1(n14814),
	.A2(n14813),
	.B(n13867),
	.C(n14812));
   NAND2xp5_ASAP7_75t_SL U13528 (.Y(n14913),
	.A(FE_OFN27200_n),
	.B(n25782));
   O2A1O1Ixp33_ASAP7_75t_SL U13529 (.Y(n24273),
	.A1(n24272),
	.A2(n24271),
	.B(n25575),
	.C(n24270));
   INVx2_ASAP7_75t_L U13530 (.Y(n16408),
	.A(FE_OFN29016_n16512));
   O2A1O1Ixp33_ASAP7_75t_SL U13532 (.Y(n26463),
	.A1(n25068),
	.A2(n25067),
	.B(n26282),
	.C(n25066));
   NAND2xp5_ASAP7_75t_L U13533 (.Y(n23724),
	.A(n23833),
	.B(n23755));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13536 (.Y(n19642),
	.A1(FE_OCPN28040_n19766),
	.A2(n23148),
	.B(n19641),
	.C(n23948));
   NAND2x1p5_ASAP7_75t_L U13537 (.Y(n16647),
	.A(FE_OCPN27635_sa10_4),
	.B(FE_OFN25959_n23011));
   NAND2xp5_ASAP7_75t_SL U13538 (.Y(n19605),
	.A(n18773),
	.B(n21157));
   AOI21x1_ASAP7_75t_SL U13539 (.Y(n23720),
	.A1(FE_OFN29076_n18540),
	.A2(n20617),
	.B(n23829));
   NOR2x1p5_ASAP7_75t_SL U13540 (.Y(n16424),
	.A(FE_OCPN29391_FE_OFN29162_sa33_2),
	.B(FE_OCPN27666_n17418));
   O2A1O1Ixp33_ASAP7_75t_R U13543 (.Y(n20819),
	.A1(n20796),
	.A2(FE_OCPN8265_n24362),
	.B(FE_OFN29075_n22745),
	.C(FE_OFN28520_n22753));
   NAND2xp5_ASAP7_75t_SL U13545 (.Y(n19901),
	.A(n17879),
	.B(n17878));
   NAND2xp5_ASAP7_75t_L U13547 (.Y(n17754),
	.A(n17753),
	.B(n17752));
   NAND2xp5_ASAP7_75t_L U13549 (.Y(n16510),
	.A(n16509),
	.B(n26294));
   NAND2x1_ASAP7_75t_SL U13550 (.Y(n14602),
	.A(n14600),
	.B(n14599));
   NAND2x1p5_ASAP7_75t_SL U13551 (.Y(n15447),
	.A(FE_OFN27115_n),
	.B(FE_OFN16459_n));
   O2A1O1Ixp33_ASAP7_75t_L U13552 (.Y(n15506),
	.A1(FE_OFN6_w3_22),
	.A2(FE_OFN25915_n15514),
	.B(n15339),
	.C(n15660));
   NAND2x1p5_ASAP7_75t_L U13553 (.Y(n15842),
	.A(FE_OFN26591_w3_3),
	.B(FE_OFN26531_n));
   NAND2xp5_ASAP7_75t_L U13554 (.Y(n15888),
	.A(w3_2_),
	.B(n25596));
   OAI21x1_ASAP7_75t_SL U13555 (.Y(n15239),
	.A1(FE_OCPN27656_w3_25),
	.A2(FE_OFN26048_w3_27),
	.B(FE_OFN27207_w3_30));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13556 (.Y(n13473),
	.A1(n15224),
	.A2(FE_OFN28455_n13348),
	.B(n13428),
	.C(n13427));
   NAND2xp5_ASAP7_75t_SL U13557 (.Y(n15560),
	.A(n15558),
	.B(n15557));
   O2A1O1Ixp33_ASAP7_75t_R U13558 (.Y(n24105),
	.A1(n26777),
	.A2(n26776),
	.B(FE_OCPN27935_n26773),
	.C(n24118));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13559 (.Y(n26576),
	.A1(n26710),
	.A2(n26709),
	.B(n26706),
	.C(n26575));
   O2A1O1Ixp33_ASAP7_75t_SRAM U13560 (.Y(n25658),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25669),
	.C(n25657));
   O2A1O1Ixp5_ASAP7_75t_L U13561 (.Y(n25312),
	.A1(n27140),
	.A2(n27139),
	.B(n27136),
	.C(FE_OFN26012_n27208));
   O2A1O1Ixp33_ASAP7_75t_SRAM U13562 (.Y(n25141),
	.A1(n25420),
	.A2(FE_OFN28561_n25419),
	.B(FE_OCPN27682_n25414),
	.C(FE_OFN25887_w3_3));
   NAND2xp5_ASAP7_75t_SL U13563 (.Y(n16392),
	.A(n20836),
	.B(n16390));
   O2A1O1Ixp33_ASAP7_75t_SL U13564 (.Y(n26700),
	.A1(n27004),
	.A2(n26702),
	.B(n26699),
	.C(n26698));
   INVx1_ASAP7_75t_SL U13567 (.Y(n26866),
	.A(FE_OCPN27283_n26867));
   NAND2x1_ASAP7_75t_SL U13568 (.Y(n19180),
	.A(n19179),
	.B(n19178));
   NAND2xp5_ASAP7_75t_L U13569 (.Y(n18507),
	.A(n21603),
	.B(n18502));
   NAND2x1p5_ASAP7_75t_L U13570 (.Y(n18364),
	.A(FE_OCPN29431_sa30_3),
	.B(FE_OFN16333_sa30_4));
   NAND2x1p5_ASAP7_75t_SL U13572 (.Y(n18582),
	.A(FE_OCPN27371_sa20_2),
	.B(FE_OCPN29380_sa20_1));
   NAND2xp5_ASAP7_75t_L U13574 (.Y(n25994),
	.A(FE_OFN16162_n25869),
	.B(FE_OCPN28137_n17170));
   NAND2x1_ASAP7_75t_SL U13576 (.Y(n17059),
	.A(sa13_4_),
	.B(n16981));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13577 (.Y(n18241),
	.A1(FE_OFN16319_n20527),
	.A2(FE_OFN28801_n16978),
	.B(n17060),
	.C(n17154));
   O2A1O1Ixp5_ASAP7_75t_SL U13578 (.Y(n20505),
	.A1(FE_OFN16162_n25869),
	.A2(n19376),
	.B(FE_OCPN28137_n17170),
	.C(n20521));
   NAND2x1_ASAP7_75t_SL U13579 (.Y(n20471),
	.A(n17637),
	.B(FE_OFN16200_sa30_2));
   NAND2x1p5_ASAP7_75t_L U13581 (.Y(n17489),
	.A(FE_OCPN27242_sa11_1),
	.B(FE_OCPN27512_sa11_2));
   NAND2x1p5_ASAP7_75t_SL U13583 (.Y(n21772),
	.A(FE_OFN28680_n),
	.B(n20739));
   NAND2xp5_ASAP7_75t_SL U13584 (.Y(n23707),
	.A(n23706),
	.B(n23705));
   NAND2xp33_ASAP7_75t_L U13585 (.Y(n23548),
	.A(sa33_6_),
	.B(n16468));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13587 (.Y(n19012),
	.A1(FE_OCPN27955_n22945),
	.A2(FE_OCPN29480_n20913),
	.B(FE_OCPN28381_n26660),
	.C(n22998));
   NAND2x1p5_ASAP7_75t_SL U13588 (.Y(n19527),
	.A(FE_OFN28764_n17928),
	.B(n17899));
   NAND2x1p5_ASAP7_75t_SL U13590 (.Y(n25350),
	.A(n16757),
	.B(FE_OFN16447_n16749));
   NAND2xp5_ASAP7_75t_SL U13594 (.Y(n20066),
	.A(n20868),
	.B(n21989));
   O2A1O1Ixp33_ASAP7_75t_L U13595 (.Y(n25238),
	.A1(n27102),
	.A2(n25240),
	.B(FE_OFN115_n27187),
	.C(n25236));
   O2A1O1Ixp5_ASAP7_75t_SL U13597 (.Y(n24211),
	.A1(n24208),
	.A2(n24207),
	.B(n26679),
	.C(n26675));
   OAI21xp5_ASAP7_75t_SL U13598 (.Y(n21491),
	.A1(FE_OCPN27951_n19098),
	.A2(n19097),
	.B(n19096));
   O2A1O1Ixp33_ASAP7_75t_SL U13599 (.Y(n14603),
	.A1(n15259),
	.A2(n14605),
	.B(n14602),
	.C(n26544));
   O2A1O1Ixp33_ASAP7_75t_SL U13600 (.Y(n14407),
	.A1(n15704),
	.A2(n14406),
	.B(n14405),
	.C(n14404));
   NAND2xp5_ASAP7_75t_R U13601 (.Y(n16023),
	.A(w3_10_),
	.B(w3_8_));
   NAND2xp5_ASAP7_75t_L U13602 (.Y(n14585),
	.A(FE_OFN16412_w3_26),
	.B(FE_OFN25880_w3_24));
   O2A1O1Ixp5_ASAP7_75t_SL U13603 (.Y(n26499),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(n26498),
	.C(n26497));
   O2A1O1Ixp33_ASAP7_75t_R U13604 (.Y(n25558),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(FE_OCPN28119_n26955),
	.C(n25570));
   O2A1O1Ixp33_ASAP7_75t_L U13605 (.Y(n25890),
	.A1(FE_OFN16158_n26959),
	.A2(n25892),
	.B(n25889),
	.C(n25895));
   NAND2xp5_ASAP7_75t_SL U13606 (.Y(n25859),
	.A(FE_OFN28615_n26191),
	.B(n25854));
   O2A1O1Ixp5_ASAP7_75t_SL U13607 (.Y(n25332),
	.A1(n27168),
	.A2(n27167),
	.B(n27163),
	.C(n26747));
   O2A1O1Ixp33_ASAP7_75t_R U13608 (.Y(n26956),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(FE_OCPN28119_n26955),
	.C(n26963));
   O2A1O1Ixp33_ASAP7_75t_L U13609 (.Y(n26325),
	.A1(n26315),
	.A2(n26314),
	.B(n26313),
	.C(n26312));
   O2A1O1Ixp5_ASAP7_75t_SL U13610 (.Y(n26213),
	.A1(n27027),
	.A2(n25701),
	.B(n25700),
	.C(n25699));
   O2A1O1Ixp33_ASAP7_75t_L U13611 (.Y(n24715),
	.A1(n17506),
	.A2(n24717),
	.B(n24714),
	.C(n24721));
   NAND2xp5_ASAP7_75t_SL U13612 (.Y(n25684),
	.A(FE_OFN28525_n25751),
	.B(n26705));
   NAND2xp5_ASAP7_75t_SL U13613 (.Y(n24573),
	.A(n25251),
	.B(n25966));
   NAND2xp5_ASAP7_75t_SL U13614 (.Y(n24194),
	.A(n16364),
	.B(n16363));
   O2A1O1Ixp5_ASAP7_75t_SL U13615 (.Y(n16486),
	.A1(n23557),
	.A2(n16485),
	.B(n26770),
	.C(n16484));
   O2A1O1Ixp33_ASAP7_75t_L U13617 (.Y(n19284),
	.A1(FE_OCPN29387_n25273),
	.A2(n25208),
	.B(n27183),
	.C(n25215));
   O2A1O1Ixp5_ASAP7_75t_L U13618 (.Y(n20181),
	.A1(FE_OCPN28196_n22547),
	.A2(n20180),
	.B(n27183),
	.C(n20179));
   NAND2xp5_ASAP7_75t_SL U13619 (.Y(n27140),
	.A(sa02_7_),
	.B(n17815));
   O2A1O1Ixp5_ASAP7_75t_SL U13620 (.Y(n19807),
	.A1(FE_OFN16202_n19806),
	.A2(n19805),
	.B(n24974),
	.C(n24677));
   O2A1O1Ixp5_ASAP7_75t_SL U13621 (.Y(n22217),
	.A1(n22216),
	.A2(n22215),
	.B(n26282),
	.C(n22214));
   O2A1O1Ixp33_ASAP7_75t_SL U13622 (.Y(n23847),
	.A1(n25639),
	.A2(n25638),
	.B(n26323),
	.C(n23846));
   NAND2xp5_ASAP7_75t_SL U13623 (.Y(n20041),
	.A(n20040),
	.B(n20039));
   NAND2xp5_ASAP7_75t_L U13624 (.Y(n25885),
	.A(n17172),
	.B(n17096));
   NAND2xp5_ASAP7_75t_SL U13625 (.Y(n20114),
	.A(n19930),
	.B(n19929));
   NAND2xp5_ASAP7_75t_R U13626 (.Y(n23467),
	.A(sa03_7_),
	.B(FE_OFN156_sa03_6));
   O2A1O1Ixp33_ASAP7_75t_SL U13629 (.Y(n19692),
	.A1(n23144),
	.A2(n19691),
	.B(n24974),
	.C(n19690));
   NAND2xp5_ASAP7_75t_SL U13630 (.Y(n24460),
	.A(n16654),
	.B(n19669));
   NAND2x1_ASAP7_75t_L U13631 (.Y(n25139),
	.A(FE_OFN59_sa10_7),
	.B(sa10_6_));
   O2A1O1Ixp5_ASAP7_75t_SL U13632 (.Y(n19157),
	.A1(n21180),
	.A2(n19156),
	.B(n26637),
	.C(n19155));
   NAND2xp33_ASAP7_75t_SL U13633 (.Y(n17506),
	.A(sa11_6_),
	.B(n19161));
   O2A1O1Ixp5_ASAP7_75t_SL U13634 (.Y(n22520),
	.A1(n22519),
	.A2(n22518),
	.B(n26082),
	.C(n22517));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13635 (.Y(n18513),
	.A1(n24798),
	.A2(n24797),
	.B(n26584),
	.C(n18512));
   NOR2x1p5_ASAP7_75t_SL U13636 (.Y(n18176),
	.A(FE_OFN28688_sa22_2),
	.B(FE_OFN29152_sa22_0));
   O2A1O1Ixp5_ASAP7_75t_SL U13637 (.Y(n22866),
	.A1(n22865),
	.A2(n22864),
	.B(n26878),
	.C(n22863));
   O2A1O1Ixp33_ASAP7_75t_SL U13638 (.Y(n26882),
	.A1(n21802),
	.A2(n18234),
	.B(n27117),
	.C(n18233));
   O2A1O1Ixp33_ASAP7_75t_L U13639 (.Y(n20645),
	.A1(FE_OFN28729_n20617),
	.A2(FE_OFN29081_n18526),
	.B(FE_OFN29112_FE_OCPN27870_n18527),
	.C(n20643));
   O2A1O1Ixp5_ASAP7_75t_SL U13640 (.Y(n18154),
	.A1(n23534),
	.A2(n18153),
	.B(n26770),
	.C(n18152));
   O2A1O1Ixp5_ASAP7_75t_SRAM U13641 (.Y(n16900),
	.A1(n24335),
	.A2(n24334),
	.B(n26770),
	.C(n24337));
   O2A1O1Ixp5_ASAP7_75t_SL U13642 (.Y(n19028),
	.A1(n26569),
	.A2(n26568),
	.B(n26567),
	.C(n19027));
   NAND2xp5_ASAP7_75t_L U13643 (.Y(n26710),
	.A(sa23_7_),
	.B(FE_OFN45_sa23_6));
   NAND2xp33_ASAP7_75t_L U13644 (.Y(n26464),
	.A(sa01_6_),
	.B(sa01_7_));
   NAND2x1p5_ASAP7_75t_R U13646 (.Y(n26607),
	.A(FE_OFN165_sa12_7),
	.B(n17915));
   NAND2xp5_ASAP7_75t_L U13647 (.Y(n25918),
	.A(FE_OCPN27541_n26748),
	.B(n25935));
   NAND2x1_ASAP7_75t_SL U13648 (.Y(n20301),
	.A(n17869),
	.B(n23640));
   O2A1O1Ixp33_ASAP7_75t_L U13649 (.Y(n17892),
	.A1(n17891),
	.A2(n17890),
	.B(n25575),
	.C(n17889));
   O2A1O1Ixp5_ASAP7_75t_SL U13651 (.Y(n20894),
	.A1(n20893),
	.A2(n20892),
	.B(n26407),
	.C(n20891));
   O2A1O1Ixp5_ASAP7_75t_SL U13652 (.Y(n25769),
	.A1(n24065),
	.A2(n24064),
	.B(n25682),
	.C(n24063));
   NAND2xp5_ASAP7_75t_L U13653 (.Y(n25509),
	.A(FE_OCPN29443_n25507),
	.B(FE_OFN28907_n26049));
   O2A1O1Ixp33_ASAP7_75t_L U13654 (.Y(n25242),
	.A1(n27168),
	.A2(n25823),
	.B(n26625),
	.C(FE_OFN28907_n26049));
   O2A1O1Ixp5_ASAP7_75t_SL U13655 (.Y(n21699),
	.A1(n21698),
	.A2(n21697),
	.B(n26323),
	.C(n21696));
   NAND2xp5_ASAP7_75t_L U13656 (.Y(n21493),
	.A(FE_OFN28499_sa00_6),
	.B(sa00_7_));
   O2A1O1Ixp5_ASAP7_75t_L U13661 (.Y(n24432),
	.A1(n24225),
	.A2(n24224),
	.B(n26282),
	.C(n24223));
   O2A1O1Ixp5_ASAP7_75t_SL U13663 (.Y(n27170),
	.A1(n27168),
	.A2(n27167),
	.B(n27166),
	.C(n27165));
   NAND2xp5_ASAP7_75t_SL U13664 (.Y(n25344),
	.A(n26052),
	.B(n25922));
   O2A1O1Ixp33_ASAP7_75t_SL U13665 (.Y(n26433),
	.A1(FE_OFN16180_n26542),
	.A2(n26431),
	.B(n26430),
	.C(n26429));
   O2A1O1Ixp33_ASAP7_75t_SRAM U13666 (.Y(n25430),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25429),
	.C(n25428));
   O2A1O1Ixp5_ASAP7_75t_R U13667 (.Y(n25673),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25671),
	.C(n25670));
   NAND2xp5_ASAP7_75t_SL U13668 (.Y(n25004),
	.A(n25000),
	.B(n24999));
   OAI21x1_ASAP7_75t_SL U13670 (.Y(n25363),
	.A1(n19750),
	.A2(n23899),
	.B(n19749));
   O2A1O1Ixp5_ASAP7_75t_SL U13672 (.Y(n24301),
	.A1(n23535),
	.A2(n16733),
	.B(n24610),
	.C(n16732));
   INVxp33_ASAP7_75t_SRAM U13674 (.Y(n27219),
	.A(w2_18_));
   O2A1O1Ixp5_ASAP7_75t_SL U13680 (.Y(n26428),
	.A1(n24624),
	.A2(n16970),
	.B(n26770),
	.C(n16969));
   OAI21x1_ASAP7_75t_SL U13683 (.Y(n26839),
	.A1(n18855),
	.A2(n23899),
	.B(n18854));
   O2A1O1Ixp33_ASAP7_75t_SL U13685 (.Y(n24418),
	.A1(n24044),
	.A2(n24043),
	.B(n26249),
	.C(n24042));
   OAI21xp5_ASAP7_75t_SL U13686 (.Y(n25495),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(FE_OCPN4698_n25497),
	.B(n25496));
   NAND2xp33_ASAP7_75t_SRAM U13690 (.Y(n24471),
	.A(FE_OFN28482_ld_r),
	.B(text_in_r_26_));
   O2A1O1Ixp33_ASAP7_75t_L U13691 (.Y(n26505),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(n27147),
	.B(FE_OCPN7556_n26504),
	.C(n26503));
   OAI21xp5_ASAP7_75t_SL U13692 (.Y(n26119),
	.A1(text_in_r_96_),
	.A2(FE_OFN28484_ld_r),
	.B(n26114));
   OAI21xp33_ASAP7_75t_L U13693 (.Y(n24757),
	.A1(n24758),
	.A2(FE_OCPN27430_n26334),
	.B(FE_OFN28489_ld_r));
   OAI21xp5_ASAP7_75t_SL U13694 (.Y(n26989),
	.A1(text_in_r_48_),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B(n26985));
   INVxp67_ASAP7_75t_SL U13696 (.Y(n26951),
	.A(w2_10_));
   OAI21xp5_ASAP7_75t_SL U13697 (.Y(n27131),
	.A1(n27133),
	.A2(n27132),
	.B(FE_OFN28484_ld_r));
   O2A1O1Ixp5_ASAP7_75t_SL U13698 (.Y(n27199),
	.A1(FE_OFN116_n27187),
	.A2(n27186),
	.B(FE_OCPN8214_n27185),
	.C(n27184));
   O2A1O1Ixp5_ASAP7_75t_SL U13699 (.Y(n25813),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OFN26024_n26115),
	.B(n25812),
	.C(n25811));
   NAND2x1_ASAP7_75t_SL U13701 (.Y(n27182),
	.A(n22538),
	.B(n22537));
   NAND2xp5_ASAP7_75t_SL U13702 (.Y(n26057),
	.A(n23862),
	.B(n23861));
   NAND2xp33_ASAP7_75t_SL U13703 (.Y(n26281),
	.A(FE_OCPN29330_n26459),
	.B(n23072));
   O2A1O1Ixp5_ASAP7_75t_SL U13705 (.Y(n27068),
	.A1(FE_OCPN28442_n27056),
	.A2(n27055),
	.B(n27054),
	.C(n27053));
   INVxp33_ASAP7_75t_SRAM U13706 (.Y(n27085),
	.A(w2_15_));
   O2A1O1Ixp5_ASAP7_75t_SL U13707 (.Y(n25481),
	.A1(FE_OCPN28100_n25470),
	.A2(n25469),
	.B(n25468),
	.C(n25467));
   O2A1O1Ixp5_ASAP7_75t_SL U13718 (.Y(n461),
	.A1(FE_OFN40_w0_19),
	.A2(text_in_r_115_),
	.B(n26232),
	.C(n26231));
   O2A1O1Ixp5_ASAP7_75t_SL U13719 (.Y(n462),
	.A1(FE_OFN25897_w3_4),
	.A2(text_in_r_4_),
	.B(n25666),
	.C(n25665));
   O2A1O1Ixp5_ASAP7_75t_SL U13722 (.Y(n432),
	.A1(FE_OCPN27985_n24831),
	.A2(text_in_r_1_),
	.B(n24851),
	.C(n24850));
   O2A1O1Ixp5_ASAP7_75t_SL U13723 (.Y(n523),
	.A1(w2_7_),
	.A2(text_in_r_39_),
	.B(n26629),
	.C(n26628));
   OAI22xp5_ASAP7_75t_L U13724 (.Y(n538),
	.A1(ld),
	.A2(n16115),
	.B1(key_55_),
	.B2(n16115));
   NAND2xp5_ASAP7_75t_SL U13726 (.Y(n649),
	.A(n16279),
	.B(n16278));
   OAI21xp5_ASAP7_75t_SL U13728 (.Y(n26392),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OCPN27274_n26394),
	.B(n26393));
   OAI22xp5_ASAP7_75t_L U13730 (.Y(n532),
	.A1(n16125),
	.A2(n16153),
	.B1(key_39_),
	.B2(n16153));
   NAND2xp5_ASAP7_75t_L U13733 (.Y(n16254),
	.A(FE_OFN28701_w3_16),
	.B(FE_OFN26021_n16253));
   OAI22xp5_ASAP7_75t_L U13734 (.Y(n613),
	.A1(ld),
	.A2(FE_OFN16361_n16263),
	.B1(key_57_),
	.B2(FE_OFN16361_n16263));
   OAI22xp33_ASAP7_75t_L U13736 (.Y(n553),
	.A1(ld),
	.A2(FE_OFN26630_n16190),
	.B1(key_61_),
	.B2(FE_OFN26630_n16190));
   O2A1O1Ixp5_ASAP7_75t_SL U13737 (.Y(n386),
	.A1(w1_17_),
	.A2(text_in_r_81_),
	.B(n26220),
	.C(n26219));
   AOI22x1_ASAP7_75t_SL U13739 (.Y(n16059),
	.A1(w1_4_),
	.A2(n14663),
	.B1(FE_OFN16273_n14664),
	.B2(n26243));
   OAI21xp5_ASAP7_75t_SL U13741 (.Y(n639),
	.A1(n16235),
	.A2(n16234),
	.B(n16233));
   OAI21xp33_ASAP7_75t_L U13742 (.Y(n16255),
	.A1(n16252),
	.A2(n16251),
	.B(n16253));
   OAI21x1_ASAP7_75t_SL U13746 (.Y(n26843),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OFN28565_n26845),
	.B(n26844));
   OAI22x1_ASAP7_75t_SL U13748 (.Y(n16151),
	.A1(w2_7_),
	.A2(n16125),
	.B1(n16152),
	.B2(n16125));
   OAI21xp5_ASAP7_75t_L U13750 (.Y(n24637),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OCPN29365_n24639),
	.B(n24638));
   OAI22xp5_ASAP7_75t_SL U13751 (.Y(n16182),
	.A1(n24236),
	.A2(n16053),
	.B1(FE_OFN16262_n16052),
	.B2(w1_6_));
   OAI22xp5_ASAP7_75t_SRAM U13752 (.Y(n577),
	.A1(ld),
	.A2(FE_OFN25975_n16217),
	.B1(key_59_),
	.B2(FE_OFN25975_n16217));
   OAI22xp5_ASAP7_75t_L U13753 (.Y(n616),
	.A1(FE_OFN21_n16125),
	.A2(n16083),
	.B1(key_32_),
	.B2(n16083));
   A2O1A1Ixp33_ASAP7_75t_SL U13754 (.Y(n16261),
	.A1(w2_24_),
	.A2(FE_OFN19_n16125),
	.B(n16258),
	.C(n16257));
   OAI21x1_ASAP7_75t_SL U13757 (.Y(n16247),
	.A1(n16243),
	.A2(n27219),
	.B(n16242));
   OAI22xp5_ASAP7_75t_SRAM U13758 (.Y(n598),
	.A1(ld),
	.A2(n16192),
	.B1(key_51_),
	.B2(n16192));
   OAI21xp5_ASAP7_75t_SL U13765 (.Y(n25930),
	.A1(text_in_r_32_),
	.A2(FE_DBTN0_ld_r),
	.B(n25926));
   OAI22xp33_ASAP7_75t_L U13766 (.Y(n574),
	.A1(FE_OFN21_n16125),
	.A2(n16214),
	.B1(key_52_),
	.B2(n16214));
   OAI21xp33_ASAP7_75t_SL U13767 (.Y(n624),
	.A1(n16212),
	.A2(n16211),
	.B(n16210));
   OAI21xp5_ASAP7_75t_L U13768 (.Y(n16233),
	.A1(FE_OFN26072_n26720),
	.A2(FE_OFN21_n16125),
	.B(n16232));
   OAI21xp5_ASAP7_75t_L U13770 (.Y(n16253),
	.A1(w2_16_),
	.A2(n16250),
	.B(n16249));
   OAI21xp5_ASAP7_75t_SL U13771 (.Y(n16257),
	.A1(ld),
	.A2(w2_24_),
	.B(n16258));
   OAI21xp5_ASAP7_75t_L U13772 (.Y(n16210),
	.A1(n16125),
	.A2(FE_OFN16184_w3_9),
	.B(n16209));
   OAI21x1_ASAP7_75t_SL U13773 (.Y(n15916),
	.A1(n15371),
	.A2(n25931),
	.B(n15370));
   OAI21xp33_ASAP7_75t_SL U13774 (.Y(n26038),
	.A1(FE_OFN16213_ld_r),
	.A2(FE_OCPN27462_n26215),
	.B(n26039));
   OAI22xp5_ASAP7_75t_L U13775 (.Y(n562),
	.A1(FE_OFN0_ld),
	.A2(n16104),
	.B1(key_53_),
	.B2(n16104));
   OAI22xp5_ASAP7_75t_SL U13777 (.Y(n535),
	.A1(ld),
	.A2(n16149),
	.B1(key_47_),
	.B2(n16149));
   OAI21xp5_ASAP7_75t_SL U13778 (.Y(n16232),
	.A1(key_20_),
	.A2(FE_OFN26_n16125),
	.B(n16231));
   OAI22xp33_ASAP7_75t_L U13779 (.Y(n529),
	.A1(ld),
	.A2(FE_OFN26154_n16132),
	.B1(key_63_),
	.B2(FE_OFN26154_n16132));
   FAx1_ASAP7_75t_SL U13781 (.SN(n25898),
	.A(FE_OCPN28054_n26501),
	.B(FE_OCPN27366_n26326),
	.CI(n25893));
   A2O1A1Ixp33_ASAP7_75t_SL U13782 (.Y(n15369),
	.A1(FE_OFN26_n16125),
	.A2(FE_OFN16276_w3_5),
	.B(n15368),
	.C(n15776));
   OAI21xp5_ASAP7_75t_SL U13783 (.Y(n16166),
	.A1(n16134),
	.A2(n25841),
	.B(n16133));
   OAI22xp5_ASAP7_75t_L U13784 (.Y(n541),
	.A1(FE_OFN21_n16125),
	.A2(n16198),
	.B1(key_62_),
	.B2(n16198));
   INVx2_ASAP7_75t_SL U13786 (.Y(n26895),
	.A(n25982));
   NAND2x1p5_ASAP7_75t_L U13788 (.Y(n16231),
	.A(FE_OFN22_n16125),
	.B(n16234));
   OAI21xp5_ASAP7_75t_SL U13789 (.Y(n16094),
	.A1(n16091),
	.A2(n25247),
	.B(n16090));
   AOI22x1_ASAP7_75t_SL U13790 (.Y(n16243),
	.A1(w1_18_),
	.A2(n16099),
	.B1(FE_OFN26541_n16100),
	.B2(n24412));
   OAI21xp5_ASAP7_75t_L U13791 (.Y(n16209),
	.A1(key_9_),
	.A2(FE_OFN25_n16125),
	.B(n16208));
   NAND2xp5_ASAP7_75t_SL U13793 (.Y(n26481),
	.A(n26742),
	.B(n26477));
   INVx1_ASAP7_75t_SL U13796 (.Y(n15267),
	.A(n15266));
   NAND2xp5_ASAP7_75t_SL U13797 (.Y(n24177),
	.A(FE_OCPN29470_n24175),
	.B(n24173));
   A2O1A1Ixp33_ASAP7_75t_SL U13798 (.Y(n24523),
	.A1(FE_OFN27069_n24478),
	.A2(n19158),
	.B(n26777),
	.C(n19157));
   OAI21xp5_ASAP7_75t_SL U13799 (.Y(n16265),
	.A1(n16225),
	.A2(n26963),
	.B(n16224));
   INVx1_ASAP7_75t_SRAM U13800 (.Y(n26330),
	.A(FE_OCPN7636_n25940));
   OAI21xp5_ASAP7_75t_SL U13801 (.Y(n16271),
	.A1(n16268),
	.A2(n27173),
	.B(n16267));
   OAI21xp5_ASAP7_75t_SL U13802 (.Y(n16148),
	.A1(n16127),
	.A2(n27085),
	.B(n16126));
   O2A1O1Ixp5_ASAP7_75t_SL U13804 (.Y(n25809),
	.A1(FE_OFN16180_n26542),
	.A2(n18158),
	.B(n25808),
	.C(n25807));
   NAND2xp33_ASAP7_75t_SRAM U13805 (.Y(n24539),
	.A(FE_OFN16263_n25976),
	.B(FE_OFN26546_n24537));
   NAND2xp5_ASAP7_75t_L U13806 (.Y(n24632),
	.A(FE_OCPN29503_n24627),
	.B(n24629));
   A2O1A1Ixp33_ASAP7_75t_SL U13807 (.Y(n24847),
	.A1(n26829),
	.A2(n25005),
	.B(n23962),
	.C(n23961));
   O2A1O1Ixp5_ASAP7_75t_SL U13809 (.Y(n26711),
	.A1(n26710),
	.A2(n26709),
	.B(n26708),
	.C(n26707));
   A2O1A1Ixp33_ASAP7_75t_L U13810 (.Y(n26586),
	.A1(n26282),
	.A2(n26250),
	.B(n25684),
	.C(n25683));
   AOI22x1_ASAP7_75t_SL U13813 (.Y(n16145),
	.A1(w1_17_),
	.A2(FE_OCPN28075_n16048),
	.B1(n16047),
	.B2(n26210));
   NAND2xp33_ASAP7_75t_SL U13814 (.Y(n25446),
	.A(FE_OFN29143_n25444),
	.B(n25697));
   NOR2x1_ASAP7_75t_L U13815 (.Y(n26363),
	.A(n27120),
	.B(FE_OCPN27641_n27121));
   NAND2xp5_ASAP7_75t_SL U13816 (.Y(n24285),
	.A(n26836),
	.B(n24282));
   A2O1A1Ixp33_ASAP7_75t_SL U13817 (.Y(n26205),
	.A1(n27216),
	.A2(n26494),
	.B(n26204),
	.C(n26203));
   AOI22x1_ASAP7_75t_SL U13818 (.Y(n16268),
	.A1(w1_8_),
	.A2(FE_OCPN28186_n16123),
	.B1(n16122),
	.B2(n26932));
   A2O1A1Ixp33_ASAP7_75t_SL U13823 (.Y(n26228),
	.A1(FE_OFN16170_n26637),
	.A2(n26226),
	.B(n26225),
	.C(n26224));
   A2O1A1Ixp33_ASAP7_75t_SL U13824 (.Y(n25343),
	.A1(FE_OFN16177_n27207),
	.A2(n26057),
	.B(n26054),
	.C(n25923));
   NAND2xp5_ASAP7_75t_SL U13826 (.Y(n26005),
	.A(FE_OFN25911_n26491),
	.B(n26190));
   NAND2xp5_ASAP7_75t_L U13827 (.Y(n26195),
	.A(FE_OFN28615_n26191),
	.B(n26190));
   A2O1A1Ixp33_ASAP7_75t_L U13830 (.Y(n24745),
	.A1(n26819),
	.A2(n26725),
	.B(n26722),
	.C(n24744));
   NAND2xp33_ASAP7_75t_SL U13831 (.Y(n25925),
	.A(FE_OFN104_n27179),
	.B(n25922));
   NAND2xp33_ASAP7_75t_L U13832 (.Y(n24343),
	.A(FE_OFN29011_n27113),
	.B(n24340));
   AOI22x1_ASAP7_75t_SL U13833 (.Y(n16179),
	.A1(w1_12_),
	.A2(FE_OFN25929_n16073),
	.B1(FE_OCPN29386_n16073),
	.B2(n25128));
   INVx1_ASAP7_75t_SL U13840 (.Y(n26190),
	.A(n26192));
   A2O1A1Ixp33_ASAP7_75t_SL U13843 (.Y(n25858),
	.A1(FE_OFN16176_n27207),
	.A2(n26196),
	.B(FE_OCPN27583_n26193),
	.C(n25857));
   A2O1A1Ixp33_ASAP7_75t_SL U13844 (.Y(n14745),
	.A1(FE_OFN16411_n15884),
	.A2(n13798),
	.B(n13797),
	.C(n13796));
   NAND2xp5_ASAP7_75t_SL U13847 (.Y(n24811),
	.A(FE_OFN27169_n26683),
	.B(n24807));
   A2O1A1Ixp33_ASAP7_75t_SL U13850 (.Y(n16073),
	.A1(FE_OFN16411_n15884),
	.A2(n14894),
	.B(n14893),
	.C(n14892));
   A2O1A1Ixp33_ASAP7_75t_SL U13853 (.Y(n16088),
	.A1(n15896),
	.A2(n15059),
	.B(n15058),
	.C(n15057));
   O2A1O1Ixp5_ASAP7_75t_SL U13856 (.Y(n22652),
	.A1(n22651),
	.A2(n22650),
	.B(n26584),
	.C(n22649));
   INVxp67_ASAP7_75t_L U13858 (.Y(n24209),
	.A(n24211));
   A2O1A1Ixp33_ASAP7_75t_SL U13860 (.Y(n13722),
	.A1(n13707),
	.A2(n13706),
	.B(n14585),
	.C(n13705));
   O2A1O1Ixp33_ASAP7_75t_SL U13861 (.Y(n26867),
	.A1(n21417),
	.A2(n26083),
	.B(n26082),
	.C(n26081));
   A2O1A1Ixp33_ASAP7_75t_SL U13864 (.Y(n16123),
	.A1(n15896),
	.A2(n15656),
	.B(n15655),
	.C(n15654));
   NAND2xp5_ASAP7_75t_L U13865 (.Y(n19147),
	.A(n19146),
	.B(FE_OCPN4686_n19142));
   NAND2xp5_ASAP7_75t_L U13868 (.Y(n19148),
	.A(n19143),
	.B(FE_OCPN4686_n19142));
   NOR3x1_ASAP7_75t_SL U13877 (.Y(n25751),
	.A(n22477),
	.B(n22476),
	.C(n22475));
   NOR3x1_ASAP7_75t_SL U13883 (.Y(n25733),
	.A(n22961),
	.B(n22960),
	.C(n22959));
   NAND2xp5_ASAP7_75t_SL U13884 (.Y(n13472),
	.A(n13471),
	.B(n13470));
   INVxp67_ASAP7_75t_SL U13886 (.Y(n14402),
	.A(n14403));
   NAND2xp33_ASAP7_75t_SL U13887 (.Y(n20322),
	.A(n20317),
	.B(n20319));
   NAND3xp33_ASAP7_75t_SL U13888 (.Y(n19375),
	.A(n24164),
	.B(n19371),
	.C(n19370));
   A2O1A1Ixp33_ASAP7_75t_SL U13889 (.Y(n25563),
	.A1(n19391),
	.A2(n19390),
	.B(n26959),
	.C(n19389));
   NAND2xp5_ASAP7_75t_SL U13891 (.Y(n23461),
	.A(n21334),
	.B(n21039));
   NAND2xp5_ASAP7_75t_L U13892 (.Y(n19735),
	.A(n19734),
	.B(n19733));
   NAND3xp33_ASAP7_75t_SL U13894 (.Y(n14467),
	.A(n14465),
	.B(n14464),
	.C(n14463));
   A2O1A1Ixp33_ASAP7_75t_SL U13895 (.Y(n15892),
	.A1(n15890),
	.A2(n15889),
	.B(FE_OFN28682_n15888),
	.C(n15887));
   NAND2xp5_ASAP7_75t_SL U13898 (.Y(n21472),
	.A(n17292),
	.B(n17291));
   O2A1O1Ixp33_ASAP7_75t_L U13904 (.Y(n14963),
	.A1(n14962),
	.A2(n14961),
	.B(n16042),
	.C(n14960));
   NAND2xp5_ASAP7_75t_SL U13905 (.Y(n19371),
	.A(n19369),
	.B(n19368));
   A2O1A1Ixp33_ASAP7_75t_L U13906 (.Y(n17232),
	.A1(n19694),
	.A2(n17215),
	.B(n25139),
	.C(n17214));
   NOR3xp33_ASAP7_75t_SL U13908 (.Y(n22154),
	.A(n22150),
	.B(n22149),
	.C(n22148));
   NOR3xp33_ASAP7_75t_SL U13909 (.Y(n19900),
	.A(n19898),
	.B(n22692),
	.C(n20335));
   NOR3xp33_ASAP7_75t_SL U13910 (.Y(n23368),
	.A(n23367),
	.B(n24545),
	.C(n23366));
   NOR3x1_ASAP7_75t_SL U13913 (.Y(n24571),
	.A(n17504),
	.B(FE_OCPN27807_n23375),
	.C(n17503));
   NOR3xp33_ASAP7_75t_SL U13919 (.Y(n25289),
	.A(n25288),
	.B(n25990),
	.C(n25287));
   NOR3x1_ASAP7_75t_SL U13920 (.Y(n17080),
	.A(n17076),
	.B(n17100),
	.C(n18918));
   INVx1_ASAP7_75t_SL U13921 (.Y(n13468),
	.A(n13465));
   NAND2xp5_ASAP7_75t_L U13922 (.Y(n17755),
	.A(n17751),
	.B(n17752));
   NOR3xp33_ASAP7_75t_SL U13923 (.Y(n23687),
	.A(n18559),
	.B(FE_OFN28921_n20660),
	.C(n20643));
   NOR3xp33_ASAP7_75t_SL U13924 (.Y(n20084),
	.A(n20082),
	.B(FE_OCPN28156_n26304),
	.C(n21990));
   NAND3xp33_ASAP7_75t_SL U13926 (.Y(n17076),
	.A(n17075),
	.B(n17074),
	.C(n20497));
   NAND3xp33_ASAP7_75t_SL U13927 (.Y(n19459),
	.A(n18050),
	.B(n18049),
	.C(n23454));
   NOR2xp33_ASAP7_75t_SL U13929 (.Y(n13756),
	.A(n15787),
	.B(n13760));
   NOR3x1_ASAP7_75t_SL U13930 (.Y(n18271),
	.A(n18270),
	.B(n18269),
	.C(n19435));
   NOR2xp33_ASAP7_75t_SL U13931 (.Y(n13763),
	.A(n13761),
	.B(n13760));
   OAI22xp33_ASAP7_75t_SL U13932 (.Y(n14888),
	.A1(n15896),
	.A2(n14887),
	.B1(n14886),
	.B2(n14887));
   NAND2xp5_ASAP7_75t_SL U13933 (.Y(n17644),
	.A(n17643),
	.B(n17642));
   NAND2xp5_ASAP7_75t_SL U13937 (.Y(n19471),
	.A(n19469),
	.B(n19468));
   NAND2xp33_ASAP7_75t_L U13938 (.Y(n20939),
	.A(n20936),
	.B(n20937));
   NOR2x1_ASAP7_75t_SL U13939 (.Y(n17429),
	.A(n16688),
	.B(n16687));
   NOR3x1_ASAP7_75t_SL U13940 (.Y(n21382),
	.A(n19203),
	.B(n21344),
	.C(n23246));
   NAND3xp33_ASAP7_75t_L U13941 (.Y(n20067),
	.A(n21933),
	.B(n16519),
	.C(n16518));
   NOR2xp33_ASAP7_75t_SL U13943 (.Y(n23003),
	.A(n23515),
	.B(n23001));
   OAI22xp33_ASAP7_75t_SL U13944 (.Y(n23004),
	.A1(FE_OFN29026_n20911),
	.A2(n22996),
	.B1(FE_OFN28752_n),
	.B2(n22996));
   NAND3xp33_ASAP7_75t_SL U13945 (.Y(n17099),
	.A(FE_OFN28913_n18247),
	.B(FE_OCPN29568_n18257),
	.C(n25882));
   NOR2xp33_ASAP7_75t_SL U13946 (.Y(n14863),
	.A(n15896),
	.B(n14887));
   NOR3x1_ASAP7_75t_SL U13948 (.Y(n26080),
	.A(n21354),
	.B(n21373),
	.C(n22511));
   NAND3x1_ASAP7_75t_SL U13949 (.Y(n19882),
	.A(n19881),
	.B(n19880),
	.C(n19879));
   NAND2xp5_ASAP7_75t_SL U13950 (.Y(n17089),
	.A(n17007),
	.B(n17006));
   NOR2xp33_ASAP7_75t_L U13951 (.Y(n16491),
	.A(n16508),
	.B(n21962));
   NAND3xp33_ASAP7_75t_SL U13952 (.Y(n23051),
	.A(n16650),
	.B(n16649),
	.C(n19689));
   NAND2xp5_ASAP7_75t_SL U13954 (.Y(n17287),
	.A(n17283),
	.B(n17284));
   NOR3xp33_ASAP7_75t_SL U13955 (.Y(n18941),
	.A(n17097),
	.B(n25885),
	.C(FE_OFN28559_n18278));
   NAND2xp5_ASAP7_75t_L U13956 (.Y(n15122),
	.A(n15121),
	.B(n15120));
   NAND2xp5_ASAP7_75t_SL U13957 (.Y(n17286),
	.A(n17285),
	.B(n17284));
   NAND3xp33_ASAP7_75t_SL U13958 (.Y(n18641),
	.A(n18639),
	.B(n21167),
	.C(n21168));
   NOR3xp33_ASAP7_75t_SL U13960 (.Y(n22646),
	.A(n18391),
	.B(n18467),
	.C(n18390));
   NAND3xp33_ASAP7_75t_L U13961 (.Y(n21302),
	.A(n21300),
	.B(n21299),
	.C(n21298));
   NAND2xp5_ASAP7_75t_SL U13962 (.Y(n18870),
	.A(n21275),
	.B(n18866));
   NAND2xp5_ASAP7_75t_L U13963 (.Y(n22027),
	.A(n22026),
	.B(n22025));
   NAND2x1_ASAP7_75t_SL U13964 (.Y(n20212),
	.A(n21002),
	.B(n20171));
   NOR2x1_ASAP7_75t_SL U13965 (.Y(n18748),
	.A(n19106),
	.B(n18741));
   NOR3xp33_ASAP7_75t_L U13966 (.Y(n16509),
	.A(n16508),
	.B(FE_OFN28549_n21934),
	.C(n16507));
   NAND3xp33_ASAP7_75t_SL U13967 (.Y(n25544),
	.A(n25995),
	.B(n18254),
	.C(n17028));
   NOR2x1_ASAP7_75t_SL U13970 (.Y(n17285),
	.A(n17245),
	.B(n19594));
   OAI22xp33_ASAP7_75t_L U13973 (.Y(n13563),
	.A1(n15188),
	.A2(n13413),
	.B1(FE_OCPN27656_w3_25),
	.B2(n13413));
   OAI22xp5_ASAP7_75t_L U13976 (.Y(n13914),
	.A1(FE_OFN28628_n15667),
	.A2(n13903),
	.B1(n14798),
	.B2(n13903));
   NAND2xp5_ASAP7_75t_L U13977 (.Y(n21380),
	.A(n21379),
	.B(n21378));
   NAND3xp33_ASAP7_75t_SL U13979 (.Y(n16322),
	.A(n20873),
	.B(n20856),
	.C(n21938));
   NAND3xp33_ASAP7_75t_SRAM U13980 (.Y(n19606),
	.A(FE_OCPN29553_n19602),
	.B(n21473),
	.C(n19601));
   NAND3xp33_ASAP7_75t_SL U13981 (.Y(n18557),
	.A(n23804),
	.B(n21638),
	.C(n23750));
   NOR3xp33_ASAP7_75t_SL U13984 (.Y(n23140),
	.A(n16645),
	.B(n17203),
	.C(n16644));
   NAND3x1_ASAP7_75t_SL U13985 (.Y(n18267),
	.A(n25994),
	.B(n24165),
	.C(n17017));
   AND3x2_ASAP7_75t_SL U13986 (.Y(n21004),
	.A(n22892),
	.B(n22891),
	.C(n19261));
   NOR3xp33_ASAP7_75t_SL U13987 (.Y(n25562),
	.A(n17105),
	.B(n19411),
	.C(n17104));
   NAND2xp33_ASAP7_75t_L U13988 (.Y(n16343),
	.A(n16359),
	.B(n18068));
   NAND2xp5_ASAP7_75t_L U13989 (.Y(n23804),
	.A(n18556),
	.B(n18555));
   OAI22xp5_ASAP7_75t_L U13990 (.Y(n14712),
	.A1(FE_OCPN29536_FE_OFN8_w3_14),
	.A2(n14098),
	.B1(FE_OCPN28296_n15386),
	.B2(n14098));
   NAND2xp5_ASAP7_75t_L U13991 (.Y(n26165),
	.A(n22021),
	.B(n18990));
   OAI22xp33_ASAP7_75t_L U13993 (.Y(n18695),
	.A1(n21553),
	.A2(n22436),
	.B1(FE_OCPN29409_n22461),
	.B2(n22436));
   NAND2xp5_ASAP7_75t_SL U13996 (.Y(n14951),
	.A(n13977),
	.B(n13976));
   NOR2x1_ASAP7_75t_L U13998 (.Y(n19201),
	.A(FE_OCPN27496_n21820),
	.B(n19198));
   OAI21xp33_ASAP7_75t_SL U13999 (.Y(n21415),
	.A1(FE_OCPN29378_n23266),
	.A2(FE_OCPN28447_n23392),
	.B(n19197));
   NAND3x1_ASAP7_75t_SL U14000 (.Y(n21875),
	.A(n19647),
	.B(n19646),
	.C(n19775));
   OAI21xp5_ASAP7_75t_L U14001 (.Y(n14429),
	.A1(n15568),
	.A2(n15808),
	.B(n14426));
   NOR2x1_ASAP7_75t_SL U14002 (.Y(n15045),
	.A(n14855),
	.B(FE_OFN28691_n13725));
   NAND2xp5_ASAP7_75t_SL U14003 (.Y(n17027),
	.A(n19372),
	.B(n17117));
   NAND2xp5_ASAP7_75t_L U14004 (.Y(n18287),
	.A(FE_OFN29035_n17116),
	.B(n18284));
   INVx2_ASAP7_75t_L U14006 (.Y(n15595),
	.A(n14417));
   OAI22xp5_ASAP7_75t_SL U14007 (.Y(n21412),
	.A1(FE_OCPN29435_n17445),
	.A2(n23262),
	.B1(FE_OCPN27730_n17464),
	.B2(n23262));
   OA21x2_ASAP7_75t_SRAM U14008 (.Y(n20855),
	.A1(n20854),
	.A2(n20853),
	.B(n25322));
   OAI22xp33_ASAP7_75t_L U14013 (.Y(n20200),
	.A1(n17757),
	.A2(n20168),
	.B1(n17808),
	.B2(n20168));
   NAND2xp5_ASAP7_75t_L U14015 (.Y(n17852),
	.A(FE_OCPN27642_n16758),
	.B(FE_OCPN28298_n));
   NAND2xp5_ASAP7_75t_L U14016 (.Y(n23501),
	.A(FE_OCPN29374_FE_OFN29191_sa23_2),
	.B(n20903));
   NAND2x1p5_ASAP7_75t_SL U14018 (.Y(n18015),
	.A(FE_OFN29123_n),
	.B(n21317));
   NOR2xp33_ASAP7_75t_L U14019 (.Y(n16495),
	.A(FE_OCPN28394_FE_OFN27043_n),
	.B(n16397));
   NOR2x1_ASAP7_75t_L U14020 (.Y(n19411),
	.A(n17002),
	.B(FE_OFN28738_n16989));
   OA21x2_ASAP7_75t_SL U14021 (.Y(n18046),
	.A1(n21304),
	.A2(n21752),
	.B(FE_OFN29158_n18860));
   OAI22xp33_ASAP7_75t_SL U14022 (.Y(n15542),
	.A1(n15541),
	.A2(n15540),
	.B1(FE_OFN26614_n),
	.B2(n15540));
   OAI22xp5_ASAP7_75t_L U14024 (.Y(n18811),
	.A1(n22392),
	.A2(n24855),
	.B1(FE_OCPN28229_n17529),
	.B2(n24855));
   NAND2xp5_ASAP7_75t_L U14027 (.Y(n14693),
	.A(FE_OFN28758_n15422),
	.B(n14157));
   NOR2xp67_ASAP7_75t_L U14030 (.Y(n22751),
	.A(n19502),
	.B(n23217));
   OAI22xp5_ASAP7_75t_L U14032 (.Y(n23176),
	.A1(n18162),
	.A2(n21117),
	.B1(n23315),
	.B2(n21117));
   OAI22xp33_ASAP7_75t_SRAM U14033 (.Y(n13452),
	.A1(FE_OFN16193_n15200),
	.A2(n13451),
	.B1(FE_OFN28604_n14534),
	.B2(n13451));
   NAND2xp5_ASAP7_75t_R U14034 (.Y(n16004),
	.A(n14695),
	.B(n15956));
   NAND2xp5_ASAP7_75t_SL U14035 (.Y(n20540),
	.A(n22256),
	.B(n20561));
   NOR2x1_ASAP7_75t_SL U14036 (.Y(n19839),
	.A(FE_OCPN27951_n19098),
	.B(n19097));
   INVx2_ASAP7_75t_SL U14037 (.Y(n21120),
	.A(n20720));
   NOR3xp33_ASAP7_75t_R U14038 (.Y(n15093),
	.A(n13725),
	.B(FE_OCPN29537_FE_OFN28699_w3_6),
	.C(n13736));
   NOR2x1p5_ASAP7_75t_L U14041 (.Y(n24694),
	.A(n18166),
	.B(n23160));
   INVx2_ASAP7_75t_SL U14042 (.Y(n18739),
	.A(n17251));
   NOR2x1_ASAP7_75t_L U14043 (.Y(n23267),
	.A(FE_OCPN27601_n17475),
	.B(n19166));
   NAND2x1p5_ASAP7_75t_SL U14044 (.Y(n17330),
	.A(FE_OFN16141_sa01_3),
	.B(n26456));
   OAI22xp33_ASAP7_75t_SL U14047 (.Y(n21425),
	.A1(n17445),
	.A2(n21860),
	.B1(FE_OCPN27562_n17447),
	.B2(n21860));
   OAI22xp5_ASAP7_75t_L U14050 (.Y(n15810),
	.A1(n15034),
	.A2(n15636),
	.B1(FE_OFN28747_n),
	.B2(n15636));
   OAI22xp33_ASAP7_75t_R U14052 (.Y(n15600),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(n15860),
	.B1(FE_OFN28732_n),
	.B2(n15860));
   NOR2x1p5_ASAP7_75t_SL U14058 (.Y(n16978),
	.A(FE_OFN28862_n),
	.B(n17103));
   NAND2xp33_ASAP7_75t_SRAM U14059 (.Y(n14945),
	.A(n15972),
	.B(FE_OFN28574_n16016));
   NAND2x1_ASAP7_75t_SL U14060 (.Y(n16000),
	.A(FE_OFN26641_w3_14),
	.B(FE_PSN8324_n15987));
   NAND2x1p5_ASAP7_75t_SL U14061 (.Y(n17251),
	.A(FE_OCPN27818_n17267),
	.B(n17265));
   NAND2x1p5_ASAP7_75t_SL U14062 (.Y(n18767),
	.A(n17265),
	.B(FE_OFN42_sa00_0));
   NAND2xp5_ASAP7_75t_SL U14064 (.Y(n17998),
	.A(FE_OCPN27726_n),
	.B(n21304));
   OAI21xp33_ASAP7_75t_SRAM U14065 (.Y(n26832),
	.A1(text_in_r_23_),
	.A2(FE_OCPN29502_w3_23),
	.B(n26830));
   NOR2x1_ASAP7_75t_SL U14066 (.Y(n19399),
	.A(FE_OFN28479_sa13_2),
	.B(n19360));
   NAND2xp5_ASAP7_75t_SL U14067 (.Y(n19981),
	.A(n19979),
	.B(FE_OFN25993_n16767));
   NOR2x1p5_ASAP7_75t_L U14069 (.Y(n17606),
	.A(FE_OCPN29431_sa30_3),
	.B(n21627));
   NAND2xp5_ASAP7_75t_SL U14070 (.Y(n26026),
	.A(FE_OFN28895_sa30_2),
	.B(n17637));
   NOR2x1_ASAP7_75t_L U14073 (.Y(n15757),
	.A(FE_OFN28701_w3_16),
	.B(n23974));
   NAND2x1p5_ASAP7_75t_L U14074 (.Y(n15969),
	.A(w3_10_),
	.B(FE_OFN25961_w3_8));
   NOR2x1p5_ASAP7_75t_SL U14075 (.Y(n25869),
	.A(FE_OFN28725_n16982),
	.B(n17065));
   NAND2xp5_ASAP7_75t_L U14076 (.Y(n15994),
	.A(n24755),
	.B(n15922));
   NOR2x1p5_ASAP7_75t_SL U14077 (.Y(n15857),
	.A(FE_OFN29052_w3_5),
	.B(FE_OCPN29500_FE_OFN28662_w3_7));
   OAI22xp33_ASAP7_75t_SRAM U14079 (.Y(n25427),
	.A1(FE_OFN16179_w3_19),
	.A2(FE_OFN28489_ld_r),
	.B1(text_in_r_19_),
	.B2(FE_OFN28489_ld_r));
   NOR3xp33_ASAP7_75t_L U14080 (.Y(n13459),
	.A(FE_OCPN29350_w3_25),
	.B(FE_OFN27206_w3_30),
	.C(n25675));
   OAI22xp33_ASAP7_75t_SRAM U14081 (.Y(n25960),
	.A1(text_in_r_21_),
	.A2(FE_OFN28489_ld_r),
	.B1(n25961),
	.B2(FE_OFN28489_ld_r));
   NOR2xp33_ASAP7_75t_SL U14082 (.Y(n18165),
	.A(sa22_3_),
	.B(n18164));
   NAND2x1_ASAP7_75t_SL U14083 (.Y(n16329),
	.A(FE_OFN26095_n16293),
	.B(FE_OFN26096_n16294));
   NAND2x2_ASAP7_75t_SL U14084 (.Y(n21818),
	.A(n21844),
	.B(FE_OCPN27241_sa11_1));
   NOR2x1_ASAP7_75t_SL U14086 (.Y(n22505),
	.A(FE_OFN138_sa11_0),
	.B(n17489));
   NOR2x1p5_ASAP7_75t_SL U14088 (.Y(n18707),
	.A(FE_OFN28672_sa01_2),
	.B(FE_OFN125_sa01_1));
   NAND2x2_ASAP7_75t_SL U14089 (.Y(n18693),
	.A(FE_OCPN27423_sa01_0),
	.B(n17359));
   NOR3x1_ASAP7_75t_SL U14090 (.Y(n25102),
	.A(n18379),
	.B(n17601),
	.C(FE_OFN16200_sa30_2));
   NOR2x1p5_ASAP7_75t_SL U14091 (.Y(n27117),
	.A(sa22_6_),
	.B(n22300));
   NOR2x1p5_ASAP7_75t_SL U14093 (.Y(n17265),
	.A(FE_OFN28744_FE_OCPN27908),
	.B(FE_OFN148_sa00_1));
   NAND2x2_ASAP7_75t_SL U14094 (.Y(n17275),
	.A(FE_OFN29172_sa00_4),
	.B(n19834));
   NAND2x1_ASAP7_75t_SL U14095 (.Y(n17744),
	.A(FE_OCPN27261_sa02_0),
	.B(n22882));
   NOR2x1p5_ASAP7_75t_SL U14098 (.Y(n18521),
	.A(FE_OCPN27557_sa20_4),
	.B(FE_OFN29150_sa20_5));
   NOR2x1p5_ASAP7_75t_SL U14099 (.Y(n17761),
	.A(n17763),
	.B(FE_OCPN27566_FE_OFN16138_sa02_5));
   NAND2x1p5_ASAP7_75t_L U14104 (.Y(n19011),
	.A(FE_OCPN27803_sa23_4),
	.B(FE_OFN27078_sa23_5));
   NAND2x1p5_ASAP7_75t_SL U14108 (.Y(n16581),
	.A(FE_OFN27196_n),
	.B(FE_OFN130_sa10_5));
   NOR2x1p5_ASAP7_75t_SL U14110 (.Y(n21327),
	.A(FE_OFN28689_sa03_5),
	.B(FE_OCPN27405_sa03_4));
   NAND2xp5_ASAP7_75t_SL U14112 (.Y(n16278),
	.A(FE_OFN28699_w3_6),
	.B(n16276));
   A2O1A1Ixp33_ASAP7_75t_SL U14114 (.Y(n524),
	.A1(n26696),
	.A2(n26695),
	.B(n26694),
	.C(n26693));
   OAI21xp5_ASAP7_75t_SL U14116 (.Y(n653),
	.A1(n16156),
	.A2(FE_OCPN29500_FE_OFN28662_w3_7),
	.B(n16155));
   NAND3xp33_ASAP7_75t_SL U14117 (.Y(n26797),
	.A(FE_OFN25881_w3_24),
	.B(n26800),
	.C(n26799));
   NAND3xp33_ASAP7_75t_SL U14119 (.Y(n26473),
	.A(n26474),
	.B(n26476),
	.C(n26475));
   A2O1A1Ixp33_ASAP7_75t_SL U14120 (.Y(n26476),
	.A1(n26472),
	.A2(FE_OFN28487_ld_r),
	.B(n26471),
	.C(n26470));
   O2A1O1Ixp5_ASAP7_75t_SL U14123 (.Y(n359),
	.A1(w1_19_),
	.A2(text_in_r_83_),
	.B(n25760),
	.C(n25759));
   A2O1A1Ixp33_ASAP7_75t_SL U14124 (.Y(n26390),
	.A1(n26769),
	.A2(n26770),
	.B(n26766),
	.C(FE_OCPN27310_n26389));
   OAI22xp33_ASAP7_75t_SL U14126 (.Y(n586),
	.A1(ld),
	.A2(n16244),
	.B1(key_50_),
	.B2(n16244));
   A2O1A1Ixp33_ASAP7_75t_SL U14127 (.Y(n25249),
	.A1(FE_OCPN28138_n26654),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B(n25245),
	.C(n25244));
   FAx1_ASAP7_75t_SL U14128 (.SN(n25984),
	.A(FE_OCPN27525_n26434),
	.B(FE_OCPN27514_n25981),
	.CI(n25980));
   NAND3xp33_ASAP7_75t_SL U14129 (.Y(n26820),
	.A(n26822),
	.B(n26823),
	.C(n26821));
   O2A1O1Ixp33_ASAP7_75t_SL U14131 (.Y(n26785),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OFN26024_n26115),
	.B(n26783),
	.C(n26782));
   NAND2xp5_ASAP7_75t_SL U14132 (.Y(n26985),
	.A(n27144),
	.B(n26986));
   OAI22xp5_ASAP7_75t_L U14133 (.Y(n592),
	.A1(ld),
	.A2(n15917),
	.B1(key_33_),
	.B2(n15917));
   A2O1A1Ixp33_ASAP7_75t_SL U14134 (.Y(n16239),
	.A1(FE_OFN28472_ld),
	.A2(FE_OFN28858_FE_OCPN27664_w3_25),
	.B(n16238),
	.C(FE_OFN25892_n16264));
   AOI22xp5_ASAP7_75t_L U14135 (.Y(n24535),
	.A1(FE_OCPN27274_n26394),
	.A2(n24531),
	.B1(FE_OFN48_w0_2),
	.B2(n24514));
   NOR3xp33_ASAP7_75t_SL U14136 (.Y(n27184),
	.A(FE_OFN116_n27187),
	.B(n27185),
	.C(n27186));
   A2O1A1Ixp33_ASAP7_75t_SL U14137 (.Y(n26414),
	.A1(n26412),
	.A2(FE_OCPN29443_n25507),
	.B(FE_OCPN7589_n26420),
	.C(n26410));
   A2O1A1Ixp33_ASAP7_75t_SL U14138 (.Y(n26851),
	.A1(n17580),
	.A2(n24830),
	.B(n24829),
	.C(n24828));
   A2O1A1Ixp33_ASAP7_75t_SL U14139 (.Y(n26658),
	.A1(FE_OCPN28138_n26654),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B(n26653),
	.C(n26652));
   INVx1_ASAP7_75t_L U14140 (.Y(n15917),
	.A(n15916));
   OAI22xp33_ASAP7_75t_L U14142 (.Y(n556),
	.A1(ld),
	.A2(n15777),
	.B1(key_37_),
	.B2(n15777));
   OAI21xp33_ASAP7_75t_L U14143 (.Y(n26947),
	.A1(FE_OFN1_ld_r),
	.A2(n27143),
	.B(n26948));
   A2O1A1Ixp33_ASAP7_75t_SL U14144 (.Y(n26043),
	.A1(FE_OCPN27462_n26215),
	.A2(FE_OFN28487_ld_r),
	.B(n26039),
	.C(n26038));
   OAI21xp5_ASAP7_75t_SL U14145 (.Y(n645),
	.A1(n15776),
	.A2(FE_OFN16276_w3_5),
	.B(n15369));
   FAx1_ASAP7_75t_SL U14148 (.SN(n26098),
	.A(FE_OFN28968_n26780),
	.B(FE_OCPN27941_n),
	.CI(n26092));
   OAI22xp33_ASAP7_75t_SL U14149 (.Y(n565),
	.A1(FE_OFN21_n16125),
	.A2(FE_OFN26121_n16107),
	.B1(key_60_),
	.B2(FE_OFN26121_n16107));
   NAND2xp5_ASAP7_75t_SL U14150 (.Y(n24525),
	.A(n24522),
	.B(FE_OFN26546_n24537));
   A2O1A1Ixp33_ASAP7_75t_SL U14151 (.Y(n27210),
	.A1(FE_OFN16177_n27207),
	.A2(n27206),
	.B(n27205),
	.C(n27204));
   FAx1_ASAP7_75t_SL U14152 (.SN(n26230),
	.A(FE_OCPN27374_n26394),
	.B(n26228),
	.CI(FE_OCPN27678_n26227));
   OAI22xp33_ASAP7_75t_L U14153 (.Y(n619),
	.A1(n16125),
	.A2(n16200),
	.B1(key_41_),
	.B2(n16200));
   A2O1A1Ixp33_ASAP7_75t_SL U14155 (.Y(n26809),
	.A1(n27062),
	.A2(n27061),
	.B(n24482),
	.C(n24481));
   A2O1A1Ixp33_ASAP7_75t_SL U14156 (.Y(n16052),
	.A1(n15271),
	.A2(n15270),
	.B(n15269),
	.C(n15268));
   NOR2xp67_ASAP7_75t_SL U14158 (.Y(n26444),
	.A(n26445),
	.B(n26443));
   NAND2xp5_ASAP7_75t_SL U14159 (.Y(n25703),
	.A(n27031),
	.B(n25704));
   FAx1_ASAP7_75t_SL U14161 (.SN(n24987),
	.A(FE_OCPN28311_n26789),
	.B(n24982),
	.CI(FE_OCPN27497_n25431));
   A2O1A1Ixp33_ASAP7_75t_SL U14162 (.Y(n24686),
	.A1(n26823),
	.A2(n26822),
	.B(FE_OCPN27505_n24684),
	.C(n24683));
   INVx1_ASAP7_75t_L U14163 (.Y(n16202),
	.A(n16201));
   FAx1_ASAP7_75t_SL U14164 (.SN(n27109),
	.A(FE_OCPN27235_n27143),
	.B(FE_OCPN29258_n27171),
	.CI(n27103));
   O2A1O1Ixp33_ASAP7_75t_SL U14165 (.Y(n25409),
	.A1(FE_PSN8314_n25722),
	.A2(n25406),
	.B(n25488),
	.C(n25405));
   O2A1O1Ixp33_ASAP7_75t_SL U14166 (.Y(n26039),
	.A1(n26037),
	.A2(n26036),
	.B(FE_OCPN8225_n26172),
	.C(n26035));
   O2A1O1Ixp5_ASAP7_75t_SL U14168 (.Y(n27083),
	.A1(n27081),
	.A2(FE_OCPN28438_n27080),
	.B(FE_OCPN27391_n27079),
	.C(n27078));
   NOR3xp33_ASAP7_75t_SL U14170 (.Y(n25482),
	.A(FE_OCPN27723_n),
	.B(n25483),
	.C(n25484));
   A2O1A1Ixp33_ASAP7_75t_SL U14173 (.Y(n26394),
	.A1(n26082),
	.A2(n24633),
	.B(n24513),
	.C(n24512));
   INVxp67_ASAP7_75t_SL U14174 (.Y(n16266),
	.A(n16265));
   AOI22x1_ASAP7_75t_SL U14177 (.Y(n15902),
	.A1(w1_2_),
	.A2(n14007),
	.B1(FE_OFN16254_n14008),
	.B2(n26185));
   XNOR2x2_ASAP7_75t_SL U14181 (.Y(n16234),
	.A(w2_20_),
	.B(n16213));
   NAND2xp33_ASAP7_75t_SL U14182 (.Y(n25522),
	.A(n26197),
	.B(n26496));
   XNOR2x2_ASAP7_75t_SL U14183 (.Y(n16119),
	.A(u0_rcon_29_),
	.B(n14823));
   A2O1A1Ixp33_ASAP7_75t_L U14184 (.Y(n24933),
	.A1(n26819),
	.A2(n26818),
	.B(n26815),
	.C(n24932));
   A2O1A1Ixp33_ASAP7_75t_L U14186 (.Y(n24115),
	.A1(n26769),
	.A2(n26770),
	.B(n26766),
	.C(FE_OFN29227_n24510));
   NAND3xp33_ASAP7_75t_SL U14187 (.Y(n24599),
	.A(n24600),
	.B(n24602),
	.C(n24601));
   NAND2xp5_ASAP7_75t_SL U14188 (.Y(n16208),
	.A(FE_OFN28462_ld),
	.B(n16211));
   NAND2x1_ASAP7_75t_L U14190 (.Y(n16203),
	.A(FE_OFN28472_ld),
	.B(n16206));
   OR2x2_ASAP7_75t_L U14192 (.Y(n26927),
	.A(FE_OFN16213_ld_r),
	.B(FE_OCPN29576_n26930));
   NAND2xp5_ASAP7_75t_SL U14194 (.Y(n24513),
	.A(FE_OCPN29503_n24627),
	.B(n24510));
   A2O1A1Ixp33_ASAP7_75t_SL U14196 (.Y(n14008),
	.A1(n15271),
	.A2(n13409),
	.B(n13408),
	.C(n13407));
   NAND2xp33_ASAP7_75t_SL U14198 (.Y(n24583),
	.A(n25167),
	.B(n24807));
   NAND2x1_ASAP7_75t_L U14200 (.Y(n25538),
	.A(FE_OFN26558_n26911),
	.B(FE_OFN16340_n26317));
   NOR2xp33_ASAP7_75t_SL U14201 (.Y(n14604),
	.A(w0_7_),
	.B(n14601));
   O2A1O1Ixp33_ASAP7_75t_SL U14203 (.Y(n15266),
	.A1(n15265),
	.A2(n15264),
	.B(n15263),
	.C(n15262));
   A2O1A1Ixp33_ASAP7_75t_SL U14207 (.Y(n26638),
	.A1(n27117),
	.A2(n27052),
	.B(n25614),
	.C(n25613));
   A2O1A1Ixp33_ASAP7_75t_SL U14208 (.Y(n16100),
	.A1(n16042),
	.A2(n15469),
	.B(n15468),
	.C(n15467));
   NAND2xp5_ASAP7_75t_SL U14209 (.Y(n24934),
	.A(n24931),
	.B(FE_OFN16271_n26814));
   AOI22x1_ASAP7_75t_SL U14210 (.Y(n15910),
	.A1(w1_3_),
	.A2(n14090),
	.B1(FE_OFN27216_n14091),
	.B2(n26578));
   A2O1A1Ixp33_ASAP7_75t_SL U14211 (.Y(n24878),
	.A1(n26819),
	.A2(FE_OCPN8227_n25950),
	.B(n25947),
	.C(n24877));
   NAND2xp5_ASAP7_75t_SL U14212 (.Y(n13626),
	.A(n13625),
	.B(n13624));
   O2A1O1Ixp33_ASAP7_75t_SL U14213 (.Y(n25124),
	.A1(FE_OFN16413_n26687),
	.A2(n26258),
	.B(n26255),
	.C(n25123));
   A2O1A1Ixp33_ASAP7_75t_SL U14214 (.Y(n15774),
	.A1(n14183),
	.A2(n14182),
	.B(n14181),
	.C(n14180));
   NAND2xp5_ASAP7_75t_SL U14215 (.Y(n13408),
	.A(n13405),
	.B(n24531));
   INVx2_ASAP7_75t_L U14216 (.Y(n25167),
	.A(FE_OCPN27825_n25169));
   O2A1O1Ixp33_ASAP7_75t_SL U14217 (.Y(n26478),
	.A1(n26542),
	.A2(n26431),
	.B(n25264),
	.C(n25263));
   NOR2xp33_ASAP7_75t_SL U14219 (.Y(n25313),
	.A(n27208),
	.B(FE_OCPN29514_n27136));
   NOR3x1_ASAP7_75t_SL U14220 (.Y(n26814),
	.A(n21080),
	.B(n21079),
	.C(n21078));
   A2O1A1Ixp33_ASAP7_75t_SL U14222 (.Y(n26440),
	.A1(n26139),
	.A2(n24214),
	.B(n24213),
	.C(n24212));
   NAND2x1_ASAP7_75t_SL U14223 (.Y(n26906),
	.A(n26902),
	.B(n26901));
   NAND2xp5_ASAP7_75t_L U14224 (.Y(n25766),
	.A(FE_OFN26148_n26245),
	.B(n25763));
   A2O1A1Ixp33_ASAP7_75t_SL U14225 (.Y(n16075),
	.A1(n16042),
	.A2(n16041),
	.B(n16040),
	.C(n16039));
   A2O1A1Ixp33_ASAP7_75t_L U14226 (.Y(n26055),
	.A1(FE_OFN16177_n27207),
	.A2(n26057),
	.B(n26054),
	.C(n26053));
   NAND2xp5_ASAP7_75t_L U14227 (.Y(n25614),
	.A(FE_OFN29224_FE_OCPN28074_n27049),
	.B(n25611));
   NAND2xp5_ASAP7_75t_L U14228 (.Y(n25177),
	.A(FE_OFN16292_n25175),
	.B(FE_OFN29141_n26574));
   A2O1A1Ixp33_ASAP7_75t_SL U14229 (.Y(n25390),
	.A1(FE_OCPN29587_n26857),
	.A2(FE_OFN29242_n26856),
	.B(n24452),
	.C(n24451));
   A2O1A1Ixp33_ASAP7_75t_SL U14231 (.Y(n25861),
	.A1(n22896),
	.A2(n21008),
	.B(n26976),
	.C(n21007));
   NAND2xp33_ASAP7_75t_SL U14233 (.Y(n26204),
	.A(w2_4_),
	.B(FE_OFN25911_n26491));
   A2O1A1Ixp33_ASAP7_75t_SL U14235 (.Y(n25165),
	.A1(n25163),
	.A2(n25162),
	.B(n26607),
	.C(n25161));
   INVx2_ASAP7_75t_SL U14236 (.Y(n26053),
	.A(n26051));
   XOR2x2_ASAP7_75t_SL U14237 (.Y(n15904),
	.A(u0_rcon_30_),
	.B(n14407));
   NAND2xp5_ASAP7_75t_L U14238 (.Y(n24213),
	.A(n24210),
	.B(n24209));
   A2O1A1Ixp33_ASAP7_75t_SL U14242 (.Y(n16045),
	.A1(n16042),
	.A2(n14661),
	.B(n14660),
	.C(n14659));
   NAND2xp5_ASAP7_75t_L U14243 (.Y(n14599),
	.A(n14598),
	.B(n14597));
   NAND2xp5_ASAP7_75t_L U14244 (.Y(n14600),
	.A(n14591),
	.B(n14597));
   A2O1A1Ixp33_ASAP7_75t_SL U14246 (.Y(n15919),
	.A1(FE_OFN16411_n15884),
	.A2(n14470),
	.B(n14469),
	.C(n14468));
   A2O1A1Ixp33_ASAP7_75t_SL U14248 (.Y(n15466),
	.A1(n15464),
	.A2(n15463),
	.B(n16023),
	.C(n15462));
   A2O1A1Ixp33_ASAP7_75t_SL U14249 (.Y(n27189),
	.A1(n23788),
	.A2(n23787),
	.B(n26517),
	.C(n23786));
   NAND2xp5_ASAP7_75t_SL U14250 (.Y(n15763),
	.A(n15762),
	.B(n15761));
   NAND2xp33_ASAP7_75t_R U14252 (.Y(n16040),
	.A(w0_16_),
	.B(n16037));
   NAND2xp5_ASAP7_75t_L U14256 (.Y(n14969),
	.A(n14966),
	.B(n26221));
   NAND2xp5_ASAP7_75t_R U14257 (.Y(n13797),
	.A(n13794),
	.B(n24495));
   NAND2xp33_ASAP7_75t_SL U14260 (.Y(n14181),
	.A(n14178),
	.B(n25616));
   NAND2xp33_ASAP7_75t_SL U14262 (.Y(n19427),
	.A(n19422),
	.B(n19421));
   A2O1A1Ixp33_ASAP7_75t_SL U14263 (.Y(n25414),
	.A1(n21521),
	.A2(n18911),
	.B(n23467),
	.C(n18910));
   O2A1O1Ixp33_ASAP7_75t_L U14264 (.Y(n22791),
	.A1(n22790),
	.A2(n22789),
	.B(n25682),
	.C(n22788));
   NOR3x1_ASAP7_75t_SL U14267 (.Y(n15462),
	.A(n15461),
	.B(n15460),
	.C(n15459));
   A2O1A1Ixp33_ASAP7_75t_SL U14268 (.Y(n26054),
	.A1(n23895),
	.A2(n23894),
	.B(n26517),
	.C(n23893));
   O2A1O1Ixp33_ASAP7_75t_L U14269 (.Y(n22912),
	.A1(n22911),
	.A2(n22910),
	.B(n27216),
	.C(n22909));
   NAND3x1_ASAP7_75t_SL U14270 (.Y(n21005),
	.A(n21004),
	.B(n21003),
	.C(FE_OCPN8255_n21002));
   NAND2xp33_ASAP7_75t_SL U14271 (.Y(n23223),
	.A(n23219),
	.B(n23221));
   OAI21xp5_ASAP7_75t_SL U14272 (.Y(n25174),
	.A1(n24404),
	.A2(n26464),
	.B(n18730));
   NAND2xp5_ASAP7_75t_L U14273 (.Y(n23222),
	.A(FE_OCPN29492_sa12_4),
	.B(n23221));
   AND2x2_ASAP7_75t_L U14274 (.Y(n23287),
	.A(n23286),
	.B(n23285));
   NAND2x1_ASAP7_75t_SL U14275 (.Y(n26818),
	.A(n21298),
	.B(n21041));
   NOR2xp67_ASAP7_75t_L U14276 (.Y(n24419),
	.A(n19307),
	.B(n19324));
   NAND2xp5_ASAP7_75t_SL U14277 (.Y(n20354),
	.A(n20322),
	.B(n20321));
   A2O1A1Ixp33_ASAP7_75t_SL U14278 (.Y(n25099),
	.A1(n26573),
	.A2(n26572),
	.B(n26571),
	.C(n19028));
   O2A1O1Ixp5_ASAP7_75t_SL U14279 (.Y(n17820),
	.A1(n25277),
	.A2(n17819),
	.B(n27183),
	.C(n17818));
   A2O1A1Ixp33_ASAP7_75t_SL U14280 (.Y(n26193),
	.A1(n23862),
	.A2(n20699),
	.B(n26517),
	.C(n20698));
   NAND2xp5_ASAP7_75t_SL U14281 (.Y(n15251),
	.A(n15250),
	.B(n15249));
   NAND2xp5_ASAP7_75t_L U14282 (.Y(n14469),
	.A(n14466),
	.B(n24320));
   NAND2x1_ASAP7_75t_SL U14283 (.Y(n24229),
	.A(n24432),
	.B(n24433));
   A2O1A1Ixp33_ASAP7_75t_SL U14284 (.Y(n13476),
	.A1(n13474),
	.A2(n13473),
	.B(n15259),
	.C(n13472));
   OR2x2_ASAP7_75t_SRAM U14286 (.Y(n24405),
	.A(n24404),
	.B(n26464));
   OAI21xp5_ASAP7_75t_SL U14287 (.Y(n25039),
	.A1(n23946),
	.A2(n23945),
	.B(n23944));
   O2A1O1Ixp5_ASAP7_75t_SL U14288 (.Y(n27136),
	.A1(n25310),
	.A2(n25309),
	.B(n27183),
	.C(n25308));
   O2A1O1Ixp5_ASAP7_75t_L U14290 (.Y(n21866),
	.A1(n21865),
	.A2(n21864),
	.B(n26082),
	.C(n21863));
   OAI21xp5_ASAP7_75t_L U14291 (.Y(n15736),
	.A1(n13875),
	.A2(FE_OFN72_n15506),
	.B(n15734));
   NAND2xp5_ASAP7_75t_SL U14292 (.Y(n22401),
	.A(n19736),
	.B(n19735));
   O2A1O1Ixp5_ASAP7_75t_SL U14294 (.Y(n20698),
	.A1(n23762),
	.A2(n20697),
	.B(n26323),
	.C(n20696));
   NAND2xp5_ASAP7_75t_SL U14295 (.Y(n13795),
	.A(n13793),
	.B(n13792));
   NAND2x1_ASAP7_75t_SL U14298 (.Y(n25442),
	.A(n20589),
	.B(n20588));
   NAND2xp5_ASAP7_75t_L U14299 (.Y(n19421),
	.A(n19420),
	.B(n19419));
   OAI21xp5_ASAP7_75t_SL U14300 (.Y(n15461),
	.A1(n15444),
	.A2(FE_OFN16348_n15949),
	.B(n15443));
   O2A1O1Ixp5_ASAP7_75t_SL U14301 (.Y(n23409),
	.A1(n23408),
	.A2(n23407),
	.B(n27062),
	.C(n23406));
   NAND2xp5_ASAP7_75t_SL U14302 (.Y(n15249),
	.A(n15248),
	.B(n15247));
   NAND2xp5_ASAP7_75t_SL U14303 (.Y(n13498),
	.A(n13494),
	.B(n13493));
   A2O1A1Ixp33_ASAP7_75t_SL U14305 (.Y(n15532),
	.A1(n15531),
	.A2(n15530),
	.B(n13901),
	.C(n15529));
   A2O1A1Ixp33_ASAP7_75t_SL U14306 (.Y(n17439),
	.A1(n17438),
	.A2(n17437),
	.B(n24331),
	.C(n17436));
   O2A1O1Ixp5_ASAP7_75t_SL U14307 (.Y(n24387),
	.A1(n23621),
	.A2(n23620),
	.B(n25682),
	.C(n23619));
   NOR3xp33_ASAP7_75t_SL U14309 (.Y(n18611),
	.A(n18563),
	.B(n23831),
	.C(n18562));
   NAND2xp5_ASAP7_75t_SL U14311 (.Y(n17683),
	.A(n17682),
	.B(n17681));
   A2O1A1Ixp33_ASAP7_75t_SL U14312 (.Y(n15529),
	.A1(n15528),
	.A2(n15527),
	.B(n15526),
	.C(n15757));
   O2A1O1Ixp5_ASAP7_75t_SL U14313 (.Y(n18730),
	.A1(n24393),
	.A2(n18729),
	.B(n26679),
	.C(n24399));
   NOR3xp33_ASAP7_75t_L U14314 (.Y(n16670),
	.A(n16636),
	.B(n16635),
	.C(n24725));
   A2O1A1Ixp33_ASAP7_75t_SL U14315 (.Y(n15136),
	.A1(n15135),
	.A2(n15134),
	.B(FE_OFN28682_n15888),
	.C(n15133));
   NAND2xp5_ASAP7_75t_L U14316 (.Y(n20588),
	.A(FE_OFN107_n22745),
	.B(FE_OFN16380_n20584));
   OAI21xp5_ASAP7_75t_SL U14317 (.Y(n15737),
	.A1(n15710),
	.A2(n15709),
	.B(n15708));
   NAND2xp5_ASAP7_75t_SL U14319 (.Y(n19235),
	.A(n19221),
	.B(n19220));
   NAND3xp33_ASAP7_75t_SL U14320 (.Y(n25884),
	.A(n25882),
	.B(n25881),
	.C(n25880));
   O2A1O1Ixp5_ASAP7_75t_SL U14321 (.Y(n26050),
	.A1(n27071),
	.A2(n25339),
	.B(n26942),
	.C(n27080));
   NOR3xp33_ASAP7_75t_L U14322 (.Y(n23351),
	.A(n23332),
	.B(n23331),
	.C(n23330));
   O2A1O1Ixp33_ASAP7_75t_L U14323 (.Y(n23350),
	.A1(n23349),
	.A2(n23348),
	.B(n26878),
	.C(n23347));
   NAND2xp5_ASAP7_75t_SL U14324 (.Y(n15443),
	.A(n15442),
	.B(n15441));
   NAND3xp33_ASAP7_75t_SL U14325 (.Y(n23521),
	.A(n23509),
	.B(n23508),
	.C(n19010));
   NAND2xp5_ASAP7_75t_SL U14326 (.Y(n21595),
	.A(n21589),
	.B(n21592));
   NAND2xp5_ASAP7_75t_SL U14329 (.Y(n21594),
	.A(n21593),
	.B(n21592));
   O2A1O1Ixp5_ASAP7_75t_SL U14331 (.Y(n15887),
	.A1(n15886),
	.A2(n15885),
	.B(n15884),
	.C(n15883));
   A2O1A1Ixp33_ASAP7_75t_L U14332 (.Y(n14401),
	.A1(n14391),
	.A2(n14390),
	.B(n13901),
	.C(n14389));
   NOR3xp33_ASAP7_75t_SL U14334 (.Y(n23674),
	.A(n20006),
	.B(n20005),
	.C(n20004));
   NAND2x1p5_ASAP7_75t_SL U14335 (.Y(n23113),
	.A(n18691),
	.B(n18690));
   NAND2xp5_ASAP7_75t_SL U14336 (.Y(n20764),
	.A(n20760),
	.B(n20761));
   NOR2x1_ASAP7_75t_L U14337 (.Y(n25065),
	.A(n21537),
	.B(n20377));
   AOI21xp5_ASAP7_75t_R U14338 (.Y(n19237),
	.A1(n21404),
	.A2(n19209),
	.B(n17506));
   NOR2xp33_ASAP7_75t_SL U14339 (.Y(n24264),
	.A(n24253),
	.B(n24252));
   NOR3xp33_ASAP7_75t_SL U14341 (.Y(n22410),
	.A(n22382),
	.B(n22381),
	.C(FE_OCPN28392_n22380));
   NAND2xp5_ASAP7_75t_SL U14342 (.Y(n21421),
	.A(n21420),
	.B(n21419));
   NAND3xp33_ASAP7_75t_SL U14343 (.Y(n22608),
	.A(n22595),
	.B(n22594),
	.C(n22593));
   NOR3x1_ASAP7_75t_L U14344 (.Y(n19070),
	.A(n17644),
	.B(n18373),
	.C(n19044));
   OA222x2_ASAP7_75t_L U14345 (.Y(n14587),
	.A1(n14586),
	.A2(n14585),
	.B1(n15199),
	.B2(n14585),
	.C1(n14584),
	.C2(n14585));
   O2A1O1Ixp5_ASAP7_75t_L U14347 (.Y(n16669),
	.A1(n16668),
	.A2(n16667),
	.B(n24974),
	.C(n16666));
   NAND2xp33_ASAP7_75t_SL U14348 (.Y(n15442),
	.A(n15436),
	.B(n15439));
   NOR3xp33_ASAP7_75t_SL U14350 (.Y(n17215),
	.A(n17199),
	.B(n23043),
	.C(n17198));
   NAND2xp33_ASAP7_75t_SL U14351 (.Y(n20940),
	.A(n20939),
	.B(n20938));
   NAND2xp5_ASAP7_75t_SL U14352 (.Y(n16716),
	.A(n16715),
	.B(n16714));
   NOR3x1_ASAP7_75t_SL U14353 (.Y(n23371),
	.A(n17459),
	.B(n23272),
	.C(n17462));
   NAND2xp5_ASAP7_75t_L U14354 (.Y(n14586),
	.A(n14570),
	.B(n14569));
   NAND2xp5_ASAP7_75t_SL U14355 (.Y(n13609),
	.A(n13608),
	.B(n13607));
   NAND2xp5_ASAP7_75t_L U14356 (.Y(n14650),
	.A(n14649),
	.B(n14648));
   NAND2xp5_ASAP7_75t_SL U14357 (.Y(n14169),
	.A(n14156),
	.B(n14155));
   NOR3x1_ASAP7_75t_L U14358 (.Y(n25823),
	.A(n18067),
	.B(n24194),
	.C(n18066));
   NAND3xp33_ASAP7_75t_SL U14359 (.Y(n19349),
	.A(n23519),
	.B(n19348),
	.C(n20943));
   NAND3xp33_ASAP7_75t_SL U14360 (.Y(n19490),
	.A(n21529),
	.B(n18898),
	.C(n21290));
   NOR3x1_ASAP7_75t_L U14361 (.Y(n22202),
	.A(n21556),
	.B(n22177),
	.C(n22176));
   OAI21xp5_ASAP7_75t_SL U14362 (.Y(n14239),
	.A1(n15639),
	.A2(n15856),
	.B(n14219));
   NOR3x1_ASAP7_75t_SL U14363 (.Y(n25847),
	.A(n16392),
	.B(n21977),
	.C(n16391));
   NOR3x1_ASAP7_75t_L U14364 (.Y(n23717),
	.A(n20632),
	.B(n23835),
	.C(n21647));
   NAND2xp5_ASAP7_75t_SL U14365 (.Y(n18691),
	.A(n18688),
	.B(n18689));
   NOR3xp33_ASAP7_75t_SL U14366 (.Y(n21573),
	.A(n21570),
	.B(n23082),
	.C(n21569));
   NAND2xp5_ASAP7_75t_SL U14367 (.Y(n23708),
	.A(n23704),
	.B(n23705));
   O2A1O1Ixp33_ASAP7_75t_L U14368 (.Y(n14389),
	.A1(n15519),
	.A2(n14388),
	.B(n13867),
	.C(n14387));
   NOR3x1_ASAP7_75t_L U14370 (.Y(n22348),
	.A(n17871),
	.B(n22704),
	.C(n17870));
   NAND2xp5_ASAP7_75t_SL U14371 (.Y(n18690),
	.A(n26997),
	.B(n18689));
   NAND2xp5_ASAP7_75t_R U14372 (.Y(n14156),
	.A(n14151),
	.B(n14153));
   NAND2xp5_ASAP7_75t_SL U14373 (.Y(n15647),
	.A(n15645),
	.B(n15644));
   OR3x1_ASAP7_75t_SL U14374 (.Y(n19341),
	.A(n19340),
	.B(n19339),
	.C(n22045));
   NOR3xp33_ASAP7_75t_SL U14375 (.Y(n23240),
	.A(n22259),
	.B(n23214),
	.C(n22258));
   NAND2xp33_ASAP7_75t_SL U14376 (.Y(n14155),
	.A(n14154),
	.B(n14153));
   OAI21xp5_ASAP7_75t_L U14377 (.Y(n14166),
	.A1(n14959),
	.A2(FE_OFN28544_n13805),
	.B(n14164));
   NAND2xp5_ASAP7_75t_SL U14378 (.Y(n14130),
	.A(n14125),
	.B(n14127));
   NAND2xp5_ASAP7_75t_L U14379 (.Y(n15231),
	.A(n15225),
	.B(n15228));
   NAND2xp5_ASAP7_75t_SL U14380 (.Y(n21457),
	.A(n17287),
	.B(n17286));
   NAND2xp5_ASAP7_75t_SL U14381 (.Y(n23082),
	.A(n21568),
	.B(n21567));
   NAND2xp5_ASAP7_75t_R U14383 (.Y(n14129),
	.A(n14128),
	.B(n14127));
   NAND3xp33_ASAP7_75t_SL U14384 (.Y(n18666),
	.A(n17378),
	.B(n17377),
	.C(n20389));
   NOR3xp33_ASAP7_75t_SL U14386 (.Y(n22389),
	.A(n17704),
	.B(n19710),
	.C(n19739));
   NOR2x1_ASAP7_75t_SL U14387 (.Y(n25223),
	.A(n17016),
	.B(n17015));
   NAND2xp5_ASAP7_75t_L U14388 (.Y(n13446),
	.A(n13436),
	.B(n13435));
   NAND2xp5_ASAP7_75t_SL U14389 (.Y(n14219),
	.A(n14218),
	.B(n14217));
   OA222x2_ASAP7_75t_SL U14390 (.Y(n16025),
	.A1(n16024),
	.A2(n16023),
	.B1(n16022),
	.B2(n16023),
	.C1(n16021),
	.C2(n16023));
   NOR2x1_ASAP7_75t_SL U14391 (.Y(n26360),
	.A(n16728),
	.B(n16727));
   NAND2xp33_ASAP7_75t_L U14392 (.Y(n24261),
	.A(n24260),
	.B(n24259));
   NOR2x1_ASAP7_75t_SL U14393 (.Y(n26549),
	.A(n22996),
	.B(n19025));
   NOR3xp33_ASAP7_75t_SL U14395 (.Y(n19348),
	.A(n19347),
	.B(n22998),
	.C(n26661));
   NAND2xp5_ASAP7_75t_SL U14396 (.Y(n20643),
	.A(n20666),
	.B(n18558));
   NOR3xp33_ASAP7_75t_L U14397 (.Y(n17480),
	.A(n26076),
	.B(n21360),
	.C(n17477));
   NOR3xp33_ASAP7_75t_L U14398 (.Y(n18781),
	.A(n18772),
	.B(n19845),
	.C(n18771));
   NAND2xp5_ASAP7_75t_L U14399 (.Y(n20296),
	.A(n20000),
	.B(n19999));
   NAND2xp5_ASAP7_75t_L U14400 (.Y(n17812),
	.A(n20143),
	.B(n17809));
   NOR3xp33_ASAP7_75t_SL U14401 (.Y(n18049),
	.A(n21753),
	.B(n21058),
	.C(n18864));
   AND2x2_ASAP7_75t_R U14402 (.Y(n20884),
	.A(n20883),
	.B(n20882));
   NOR3xp33_ASAP7_75t_SL U14403 (.Y(n18898),
	.A(n18893),
	.B(n23431),
	.C(n24243));
   NOR2xp33_ASAP7_75t_SL U14404 (.Y(n24587),
	.A(n22230),
	.B(n22229));
   NAND2x1p5_ASAP7_75t_L U14405 (.Y(n26661),
	.A(n19346),
	.B(n19345));
   NAND2xp5_ASAP7_75t_SL U14406 (.Y(n19893),
	.A(n16817),
	.B(n20333));
   NAND3xp33_ASAP7_75t_SL U14407 (.Y(n17354),
	.A(n21534),
	.B(n20367),
	.C(n17351));
   NOR3xp33_ASAP7_75t_SL U14408 (.Y(n17377),
	.A(n17376),
	.B(n21548),
	.C(n22453));
   NAND2xp33_ASAP7_75t_SL U14409 (.Y(n17944),
	.A(n17940),
	.B(n17941));
   NAND2xp5_ASAP7_75t_SL U14410 (.Y(n20035),
	.A(n20032),
	.B(n20031));
   NOR3xp33_ASAP7_75t_SL U14411 (.Y(n18558),
	.A(n18557),
	.B(n23835),
	.C(n21673));
   OR2x2_ASAP7_75t_SRAM U14412 (.Y(n22081),
	.A(FE_OCPN29436_n22080),
	.B(FE_OCPN27685_n26968));
   NOR2x1_ASAP7_75t_SL U14413 (.Y(n21567),
	.A(n26461),
	.B(n21566));
   NAND3xp33_ASAP7_75t_SL U14414 (.Y(n21354),
	.A(FE_OCPN29416_n22516),
	.B(n21353),
	.C(n21410));
   NAND2xp33_ASAP7_75t_L U14415 (.Y(n15890),
	.A(n15821),
	.B(n15820));
   NAND2xp5_ASAP7_75t_SL U14416 (.Y(n14164),
	.A(n14163),
	.B(n14162));
   AND3x1_ASAP7_75t_SL U14418 (.Y(n14127),
	.A(n14693),
	.B(n14124),
	.C(n14123));
   NOR2xp33_ASAP7_75t_R U14419 (.Y(n14527),
	.A(FE_OFN16145_n15214),
	.B(n14525));
   NAND3x1_ASAP7_75t_SL U14420 (.Y(n18771),
	.A(n17299),
	.B(n21157),
	.C(n19833));
   AND2x2_ASAP7_75t_SL U14421 (.Y(n23502),
	.A(n23517),
	.B(n23501));
   AND2x2_ASAP7_75t_SRAM U14422 (.Y(n20667),
	.A(n23710),
	.B(n23766));
   NAND2x1_ASAP7_75t_SL U14423 (.Y(n23710),
	.A(n18587),
	.B(n18586));
   NOR2x1p5_ASAP7_75t_L U14424 (.Y(n26151),
	.A(n22033),
	.B(n19333));
   NOR3xp33_ASAP7_75t_SL U14425 (.Y(n24647),
	.A(n17554),
	.B(n20104),
	.C(FE_OCPN27937_n18841));
   NAND2x1_ASAP7_75t_L U14426 (.Y(n20810),
	.A(n20550),
	.B(n20549));
   NAND2xp5_ASAP7_75t_L U14427 (.Y(n17961),
	.A(n17960),
	.B(n17959));
   NAND2xp5_ASAP7_75t_SL U14428 (.Y(n24079),
	.A(n17509),
	.B(FE_OCPN28417_n21396));
   OAI22xp5_ASAP7_75t_L U14429 (.Y(n14700),
	.A1(n15380),
	.A2(n14699),
	.B1(FE_PSN8271_n15924),
	.B2(n14699));
   NOR3xp33_ASAP7_75t_SL U14430 (.Y(n21353),
	.A(n24562),
	.B(n21848),
	.C(n21350));
   NAND2xp5_ASAP7_75t_L U14431 (.Y(n21381),
	.A(n21376),
	.B(n21378));
   NOR2x1_ASAP7_75t_SL U14433 (.Y(n16817),
	.A(n23643),
	.B(n20344));
   NOR2x1_ASAP7_75t_L U14435 (.Y(n22244),
	.A(n23581),
	.B(n22259));
   NAND2xp5_ASAP7_75t_L U14436 (.Y(n20572),
	.A(n17914),
	.B(n17913));
   NAND2xp5_ASAP7_75t_L U14437 (.Y(n14296),
	.A(n14291),
	.B(n14293));
   NAND2xp5_ASAP7_75t_SL U14438 (.Y(n19654),
	.A(n19652),
	.B(n19651));
   NOR3xp33_ASAP7_75t_R U14439 (.Y(n21299),
	.A(n21518),
	.B(n21707),
	.C(n21297));
   NOR2x1_ASAP7_75t_SL U14441 (.Y(n18747),
	.A(n18757),
	.B(n19844));
   NAND2xp33_ASAP7_75t_SL U14442 (.Y(n14123),
	.A(n14122),
	.B(n14121));
   NAND2xp33_ASAP7_75t_SL U14445 (.Y(n20628),
	.A(n20625),
	.B(n23882));
   OAI21xp5_ASAP7_75t_SL U14446 (.Y(n15519),
	.A1(n13875),
	.A2(n14368),
	.B(n14367));
   OA21x2_ASAP7_75t_L U14447 (.Y(n18874),
	.A1(n23431),
	.A2(n21525),
	.B(FE_OCPN27405_sa03_4));
   NAND2xp33_ASAP7_75t_L U14448 (.Y(n14525),
	.A(n14518),
	.B(n14517));
   NAND2xp5_ASAP7_75t_SL U14449 (.Y(n20138),
	.A(n17789),
	.B(n19257));
   NAND2xp33_ASAP7_75t_SL U14450 (.Y(n20627),
	.A(n20626),
	.B(n23882));
   NAND2x1_ASAP7_75t_SL U14451 (.Y(n23480),
	.A(n19018),
	.B(n19017));
   NAND2xp5_ASAP7_75t_SL U14452 (.Y(n21232),
	.A(n21644),
	.B(n21638));
   NOR3xp33_ASAP7_75t_SL U14453 (.Y(n24041),
	.A(n20252),
	.B(n20251),
	.C(FE_OFN27046_n22024));
   NOR2xp33_ASAP7_75t_SL U14454 (.Y(n18370),
	.A(n18369),
	.B(n20438));
   OR3x1_ASAP7_75t_L U14455 (.Y(n13892),
	.A(n15698),
	.B(FE_OFN28909_w3_23),
	.C(FE_OCPN4685_n15658));
   NAND2xp33_ASAP7_75t_SL U14456 (.Y(n16387),
	.A(n16291),
	.B(n20034));
   OR2x2_ASAP7_75t_L U14457 (.Y(n13482),
	.A(n13481),
	.B(FE_OFN28453_n13348));
   AND2x2_ASAP7_75t_R U14458 (.Y(n24185),
	.A(n25815),
	.B(n24182));
   NAND3x1_ASAP7_75t_SL U14460 (.Y(n18745),
	.A(n18744),
	.B(n19602),
	.C(n18743));
   NAND2xp5_ASAP7_75t_R U14461 (.Y(n19306),
	.A(n19344),
	.B(n22986));
   NAND2x1_ASAP7_75t_SL U14463 (.Y(n23498),
	.A(n20258),
	.B(n20257));
   NOR2xp33_ASAP7_75t_L U14464 (.Y(n19261),
	.A(n22872),
	.B(n22871));
   OAI21x1_ASAP7_75t_SL U14465 (.Y(n22899),
	.A1(FE_OCPN29533_n26971),
	.A2(FE_OFN27058_n22094),
	.B(n22070));
   NOR2x2_ASAP7_75t_L U14466 (.Y(n22060),
	.A(FE_OFN28703_FE_OCPN27740_sa02_4),
	.B(n22903));
   OA21x2_ASAP7_75t_SRAM U14467 (.Y(n14019),
	.A1(FE_OFN27214_w3_17),
	.A2(FE_OFN27074_n13868),
	.B(n14018));
   NOR2xp33_ASAP7_75t_L U14468 (.Y(n16598),
	.A(FE_OCPN5015_n23031),
	.B(n21906));
   NAND2xp5_ASAP7_75t_L U14469 (.Y(n17203),
	.A(n19775),
	.B(n19777));
   AND3x1_ASAP7_75t_R U14471 (.Y(n21857),
	.A(n23288),
	.B(n21856),
	.C(n21855));
   OA21x2_ASAP7_75t_SRAM U14472 (.Y(n17122),
	.A1(n17121),
	.A2(FE_OCPN28204_n20526),
	.B(n17145));
   NAND2xp5_ASAP7_75t_SL U14473 (.Y(n17105),
	.A(n17046),
	.B(n25995));
   NAND2x1_ASAP7_75t_L U14474 (.Y(n20364),
	.A(n20359),
	.B(n20361));
   NAND2x1_ASAP7_75t_L U14475 (.Y(n20363),
	.A(n20362),
	.B(n20361));
   NAND2xp5_ASAP7_75t_L U14478 (.Y(n19017),
	.A(n22934),
	.B(n19016));
   NOR2x1_ASAP7_75t_SL U14479 (.Y(n19204),
	.A(FE_OCPN28082_n21860),
	.B(n17456));
   NOR2x1p5_ASAP7_75t_SL U14480 (.Y(n25063),
	.A(n23099),
	.B(n21546));
   OA21x2_ASAP7_75t_L U14481 (.Y(n21029),
	.A1(FE_OCPN28184_n18020),
	.A2(FE_PSN8319_n21725),
	.B(FE_OFN28608_n21027));
   NOR2x1_ASAP7_75t_SL U14482 (.Y(n21014),
	.A(FE_OCPN27611_n23426),
	.B(n21728));
   OAI222xp33_ASAP7_75t_L U14484 (.Y(n14636),
	.A1(n13844),
	.A2(n14635),
	.B1(FE_PSN8324_n15987),
	.B2(n14635),
	.C1(FE_OFN26641_w3_14),
	.C2(n14635));
   OR3x1_ASAP7_75t_R U14488 (.Y(n14069),
	.A(n14303),
	.B(FE_OFN28_w3_23),
	.C(n15658));
   NOR2xp33_ASAP7_75t_L U14489 (.Y(n14612),
	.A(n14632),
	.B(n13851));
   OAI222xp33_ASAP7_75t_SRAM U14490 (.Y(n14624),
	.A1(FE_OFN26634_w3_14),
	.A2(n14686),
	.B1(FE_OFN26131_n15376),
	.B2(n14686),
	.C1(FE_OCPN28407_FE_OFN16433_w3_11),
	.C2(n14686));
   AND3x2_ASAP7_75t_SL U14491 (.Y(n17989),
	.A(FE_OCPN28001_n21310),
	.B(n21317),
	.C(FE_OCPN27405_sa03_4));
   OAI21xp5_ASAP7_75t_L U14492 (.Y(n15217),
	.A1(FE_OFN27210_w3_30),
	.A2(n14479),
	.B(FE_OFN28604_n14534));
   OA21x2_ASAP7_75t_SRAM U14494 (.Y(n17534),
	.A1(n19938),
	.A2(n19932),
	.B(n19725));
   OR3x1_ASAP7_75t_SRAM U14495 (.Y(n15313),
	.A(n15312),
	.B(FE_OFN28909_w3_23),
	.C(FE_OFN29192_n13870));
   OAI22xp33_ASAP7_75t_SRAM U14496 (.Y(n15846),
	.A1(n15787),
	.A2(n15844),
	.B1(n15843),
	.B2(n15844));
   NOR3xp33_ASAP7_75t_L U14497 (.Y(n21572),
	.A(n26460),
	.B(n20391),
	.C(n22584));
   OR2x2_ASAP7_75t_SRAM U14499 (.Y(n18845),
	.A(n17527),
	.B(n18846));
   OAI21xp33_ASAP7_75t_SL U14500 (.Y(n14452),
	.A1(n14448),
	.A2(FE_OFN28792_n15787),
	.B(n15002));
   NAND2xp5_ASAP7_75t_L U14501 (.Y(n14450),
	.A(n14449),
	.B(n15851));
   OA21x2_ASAP7_75t_L U14503 (.Y(n17252),
	.A1(FE_OCPN27679_n18631),
	.A2(n18776),
	.B(n17271));
   INVxp67_ASAP7_75t_L U14504 (.Y(n16342),
	.A(n16341));
   NOR2x1p5_ASAP7_75t_L U14505 (.Y(n22838),
	.A(FE_OFN26548_n18206),
	.B(n21770));
   OAI22xp5_ASAP7_75t_SL U14508 (.Y(n23773),
	.A1(FE_OCPN27715_n23875),
	.A2(FE_OCPN29567_n23806),
	.B1(n20617),
	.B2(FE_OCPN29567_n23806));
   OA21x2_ASAP7_75t_R U14509 (.Y(n15720),
	.A1(FE_OFN26535_w3_19),
	.A2(FE_OFN28551_FE_OFN26114_n),
	.B(n15719));
   OA21x2_ASAP7_75t_SRAM U14511 (.Y(n13767),
	.A1(n15028),
	.A2(n15809),
	.B(FE_OFN29052_w3_5));
   OA21x2_ASAP7_75t_SL U14512 (.Y(n17387),
	.A1(n21553),
	.A2(n27006),
	.B(FE_OCPN27887_n17331));
   NOR2xp33_ASAP7_75t_L U14513 (.Y(n14630),
	.A(n14912),
	.B(n14957));
   OA21x2_ASAP7_75t_L U14516 (.Y(n14061),
	.A1(FE_OFN26535_w3_19),
	.A2(FE_OFN27151_n),
	.B(n14276));
   NOR2x1_ASAP7_75t_SL U14517 (.Y(n15124),
	.A(n15028),
	.B(n13725));
   NOR2x1_ASAP7_75t_L U14518 (.Y(n14157),
	.A(n14941),
	.B(n14897));
   OA21x2_ASAP7_75t_SRAM U14519 (.Y(n13957),
	.A1(FE_OFN28884_n),
	.A2(FE_OFN28856_n15450),
	.B(FE_OFN25920_n15995));
   OR3x1_ASAP7_75t_SRAM U14521 (.Y(n15334),
	.A(n15658),
	.B(FE_OFN28_w3_23),
	.C(FE_OFN28769_n15478));
   NAND2x1p5_ASAP7_75t_SL U14522 (.Y(n23871),
	.A(FE_OFN29140_n18527),
	.B(n20617));
   OA21x2_ASAP7_75t_SL U14524 (.Y(n18580),
	.A1(FE_OFN29081_n18526),
	.A2(n18548),
	.B(FE_OCPN28163_FE_OFN99_sa20_5));
   NAND2x1_ASAP7_75t_SL U14525 (.Y(n21239),
	.A(FE_OFN29140_n18527),
	.B(FE_OFN28986_n18597));
   OR3x1_ASAP7_75t_SRAM U14526 (.Y(n13889),
	.A(FE_OFN29192_n13870),
	.B(FE_OFN28909_w3_23),
	.C(n13916));
   NOR3x2_ASAP7_75t_SL U14527 (.Y(n22533),
	.A(n20195),
	.B(FE_OFN29210_FE_OCPN27261_sa02_0),
	.C(FE_OFN29049_n17756));
   NOR2x1_ASAP7_75t_L U14528 (.Y(n16551),
	.A(n16552),
	.B(n16610));
   NAND2xp5_ASAP7_75t_L U14529 (.Y(n14944),
	.A(n15993),
	.B(FE_OFN28574_n16016));
   NOR2x1p5_ASAP7_75t_SL U14532 (.Y(n17527),
	.A(FE_OCPN29420_FE_OFN16128_sa32_2),
	.B(n18832));
   NAND2x1_ASAP7_75t_SL U14533 (.Y(n15719),
	.A(FE_OCPN29578_FE_OFN27214_w3_17),
	.B(FE_OCPN27928_FE_OFN4_w3_22));
   NAND2x2_ASAP7_75t_SL U14534 (.Y(n20195),
	.A(n17763),
	.B(n20993));
   NOR2x1p5_ASAP7_75t_SL U14535 (.Y(n16427),
	.A(FE_OFN25938_sa33_3),
	.B(n23556));
   NAND2xp5_ASAP7_75t_SL U14537 (.Y(n22526),
	.A(n17760),
	.B(n17742));
   NAND2x1_ASAP7_75t_L U14539 (.Y(n19677),
	.A(n16547),
	.B(FE_OFN28916_sa10_4));
   NAND2xp5_ASAP7_75t_L U14540 (.Y(n21845),
	.A(FE_OCPN29504_sa11_4),
	.B(n17452));
   NAND2x1p5_ASAP7_75t_SL U14541 (.Y(n13725),
	.A(FE_OFN25897_w3_4),
	.B(n15857));
   NAND2x1p5_ASAP7_75t_SL U14542 (.Y(n16989),
	.A(FE_OFN28478_sa13_2),
	.B(n16988));
   INVx2_ASAP7_75t_R U14543 (.Y(n26679),
	.A(n27015));
   OAI22xp33_ASAP7_75t_R U14544 (.Y(n16003),
	.A1(FE_OFN29125_n),
	.A2(n15998),
	.B1(FE_OCPN29508_FE_OFN16184_w3_9),
	.B2(n15998));
   NOR2x1p5_ASAP7_75t_L U14546 (.Y(n20490),
	.A(FE_OFN28775_n16992),
	.B(FE_OCPN27836_n16976));
   NAND2x1_ASAP7_75t_SL U14548 (.Y(n23306),
	.A(n21084),
	.B(n18164));
   OAI21xp33_ASAP7_75t_SRAM U14550 (.Y(n24756),
	.A1(text_in_r_12_),
	.A2(FE_OCPN29520_n24755),
	.B(n24754));
   OAI21xp33_ASAP7_75t_SRAM U14551 (.Y(n25962),
	.A1(text_in_r_21_),
	.A2(n25961),
	.B(n25960));
   NOR2x1p5_ASAP7_75t_SL U14552 (.Y(n14941),
	.A(FE_OFN26641_w3_14),
	.B(n15447));
   OR2x2_ASAP7_75t_L U14553 (.Y(n16776),
	.A(FE_OCPN29580_n),
	.B(FE_OCPN27553_n19975));
   NOR2xp33_ASAP7_75t_SL U14554 (.Y(n15896),
	.A(w3_2_),
	.B(n25596));
   NAND2x1_ASAP7_75t_SL U14555 (.Y(n18019),
	.A(FE_OCPN29349_FE_OCPN27405_sa03_4),
	.B(n21310));
   NAND2x1p5_ASAP7_75t_SL U14556 (.Y(n15987),
	.A(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(FE_OCPN28408_FE_OFN16433_w3_11));
   NOR2x1p5_ASAP7_75t_L U14557 (.Y(n18045),
	.A(FE_OFN141_sa03_1),
	.B(FE_OFN29199_FE_OCPN27726_n));
   NOR2x2_ASAP7_75t_SL U14558 (.Y(n18159),
	.A(FE_OFN28688_sa22_2),
	.B(n22310));
   NOR2x1p5_ASAP7_75t_SL U14559 (.Y(n17995),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2),
	.B(FE_OFN28523_sa03_1));
   NAND2x1_ASAP7_75t_SL U14560 (.Y(n16394),
	.A(FE_OFN28669_sa31_5),
	.B(FE_OFN26595_sa31_4));
   NAND3xp33_ASAP7_75t_L U14561 (.Y(n13348),
	.A(FE_OFN27130_w3_28),
	.B(FE_OCPN29428_FE_OFN27131_w3_29),
	.C(FE_OCPN28096_w3_31));
   NOR2x1p5_ASAP7_75t_L U14562 (.Y(n20256),
	.A(FE_OFN27078_sa23_5),
	.B(FE_OCPN27577_sa23_4));
   NOR2x1_ASAP7_75t_SL U14563 (.Y(n17254),
	.A(FE_OFN29249_n),
	.B(n17298));
   NOR2x1_ASAP7_75t_L U14564 (.Y(n17553),
	.A(FE_OFN28696_sa32_4),
	.B(FE_OFN28707_n));
   INVx2_ASAP7_75t_L U14565 (.Y(n16790),
	.A(FE_OCPN27246_n22663));
   NOR2x1p5_ASAP7_75t_SL U14566 (.Y(n16418),
	.A(FE_OCPN29391_FE_OFN29162_sa33_2),
	.B(n16875));
   INVx2_ASAP7_75t_SL U14568 (.Y(n15259),
	.A(n13634));
   NAND2x1p5_ASAP7_75t_SL U14569 (.Y(n16992),
	.A(FE_OCPN29351_FE_OFN26116_sa13_1),
	.B(n20514));
   NAND2x1p5_ASAP7_75t_SL U14570 (.Y(n17679),
	.A(FE_OCPN27499_FE_OFN16151_sa32_5),
	.B(FE_OFN29235_n));
   NOR2x1p5_ASAP7_75t_SL U14571 (.Y(n15667),
	.A(w3_21_),
	.B(FE_OFN37_w3_23));
   NAND2xp5_ASAP7_75t_SL U14572 (.Y(n25091),
	.A(FE_OCPN29373_FE_OFN29191_sa23_2),
	.B(n18970));
   NOR2x1_ASAP7_75t_L U14576 (.Y(n15455),
	.A(FE_OCPN29534_FE_OFN8_w3_14),
	.B(FE_OCPN29508_FE_OFN16184_w3_9));
   NOR2x1p5_ASAP7_75t_SL U14577 (.Y(n16417),
	.A(FE_OFN28694_sa33_4),
	.B(FE_OFN28679_sa33_5));
   NOR3x2_ASAP7_75t_SL U14578 (.Y(n23336),
	.A(FE_OFN55_sa22_5),
	.B(FE_OFN16135_sa22_4),
	.C(FE_OFN26136_sa22_3));
   NAND2xp5_ASAP7_75t_L U14579 (.Y(n17756),
	.A(FE_OFN16234_sa02_2),
	.B(sa02_1_));
   INVxp33_ASAP7_75t_SRAM U14580 (.Y(n13225),
	.A(text_in_r_49_));
   NAND2x1_ASAP7_75t_SL U14590 (.Y(n17345),
	.A(FE_OFN28672_sa01_2),
	.B(sa01_1_));
   INVxp33_ASAP7_75t_SRAM U14592 (.Y(n13051),
	.A(text_in_r_39_));
   INVxp33_ASAP7_75t_SRAM U14593 (.Y(n13215),
	.A(text_in_r_83_));
   NAND2xp5_ASAP7_75t_SL U14594 (.Y(n13726),
	.A(w3_4_),
	.B(w3_5_));
   A2O1A1Ixp33_ASAP7_75t_SL U14598 (.Y(n355),
	.A1(n26438),
	.A2(n26437),
	.B(n26436),
	.C(n26435));
   A2O1A1Ixp33_ASAP7_75t_SL U14599 (.Y(n474),
	.A1(n25965),
	.A2(n25964),
	.B(n25963),
	.C(n25962));
   NAND3xp33_ASAP7_75t_SL U14601 (.Y(n26435),
	.A(n26436),
	.B(n26438),
	.C(n26437));
   OAI21xp33_ASAP7_75t_SRAM U14602 (.Y(n567),
	.A1(key_68_),
	.A2(FE_OFN25_n16125),
	.B(n14665));
   A2O1A1Ixp33_ASAP7_75t_SL U14603 (.Y(n445),
	.A1(n24690),
	.A2(n24689),
	.B(FE_OFN27209_w3_30),
	.C(n24687));
   NAND3xp33_ASAP7_75t_SL U14604 (.Y(n26846),
	.A(FE_OFN25961_w3_8),
	.B(n26849),
	.C(n26848));
   NAND3xp33_ASAP7_75t_SL U14605 (.Y(n26918),
	.A(n26919),
	.B(n26921),
	.C(n26920));
   NOR2xp67_ASAP7_75t_SL U14606 (.Y(n25663),
	.A(n25662),
	.B(n25664));
   OAI21xp33_ASAP7_75t_R U14608 (.Y(n543),
	.A1(key_70_),
	.A2(FE_OFN25_n16125),
	.B(n16054));
   A2O1A1Ixp33_ASAP7_75t_SL U14609 (.Y(n427),
	.A1(n27175),
	.A2(n27174),
	.B(n27173),
	.C(n27172));
   NAND2xp5_ASAP7_75t_SL U14611 (.Y(n623),
	.A(n16255),
	.B(n16254));
   A2O1A1Ixp33_ASAP7_75t_SL U14612 (.Y(n507),
	.A1(n25249),
	.A2(n25248),
	.B(n25247),
	.C(n25246));
   A2O1A1Ixp33_ASAP7_75t_SL U14613 (.Y(n487),
	.A1(n27199),
	.A2(n27198),
	.B(n27197),
	.C(n27196));
   A2O1A1Ixp33_ASAP7_75t_SL U14614 (.Y(n466),
	.A1(n27162),
	.A2(n27161),
	.B(n27160),
	.C(n27159));
   A2O1A1Ixp33_ASAP7_75t_SL U14615 (.Y(n16155),
	.A1(FE_OFN26_n16125),
	.A2(FE_OCPN29500_FE_OFN28662_w3_7),
	.B(n16154),
	.C(n16156));
   O2A1O1Ixp5_ASAP7_75t_SL U14616 (.Y(n26548),
	.A1(FE_OCPN5056_n26535),
	.A2(n26534),
	.B(n26533),
	.C(n26532));
   NAND3xp33_ASAP7_75t_SL U14617 (.Y(n25781),
	.A(FE_OFN26163_w3_13),
	.B(n25784),
	.C(n25783));
   INVx1_ASAP7_75t_SL U14618 (.Y(n26388),
	.A(FE_OCPN27310_n26389));
   NAND3xp33_ASAP7_75t_SL U14619 (.Y(n26610),
	.A(n26611),
	.B(n26613),
	.C(n26612));
   OAI21xp33_ASAP7_75t_SRAM U14620 (.Y(n600),
	.A1(key_88_),
	.A2(FE_OFN19_n16125),
	.B(n16165));
   NAND3xp33_ASAP7_75t_SL U14621 (.Y(n27172),
	.A(n27173),
	.B(n27175),
	.C(n27174));
   O2A1O1Ixp5_ASAP7_75t_SL U14622 (.Y(n25652),
	.A1(FE_OCPN29515_n27136),
	.A2(n25626),
	.B(n25625),
	.C(n25624));
   NOR2xp33_ASAP7_75t_SL U14623 (.Y(n25153),
	.A(n25152),
	.B(n25154));
   NAND3xp33_ASAP7_75t_SL U14624 (.Y(n26759),
	.A(n26760),
	.B(n26762),
	.C(n26761));
   NAND3xp33_ASAP7_75t_SL U14625 (.Y(n24494),
	.A(n24495),
	.B(n24497),
	.C(n24496));
   OAI21xp33_ASAP7_75t_SRAM U14626 (.Y(n542),
	.A1(key_102_),
	.A2(FE_OFN28472_ld),
	.B(n15272));
   NAND3xp33_ASAP7_75t_SL U14629 (.Y(n25246),
	.A(n25247),
	.B(n25249),
	.C(n25248));
   OAI21xp33_ASAP7_75t_SL U14630 (.Y(n635),
	.A1(n16247),
	.A2(FE_OFN16421_n23974),
	.B(n16246));
   NAND3xp33_ASAP7_75t_SL U14631 (.Y(n26354),
	.A(n26355),
	.B(n26357),
	.C(n26356));
   OAI21xp5_ASAP7_75t_SL U14632 (.Y(n638),
	.A1(FE_OFN16287_n16230),
	.A2(FE_OFN28890_n),
	.B(n16229));
   NAND3xp33_ASAP7_75t_SL U14634 (.Y(n26286),
	.A(n26287),
	.B(n26289),
	.C(n26288));
   OAI21xp5_ASAP7_75t_SL U14635 (.Y(n26421),
	.A1(FE_OFN1_ld_r),
	.A2(FE_OCPN5088_n27079),
	.B(n26422));
   OAI21xp5_ASAP7_75t_SL U14636 (.Y(n26740),
	.A1(FE_OFN2_ld_r),
	.A2(n26742),
	.B(n26741));
   AOI21x1_ASAP7_75t_SL U14637 (.Y(n27223),
	.A1(FE_OCPN29287_n27210),
	.A2(n25311),
	.B(n27209));
   NOR3xp33_ASAP7_75t_SL U14638 (.Y(n25705),
	.A(n25707),
	.B(w1_0_),
	.C(n25706));
   OAI21xp33_ASAP7_75t_SRAM U14640 (.Y(n612),
	.A1(key_89_),
	.A2(FE_OFN22_n16125),
	.B(n16140));
   NOR3xp33_ASAP7_75t_SL U14641 (.Y(n25928),
	.A(n25930),
	.B(w2_0_),
	.C(n25929));
   NAND3xp33_ASAP7_75t_L U14642 (.Y(n26931),
	.A(n26932),
	.B(n26934),
	.C(n26933));
   A2O1A1Ixp33_ASAP7_75t_SL U14643 (.Y(n27175),
	.A1(n27171),
	.A2(FE_OFN16215_ld_r),
	.B(n27170),
	.C(n27169));
   NAND3xp33_ASAP7_75t_SL U14644 (.Y(n26655),
	.A(n26656),
	.B(n26658),
	.C(n26657));
   OAI21xp33_ASAP7_75t_SRAM U14645 (.Y(n566),
	.A1(key_100_),
	.A2(FE_OFN28472_ld),
	.B(n13635));
   OAI21xp5_ASAP7_75t_SL U14647 (.Y(n26916),
	.A1(FE_OFN1_ld_r),
	.A2(FE_OCPN27442_n27202),
	.B(n26917));
   OAI21xp33_ASAP7_75t_SRAM U14648 (.Y(n531),
	.A1(key_71_),
	.A2(FE_OFN28463_ld),
	.B(n15772));
   OAI21xp33_ASAP7_75t_SRAM U14649 (.Y(n552),
	.A1(key_93_),
	.A2(FE_OFN22_n16125),
	.B(n16121));
   O2A1O1Ixp5_ASAP7_75t_SL U14650 (.Y(n26189),
	.A1(n26178),
	.A2(n26177),
	.B(n26176),
	.C(n26175));
   OAI21xp5_ASAP7_75t_SL U14651 (.Y(n26807),
	.A1(FE_OFN2_ld_r),
	.A2(n26809),
	.B(n26808));
   O2A1O1Ixp5_ASAP7_75t_SL U14652 (.Y(n26264),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(FE_OCPN27519_n25407),
	.B(n26263),
	.C(n26262));
   O2A1O1Ixp33_ASAP7_75t_SL U14653 (.Y(n26219),
	.A1(FE_OFN16214_ld_r),
	.A2(n26218),
	.B(n26217),
	.C(n26216));
   O2A1O1Ixp5_ASAP7_75t_SL U14654 (.Y(n25426),
	.A1(FE_OFN16214_ld_r),
	.A2(n26732),
	.B(n25425),
	.C(n25424));
   A2O1A1Ixp33_ASAP7_75t_SL U14655 (.Y(n519),
	.A1(FE_OCPN27430_n26334),
	.A2(n24758),
	.B(n24757),
	.C(n24756));
   OAI21xp5_ASAP7_75t_L U14656 (.Y(n26020),
	.A1(n26021),
	.A2(FE_OCPN7605_n26234),
	.B(FE_OFN16215_ld_r));
   OAI21xp33_ASAP7_75t_SL U14658 (.Y(n629),
	.A1(n16050),
	.A2(n25140),
	.B(n15912));
   OAI21xp5_ASAP7_75t_SL U14660 (.Y(n631),
	.A1(FE_OCPN29371_n16191),
	.A2(FE_OFN29087_n),
	.B(n16177));
   NOR3xp33_ASAP7_75t_SL U14661 (.Y(n26175),
	.A(n26178),
	.B(n26176),
	.C(n26177));
   NAND2xp5_ASAP7_75t_L U14662 (.Y(n25949),
	.A(FE_OFN16322_n25946),
	.B(FE_OCPN27535_n));
   OAI21xp5_ASAP7_75t_SL U14663 (.Y(n24492),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OCPN27379_n26809),
	.B(n24493));
   OAI21xp33_ASAP7_75t_SRAM U14664 (.Y(n576),
	.A1(key_91_),
	.A2(FE_OFN22_n16125),
	.B(n16137));
   OAI21xp33_ASAP7_75t_R U14665 (.Y(n585),
	.A1(key_82_),
	.A2(FE_OFN27_n16125),
	.B(n16101));
   OAI21xp33_ASAP7_75t_SRAM U14666 (.Y(n530),
	.A1(key_103_),
	.A2(FE_OFN28472_ld),
	.B(n14606));
   OAI21xp33_ASAP7_75t_R U14667 (.Y(n579),
	.A1(key_66_),
	.A2(FE_OFN25_n16125),
	.B(n14009));
   A2O1A1Ixp33_ASAP7_75t_L U14669 (.Y(n25981),
	.A1(n27127),
	.A2(FE_OCPN7622_n24526),
	.B(n24525),
	.C(n24524));
   OAI21xp5_ASAP7_75t_SL U14670 (.Y(n26757),
	.A1(FE_OFN1_ld_r),
	.A2(n27142),
	.B(n26758));
   OAI22xp5_ASAP7_75t_L U14671 (.Y(n604),
	.A1(ld),
	.A2(FE_OFN16360_n16051),
	.B1(key_35_),
	.B2(FE_OFN16360_n16051));
   OAI21xp33_ASAP7_75t_SRAM U14672 (.Y(n588),
	.A1(key_90_),
	.A2(FE_OFN22_n16125),
	.B(n16067));
   NOR2xp67_ASAP7_75t_SL U14674 (.Y(n26590),
	.A(n27031),
	.B(n26591));
   OAI21xp33_ASAP7_75t_SRAM U14676 (.Y(n591),
	.A1(key_65_),
	.A2(FE_OFN28463_ld),
	.B(n14012));
   OAI21xp5_ASAP7_75t_SL U14678 (.Y(n26337),
	.A1(FE_OFN28482_ld_r),
	.A2(FE_OCPN27534_n),
	.B(n26338));
   OAI21xp5_ASAP7_75t_SL U14679 (.Y(n636),
	.A1(n16222),
	.A2(n25051),
	.B(n16221));
   OAI21xp33_ASAP7_75t_SRAM U14680 (.Y(n611),
	.A1(key_121_),
	.A2(FE_OFN28468_ld),
	.B(n15769));
   OAI21xp33_ASAP7_75t_SRAM U14681 (.Y(n621),
	.A1(key_80_),
	.A2(FE_OFN28462_ld),
	.B(n16077));
   NAND2xp5_ASAP7_75t_L U14682 (.Y(n26487),
	.A(n26892),
	.B(n26484));
   OAI21xp5_ASAP7_75t_SL U14683 (.Y(n26237),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(FE_OCPN28138_n26654),
	.B(n26238));
   OAI21xp33_ASAP7_75t_SRAM U14684 (.Y(n551),
	.A1(key_125_),
	.A2(FE_OFN28468_ld),
	.B(n14824));
   A2O1A1Ixp33_ASAP7_75t_SL U14685 (.Y(n26676),
	.A1(n26679),
	.A2(n26678),
	.B(FE_OCPN28279_n),
	.C(n26674));
   OAI21xp33_ASAP7_75t_SRAM U14688 (.Y(n549),
	.A1(key_86_),
	.A2(FE_OFN27_n16125),
	.B(n15775));
   FAx1_ASAP7_75t_SL U14689 (.SN(n26207),
	.A(FE_OCPN27363_n26649),
	.B(FE_OCPN27271_n26961),
	.CI(n26205));
   OAI21xp33_ASAP7_75t_L U14691 (.Y(n558),
	.A1(key_78_),
	.A2(FE_OFN25_n16125),
	.B(n14746));
   OAI21xp5_ASAP7_75t_SL U14692 (.Y(n643),
	.A1(n16110),
	.A2(n25961),
	.B(n16109));
   AOI22xp5_ASAP7_75t_SL U14693 (.Y(n24910),
	.A1(n26349),
	.A2(n24913),
	.B1(FE_OFN26531_n),
	.B2(n24907));
   OAI21xp5_ASAP7_75t_SL U14694 (.Y(n26283),
	.A1(FE_OFN16213_ld_r),
	.A2(n26285),
	.B(n26284));
   O2A1O1Ixp33_ASAP7_75t_SL U14695 (.Y(n25245),
	.A1(n27168),
	.A2(FE_OFN28500_FE_OCPN5078_n25823),
	.B(n25243),
	.C(n25242));
   OAI21xp33_ASAP7_75t_SRAM U14697 (.Y(n597),
	.A1(key_83_),
	.A2(FE_OFN27_n16125),
	.B(n16064));
   OAI21xp33_ASAP7_75t_SRAM U14698 (.Y(n609),
	.A1(key_81_),
	.A2(FE_OFN28462_ld),
	.B(n16049));
   OAI21xp33_ASAP7_75t_SRAM U14699 (.Y(n528),
	.A1(key_95_),
	.A2(FE_OFN22_n16125),
	.B(n16057));
   A2O1A1Ixp33_ASAP7_75t_SL U14700 (.Y(n26961),
	.A1(n26942),
	.A2(n26201),
	.B(n26200),
	.C(n26199));
   NAND3xp33_ASAP7_75t_SL U14702 (.Y(n24107),
	.A(n24108),
	.B(FE_OFN16263_n25976),
	.C(n24109));
   OAI21xp33_ASAP7_75t_SRAM U14703 (.Y(n573),
	.A1(key_84_),
	.A2(FE_OFN27_n16125),
	.B(n16046));
   INVx1_ASAP7_75t_SL U14704 (.Y(n24825),
	.A(n24827));
   OAI21xp33_ASAP7_75t_SRAM U14705 (.Y(n534),
	.A1(key_79_),
	.A2(FE_OFN25_n16125),
	.B(n15900));
   OAI21xp33_ASAP7_75t_SRAM U14707 (.Y(n615),
	.A1(key_64_),
	.A2(FE_OFN25_n16125),
	.B(n14473));
   OAI21xp33_ASAP7_75t_SRAM U14708 (.Y(n587),
	.A1(key_122_),
	.A2(FE_OFN28468_ld),
	.B(n14329));
   OAI21xp33_ASAP7_75t_SRAM U14709 (.Y(n614),
	.A1(key_96_),
	.A2(FE_OFN28472_ld),
	.B(n13724));
   A2O1A1Ixp33_ASAP7_75t_SL U14710 (.Y(n26674),
	.A1(n26679),
	.A2(n25172),
	.B(n25171),
	.C(n25170));
   OAI21xp33_ASAP7_75t_SRAM U14711 (.Y(n620),
	.A1(key_112_),
	.A2(FE_OFN28462_ld),
	.B(n16043));
   OAI21xp33_ASAP7_75t_SRAM U14712 (.Y(n575),
	.A1(key_123_),
	.A2(FE_OFN28461_ld),
	.B(n15365));
   O2A1O1Ixp5_ASAP7_75t_SL U14714 (.Y(n26326),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(n25863),
	.C(n25862));
   OAI21xp33_ASAP7_75t_SRAM U14715 (.Y(n555),
	.A1(key_69_),
	.A2(FE_OFN28462_ld),
	.B(n14006));
   OAI21xp5_ASAP7_75t_SL U14716 (.Y(n16215),
	.A1(ld),
	.A2(w2_27_),
	.B(n16216));
   A2O1A1Ixp33_ASAP7_75t_SL U14717 (.Y(n26527),
	.A1(n27127),
	.A2(n25255),
	.B(n24573),
	.C(n24572));
   OAI21xp33_ASAP7_75t_SRAM U14718 (.Y(n564),
	.A1(key_92_),
	.A2(FE_OFN22_n16125),
	.B(n15908));
   A2O1A1Ixp33_ASAP7_75t_SL U14719 (.Y(n15268),
	.A1(n15270),
	.A2(n15271),
	.B(n15267),
	.C(n24506));
   OAI21xp33_ASAP7_75t_SRAM U14720 (.Y(n584),
	.A1(key_114_),
	.A2(FE_OFN26_n16125),
	.B(n15470));
   A2O1A1Ixp33_ASAP7_75t_L U14721 (.Y(n27157),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(n26366),
	.C(n26365));
   INVxp33_ASAP7_75t_SRAM U14722 (.Y(n26218),
	.A(FE_OCPN27884_n26717));
   OAI21xp33_ASAP7_75t_SRAM U14723 (.Y(n606),
	.A1(key_77_),
	.A2(FE_OFN25_n16125),
	.B(n16098));
   NAND2xp5_ASAP7_75t_L U14724 (.Y(n24482),
	.A(n27057),
	.B(FE_OFN29181_n24479));
   OAI21xp33_ASAP7_75t_SRAM U14725 (.Y(n603),
	.A1(key_67_),
	.A2(FE_OFN28463_ld),
	.B(n14092));
   OAI21xp33_ASAP7_75t_SRAM U14726 (.Y(n618),
	.A1(key_73_),
	.A2(FE_OFN28462_ld),
	.B(n15920));
   AOI22xp5_ASAP7_75t_L U14727 (.Y(n24240),
	.A1(FE_OFN29037_n),
	.A2(n24236),
	.B1(w1_6_),
	.B2(FE_OFN161_n26440));
   OAI21xp33_ASAP7_75t_R U14728 (.Y(n582),
	.A1(key_74_),
	.A2(FE_OFN25_n16125),
	.B(n16089));
   NOR3xp33_ASAP7_75t_SL U14729 (.Y(n25919),
	.A(FE_OCPN27522_n25921),
	.B(n27171),
	.C(n25920));
   NOR3xp33_ASAP7_75t_SL U14730 (.Y(n25405),
	.A(FE_PSN8314_n25722),
	.B(n25488),
	.C(n25406));
   NAND2xp5_ASAP7_75t_SL U14731 (.Y(n25365),
	.A(n25361),
	.B(n25360));
   FAx1_ASAP7_75t_SL U14732 (.SN(n26716),
	.A(n26713),
	.B(FE_OCPN27922_n26712),
	.CI(n26711));
   A2O1A1Ixp33_ASAP7_75t_SL U14733 (.Y(n26728),
	.A1(n22405),
	.A2(n24930),
	.B(n24929),
	.C(n24928));
   A2O1A1Ixp33_ASAP7_75t_SL U14734 (.Y(n25407),
	.A1(n26679),
	.A2(n25172),
	.B(n24583),
	.C(n24582));
   OAI21xp33_ASAP7_75t_SRAM U14735 (.Y(n540),
	.A1(key_94_),
	.A2(FE_OFN28472_ld),
	.B(n15905));
   NAND2xp5_ASAP7_75t_SL U14736 (.Y(n25801),
	.A(FE_OFN29024_n),
	.B(n25798));
   OAI21xp33_ASAP7_75t_R U14738 (.Y(n570),
	.A1(key_76_),
	.A2(FE_OFN25_n16125),
	.B(n16074));
   O2A1O1Ixp33_ASAP7_75t_SL U14739 (.Y(n26128),
	.A1(FE_OFN16180_n26542),
	.A2(n26127),
	.B(n26126),
	.C(n26125));
   NAND2xp5_ASAP7_75t_SL U14740 (.Y(n26200),
	.A(n26197),
	.B(n26507));
   OAI21xp33_ASAP7_75t_SRAM U14741 (.Y(n539),
	.A1(key_126_),
	.A2(FE_OFN28467_ld),
	.B(n14409));
   INVxp67_ASAP7_75t_L U14743 (.Y(n27200),
	.A(n27202));
   AOI22x1_ASAP7_75t_SL U14744 (.Y(n16091),
	.A1(w1_14_),
	.A2(FE_OFN27218_n14745),
	.B1(n14744),
	.B2(n25499));
   A2O1A1Ixp33_ASAP7_75t_SL U14745 (.Y(n26215),
	.A1(FE_OFN16169_n26567),
	.A2(FE_OFN28506_n26996),
	.B(n25450),
	.C(n25449));
   OAI21xp33_ASAP7_75t_SRAM U14746 (.Y(n546),
	.A1(key_75_),
	.A2(FE_OFN28464_ld),
	.B(n16118));
   O2A1O1Ixp33_ASAP7_75t_L U14747 (.Y(n26778),
	.A1(n26777),
	.A2(n26776),
	.B(n26775),
	.C(n26774));
   NAND3xp33_ASAP7_75t_SL U14748 (.Y(n26648),
	.A(FE_OCPN29471_n24175),
	.B(n26651),
	.C(n26649));
   NAND3xp33_ASAP7_75t_SL U14750 (.Y(n24386),
	.A(n25688),
	.B(n24388),
	.C(n24387));
   NAND2xp33_ASAP7_75t_L U14751 (.Y(n26752),
	.A(FE_OCPN27541_n26748),
	.B(n26747));
   NAND2xp5_ASAP7_75t_SL U14752 (.Y(n25973),
	.A(n26477),
	.B(n25970));
   XNOR2x2_ASAP7_75t_SL U14753 (.Y(n16138),
	.A(u0_rcon_25_),
	.B(n15768));
   A2O1A1Ixp33_ASAP7_75t_SL U14754 (.Y(n24684),
	.A1(n26819),
	.A2(FE_OCPN8227_n25950),
	.B(n24009),
	.C(n24008));
   OAI21xp33_ASAP7_75t_SRAM U14755 (.Y(n561),
	.A1(key_85_),
	.A2(FE_OFN27_n16125),
	.B(n14827));
   A2O1A1Ixp33_ASAP7_75t_SL U14756 (.Y(n24631),
	.A1(n26082),
	.A2(n24633),
	.B(n24630),
	.C(FE_OFN117_n24628));
   OAI21xp33_ASAP7_75t_SRAM U14757 (.Y(n590),
	.A1(key_97_),
	.A2(FE_OFN28471_ld),
	.B(n13480));
   NAND2xp5_ASAP7_75t_SL U14759 (.Y(n25171),
	.A(n25167),
	.B(n25166));
   NAND2xp5_ASAP7_75t_L U14762 (.Y(n24929),
	.A(FE_OCPN29539_n24927),
	.B(n24924));
   OAI21xp33_ASAP7_75t_SRAM U14764 (.Y(n602),
	.A1(key_99_),
	.A2(FE_OFN28471_ld),
	.B(n13549));
   INVx2_ASAP7_75t_SL U14765 (.Y(n26507),
	.A(n26508));
   NOR2xp33_ASAP7_75t_SL U14766 (.Y(n25333),
	.A(n26749),
	.B(FE_OFN26650_n27164));
   NOR3xp33_ASAP7_75t_SL U14768 (.Y(n24197),
	.A(FE_OCPN5077_n25855),
	.B(n24198),
	.C(n25856));
   OAI21xp33_ASAP7_75t_SRAM U14769 (.Y(n605),
	.A1(key_109_),
	.A2(FE_OFN26_n16125),
	.B(n15143));
   A2O1A1Ixp33_ASAP7_75t_SL U14770 (.Y(n27079),
	.A1(FE_OFN16176_n27207),
	.A2(n27192),
	.B(n25829),
	.C(n25828));
   A2O1A1Ixp33_ASAP7_75t_L U14771 (.Y(n24008),
	.A1(n26819),
	.A2(FE_OCPN8227_n25950),
	.B(n25947),
	.C(n24007));
   INVx1_ASAP7_75t_SL U14773 (.Y(n16076),
	.A(n16075));
   A2O1A1Ixp33_ASAP7_75t_L U14775 (.Y(n25940),
	.A1(n27183),
	.A2(n27182),
	.B(n25925),
	.C(n25924));
   NOR2xp33_ASAP7_75t_L U14776 (.Y(n25863),
	.A(n26508),
	.B(n26954));
   NAND2xp5_ASAP7_75t_L U14777 (.Y(n25724),
	.A(FE_OCPN29457_n25722),
	.B(n25719));
   A2O1A1Ixp33_ASAP7_75t_SL U14779 (.Y(n13630),
	.A1(n13628),
	.A2(n13627),
	.B(n13689),
	.C(n13626));
   NOR2xp33_ASAP7_75t_R U14780 (.Y(n26775),
	.A(w0_3_),
	.B(n26771));
   A2O1A1Ixp33_ASAP7_75t_SL U14781 (.Y(n26172),
	.A1(n26139),
	.A2(n25178),
	.B(n25177),
	.C(n25176));
   OAI21xp33_ASAP7_75t_SRAM U14782 (.Y(n596),
	.A1(key_115_),
	.A2(FE_OFN22_n16125),
	.B(n14972));
   O2A1O1Ixp33_ASAP7_75t_SL U14784 (.Y(n25755),
	.A1(FE_OFN16413_n26687),
	.A2(n26258),
	.B(n25125),
	.C(n25124));
   XNOR2x2_ASAP7_75t_SL U14785 (.Y(n16080),
	.A(w1_0_),
	.B(n13723));
   OAI21xp33_ASAP7_75t_SRAM U14787 (.Y(n537),
	.A1(key_87_),
	.A2(FE_OFN28462_ld),
	.B(n14975));
   O2A1O1Ixp5_ASAP7_75t_SL U14788 (.Y(n26049),
	.A1(n27102),
	.A2(n25240),
	.B(n25239),
	.C(n25238));
   A2O1A1Ixp33_ASAP7_75t_L U14789 (.Y(n26845),
	.A1(n26857),
	.A2(n26793),
	.B(n25009),
	.C(n25008));
   NOR2xp33_ASAP7_75t_SL U14790 (.Y(n24981),
	.A(FE_OFN28582_n25657),
	.B(n25132));
   A2O1A1Ixp33_ASAP7_75t_SL U14791 (.Y(n26780),
	.A1(FE_OFN16170_n26637),
	.A2(n26226),
	.B(n26086),
	.C(n26085));
   NAND2xp5_ASAP7_75t_L U14795 (.Y(n26086),
	.A(FE_OCPN27394_n26223),
	.B(n26866));
   A2O1A1Ixp33_ASAP7_75t_SL U14797 (.Y(n24384),
	.A1(n25736),
	.A2(n26249),
	.B(n26178),
	.C(n24383));
   A2O1A1Ixp33_ASAP7_75t_SL U14798 (.Y(n15262),
	.A1(n15261),
	.A2(n15260),
	.B(n15259),
	.C(n15258));
   OAI21xp33_ASAP7_75t_SRAM U14799 (.Y(n581),
	.A1(key_106_),
	.A2(FE_OFN26_n16125),
	.B(n15060));
   INVx1_ASAP7_75t_L U14800 (.Y(n16122),
	.A(FE_OCPN28186_n16123));
   OAI21xp33_ASAP7_75t_SRAM U14802 (.Y(n560),
	.A1(key_117_),
	.A2(FE_OFN26_n16125),
	.B(n14003));
   A2O1A1Ixp33_ASAP7_75t_SL U14804 (.Y(n26922),
	.A1(FE_OFN16169_n26567),
	.A2(n24812),
	.B(n24811),
	.C(n24810));
   OAI21xp33_ASAP7_75t_SRAM U14805 (.Y(n545),
	.A1(key_107_),
	.A2(FE_OFN28460_ld),
	.B(n15897));
   AOI22xp5_ASAP7_75t_SL U14806 (.Y(n16219),
	.A1(w1_10_),
	.A2(n16088),
	.B1(n16087),
	.B2(n26041));
   A2O1A1Ixp33_ASAP7_75t_L U14807 (.Y(n24818),
	.A1(FE_OCPN5172_n26281),
	.A2(n26282),
	.B(FE_OFN27123_n26275),
	.C(n24817));
   A2O1A1Ixp33_ASAP7_75t_SL U14809 (.Y(n27121),
	.A1(n23567),
	.A2(n23566),
	.B(n24331),
	.C(n23565));
   A2O1A1Ixp33_ASAP7_75t_SL U14812 (.Y(n25357),
	.A1(n22350),
	.A2(n20354),
	.B(n24263),
	.C(n20353));
   O2A1O1Ixp5_ASAP7_75t_SL U14813 (.Y(n26773),
	.A1(n24518),
	.A2(n24104),
	.B(n27127),
	.C(n24103));
   A2O1A1Ixp33_ASAP7_75t_L U14814 (.Y(n26616),
	.A1(n27183),
	.A2(n27182),
	.B(n27177),
	.C(w2_7_));
   O2A1O1Ixp33_ASAP7_75t_SL U14815 (.Y(n25263),
	.A1(n26542),
	.A2(n26431),
	.B(n26428),
	.C(n25262));
   A2O1A1Ixp33_ASAP7_75t_SL U14816 (.Y(n25462),
	.A1(n23469),
	.A2(n23468),
	.B(n23467),
	.C(n23466));
   A2O1A1Ixp33_ASAP7_75t_SL U14818 (.Y(n25250),
	.A1(n24303),
	.A2(n24302),
	.B(n26542),
	.C(n24301));
   O2A1O1Ixp5_ASAP7_75t_SL U14821 (.Y(n26317),
	.A1(n25536),
	.A2(n25535),
	.B(n27216),
	.C(n27212));
   A2O1A1Ixp33_ASAP7_75t_SL U14822 (.Y(n25176),
	.A1(n26139),
	.A2(n25178),
	.B(n25748),
	.C(n26574));
   A2O1A1Ixp33_ASAP7_75t_SL U14824 (.Y(n16063),
	.A1(n14971),
	.A2(n14970),
	.B(n14969),
	.C(n14968));
   A2O1A1Ixp33_ASAP7_75t_SL U14825 (.Y(n24175),
	.A1(n25299),
	.A2(n22913),
	.B(n26976),
	.C(n22912));
   A2O1A1Ixp33_ASAP7_75t_SL U14826 (.Y(n16048),
	.A1(n16042),
	.A2(n14742),
	.B(n14741),
	.C(n14740));
   OAI21xp33_ASAP7_75t_SRAM U14827 (.Y(n536),
	.A1(key_119_),
	.A2(FE_OFN22_n16125),
	.B(n13866));
   A2O1A1Ixp33_ASAP7_75t_L U14828 (.Y(n14005),
	.A1(n13595),
	.A2(n13333),
	.B(n13332),
	.C(n13331));
   NOR3xp33_ASAP7_75t_SL U14829 (.Y(n13720),
	.A(n13722),
	.B(w0_0_),
	.C(n13721));
   O2A1O1Ixp5_ASAP7_75t_SL U14830 (.Y(n24977),
	.A1(n24976),
	.A2(n24975),
	.B(n24974),
	.C(n24973));
   A2O1A1Ixp33_ASAP7_75t_SL U14831 (.Y(n26369),
	.A1(n21435),
	.A2(n21434),
	.B(n26078),
	.C(n21433));
   A2O1A1Ixp33_ASAP7_75t_SL U14835 (.Y(n26528),
	.A1(n22276),
	.A2(n21811),
	.B(n23345),
	.C(n21810));
   A2O1A1Ixp33_ASAP7_75t_L U14836 (.Y(n16039),
	.A1(n16041),
	.A2(n16042),
	.B(n16038),
	.C(n26486));
   A2O1A1Ixp33_ASAP7_75t_SL U14837 (.Y(n26938),
	.A1(n21999),
	.A2(n21998),
	.B(n26315),
	.C(n21997));
   INVxp67_ASAP7_75t_L U14842 (.Y(n24931),
	.A(n24932));
   NAND2xp5_ASAP7_75t_SL U14843 (.Y(n14247),
	.A(n14244),
	.B(n26272));
   O2A1O1Ixp5_ASAP7_75t_SL U14846 (.Y(n24904),
	.A1(n24901),
	.A2(n24900),
	.B(n26857),
	.C(n24899));
   A2O1A1Ixp33_ASAP7_75t_SL U14847 (.Y(n15140),
	.A1(FE_OFN16411_n15884),
	.A2(n15142),
	.B(n15139),
	.C(w0_13_));
   NAND2xp5_ASAP7_75t_SL U14848 (.Y(n24973),
	.A(n24972),
	.B(n24971));
   INVx1_ASAP7_75t_SL U14849 (.Y(n25262),
	.A(n25261));
   A2O1A1Ixp33_ASAP7_75t_SL U14850 (.Y(n27179),
	.A1(n22573),
	.A2(n22572),
	.B(n27140),
	.C(n22571));
   OAI21xp5_ASAP7_75t_SL U14852 (.Y(n15256),
	.A1(n15253),
	.A2(n15252),
	.B(n15251));
   NOR2x1_ASAP7_75t_SL U14854 (.Y(n25418),
	.A(FE_OFN16179_w3_19),
	.B(FE_OFN28902_n25414));
   OA21x2_ASAP7_75t_SL U14855 (.Y(n24420),
	.A1(n24419),
	.A2(n26710),
	.B(n24418));
   AND2x2_ASAP7_75t_SL U14856 (.Y(n13622),
	.A(n13619),
	.B(n13618));
   NAND2xp5_ASAP7_75t_L U14857 (.Y(n23970),
	.A(n23965),
	.B(n23966));
   NAND2xp5_ASAP7_75t_SL U14858 (.Y(n21056),
	.A(n21055),
	.B(n21054));
   A2O1A1Ixp33_ASAP7_75t_SL U14859 (.Y(n13796),
	.A1(FE_OFN16411_n15884),
	.A2(n13798),
	.B(n13795),
	.C(w0_14_));
   O2A1O1Ixp5_ASAP7_75t_SL U14860 (.Y(n24803),
	.A1(FE_OCPN5109_n26551),
	.A2(n24777),
	.B(n26567),
	.C(FE_OCPN27507_n25695));
   O2A1O1Ixp5_ASAP7_75t_SL U14861 (.Y(n21810),
	.A1(n22308),
	.A2(n21809),
	.B(n26878),
	.C(n21808));
   A2O1A1Ixp33_ASAP7_75t_SL U14862 (.Y(n26491),
	.A1(n20183),
	.A2(n20182),
	.B(n26976),
	.C(n20181));
   NAND3xp33_ASAP7_75t_SL U14863 (.Y(n24005),
	.A(n23991),
	.B(n23990),
	.C(n23989));
   AOI21x1_ASAP7_75t_SL U14864 (.Y(n24932),
	.A1(n26857),
	.A2(n26856),
	.B(n26853));
   NAND2xp5_ASAP7_75t_SL U14866 (.Y(n21054),
	.A(n21053),
	.B(n21052));
   A2O1A1Ixp33_ASAP7_75t_SL U14867 (.Y(n24750),
	.A1(n19888),
	.A2(n16827),
	.B(n24263),
	.C(n16826));
   O2A1O1Ixp5_ASAP7_75t_SL U14868 (.Y(n27094),
	.A1(FE_OCPN28115_n25293),
	.A2(n25292),
	.B(n26915),
	.C(n25291));
   O2A1O1Ixp5_ASAP7_75t_SL U14870 (.Y(n25232),
	.A1(n25231),
	.A2(n25230),
	.B(n26915),
	.C(n25229));
   NAND2xp5_ASAP7_75t_L U14872 (.Y(n21055),
	.A(n21050),
	.B(n21052));
   A2O1A1Ixp33_ASAP7_75t_SL U14873 (.Y(n27020),
	.A1(n23480),
	.A2(n22055),
	.B(n26710),
	.C(n22054));
   A2O1A1Ixp33_ASAP7_75t_SL U14874 (.Y(n27203),
	.A1(n25628),
	.A2(n23736),
	.B(n26517),
	.C(n23735));
   NOR2x1_ASAP7_75t_L U14875 (.Y(n18155),
	.A(n18127),
	.B(n18126));
   NAND2x1p5_ASAP7_75t_SL U14876 (.Y(n26404),
	.A(n20042),
	.B(n20041));
   A2O1A1Ixp33_ASAP7_75t_SL U14878 (.Y(n16732),
	.A1(n16742),
	.A2(n16741),
	.B(n24331),
	.C(n16731));
   NAND2xp33_ASAP7_75t_L U14879 (.Y(n24109),
	.A(n27117),
	.B(FE_OFN28690_n25979));
   A2O1A1Ixp33_ASAP7_75t_SL U14881 (.Y(n25556),
	.A1(n25555),
	.A2(n25554),
	.B(n27095),
	.C(n25553));
   NOR2x1_ASAP7_75t_SL U14882 (.Y(n24809),
	.A(n26441),
	.B(n26442));
   A2O1A1Ixp33_ASAP7_75t_L U14884 (.Y(n14968),
	.A1(n14971),
	.A2(n14970),
	.B(n14967),
	.C(w0_19_));
   NAND3xp33_ASAP7_75t_SL U14885 (.Y(n22650),
	.A(n22639),
	.B(n22638),
	.C(n25121));
   A2O1A1Ixp33_ASAP7_75t_SL U14886 (.Y(n25956),
	.A1(n23674),
	.A2(n23673),
	.B(n24263),
	.C(n23672));
   NAND2x1p5_ASAP7_75t_SL U14887 (.Y(n24449),
	.A(n24274),
	.B(n24273));
   O2A1O1Ixp33_ASAP7_75t_SL U14888 (.Y(n20948),
	.A1(n20947),
	.A2(n20946),
	.B(n26249),
	.C(n20945));
   NOR2xp33_ASAP7_75t_SL U14889 (.Y(n14598),
	.A(n14596),
	.B(n14595));
   NAND2xp5_ASAP7_75t_SL U14890 (.Y(n23202),
	.A(n23181),
	.B(n23180));
   A2O1A1Ixp33_ASAP7_75t_SL U14891 (.Y(n26002),
	.A1(n26001),
	.A2(n26000),
	.B(n26959),
	.C(n25999));
   NAND3xp33_ASAP7_75t_L U14892 (.Y(n19324),
	.A(n19323),
	.B(n22007),
	.C(n19322));
   OAI222xp33_ASAP7_75t_L U14893 (.Y(n20535),
	.A1(n20531),
	.A2(n27102),
	.B1(n20520),
	.B2(n27102),
	.C1(n20519),
	.C2(n27102));
   NOR2x1_ASAP7_75t_L U14894 (.Y(n21003),
	.A(n21001),
	.B(n21000));
   NAND2xp33_ASAP7_75t_SL U14895 (.Y(n13617),
	.A(n13611),
	.B(n13614));
   A2O1A1Ixp33_ASAP7_75t_SL U14896 (.Y(n25340),
	.A1(n26045),
	.A2(n26044),
	.B(n27168),
	.C(n26050));
   NAND2xp33_ASAP7_75t_SL U14899 (.Y(n13616),
	.A(n13615),
	.B(n13614));
   NAND2xp33_ASAP7_75t_SL U14900 (.Y(n13367),
	.A(n13366),
	.B(n13365));
   A2O1A1Ixp33_ASAP7_75t_SL U14902 (.Y(n25485),
	.A1(n22266),
	.A2(n22265),
	.B(n24377),
	.C(n22264));
   A2O1A1Ixp33_ASAP7_75t_L U14903 (.Y(n14468),
	.A1(FE_OFN16411_n15884),
	.A2(n14470),
	.B(n14467),
	.C(w0_9_));
   NOR2xp67_ASAP7_75t_L U14904 (.Y(n15138),
	.A(n15137),
	.B(n15136));
   A2O1A1Ixp33_ASAP7_75t_SL U14905 (.Y(n14891),
	.A1(n14890),
	.A2(n14889),
	.B(FE_OFN28682_n15888),
	.C(n14888));
   NAND2xp5_ASAP7_75t_SL U14906 (.Y(n22896),
	.A(n20977),
	.B(n20976));
   OAI21xp5_ASAP7_75t_SL U14907 (.Y(n21954),
	.A1(n21953),
	.A2(n26315),
	.B(n21952));
   O2A1O1Ixp33_ASAP7_75t_L U14908 (.Y(n19619),
	.A1(n19618),
	.A2(n19617),
	.B(n26637),
	.C(n19616));
   A2O1A1Ixp33_ASAP7_75t_SL U14909 (.Y(n14967),
	.A1(n14965),
	.A2(n14964),
	.B(n15969),
	.C(n14963));
   NAND2xp33_ASAP7_75t_SL U14910 (.Y(n23180),
	.A(n23179),
	.B(n23178));
   NOR3xp33_ASAP7_75t_SL U14911 (.Y(n26572),
	.A(n18999),
	.B(n19331),
	.C(n18998));
   O2A1O1Ixp33_ASAP7_75t_SL U14912 (.Y(n25999),
	.A1(n25885),
	.A2(n25884),
	.B(n26915),
	.C(n25883));
   NAND3xp33_ASAP7_75t_SL U14913 (.Y(n25824),
	.A(n24191),
	.B(n18099),
	.C(n18098));
   NAND2xp5_ASAP7_75t_SL U14914 (.Y(n20042),
	.A(n20038),
	.B(n20039));
   A2O1A1Ixp33_ASAP7_75t_SL U14915 (.Y(n26853),
	.A1(n19683),
	.A2(n16670),
	.B(n24978),
	.C(n16669));
   NAND3xp33_ASAP7_75t_R U14916 (.Y(n18234),
	.A(n18212),
	.B(n18211),
	.C(n23175));
   NOR2xp33_ASAP7_75t_SL U14918 (.Y(n14319),
	.A(n14308),
	.B(n13901));
   NOR2xp33_ASAP7_75t_SL U14919 (.Y(n20448),
	.A(n24762),
	.B(n20445));
   NAND2xp33_ASAP7_75t_SRAM U14921 (.Y(n26109),
	.A(n26108),
	.B(FE_OFN163_sa00_7));
   NAND2xp5_ASAP7_75t_L U14922 (.Y(n20976),
	.A(n20975),
	.B(n20974));
   NAND2xp33_ASAP7_75t_SL U14924 (.Y(n20977),
	.A(n20972),
	.B(n20974));
   NAND2xp5_ASAP7_75t_L U14925 (.Y(n19323),
	.A(n19320),
	.B(n19319));
   OAI222xp33_ASAP7_75t_SRAM U14926 (.Y(n26682),
	.A1(n26671),
	.A2(n27027),
	.B1(n26670),
	.B2(n27027),
	.C1(n26669),
	.C2(n27027));
   NAND3xp33_ASAP7_75t_SL U14927 (.Y(n21423),
	.A(n25792),
	.B(n21421),
	.C(FE_OCPN29554_n22507));
   O2A1O1Ixp5_ASAP7_75t_SL U14928 (.Y(n27014),
	.A1(n22609),
	.A2(n22608),
	.B(n26282),
	.C(n22607));
   NOR2xp33_ASAP7_75t_SL U14929 (.Y(n13366),
	.A(n13364),
	.B(n13363));
   NAND2xp5_ASAP7_75t_SL U14930 (.Y(n15734),
	.A(n15733),
	.B(n15732));
   OAI21xp5_ASAP7_75t_L U14931 (.Y(n25305),
	.A1(n25304),
	.A2(n25303),
	.B(n27216));
   NOR2xp33_ASAP7_75t_SL U14932 (.Y(n13362),
	.A(FE_OFN28929_n15182),
	.B(n13363));
   NAND3xp33_ASAP7_75t_SL U14933 (.Y(n18113),
	.A(n18106),
	.B(n18446),
	.C(n18105));
   NAND2xp5_ASAP7_75t_R U14934 (.Y(n13765),
	.A(n13756),
	.B(n13762));
   NAND2xp33_ASAP7_75t_L U14935 (.Y(n13493),
	.A(n13492),
	.B(n13491));
   NAND2xp5_ASAP7_75t_R U14936 (.Y(n13764),
	.A(n13763),
	.B(n13762));
   NOR3xp33_ASAP7_75t_SL U14937 (.Y(n16524),
	.A(n16522),
	.B(n18095),
	.C(n16521));
   A2O1A1Ixp33_ASAP7_75t_SL U14938 (.Y(n13999),
	.A1(n13997),
	.A2(n13996),
	.B(n16023),
	.C(n13995));
   A2O1A1Ixp33_ASAP7_75t_SL U14939 (.Y(n23406),
	.A1(n23405),
	.A2(n23404),
	.B(n26078),
	.C(n23403));
   NAND2xp33_ASAP7_75t_SL U14940 (.Y(n25292),
	.A(n25290),
	.B(n25289));
   OR3x1_ASAP7_75t_L U14941 (.Y(n20752),
	.A(n22856),
	.B(n20748),
	.C(n21779));
   NAND3xp33_ASAP7_75t_SL U14943 (.Y(n25117),
	.A(n25115),
	.B(n25114),
	.C(n25113));
   NAND2xp33_ASAP7_75t_L U14944 (.Y(n14889),
	.A(n14885),
	.B(n14884));
   NAND2xp33_ASAP7_75t_SL U14946 (.Y(n14877),
	.A(n14876),
	.B(n14875));
   NAND2xp5_ASAP7_75t_SL U14947 (.Y(n23018),
	.A(n21881),
	.B(n21880));
   NAND3xp33_ASAP7_75t_SL U14948 (.Y(n26856),
	.A(n16628),
	.B(n16627),
	.C(n19694));
   OAI21xp5_ASAP7_75t_L U14949 (.Y(n14822),
	.A1(n15506),
	.A2(FE_OCPN8264_n13890),
	.B(n14763));
   AND2x2_ASAP7_75t_SRAM U14950 (.Y(n19247),
	.A(n19246),
	.B(n25213));
   NOR3x1_ASAP7_75t_SL U14952 (.Y(n19141),
	.A(n18769),
	.B(n18768),
	.C(n24096));
   NOR3xp33_ASAP7_75t_SL U14953 (.Y(n19477),
	.A(n19474),
	.B(n19473),
	.C(n23423));
   NOR3xp33_ASAP7_75t_L U14955 (.Y(n19859),
	.A(n19830),
	.B(n24478),
	.C(n19829));
   AO21x1_ASAP7_75t_L U14956 (.Y(n23808),
	.A1(n25642),
	.A2(n25643),
	.B(n25641));
   NAND2xp5_ASAP7_75t_SL U14957 (.Y(n20763),
	.A(n20762),
	.B(n20761));
   A2O1A1Ixp33_ASAP7_75t_L U14958 (.Y(n14465),
	.A1(n14438),
	.A2(n14437),
	.B(n14436),
	.C(n15896));
   NAND2xp33_ASAP7_75t_L U14959 (.Y(n19583),
	.A(n19582),
	.B(n19581));
   NOR2xp33_ASAP7_75t_L U14960 (.Y(n19112),
	.A(n24344),
	.B(n19105));
   NAND3xp33_ASAP7_75t_L U14961 (.Y(n21955),
	.A(n20855),
	.B(n21931),
	.C(n21992));
   NAND2xp5_ASAP7_75t_L U14962 (.Y(n19221),
	.A(n19216),
	.B(n19218));
   NAND2xp5_ASAP7_75t_SL U14963 (.Y(n19220),
	.A(n19219),
	.B(n19218));
   O2A1O1Ixp33_ASAP7_75t_L U14964 (.Y(n13995),
	.A1(n13994),
	.A2(n13993),
	.B(n16042),
	.C(n13992));
   NOR3xp33_ASAP7_75t_SL U14965 (.Y(n21132),
	.A(n21131),
	.B(n21130),
	.C(FE_OFN26009_n18213));
   AND2x2_ASAP7_75t_SRAM U14966 (.Y(n22707),
	.A(n22706),
	.B(n22705));
   NOR3x1_ASAP7_75t_SL U14968 (.Y(n22957),
	.A(n18997),
	.B(n19306),
	.C(n18996));
   NAND2xp5_ASAP7_75t_L U14969 (.Y(n25339),
	.A(n25338),
	.B(n25337));
   NAND2xp5_ASAP7_75t_L U14970 (.Y(n15732),
	.A(n15731),
	.B(n15730));
   NAND2xp5_ASAP7_75t_L U14971 (.Y(n15733),
	.A(n15727),
	.B(n15730));
   NAND2x1_ASAP7_75t_SL U14972 (.Y(n20997),
	.A(n17755),
	.B(n17754));
   NOR3x1_ASAP7_75t_SL U14973 (.Y(n25881),
	.A(n18916),
	.B(n19411),
	.C(n25199));
   OAI21xp33_ASAP7_75t_SL U14975 (.Y(n14285),
	.A1(n13875),
	.A2(n15520),
	.B(n14284));
   NOR3x1_ASAP7_75t_SL U14976 (.Y(n18962),
	.A(n18961),
	.B(n25293),
	.C(n18960));
   NOR3xp33_ASAP7_75t_L U14978 (.Y(n22792),
	.A(n22757),
	.B(n22756),
	.C(n23237));
   NAND2xp5_ASAP7_75t_L U14979 (.Y(n17368),
	.A(n17362),
	.B(n17361));
   NAND2xp5_ASAP7_75t_SL U14980 (.Y(n20468),
	.A(n20465),
	.B(n20464));
   OAI222xp33_ASAP7_75t_L U14981 (.Y(n17982),
	.A1(n20572),
	.A2(n26607),
	.B1(n17938),
	.B2(n26607),
	.C1(n17937),
	.C2(n26607));
   NOR3x1_ASAP7_75t_L U14982 (.Y(n23175),
	.A(n18210),
	.B(n21799),
	.C(n18209));
   NOR3xp33_ASAP7_75t_SL U14983 (.Y(n18737),
	.A(n18735),
	.B(n18734),
	.C(n24094));
   OR3x1_ASAP7_75t_L U14984 (.Y(n19640),
	.A(n19639),
	.B(n19638),
	.C(FE_OCPN5156_n23958));
   NAND3xp33_ASAP7_75t_SL U14985 (.Y(n18997),
	.A(n18995),
	.B(n23483),
	.C(n22018));
   NAND3xp33_ASAP7_75t_L U14986 (.Y(n22556),
	.A(n22555),
	.B(n22554),
	.C(n22553));
   NOR2xp33_ASAP7_75t_L U14987 (.Y(n14876),
	.A(n14886),
	.B(n14887));
   NOR3x1_ASAP7_75t_L U14988 (.Y(n22036),
	.A(n22035),
	.B(FE_OCPN28086_n22034),
	.C(n22033));
   NAND2x1p5_ASAP7_75t_SL U14989 (.Y(n23460),
	.A(n21711),
	.B(n18022));
   NAND2xp33_ASAP7_75t_L U14990 (.Y(n19582),
	.A(n19577),
	.B(n19579));
   NAND3xp33_ASAP7_75t_SL U14991 (.Y(n18783),
	.A(n18762),
	.B(n18761),
	.C(n19812));
   NAND2xp33_ASAP7_75t_L U14992 (.Y(n19581),
	.A(n19580),
	.B(n19579));
   NAND2xp5_ASAP7_75t_R U14993 (.Y(n17361),
	.A(n17360),
	.B(n23088));
   NOR2xp33_ASAP7_75t_SL U14994 (.Y(n22593),
	.A(n23060),
	.B(n22185));
   NOR3xp33_ASAP7_75t_L U14995 (.Y(n18542),
	.A(n18539),
	.B(n23698),
	.C(n18538));
   NOR2xp33_ASAP7_75t_SL U14996 (.Y(n17101),
	.A(n17100),
	.B(n17099));
   NAND2xp5_ASAP7_75t_SL U14999 (.Y(n23334),
	.A(n20712),
	.B(n20711));
   AND2x2_ASAP7_75t_L U15000 (.Y(n23339),
	.A(n23338),
	.B(n23337));
   NOR3xp33_ASAP7_75t_L U15002 (.Y(n24568),
	.A(n24563),
	.B(FE_PSN8302_n24562),
	.C(n24561));
   A2O1A1Ixp33_ASAP7_75t_L U15003 (.Y(n13465),
	.A1(n13464),
	.A2(n13463),
	.B(n14585),
	.C(n13462));
   NOR3x1_ASAP7_75t_SL U15004 (.Y(n19883),
	.A(n19882),
	.B(n19968),
	.C(n22349));
   INVxp67_ASAP7_75t_L U15005 (.Y(n16511),
	.A(n16510));
   AND3x1_ASAP7_75t_L U15006 (.Y(n21404),
	.A(n21382),
	.B(n19205),
	.C(n19204));
   NAND3xp33_ASAP7_75t_L U15008 (.Y(n26075),
	.A(n26073),
	.B(n26072),
	.C(n26071));
   NAND2xp5_ASAP7_75t_SL U15009 (.Y(n15232),
	.A(n15231),
	.B(n15230));
   NAND2xp5_ASAP7_75t_L U15010 (.Y(n20006),
	.A(n20003),
	.B(n23650));
   AND2x2_ASAP7_75t_R U15011 (.Y(n17688),
	.A(n17687),
	.B(n17686));
   NAND3xp33_ASAP7_75t_L U15012 (.Y(n24611),
	.A(n18447),
	.B(n18446),
	.C(n18445));
   NAND2x1_ASAP7_75t_SL U15013 (.Y(n24953),
	.A(n16572),
	.B(n16571));
   NOR3xp33_ASAP7_75t_SL U15014 (.Y(n18423),
	.A(n18419),
	.B(n23544),
	.C(FE_OFN16218_n18418));
   OAI222xp33_ASAP7_75t_L U15015 (.Y(n17440),
	.A1(n17423),
	.A2(n26542),
	.B1(n17422),
	.B2(n26542),
	.C1(n17421),
	.C2(n26542));
   NAND2xp5_ASAP7_75t_SL U15016 (.Y(n19637),
	.A(n16561),
	.B(n16560));
   NOR3x1_ASAP7_75t_SL U15017 (.Y(n19782),
	.A(n23051),
	.B(n21906),
	.C(n16651));
   NAND2xp33_ASAP7_75t_SL U15018 (.Y(n14648),
	.A(n14647),
	.B(n14643));
   NAND2xp33_ASAP7_75t_R U15019 (.Y(n23469),
	.A(n23437),
	.B(n23436));
   OR3x1_ASAP7_75t_SL U15020 (.Y(n18385),
	.A(n22645),
	.B(n18372),
	.C(n18371));
   NAND2xp33_ASAP7_75t_SL U15021 (.Y(n13608),
	.A(n13603),
	.B(n13605));
   NOR2x1_ASAP7_75t_SL U15022 (.Y(n18022),
	.A(n18859),
	.B(n18021));
   NOR3xp33_ASAP7_75t_SL U15023 (.Y(n20604),
	.A(n20601),
	.B(n23581),
	.C(n22258));
   OAI21xp33_ASAP7_75t_SL U15026 (.Y(n21990),
	.A1(FE_OCPN29483_FE_OFN26014_sa31_3),
	.A2(n20081),
	.B(n20080));
   NOR3xp33_ASAP7_75t_L U15027 (.Y(n18447),
	.A(n18444),
	.B(FE_OFN27090_n23558),
	.C(n18443));
   NOR3xp33_ASAP7_75t_SL U15028 (.Y(n17304),
	.A(n18771),
	.B(n26101),
	.C(n19578));
   NOR2xp33_ASAP7_75t_SL U15029 (.Y(n21488),
	.A(n18623),
	.B(n17270));
   NAND2x1p5_ASAP7_75t_SL U15030 (.Y(n24172),
	.A(n17158),
	.B(n17157));
   OR2x2_ASAP7_75t_SL U15031 (.Y(n19307),
	.A(n19306),
	.B(n19305));
   OAI21xp33_ASAP7_75t_L U15033 (.Y(n14470),
	.A1(FE_OFN26084_n15106),
	.A2(n15610),
	.B(n14421));
   NAND2xp5_ASAP7_75t_SL U15034 (.Y(n15126),
	.A(n15123),
	.B(n15122));
   NAND2xp5_ASAP7_75t_L U15035 (.Y(n16714),
	.A(n16713),
	.B(n16870));
   NAND2xp5_ASAP7_75t_L U15036 (.Y(n16715),
	.A(n16712),
	.B(n16870));
   NAND2xp5_ASAP7_75t_SL U15037 (.Y(n17293),
	.A(n17281),
	.B(n17280));
   NAND2xp5_ASAP7_75t_L U15039 (.Y(n20712),
	.A(n20708),
	.B(n20709));
   NAND2xp5_ASAP7_75t_L U15040 (.Y(n20711),
	.A(n20710),
	.B(n20709));
   NAND3xp33_ASAP7_75t_SL U15041 (.Y(n18270),
	.A(n18268),
	.B(n20509),
	.C(n25227));
   NAND3xp33_ASAP7_75t_SL U15042 (.Y(n20165),
	.A(n20164),
	.B(n22902),
	.C(n22084));
   NOR3x1_ASAP7_75t_SL U15043 (.Y(n18763),
	.A(n18641),
	.B(n19586),
	.C(n24089));
   AND2x2_ASAP7_75t_R U15045 (.Y(n22181),
	.A(n22180),
	.B(n22179));
   NOR2x1_ASAP7_75t_L U15046 (.Y(n19370),
	.A(n18276),
	.B(n18275));
   NAND2xp5_ASAP7_75t_SL U15048 (.Y(n21556),
	.A(n21554),
	.B(n22468));
   AND2x2_ASAP7_75t_SRAM U15049 (.Y(n22246),
	.A(n22245),
	.B(n23227));
   NOR3xp33_ASAP7_75t_L U15050 (.Y(n26079),
	.A(n21361),
	.B(n21360),
	.C(n21359));
   NAND2xp5_ASAP7_75t_SL U15051 (.Y(n20804),
	.A(n20803),
	.B(n20802));
   NOR3xp33_ASAP7_75t_SRAM U15052 (.Y(n22409),
	.A(n22385),
	.B(n22384),
	.C(n22383));
   NOR3xp33_ASAP7_75t_SL U15053 (.Y(n20164),
	.A(n20163),
	.B(FE_OCPN27652_n20176),
	.C(n20162));
   NAND2x1_ASAP7_75t_SL U15054 (.Y(n16728),
	.A(n17412),
	.B(n16722));
   NOR3xp33_ASAP7_75t_SL U15055 (.Y(n18224),
	.A(n18218),
	.B(n23164),
	.C(n18217));
   NAND2xp5_ASAP7_75t_SL U15057 (.Y(n23544),
	.A(n18125),
	.B(n16888));
   AND2x2_ASAP7_75t_L U15058 (.Y(n19667),
	.A(n19666),
	.B(n24669));
   NOR3xp33_ASAP7_75t_SL U15059 (.Y(n17049),
	.A(n17047),
	.B(n17105),
	.C(n17165));
   AND3x1_ASAP7_75t_SL U15060 (.Y(n16571),
	.A(n16570),
	.B(n16569),
	.C(n16661));
   NAND3xp33_ASAP7_75t_SL U15061 (.Y(n23376),
	.A(n22495),
	.B(n21841),
	.C(n21840));
   NAND3xp33_ASAP7_75t_SL U15062 (.Y(n17016),
	.A(n17162),
	.B(n19424),
	.C(n17014));
   NAND2x1_ASAP7_75t_SL U15063 (.Y(n17158),
	.A(n17153),
	.B(n17155));
   NAND2x1_ASAP7_75t_SL U15064 (.Y(n17157),
	.A(n17156),
	.B(n17155));
   NAND2xp5_ASAP7_75t_SL U15066 (.Y(n17341),
	.A(n17340),
	.B(n17339));
   NOR3xp33_ASAP7_75t_SL U15067 (.Y(n16590),
	.A(n24742),
	.B(n23995),
	.C(n17186));
   NOR3xp33_ASAP7_75t_SRAM U15068 (.Y(n21494),
	.A(n21466),
	.B(n21465),
	.C(n21464));
   NAND2xp5_ASAP7_75t_SL U15069 (.Y(n19078),
	.A(n18378),
	.B(n18377));
   NAND2xp33_ASAP7_75t_L U15070 (.Y(n13983),
	.A(n13979),
	.B(n13980));
   NAND2xp33_ASAP7_75t_L U15071 (.Y(n13982),
	.A(n13981),
	.B(n13980));
   AND3x1_ASAP7_75t_L U15072 (.Y(n23873),
	.A(n23872),
	.B(n23871),
	.C(n23870));
   NAND2x1_ASAP7_75t_SL U15074 (.Y(n22859),
	.A(n18207),
	.B(n20772));
   NAND2xp5_ASAP7_75t_L U15075 (.Y(n19852),
	.A(FE_OCPN27908_FE_OFN16156_sa00_2),
	.B(n19851));
   NAND2xp5_ASAP7_75t_SL U15076 (.Y(n18021),
	.A(n19485),
	.B(n18900));
   NAND2xp33_ASAP7_75t_SL U15077 (.Y(n22028),
	.A(FE_OFN28581_n23491),
	.B(n22025));
   NOR3xp33_ASAP7_75t_L U15078 (.Y(n18422),
	.A(n23534),
	.B(n18421),
	.C(n18420));
   NOR3xp33_ASAP7_75t_SL U15079 (.Y(n16364),
	.A(n20893),
	.B(n16361),
	.C(n16360));
   NAND2xp5_ASAP7_75t_L U15080 (.Y(n19270),
	.A(n19268),
	.B(n19267));
   NOR3x1_ASAP7_75t_L U15081 (.Y(n17423),
	.A(n16938),
	.B(n16937),
	.C(n16936));
   NAND2xp33_ASAP7_75t_SL U15082 (.Y(n16862),
	.A(n16861),
	.B(FE_OFN79_n16857));
   NAND3x1_ASAP7_75t_SL U15083 (.Y(n19203),
	.A(n19202),
	.B(n19201),
	.C(n23397));
   OA21x2_ASAP7_75t_L U15084 (.Y(n14153),
	.A1(FE_OFN28898_n13805),
	.A2(n14150),
	.B(n14149));
   NAND2xp33_ASAP7_75t_SL U15085 (.Y(n16863),
	.A(n16858),
	.B(FE_OFN79_n16857));
   NAND3xp33_ASAP7_75t_SL U15086 (.Y(n19990),
	.A(n19989),
	.B(n20323),
	.C(n19988));
   NAND2xp33_ASAP7_75t_L U15087 (.Y(n19999),
	.A(n19998),
	.B(n19997));
   NAND2xp5_ASAP7_75t_L U15088 (.Y(n15230),
	.A(n15229),
	.B(n15228));
   NAND2xp33_ASAP7_75t_L U15089 (.Y(n15644),
	.A(n15643),
	.B(n15642));
   NAND2xp33_ASAP7_75t_L U15090 (.Y(n20000),
	.A(n19996),
	.B(n19997));
   NAND2xp33_ASAP7_75t_R U15091 (.Y(n14554),
	.A(n14553),
	.B(n14552));
   AND2x2_ASAP7_75t_SRAM U15092 (.Y(n19213),
	.A(n19212),
	.B(n19211));
   NAND2xp5_ASAP7_75t_L U15093 (.Y(n17868),
	.A(n17867),
	.B(n17866));
   NAND2xp33_ASAP7_75t_L U15094 (.Y(n14555),
	.A(n14549),
	.B(n14552));
   NOR2xp33_ASAP7_75t_R U15095 (.Y(n13979),
	.A(n14928),
	.B(n14951));
   NAND2xp33_ASAP7_75t_L U15096 (.Y(n15645),
	.A(n15634),
	.B(n15633));
   NOR3xp33_ASAP7_75t_SL U15097 (.Y(n20564),
	.A(n20563),
	.B(n22239),
	.C(n20562));
   OR3x1_ASAP7_75t_L U15098 (.Y(n15590),
	.A(n13726),
	.B(FE_OFN28662_w3_7),
	.C(n15589));
   NAND2xp5_ASAP7_75t_L U15099 (.Y(n14149),
	.A(n14148),
	.B(n14147));
   NOR3xp33_ASAP7_75t_L U15100 (.Y(n14637),
	.A(n14633),
	.B(n14632),
	.C(n14631));
   NAND2xp5_ASAP7_75t_L U15101 (.Y(n16699),
	.A(n16697),
	.B(n16696));
   NOR2xp33_ASAP7_75t_L U15102 (.Y(n14432),
	.A(n14430),
	.B(n14429));
   NOR2xp33_ASAP7_75t_L U15103 (.Y(n14428),
	.A(n15128),
	.B(n14429));
   NAND2xp5_ASAP7_75t_L U15104 (.Y(n14295),
	.A(n14294),
	.B(n14293));
   NAND3xp33_ASAP7_75t_SL U15105 (.Y(n17457),
	.A(n21393),
	.B(n17508),
	.C(n19204));
   NOR3x1_ASAP7_75t_L U15106 (.Y(n16722),
	.A(n16721),
	.B(n18415),
	.C(n16720));
   NAND2xp5_ASAP7_75t_R U15108 (.Y(n18780),
	.A(n18779),
	.B(n18778));
   NAND2xp5_ASAP7_75t_L U15109 (.Y(n18928),
	.A(n18925),
	.B(n18924));
   NAND2xp5_ASAP7_75t_L U15110 (.Y(n18377),
	.A(n18376),
	.B(n18375));
   NAND2xp5_ASAP7_75t_SL U15111 (.Y(n18378),
	.A(n18374),
	.B(n18375));
   NOR3xp33_ASAP7_75t_SL U15112 (.Y(n19082),
	.A(n18507),
	.B(n18506),
	.C(n22122));
   OR3x1_ASAP7_75t_L U15113 (.Y(n17477),
	.A(n17476),
	.B(FE_OFN114_n22512),
	.C(n21822));
   AND2x2_ASAP7_75t_SRAM U15114 (.Y(n23954),
	.A(n23953),
	.B(n23952));
   NAND2x1p5_ASAP7_75t_SL U15115 (.Y(n25064),
	.A(n20364),
	.B(n20363));
   NAND2xp5_ASAP7_75t_L U15116 (.Y(n21570),
	.A(n21559),
	.B(n21558));
   NAND2xp5_ASAP7_75t_L U15117 (.Y(n18702),
	.A(n18701),
	.B(n18700));
   NAND2xp5_ASAP7_75t_L U15118 (.Y(n18703),
	.A(n18699),
	.B(n18700));
   OAI21xp33_ASAP7_75t_R U15120 (.Y(n22437),
	.A1(FE_OCPN29320_n22461),
	.A2(FE_OCPN27399_n22598),
	.B(n26453));
   NAND2xp33_ASAP7_75t_SL U15121 (.Y(n17866),
	.A(n17865),
	.B(n22697));
   NAND2xp5_ASAP7_75t_SL U15122 (.Y(n18741),
	.A(n19601),
	.B(n18740));
   NAND2xp33_ASAP7_75t_SL U15123 (.Y(n17867),
	.A(n17864),
	.B(n22697));
   AND2x2_ASAP7_75t_L U15124 (.Y(n23729),
	.A(n23728),
	.B(n23727));
   NAND2xp33_ASAP7_75t_SL U15125 (.Y(n19989),
	.A(n19987),
	.B(n19986));
   NOR2xp33_ASAP7_75t_SL U15126 (.Y(n16772),
	.A(n22679),
	.B(n25581));
   AND2x2_ASAP7_75t_R U15127 (.Y(n19520),
	.A(n19519),
	.B(n19518));
   NOR2xp33_ASAP7_75t_SRAM U15128 (.Y(n17937),
	.A(n22752),
	.B(n17936));
   OR3x1_ASAP7_75t_L U15129 (.Y(n20748),
	.A(FE_OCPN5182_n21090),
	.B(n21130),
	.C(n20746));
   NAND2xp5_ASAP7_75t_SL U15131 (.Y(n24894),
	.A(n16598),
	.B(n23950));
   NOR2xp67_ASAP7_75t_L U15132 (.Y(n18887),
	.A(n17989),
	.B(n21043));
   NAND2xp5_ASAP7_75t_L U15133 (.Y(n18959),
	.A(n18958),
	.B(n18957));
   OR3x1_ASAP7_75t_SL U15135 (.Y(n18902),
	.A(n18901),
	.B(n21504),
	.C(n21751));
   NOR2xp33_ASAP7_75t_SRAM U15137 (.Y(n21777),
	.A(n21771),
	.B(n23309));
   NAND2xp33_ASAP7_75t_SL U15138 (.Y(n20621),
	.A(n20620),
	.B(n20619));
   NOR2x1_ASAP7_75t_L U15139 (.Y(n21168),
	.A(n19090),
	.B(n18638));
   NAND2xp5_ASAP7_75t_L U15140 (.Y(n20622),
	.A(n20618),
	.B(n20619));
   NAND2x1_ASAP7_75t_L U15141 (.Y(n19181),
	.A(n19177),
	.B(n19178));
   NAND2xp5_ASAP7_75t_SL U15142 (.Y(n17014),
	.A(n17013),
	.B(n17012));
   NAND3xp33_ASAP7_75t_SL U15143 (.Y(n19404),
	.A(FE_OCPN29568_n18257),
	.B(n25872),
	.C(n16990));
   AND3x4_ASAP7_75t_SL U15144 (.Y(n17155),
	.A(n17152),
	.B(n20505),
	.C(n19386));
   NOR3xp33_ASAP7_75t_L U15145 (.Y(n16324),
	.A(n16323),
	.B(n20833),
	.C(n21929));
   NAND2xp33_ASAP7_75t_SRAM U15146 (.Y(n18958),
	.A(n18953),
	.B(n18955));
   NAND2xp33_ASAP7_75t_SRAM U15147 (.Y(n18957),
	.A(n18956),
	.B(n18955));
   OAI21x1_ASAP7_75t_SL U15148 (.Y(n23309),
	.A1(n18178),
	.A2(n23160),
	.B(n21120));
   NAND2xp33_ASAP7_75t_SRAM U15149 (.Y(n17503),
	.A(n23250),
	.B(n19210));
   NOR2x1_ASAP7_75t_SL U15150 (.Y(n23397),
	.A(n19200),
	.B(n19199));
   NOR3xp33_ASAP7_75t_SL U15151 (.Y(n17509),
	.A(n23366),
	.B(n23247),
	.C(n21837));
   NAND3xp33_ASAP7_75t_SL U15153 (.Y(n16721),
	.A(n16945),
	.B(n18446),
	.C(n16719));
   NAND2xp5_ASAP7_75t_R U15154 (.Y(n19333),
	.A(n19332),
	.B(n22986));
   NAND2xp5_ASAP7_75t_SL U15155 (.Y(n21465),
	.A(n17255),
	.B(n21468));
   AND3x1_ASAP7_75t_SRAM U15156 (.Y(n22485),
	.A(n26064),
	.B(n23254),
	.C(n22484));
   OAI21xp5_ASAP7_75t_SL U15157 (.Y(n21125),
	.A1(FE_PSN8294_n22310),
	.A2(n21770),
	.B(n21124));
   NAND3xp33_ASAP7_75t_SL U15158 (.Y(n18457),
	.A(n26025),
	.B(n18498),
	.C(n18455));
   NAND2xp33_ASAP7_75t_R U15159 (.Y(n18112),
	.A(n18111),
	.B(n18110));
   NAND2xp5_ASAP7_75t_SL U15160 (.Y(n19385),
	.A(FE_OFN29173_n),
	.B(n17078));
   AND2x2_ASAP7_75t_R U15161 (.Y(n15247),
	.A(n15243),
	.B(n15242));
   OA21x2_ASAP7_75t_SRAM U15162 (.Y(n20226),
	.A1(n22010),
	.A2(FE_OCPN27288_n25091),
	.B(n20225));
   NOR3x1_ASAP7_75t_SL U15163 (.Y(n16589),
	.A(n23043),
	.B(n23141),
	.C(n23044));
   AND2x2_ASAP7_75t_SRAM U15164 (.Y(n23458),
	.A(n23457),
	.B(n23456));
   OR2x2_ASAP7_75t_SRAM U15165 (.Y(n18200),
	.A(n18199),
	.B(n23161));
   OA21x2_ASAP7_75t_SRAM U15167 (.Y(n18167),
	.A1(n23303),
	.A2(n18166),
	.B(n21124));
   NAND2xp5_ASAP7_75t_R U15168 (.Y(n19018),
	.A(n19015),
	.B(n19016));
   OA21x2_ASAP7_75t_SRAM U15169 (.Y(n22851),
	.A1(n18162),
	.A2(FE_OFN29195_n22850),
	.B(FE_OCPN27979_FE_OFN16147_sa22_1));
   AND3x1_ASAP7_75t_SL U15170 (.Y(n19010),
	.A(n22046),
	.B(n23476),
	.C(n19009));
   NOR3xp33_ASAP7_75t_SL U15171 (.Y(n20960),
	.A(n19258),
	.B(n22881),
	.C(n22539));
   NAND2xp33_ASAP7_75t_SRAM U15172 (.Y(n18444),
	.A(n18442),
	.B(n18441));
   NAND2xp5_ASAP7_75t_L U15173 (.Y(n19987),
	.A(n19984),
	.B(n19983));
   NOR3xp33_ASAP7_75t_SRAM U15174 (.Y(n16363),
	.A(n18084),
	.B(n16496),
	.C(n16362));
   OR3x1_ASAP7_75t_SRAM U15175 (.Y(n18066),
	.A(n18065),
	.B(n18071),
	.C(n20068));
   AND3x1_ASAP7_75t_L U15176 (.Y(n17775),
	.A(n20204),
	.B(n22891),
	.C(n17774));
   OA222x2_ASAP7_75t_SRAM U15177 (.Y(n13287),
	.A1(n13596),
	.A2(n13286),
	.B1(n15255),
	.B2(n13286),
	.C1(FE_OFN16437_n),
	.C2(n13286));
   OA21x2_ASAP7_75t_R U15178 (.Y(n15284),
	.A1(n15283),
	.A2(n14289),
	.B(n15282));
   AND2x2_ASAP7_75t_SRAM U15179 (.Y(n19628),
	.A(n19627),
	.B(FE_OFN28596_n23948));
   AND2x2_ASAP7_75t_R U15180 (.Y(n15037),
	.A(n15108),
	.B(n15036));
   OA21x2_ASAP7_75t_L U15181 (.Y(n15849),
	.A1(n15639),
	.A2(n15847),
	.B(n15846));
   NAND2xp5_ASAP7_75t_SL U15182 (.Y(n17854),
	.A(n16807),
	.B(n22343));
   OA21x2_ASAP7_75t_SRAM U15183 (.Y(n15515),
	.A1(FE_OFN16352_n14289),
	.A2(n15714),
	.B(n15513));
   OA21x2_ASAP7_75t_L U15184 (.Y(n20963),
	.A1(FE_OCPN7645_n20962),
	.A2(FE_OCPN29545_n22529),
	.B(n22110));
   NAND2xp33_ASAP7_75t_SRAM U15185 (.Y(n13761),
	.A(n13759),
	.B(n13758));
   OA21x2_ASAP7_75t_SRAM U15186 (.Y(n20566),
	.A1(n23217),
	.A2(n23215),
	.B(n24056));
   NOR2x1_ASAP7_75t_SL U15188 (.Y(n16895),
	.A(n17407),
	.B(n16449));
   NAND3xp33_ASAP7_75t_R U15189 (.Y(n14625),
	.A(n14624),
	.B(n15431),
	.C(n14623));
   OA21x2_ASAP7_75t_R U15190 (.Y(n14454),
	.A1(n15567),
	.A2(n15808),
	.B(n14450));
   OA21x2_ASAP7_75t_L U15191 (.Y(n14616),
	.A1(n15447),
	.A2(FE_OCPN29570_n15423),
	.B(n14612));
   NAND2x1_ASAP7_75t_L U15192 (.Y(n19647),
	.A(n24955),
	.B(n19787));
   OA21x2_ASAP7_75t_SRAM U15193 (.Y(n23630),
	.A1(FE_OFN16267_sa21_4),
	.A2(n23628),
	.B(n23627));
   NOR2xp33_ASAP7_75t_L U15194 (.Y(n16654),
	.A(n23131),
	.B(n16653));
   OAI21xp5_ASAP7_75t_SL U15195 (.Y(n23385),
	.A1(FE_OCPN27229_sa11_2),
	.A2(FE_OCPN27848_n23255),
	.B(n19164));
   NAND2x1_ASAP7_75t_SL U15196 (.Y(n17201),
	.A(n19787),
	.B(n16542));
   OA21x2_ASAP7_75t_R U15199 (.Y(n18579),
	.A1(n23677),
	.A2(FE_OFN28815_n18523),
	.B(n21665));
   NAND2xp5_ASAP7_75t_SL U15200 (.Y(n13359),
	.A(n15182),
	.B(FE_OFN27207_w3_30));
   NOR2x1p5_ASAP7_75t_SL U15201 (.Y(n17297),
	.A(n19097),
	.B(n17275));
   OR3x1_ASAP7_75t_SRAM U15205 (.Y(n14750),
	.A(n14749),
	.B(FE_OFN28977_n),
	.C(FE_OFN28683_w3_21));
   AND2x2_ASAP7_75t_SRAM U15206 (.Y(n23280),
	.A(n23279),
	.B(n23278));
   NAND2x1_ASAP7_75t_SL U15207 (.Y(n19775),
	.A(FE_OFN28749_n),
	.B(n16551));
   NOR2xp33_ASAP7_75t_SRAM U15208 (.Y(n19734),
	.A(n17529),
	.B(n19732));
   AND3x1_ASAP7_75t_SL U15209 (.Y(n17874),
	.A(n25350),
	.B(n19973),
	.C(n17873));
   NAND2x1p5_ASAP7_75t_L U15210 (.Y(n24567),
	.A(FE_OFN29171_n17510),
	.B(FE_OFN29061_n22505));
   OA21x2_ASAP7_75t_SRAM U15211 (.Y(n13895),
	.A1(n15339),
	.A2(FE_OFN16210_n13876),
	.B(n14351));
   OR2x2_ASAP7_75t_R U15212 (.Y(n21031),
	.A(FE_OCPN27483_FE_OFN16132_sa03_5),
	.B(n23443));
   OA21x2_ASAP7_75t_SRAM U15213 (.Y(n17058),
	.A1(FE_OCPN28204_n20526),
	.A2(n17115),
	.B(n27089));
   AND2x2_ASAP7_75t_L U15214 (.Y(n18215),
	.A(n18214),
	.B(n18213));
   AND2x2_ASAP7_75t_R U15215 (.Y(n14017),
	.A(n14016),
	.B(FE_OFN28600_n14289));
   NAND2xp5_ASAP7_75t_SL U15216 (.Y(n16998),
	.A(n25988),
	.B(n17077));
   OA21x2_ASAP7_75t_SRAM U15217 (.Y(n13835),
	.A1(n15402),
	.A2(FE_OFN29018_n15921),
	.B(n13834));
   OA21x2_ASAP7_75t_SRAM U15218 (.Y(n23952),
	.A1(FE_OFN130_sa10_5),
	.A2(n23951),
	.B(n23950));
   OA21x2_ASAP7_75t_R U15219 (.Y(n13967),
	.A1(n15455),
	.A2(n15445),
	.B(n13966));
   OR2x2_ASAP7_75t_SRAM U15220 (.Y(n18848),
	.A(n18847),
	.B(n18846));
   OA21x2_ASAP7_75t_L U15221 (.Y(n14643),
	.A1(n15958),
	.A2(n14642),
	.B(n14641));
   OA21x2_ASAP7_75t_R U15222 (.Y(n13828),
	.A1(n14915),
	.A2(FE_OFN112_n15994),
	.B(n13827));
   OA21x2_ASAP7_75t_SRAM U15223 (.Y(n16675),
	.A1(n16429),
	.A2(n16947),
	.B(n16724));
   NAND2xp5_ASAP7_75t_L U15224 (.Y(n13977),
	.A(n14906),
	.B(n14112));
   OR2x2_ASAP7_75t_SRAM U15225 (.Y(n22482),
	.A(n17473),
	.B(n23374));
   OR2x2_ASAP7_75t_SRAM U15227 (.Y(n22492),
	.A(FE_OCPN28038_n23252),
	.B(n23375));
   NAND2xp33_ASAP7_75t_SL U15228 (.Y(n14148),
	.A(n14144),
	.B(n14145));
   OR2x2_ASAP7_75t_R U15229 (.Y(n20231),
	.A(FE_OCPN29480_n20913),
	.B(n20928));
   OA21x2_ASAP7_75t_SRAM U15230 (.Y(n19038),
	.A1(FE_OFN28901_sa30_4),
	.A2(n19037),
	.B(n17618));
   NAND2x1_ASAP7_75t_L U15231 (.Y(n18721),
	.A(FE_OCPN29408_n22461),
	.B(n17321));
   INVx1_ASAP7_75t_L U15232 (.Y(n19016),
	.A(n20260));
   OA21x2_ASAP7_75t_SL U15234 (.Y(n13660),
	.A1(n14593),
	.A2(n13658),
	.B(n15156));
   OA21x2_ASAP7_75t_SRAM U15235 (.Y(n13426),
	.A1(FE_OFN25966_n13646),
	.A2(n13649),
	.B(n13692));
   OR2x2_ASAP7_75t_R U15236 (.Y(n17369),
	.A(FE_OCPN29320_n22461),
	.B(FE_OFN25878_n17329));
   OA21x2_ASAP7_75t_SRAM U15237 (.Y(n20914),
	.A1(n20920),
	.A2(n20913),
	.B(n25713));
   OA21x2_ASAP7_75t_R U15238 (.Y(n19337),
	.A1(n19019),
	.A2(n20251),
	.B(FE_OFN27078_sa23_5));
   NAND2x1p5_ASAP7_75t_SL U15239 (.Y(n23372),
	.A(n17446),
	.B(n21365));
   OA21x2_ASAP7_75t_L U15240 (.Y(n19174),
	.A1(FE_OCPN28447_n23392),
	.A2(FE_OCPN29378_n23266),
	.B(n19173));
   INVxp33_ASAP7_75t_L U15241 (.Y(n18502),
	.A(n25083));
   OA21x2_ASAP7_75t_SRAM U15242 (.Y(n20472),
	.A1(FE_OCPN27428_n26027),
	.A2(n20471),
	.B(FE_OFN28513_n20470));
   OA21x2_ASAP7_75t_L U15243 (.Y(n19983),
	.A1(n19982),
	.A2(n16762),
	.B(n19981));
   NAND2x1_ASAP7_75t_L U15245 (.Y(n16406),
	.A(n16303),
	.B(n21989));
   NAND2xp5_ASAP7_75t_SL U15246 (.Y(n21936),
	.A(n16299),
	.B(n16348));
   NAND2xp5_ASAP7_75t_R U15247 (.Y(n15693),
	.A(n15528),
	.B(n14276));
   OA21x2_ASAP7_75t_L U15249 (.Y(n22819),
	.A1(n23303),
	.A2(n18166),
	.B(FE_OFN28939_n21129));
   NOR2xp33_ASAP7_75t_SL U15251 (.Y(n14837),
	.A(FE_OFN28792_n15787),
	.B(n15851));
   OR2x2_ASAP7_75t_SRAM U15252 (.Y(n14857),
	.A(FE_OFN26084_n15106),
	.B(n15817));
   NAND2xp33_ASAP7_75t_SRAM U15253 (.Y(n13759),
	.A(n15028),
	.B(n13757));
   OR2x2_ASAP7_75t_SRAM U15254 (.Y(n13908),
	.A(n15534),
	.B(n14315));
   NAND2xp5_ASAP7_75t_L U15255 (.Y(n16588),
	.A(n19630),
	.B(n16597));
   NAND2xp5_ASAP7_75t_L U15256 (.Y(n20795),
	.A(n22745),
	.B(n22742));
   OA21x2_ASAP7_75t_SRAM U15257 (.Y(n14977),
	.A1(FE_OFN28695_n),
	.A2(n14986),
	.B(n13771));
   INVx3_ASAP7_75t_SL U15258 (.Y(n19787),
	.A(n16564));
   NOR3x1_ASAP7_75t_SL U15259 (.Y(n21677),
	.A(n20623),
	.B(FE_OCPN27532_n21643),
	.C(n21642));
   NOR2xp33_ASAP7_75t_L U15260 (.Y(n18333),
	.A(n17679),
	.B(n19721));
   NOR2xp33_ASAP7_75t_L U15261 (.Y(n18073),
	.A(FE_OCPN29482_FE_OFN26014_sa31_3),
	.B(n16296));
   OAI22xp33_ASAP7_75t_SRAM U15263 (.Y(n20331),
	.A1(FE_OCPN28298_n),
	.A2(n20325),
	.B1(FE_OCPN27690_n16757),
	.B2(n20325));
   NOR2x1p5_ASAP7_75t_L U15265 (.Y(n17444),
	.A(FE_OCPN27365_sa11_4),
	.B(n23393));
   NOR3xp33_ASAP7_75t_SL U15266 (.Y(n20583),
	.A(n17916),
	.B(FE_OCPN29477_sa12_5),
	.C(n19527));
   NAND2x1p5_ASAP7_75t_SL U15268 (.Y(n15808),
	.A(n15857),
	.B(FE_OFN25900_w3_4));
   NAND2x1p5_ASAP7_75t_SL U15269 (.Y(n18011),
	.A(FE_OCPN29349_FE_OCPN27405_sa03_4),
	.B(n21318));
   OAI21xp5_ASAP7_75t_SL U15270 (.Y(n13288),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OCPN27656_w3_25),
	.B(n15183));
   NAND2x1_ASAP7_75t_SL U15272 (.Y(n20561),
	.A(n17898),
	.B(n22745));
   NAND2xp33_ASAP7_75t_SRAM U15274 (.Y(n22555),
	.A(n17757),
	.B(n17761));
   NOR2xp33_ASAP7_75t_SL U15275 (.Y(n16306),
	.A(FE_OFN29117_n),
	.B(n16408));
   OR2x2_ASAP7_75t_SRAM U15276 (.Y(n15988),
	.A(FE_OFN26007_n16010),
	.B(n15987));
   NAND2x1p5_ASAP7_75t_SL U15277 (.Y(n16874),
	.A(FE_OCPN29487_FE_OFN28694_sa33_4),
	.B(n16909));
   NAND2xp5_ASAP7_75t_SL U15278 (.Y(n24866),
	.A(n17529),
	.B(n17546));
   OR3x1_ASAP7_75t_SRAM U15279 (.Y(n20727),
	.A(FE_OFN26133_sa22_3),
	.B(FE_OFN28680_n),
	.C(n20753));
   NOR2xp33_ASAP7_75t_SRAM U15280 (.Y(n14100),
	.A(FE_OFN27115_n),
	.B(FE_OFN109_n15994));
   NAND2x1p5_ASAP7_75t_SL U15281 (.Y(n16429),
	.A(n16689),
	.B(FE_OCPN27568_sa33_3));
   NAND2xp5_ASAP7_75t_L U15282 (.Y(n17042),
	.A(n16988),
	.B(FE_OFN28479_sa13_2));
   NOR2x1p5_ASAP7_75t_SL U15283 (.Y(n16542),
	.A(FE_OCPN27636_sa10_4),
	.B(n16594));
   NAND2x1p5_ASAP7_75t_SL U15284 (.Y(n16610),
	.A(FE_OCPN27636_sa10_4),
	.B(n16547));
   INVx3_ASAP7_75t_SL U15285 (.Y(n16648),
	.A(n17223));
   OR2x2_ASAP7_75t_SRAM U15286 (.Y(n15086),
	.A(n15601),
	.B(FE_OFN26084_n15106));
   NAND2x1p5_ASAP7_75t_SL U15287 (.Y(n16436),
	.A(FE_OFN28727_sa33_1),
	.B(n16831));
   OA21x2_ASAP7_75t_SRAM U15288 (.Y(n13437),
	.A1(FE_OFN27207_w3_30),
	.A2(n15183),
	.B(n15224));
   NAND2x1p5_ASAP7_75t_SL U15289 (.Y(n22461),
	.A(n18707),
	.B(FE_OCPN27810_n));
   NOR2x1_ASAP7_75t_L U15291 (.Y(n23996),
	.A(n16594),
	.B(n19789));
   NAND2x1_ASAP7_75t_SL U15293 (.Y(n13730),
	.A(FE_OFN29052_w3_5),
	.B(FE_OFN25900_w3_4));
   NAND2xp5_ASAP7_75t_L U15295 (.Y(n25585),
	.A(sa21_6_),
	.B(FE_OFN167_sa21_7));
   NAND2xp5_ASAP7_75t_L U15296 (.Y(n26777),
	.A(sa00_7_),
	.B(n17305));
   NAND2xp5_ASAP7_75t_L U15297 (.Y(n13689),
	.A(w3_24_),
	.B(n24470));
   INVx1_ASAP7_75t_R U15298 (.Y(n15271),
	.A(n14585));
   INVx1_ASAP7_75t_SL U15299 (.Y(n15156),
	.A(n13551));
   NAND2x1p5_ASAP7_75t_R U15301 (.Y(n17584),
	.A(n17732),
	.B(n25034));
   NAND2x1_ASAP7_75t_L U15302 (.Y(n26315),
	.A(FE_OFN16197_sa31_6),
	.B(n16344));
   NOR2xp67_ASAP7_75t_L U15303 (.Y(n17580),
	.A(n17732),
	.B(n25034));
   NOR2x1p5_ASAP7_75t_SL U15304 (.Y(n24181),
	.A(FE_OFN26629_sa31_4),
	.B(FE_OFN26107_sa31_5));
   NOR2x1_ASAP7_75t_L U15305 (.Y(n26829),
	.A(sa21_6_),
	.B(FE_OFN167_sa21_7));
   NAND2xp5_ASAP7_75t_L U15306 (.Y(n26889),
	.A(sa22_6_),
	.B(n22300));
   NAND2xp5_ASAP7_75t_L U15307 (.Y(n26346),
	.A(FE_OFN25946_sa32_6),
	.B(FE_OFN25997_n));
   NAND2x1p5_ASAP7_75t_SL U15308 (.Y(n21355),
	.A(n19170),
	.B(n17451));
   NAND2x1_ASAP7_75t_R U15309 (.Y(n17463),
	.A(FE_OFN150_sa11_7),
	.B(n21340));
   NAND2xp5_ASAP7_75t_L U15310 (.Y(n15704),
	.A(FE_OFN28701_w3_16),
	.B(n23974));
   NAND2xp5_ASAP7_75t_R U15311 (.Y(n26571),
	.A(FE_OFN45_sa23_6),
	.B(FE_OFN162_sa23_7));
   NOR2x1_ASAP7_75t_L U15312 (.Y(n17452),
	.A(n19170),
	.B(FE_OFN26005_n17451));
   NAND2x1p5_ASAP7_75t_L U15313 (.Y(n15694),
	.A(FE_OFN27096_n),
	.B(FE_PSN8292_FE_OFN26041_w3_17));
   NAND2x1p5_ASAP7_75t_SL U15315 (.Y(n19509),
	.A(FE_OCPN29453_sa12_4),
	.B(FE_OFN28676_sa12_5));
   NAND2xp33_ASAP7_75t_SRAM U15317 (.Y(n16235),
	.A(FE_OFN28713_n),
	.B(FE_OFN26_n16125));
   NOR2x1_ASAP7_75t_L U15318 (.Y(n26857),
	.A(sa10_6_),
	.B(n16563));
   NAND2xp33_ASAP7_75t_SRAM U15319 (.Y(n16212),
	.A(FE_OFN25_n16125),
	.B(FE_OFN16459_n));
   NAND2xp5_ASAP7_75t_L U15320 (.Y(n24800),
	.A(sa30_6_),
	.B(n19060));
   NAND2xp5_ASAP7_75t_R U15321 (.Y(n25420),
	.A(sa03_6_),
	.B(FE_OFN118_sa03_7));
   NAND2xp5_ASAP7_75t_L U15322 (.Y(n26687),
	.A(FE_OFN28480_sa30_7),
	.B(n17629));
   NAND2x1p5_ASAP7_75t_SL U15323 (.Y(n19502),
	.A(n22721),
	.B(n22776));
   NAND2xp33_ASAP7_75t_L U15324 (.Y(n25641),
	.A(sa20_7_),
	.B(n24154));
   NAND2xp33_ASAP7_75t_L U15325 (.Y(n27027),
	.A(sa23_7_),
	.B(n26562));
   NAND2x1p5_ASAP7_75t_R U15326 (.Y(n15238),
	.A(FE_OFN16412_w3_26),
	.B(FE_OFN16159_w3_24));
   NOR2xp33_ASAP7_75t_L U15327 (.Y(n27207),
	.A(sa20_7_),
	.B(n24154));
   NAND2xp33_ASAP7_75t_L U15329 (.Y(n24978),
	.A(sa10_6_),
	.B(n16563));
   NAND2xp5_ASAP7_75t_L U15330 (.Y(n27095),
	.A(n19359),
	.B(FE_OFN127_sa13_7));
   NOR2xp67_ASAP7_75t_L U15331 (.Y(n27183),
	.A(sa02_7_),
	.B(n17815));
   NOR2x1_ASAP7_75t_L U15332 (.Y(n26139),
	.A(FE_OFN165_sa12_7),
	.B(n17915));
   NAND2x1_ASAP7_75t_SL U15333 (.Y(n15183),
	.A(n25675),
	.B(w3_25_));
   AND2x2_ASAP7_75t_SRAM U15334 (.Y(n13007),
	.A(n16281),
	.B(n13006));
   NAND2x1_ASAP7_75t_R U15335 (.Y(n26542),
	.A(FE_OFN90_sa33_7),
	.B(FE_OFN174_sa33_6));
   NOR2x1_ASAP7_75t_L U15336 (.Y(n26942),
	.A(FE_OFN16197_sa31_6),
	.B(n16344));
   INVxp67_ASAP7_75t_SRAM U15337 (.Y(n25247),
	.A(w2_14_));
   NAND2xp33_ASAP7_75t_L U15339 (.Y(n15881),
	.A(w3_0_),
	.B(w3_2_));
   NAND2xp5_ASAP7_75t_R U15340 (.Y(n13901),
	.A(FE_OFN28701_w3_16),
	.B(FE_OFN50_w3_18));
   NOR2x1p5_ASAP7_75t_L U15342 (.Y(n13867),
	.A(FE_OFN28701_w3_16),
	.B(FE_OFN50_w3_18));
   INVx1_ASAP7_75t_R U15343 (.Y(n25051),
	.A(w3_10_));
   NOR2xp33_ASAP7_75t_SL U15345 (.Y(n13551),
	.A(FE_OFN27210_w3_30),
	.B(FE_OCPN27656_w3_25));
   NAND2x1_ASAP7_75t_L U15346 (.Y(n15423),
	.A(FE_OCPN28402_w3_13),
	.B(n24755));
   NOR2xp67_ASAP7_75t_L U15349 (.Y(n26249),
	.A(sa23_7_),
	.B(sa23_6_));
   NOR3xp33_ASAP7_75t_SL U15350 (.Y(n23359),
	.A(sa11_2_),
	.B(FE_OCPN27242_sa11_1),
	.C(FE_OFN28507_sa11_0));
   NOR2x1p5_ASAP7_75t_R U15351 (.Y(n27216),
	.A(FE_OFN68_sa02_6),
	.B(sa02_7_));
   NAND2x1p5_ASAP7_75t_L U15352 (.Y(n27168),
	.A(n16377),
	.B(sa31_7_));
   NOR2x1_ASAP7_75t_L U15353 (.Y(n26282),
	.A(sa01_6_),
	.B(sa01_7_));
   NAND2xp33_ASAP7_75t_SL U15354 (.Y(n26078),
	.A(sa11_6_),
	.B(sa11_7_));
   NOR2x1_ASAP7_75t_L U15355 (.Y(n27127),
	.A(FE_OFN28499_sa00_6),
	.B(sa00_7_));
   NOR2x1p5_ASAP7_75t_L U15356 (.Y(n26915),
	.A(FE_OFN128_sa13_7),
	.B(n19359));
   NOR2x1p5_ASAP7_75t_SL U15357 (.Y(n20739),
	.A(FE_OFN16135_sa22_4),
	.B(FE_OFN26136_sa22_3));
   NAND2x1p5_ASAP7_75t_SL U15358 (.Y(n17065),
	.A(FE_OFN16444_sa13_1),
	.B(FE_OFN28478_sa13_2));
   NOR2x1_ASAP7_75t_L U15359 (.Y(n26819),
	.A(sa03_6_),
	.B(sa03_7_));
   NAND2xp5_ASAP7_75t_L U15360 (.Y(n24331),
	.A(sa33_6_),
	.B(FE_OFN90_sa33_7));
   NAND2xp5_ASAP7_75t_L U15361 (.Y(n26976),
	.A(sa02_6_),
	.B(sa02_7_));
   NAND2xp5_ASAP7_75t_L U15362 (.Y(n23899),
	.A(n17732),
	.B(FE_OFN25946_sa32_6));
   NAND2xp33_ASAP7_75t_L U15363 (.Y(n23945),
	.A(sa03_6_),
	.B(sa03_7_));
   NAND2xp33_ASAP7_75t_L U15367 (.Y(n24263),
	.A(sa21_6_),
	.B(sa21_7_));
   NAND2xp33_ASAP7_75t_L U15368 (.Y(n26517),
	.A(sa20_6_),
	.B(sa20_7_));
   NAND2xp33_ASAP7_75t_L U15369 (.Y(n23345),
	.A(sa22_6_),
	.B(sa22_7_));
   NAND2x1_ASAP7_75t_L U15370 (.Y(n24377),
	.A(FE_OFN175_sa12_6),
	.B(FE_OFN165_sa12_7));
   INVxp67_ASAP7_75t_SRAM U15371 (.Y(n27195),
	.A(w2_23_));
   NOR2x1_ASAP7_75t_L U15373 (.Y(n26584),
	.A(sa30_6_),
	.B(FE_OFN28480_sa30_7));
   NOR2x1_ASAP7_75t_L U15374 (.Y(n22405),
	.A(n17732),
	.B(FE_OFN25946_sa32_6));
   NAND2xp5_ASAP7_75t_L U15375 (.Y(n26926),
	.A(sa30_6_),
	.B(FE_OFN28480_sa30_7));
   INVxp67_ASAP7_75t_SRAM U15376 (.Y(n26416),
	.A(w2_13_));
   A2O1A1Ixp33_ASAP7_75t_L U15377 (.Y(n17772),
	.A1(n20982),
	.A2(n22528),
	.B(n20206),
	.C(FE_OFN28812_FE_OCPN27261_sa02_0));
   A2O1A1Ixp33_ASAP7_75t_R U15378 (.Y(n25302),
	.A1(FE_OFN28595_n20189),
	.A2(n22528),
	.B(n25528),
	.C(n22528));
   A2O1A1Ixp33_ASAP7_75t_SRAM U15379 (.Y(n22530),
	.A1(n22529),
	.A2(n22528),
	.B(FE_OFN27202_n),
	.C(n22528));
   NAND2xp5_ASAP7_75t_L U15380 (.Y(n26792),
	.A(FE_OFN16283_n26788),
	.B(FE_OCPN27435_n26790));
   NAND2xp5_ASAP7_75t_L U15381 (.Y(n25450),
	.A(n27023),
	.B(n25447));
   OAI21xp5_ASAP7_75t_SL U15382 (.Y(n27169),
	.A1(FE_OFN1_ld_r),
	.A2(n27171),
	.B(n27170));
   NOR2x1_ASAP7_75t_SL U15384 (.Y(n27208),
	.A(n25295),
	.B(n25294));
   OAI21x1_ASAP7_75t_L U15385 (.Y(n27197),
	.A1(n27199),
	.A2(n27198),
	.B(FE_OFN16_FE_DBTN0_ld_r));
   INVxp67_ASAP7_75t_SL U15386 (.Y(n24651),
	.A(n24652));
   O2A1O1Ixp33_ASAP7_75t_SL U15388 (.Y(n25431),
	.A1(n25139),
	.A2(FE_OCPN29562_n25138),
	.B(n24981),
	.C(n24980));
   O2A1O1Ixp5_ASAP7_75t_SL U15389 (.Y(n23735),
	.A1(n23734),
	.A2(n23733),
	.B(n26323),
	.C(n23732));
   NOR2x1_ASAP7_75t_L U15390 (.Y(n15290),
	.A(n15341),
	.B(n13890));
   NOR3x1_ASAP7_75t_SL U15391 (.Y(n21017),
	.A(FE_OCPN27675_n17986),
	.B(FE_OCPN27990_FE_OFN16132_sa03_5),
	.C(n18029));
   NOR3x1_ASAP7_75t_SL U15392 (.Y(n26721),
	.A(n21761),
	.B(n21760),
	.C(n21759));
   NAND2xp5_ASAP7_75t_L U15394 (.Y(n16976),
	.A(FE_OFN28979_n),
	.B(n16975));
   OAI21xp5_ASAP7_75t_SL U15395 (.Y(n24685),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27375_n26860),
	.B(n24686));
   NAND2xp5_ASAP7_75t_L U15396 (.Y(n24009),
	.A(FE_OFN16322_n25946),
	.B(n24006));
   OAI21xp5_ASAP7_75t_L U15397 (.Y(n26858),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27375_n26860),
	.B(n26859));
   O2A1O1Ixp33_ASAP7_75t_SRAM U15398 (.Y(n23867),
	.A1(FE_OCPN27896_n18583),
	.A2(n18521),
	.B(n23869),
	.C(n23866));
   NOR3xp33_ASAP7_75t_SL U15400 (.Y(n16447),
	.A(FE_OFN28727_sa33_1),
	.B(FE_OFN29163_sa33_2),
	.C(FE_OFN29134_sa33_0));
   O2A1O1Ixp33_ASAP7_75t_L U15401 (.Y(n26125),
	.A1(FE_OFN16180_n26542),
	.A2(n26127),
	.B(n26124),
	.C(n26130));
   NAND2xp5_ASAP7_75t_L U15402 (.Y(n26940),
	.A(n26936),
	.B(n26935));
   O2A1O1Ixp33_ASAP7_75t_SL U15403 (.Y(n22983),
	.A1(FE_OCPN28381_n26660),
	.A2(n19000),
	.B(FE_OFN16248_n20235),
	.C(n22981));
   O2A1O1Ixp33_ASAP7_75t_SRAM U15404 (.Y(n21095),
	.A1(FE_RN_0_0),
	.A2(n23322),
	.B(FE_OFN28798_FE_OCPN27947_n18177),
	.C(n22281));
   O2A1O1Ixp33_ASAP7_75t_SL U15405 (.Y(n25372),
	.A1(FE_OCPN28100_n25470),
	.A2(n25469),
	.B(n26349),
	.C(n25370));
   O2A1O1Ixp33_ASAP7_75t_L U15406 (.Y(n26353),
	.A1(FE_OCPN27491_n26351),
	.A2(n26350),
	.B(n26349),
	.C(n26348));
   OAI21xp5_ASAP7_75t_SL U15407 (.Y(n26144),
	.A1(FE_OCPN7609_n26145),
	.A2(FE_OCPN29382_n26674),
	.B(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U15408 (.Y(n26788),
	.A1(n26819),
	.A2(n26818),
	.B(n24934),
	.C(n24933));
   NAND2x1_ASAP7_75t_SL U15409 (.Y(n16556),
	.A(FE_OCPN28053_sa10_1),
	.B(FE_OCPN28145_n16535));
   NAND2xp33_ASAP7_75t_L U15410 (.Y(n15269),
	.A(w0_6_),
	.B(n15266));
   A2O1A1Ixp33_ASAP7_75t_SL U15411 (.Y(n26334),
	.A1(n26819),
	.A2(n26725),
	.B(n24746),
	.C(n24745));
   NOR2xp67_ASAP7_75t_SL U15412 (.Y(n23491),
	.A(FE_OCPN27803_sa23_4),
	.B(n22971));
   NOR2x1p5_ASAP7_75t_SL U15414 (.Y(n19000),
	.A(FE_OFN27126_sa23_3),
	.B(n19011));
   OA21x2_ASAP7_75t_R U15415 (.Y(n13684),
	.A1(n14479),
	.A2(n15203),
	.B(n13682));
   NOR3x2_ASAP7_75t_SL U15416 (.Y(n16771),
	.A(FE_OFN28903_sa21_0),
	.B(FE_OCPN27327_sa21_2),
	.C(FE_OCPN29497_sa21_1));
   O2A1O1Ixp5_ASAP7_75t_L U15417 (.Y(n22054),
	.A1(n23522),
	.A2(n22053),
	.B(n26249),
	.C(n22052));
   NOR3x1_ASAP7_75t_SL U15420 (.Y(n22197),
	.A(FE_OFN28718_sa01_1),
	.B(FE_OCPN27423_sa01_0),
	.C(FE_OFN28672_sa01_2));
   OAI22xp5_ASAP7_75t_L U15421 (.Y(n23243),
	.A1(n25682),
	.A2(n25158),
	.B1(n25164),
	.B2(n25158));
   O2A1O1Ixp33_ASAP7_75t_SRAM U15422 (.Y(n16628),
	.A1(n23980),
	.A2(n24959),
	.B(n23148),
	.C(n23043));
   O2A1O1Ixp5_ASAP7_75t_SL U15425 (.Y(n26726),
	.A1(n25139),
	.A2(FE_OCPN29562_n25138),
	.B(n25137),
	.C(n25136));
   O2A1O1Ixp33_ASAP7_75t_L U15426 (.Y(n25136),
	.A1(n25139),
	.A2(n25138),
	.B(FE_OCPN5112_n25135),
	.C(n25134));
   NAND2x1_ASAP7_75t_SL U15427 (.Y(n22329),
	.A(FE_OFN25989_sa21_4),
	.B(FE_OFN28985_sa21_5));
   NAND2xp5_ASAP7_75t_L U15428 (.Y(n24819),
	.A(n24816),
	.B(FE_OFN25939_n26275));
   A2O1A1Ixp33_ASAP7_75t_SL U15429 (.Y(n24275),
	.A1(n17580),
	.A2(n24830),
	.B(FE_OCPN27491_n26351),
	.C(n24450));
   A2O1A1Ixp33_ASAP7_75t_L U15430 (.Y(n27180),
	.A1(n27183),
	.A2(n27182),
	.B(n27177),
	.C(n27178));
   A2O1A1Ixp33_ASAP7_75t_SL U15431 (.Y(n27187),
	.A1(n25234),
	.A2(n25233),
	.B(n26959),
	.C(n25232));
   O2A1O1Ixp33_ASAP7_75t_SRAM U15432 (.Y(n17768),
	.A1(n17763),
	.A2(FE_OFN28665_FE_OCPN27566),
	.B(n17760),
	.C(FE_OFN29184_n17744));
   O2A1O1Ixp33_ASAP7_75t_SL U15433 (.Y(n20965),
	.A1(FE_OFN28704_FE_OCPN27740_sa02_4),
	.A2(FE_OFN28961_n17744),
	.B(n20961),
	.C(FE_OFN28730_FE_OCPN28416_sa02_3));
   NAND2xp5_ASAP7_75t_SL U15434 (.Y(n24427),
	.A(n26134),
	.B(FE_OCPN27806_n25497));
   A2O1A1Ixp33_ASAP7_75t_SL U15435 (.Y(n24426),
	.A1(n26139),
	.A2(n26138),
	.B(n26135),
	.C(n25497));
   NOR2x1p5_ASAP7_75t_SL U15436 (.Y(n21084),
	.A(FE_OFN16135_sa22_4),
	.B(FE_OFN26133_sa22_3));
   OAI21xp33_ASAP7_75t_L U15438 (.Y(n27097),
	.A1(n27096),
	.A2(n27095),
	.B(FE_OCPN8208_n27094));
   OAI21xp5_ASAP7_75t_SL U15439 (.Y(n25294),
	.A1(n27101),
	.A2(n27102),
	.B(n27094));
   OAI22xp33_ASAP7_75t_SL U15440 (.Y(n544),
	.A1(FE_OFN21_n16125),
	.A2(FE_OFN28964_n16273),
	.B1(key_38_),
	.B2(FE_OFN28964_n16273));
   NAND2x1_ASAP7_75t_SL U15441 (.Y(n19275),
	.A(FE_OCPN27261_sa02_0),
	.B(n17799));
   NOR2x1_ASAP7_75t_L U15442 (.Y(n26972),
	.A(FE_OFN28941_sa02_2),
	.B(n22103));
   NAND3xp33_ASAP7_75t_L U15443 (.Y(n22175),
	.A(n17359),
	.B(n17317),
	.C(FE_OCPN29429_FE_OFN16141_sa01_3));
   NOR2xp33_ASAP7_75t_SL U15444 (.Y(n19470),
	.A(n21740),
	.B(n24243));
   NAND3xp33_ASAP7_75t_SL U15445 (.Y(n18774),
	.A(FE_OCPN29302_sa00_4),
	.B(FE_OCPN29260_sa00_5),
	.C(FE_OFN29249_n));
   NAND2xp5_ASAP7_75t_L U15446 (.Y(n18642),
	.A(FE_OCPN29385_n),
	.B(n17252));
   NAND2xp5_ASAP7_75t_SL U15447 (.Y(n20961),
	.A(FE_OFN25998_n17781),
	.B(FE_OCPN8230_n20993));
   NAND2x1p5_ASAP7_75t_L U15448 (.Y(n22069),
	.A(FE_OFN28812_FE_OCPN27261_sa02_0),
	.B(n20129));
   NOR2xp33_ASAP7_75t_L U15449 (.Y(n22077),
	.A(n20186),
	.B(n26972));
   NAND2x1p5_ASAP7_75t_SL U15451 (.Y(n17996),
	.A(FE_OFN29123_n),
	.B(n21327));
   NOR2xp33_ASAP7_75t_R U15452 (.Y(n23134),
	.A(FE_OCPN5015_n23031),
	.B(n19774));
   NOR2x1_ASAP7_75t_SL U15453 (.Y(n17637),
	.A(FE_OFN16247_sa30_1),
	.B(FE_OFN28925_sa30_0));
   NAND2xp5_ASAP7_75t_SL U15454 (.Y(n23249),
	.A(n21366),
	.B(n19162));
   NOR3x1_ASAP7_75t_L U15455 (.Y(n21586),
	.A(n20471),
	.B(FE_OCPN29432_sa30_3),
	.C(FE_OCPN27971_n21627));
   NAND2x1p5_ASAP7_75t_SL U15457 (.Y(n23752),
	.A(FE_OFN29112_FE_OCPN27870_n18527),
	.B(FE_OCPN27606_n23869));
   NAND2xp5_ASAP7_75t_SL U15458 (.Y(n23766),
	.A(FE_OFN29081_n18526),
	.B(FE_OFN16295_n23837));
   NOR3xp33_ASAP7_75t_L U15459 (.Y(n16475),
	.A(n17398),
	.B(n16472),
	.C(n23558));
   NOR2x1_ASAP7_75t_L U15460 (.Y(n16698),
	.A(n24328),
	.B(FE_OCPN27593_n16908));
   NOR2x1_ASAP7_75t_SL U15461 (.Y(n19313),
	.A(FE_OFN27126_sa23_3),
	.B(n18989));
   NOR2xp67_ASAP7_75t_L U15462 (.Y(n23060),
	.A(FE_OFN16141_sa01_3),
	.B(n18719));
   NAND2xp5_ASAP7_75t_R U15463 (.Y(n18719),
	.A(n26456),
	.B(n18671));
   NOR3xp33_ASAP7_75t_L U15464 (.Y(n23573),
	.A(n22223),
	.B(FE_OFN25908_sa12_2),
	.C(FE_OCPN27253_n17923));
   NAND2x1_ASAP7_75t_SL U15465 (.Y(n22336),
	.A(n22665),
	.B(n22354));
   NOR2xp33_ASAP7_75t_L U15466 (.Y(n16503),
	.A(n25319),
	.B(FE_OFN26550_n16331));
   O2A1O1Ixp5_ASAP7_75t_L U15467 (.Y(n24805),
	.A1(n26926),
	.A2(n26995),
	.B(n26992),
	.C(FE_OFN16297_n24803));
   A2O1A1Ixp33_ASAP7_75t_SL U15468 (.Y(n26194),
	.A1(FE_OFN16176_n27207),
	.A2(n26196),
	.B(FE_OCPN27583_n26193),
	.C(n26192));
   OAI21xp5_ASAP7_75t_L U15470 (.Y(n25553),
	.A1(FE_OFN28622_n25870),
	.A2(n25552),
	.B(n26915));
   NAND3xp33_ASAP7_75t_SL U15471 (.Y(n25552),
	.A(n25551),
	.B(n25550),
	.C(n25549));
   NAND2xp33_ASAP7_75t_SL U15472 (.Y(n19929),
	.A(n19928),
	.B(n19927));
   NAND2xp5_ASAP7_75t_L U15473 (.Y(n19930),
	.A(n19925),
	.B(n19927));
   NOR2xp33_ASAP7_75t_SRAM U15474 (.Y(n19928),
	.A(n17525),
	.B(n19926));
   NAND3x2_ASAP7_75t_SL U15475 (.Y(n21725),
	.A(FE_OCPN29349_FE_OCPN27405_sa03_4),
	.B(FE_OFN21730_sa03_3),
	.C(FE_OFN29179_n));
   NAND3xp33_ASAP7_75t_SL U15477 (.Y(n24551),
	.A(n24567),
	.B(n23249),
	.C(n22514));
   INVxp33_ASAP7_75t_L U15478 (.Y(n21340),
	.A(sa11_6_));
   NOR2xp33_ASAP7_75t_SL U15479 (.Y(n22806),
	.A(n23168),
	.B(n18231));
   NOR3xp33_ASAP7_75t_L U15480 (.Y(n22868),
	.A(n22843),
	.B(n22273),
	.C(n22292));
   NOR3xp33_ASAP7_75t_SL U15481 (.Y(n25093),
	.A(n20913),
	.B(FE_OFN27126_sa23_3),
	.C(n19011));
   NAND3xp33_ASAP7_75t_SL U15483 (.Y(n22375),
	.A(n17577),
	.B(n17576),
	.C(n19916));
   OAI21xp33_ASAP7_75t_L U15484 (.Y(n17572),
	.A1(n18828),
	.A2(FE_OFN26577_n),
	.B(n17697));
   NAND3xp33_ASAP7_75t_L U15485 (.Y(n22374),
	.A(n18304),
	.B(n18329),
	.C(n18833));
   NOR2xp33_ASAP7_75t_SL U15486 (.Y(n18304),
	.A(n20095),
	.B(n18303));
   NOR2xp33_ASAP7_75t_L U15488 (.Y(n24920),
	.A(FE_OFN28539_n22336),
	.B(n22335));
   OAI21xp5_ASAP7_75t_R U15489 (.Y(n24502),
	.A1(n24348),
	.A2(n24347),
	.B(n26637));
   NAND3xp33_ASAP7_75t_SRAM U15490 (.Y(n24347),
	.A(n24346),
	.B(n24345),
	.C(n25258));
   INVxp67_ASAP7_75t_SL U15491 (.Y(n24282),
	.A(n24283));
   OAI21xp33_ASAP7_75t_L U15493 (.Y(n24096),
	.A1(FE_OCPN27968_n21154),
	.A2(FE_OCPN29415_n17237),
	.B(n21441));
   NAND2x1p5_ASAP7_75t_L U15494 (.Y(n23819),
	.A(FE_OCPN29380_sa20_1),
	.B(FE_OCPN28223_FE_OFN27219_n18522));
   NAND2x1p5_ASAP7_75t_SL U15495 (.Y(n25092),
	.A(FE_OCPN27881_FE_OFN27126_sa23_3),
	.B(n20256));
   NAND2xp5_ASAP7_75t_L U15496 (.Y(n23215),
	.A(n17953),
	.B(FE_OFN27070_n));
   NOR3x1_ASAP7_75t_R U15498 (.Y(n23603),
	.A(FE_OFN27070_n),
	.B(FE_OFN28764_n17928),
	.C(FE_OFN28476_sa12_0));
   NAND3xp33_ASAP7_75t_L U15499 (.Y(n19425),
	.A(FE_OCPN28212_n16980),
	.B(FE_OCPN28121_n16975),
	.C(FE_OFN28491_sa13_3));
   NOR3x2_ASAP7_75t_SL U15500 (.Y(n19710),
	.A(n18828),
	.B(FE_OCPN29419_FE_OFN16128_sa32_2),
	.C(n17566));
   NAND2x1p5_ASAP7_75t_L U15501 (.Y(n22690),
	.A(FE_OFN27157_n23928),
	.B(FE_OCPN28299_n));
   NAND3xp33_ASAP7_75t_SL U15502 (.Y(n23626),
	.A(FE_OCPN27631_n16774),
	.B(FE_OFN16153_n16747),
	.C(FE_OFN29066_FE_OCPN27328_sa21_2));
   NAND2xp5_ASAP7_75t_SL U15503 (.Y(n23012),
	.A(n19756),
	.B(FE_OCPN28323_FE_OFN16427_sa10_3));
   NOR3x1_ASAP7_75t_SL U15504 (.Y(n15380),
	.A(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(FE_OCPN29536_FE_OFN8_w3_14),
	.C(FE_OCPN28407_FE_OFN16433_w3_11));
   NOR2x1_ASAP7_75t_L U15505 (.Y(n24617),
	.A(n16925),
	.B(FE_OCPN27460_n16913));
   NAND3xp33_ASAP7_75t_L U15506 (.Y(n26899),
	.A(n25637),
	.B(n25636),
	.C(n25635));
   NOR2x1_ASAP7_75t_SL U15508 (.Y(n24565),
	.A(FE_OCPN27866_n),
	.B(n23381));
   NAND2xp5_ASAP7_75t_SL U15509 (.Y(n18091),
	.A(n18075),
	.B(n18074));
   NOR2xp33_ASAP7_75t_SL U15510 (.Y(n18075),
	.A(n18072),
	.B(n18071));
   NOR2xp33_ASAP7_75t_SRAM U15511 (.Y(n18074),
	.A(n20876),
	.B(n18073));
   NAND3xp33_ASAP7_75t_L U15512 (.Y(n23328),
	.A(FE_OFN26528_n23302),
	.B(n18176),
	.C(FE_OCPN27979_FE_OFN16147_sa22_1));
   NAND2xp5_ASAP7_75t_SL U15513 (.Y(n19424),
	.A(n19376),
	.B(FE_OCPN28137_n17170));
   NOR3x1_ASAP7_75t_L U15514 (.Y(n19739),
	.A(n25029),
	.B(FE_OFN27148_sa32_3),
	.C(FE_OCPN29579_n18837));
   NAND2x1_ASAP7_75t_L U15516 (.Y(n16564),
	.A(n16597),
	.B(FE_OFN26039_sa10_2));
   NAND3xp33_ASAP7_75t_L U15518 (.Y(n22183),
	.A(n17359),
	.B(n17329),
	.C(FE_OCPN27423_sa01_0));
   INVx1_ASAP7_75t_SL U15519 (.Y(n22191),
	.A(n20409));
   NOR3xp33_ASAP7_75t_SL U15520 (.Y(n21551),
	.A(n17326),
	.B(FE_OFN16141_sa01_3),
	.C(FE_OCPN28217_sa01_5));
   OAI22xp5_ASAP7_75t_L U15521 (.Y(n18620),
	.A1(FE_OFN16216_n19573),
	.A2(n19818),
	.B1(FE_OCPN28389_n21479),
	.B2(n19818));
   NOR2x1p5_ASAP7_75t_SL U15522 (.Y(n23775),
	.A(n18544),
	.B(FE_OFN28815_n18523));
   NAND2xp33_ASAP7_75t_SRAM U15523 (.Y(n23793),
	.A(n18583),
	.B(FE_OCPN27606_n23869));
   NOR2x1_ASAP7_75t_L U15524 (.Y(n23496),
	.A(n22010),
	.B(FE_OFN25889_n20913));
   NOR2xp33_ASAP7_75t_SL U15525 (.Y(n20324),
	.A(n19871),
	.B(n16798));
   NAND3xp33_ASAP7_75t_SL U15527 (.Y(n19951),
	.A(n19911),
	.B(n19938),
	.C(FE_OCPN29404_FE_OFN27148_sa32_3));
   NOR2x1_ASAP7_75t_SL U15528 (.Y(n18847),
	.A(FE_OCPN28245_n),
	.B(n17679));
   NAND2x1_ASAP7_75t_SL U15529 (.Y(n23412),
	.A(n18880),
	.B(n21064));
   NAND2x1p5_ASAP7_75t_L U15530 (.Y(n21718),
	.A(FE_OCPN27617_n18016),
	.B(n21738));
   NOR2x1_ASAP7_75t_L U15531 (.Y(n23450),
	.A(n17993),
	.B(n18015));
   NOR3xp33_ASAP7_75t_SL U15532 (.Y(n21158),
	.A(n18624),
	.B(n18623),
	.C(n18628));
   NOR2xp33_ASAP7_75t_L U15533 (.Y(n21155),
	.A(n18776),
	.B(n19129));
   NAND2xp5_ASAP7_75t_SL U15534 (.Y(n18766),
	.A(FE_OCPN29295_n18739),
	.B(n17245));
   NAND2xp5_ASAP7_75t_L U15535 (.Y(n19572),
	.A(FE_OFN28796_n17301),
	.B(n17271));
   NAND2xp5_ASAP7_75t_L U15536 (.Y(n19811),
	.A(FE_PSN8282_n21154),
	.B(FE_OCPN28389_n21479));
   NOR3x1_ASAP7_75t_SL U15537 (.Y(n22894),
	.A(FE_OFN27058_n22094),
	.B(FE_OFN28665_FE_OCPN27566),
	.C(n17771));
   NOR3xp33_ASAP7_75t_L U15538 (.Y(n20132),
	.A(n17765),
	.B(FE_OFN29102_FE_OCPN27261_sa02_0),
	.C(FE_OFN29148_n));
   NOR3xp33_ASAP7_75t_SL U15539 (.Y(n20176),
	.A(FE_OCPN29341_FE_OFN29148_n),
	.B(FE_OCPN27261_sa02_0),
	.C(n20962));
   NOR3x1_ASAP7_75t_L U15540 (.Y(n22888),
	.A(FE_OCPN27585_sa02_1),
	.B(FE_OCPN27261_sa02_0),
	.C(FE_OFN16234_sa02_2));
   NOR3xp33_ASAP7_75t_SL U15542 (.Y(n19461),
	.A(n17996),
	.B(FE_OCPN29451_n),
	.C(n18040));
   NAND2xp33_ASAP7_75t_SL U15543 (.Y(n19481),
	.A(n19464),
	.B(n18012));
   OAI21xp33_ASAP7_75t_L U15544 (.Y(n23420),
	.A1(FE_OFN29109_n),
	.A2(n19489),
	.B(n19488));
   NOR3xp33_ASAP7_75t_R U15545 (.Y(n19488),
	.A(n23443),
	.B(FE_OCPN29327_n21017),
	.C(n18008));
   NOR2x1_ASAP7_75t_L U15546 (.Y(n21278),
	.A(FE_OFN26581_n21317),
	.B(n21706));
   OAI22xp5_ASAP7_75t_L U15547 (.Y(n21279),
	.A1(FE_OCPN27998_n18019),
	.A2(FE_OCPN28184_n18020),
	.B1(n17996),
	.B2(FE_OCPN28184_n18020));
   NOR3x1_ASAP7_75t_SL U15548 (.Y(n21295),
	.A(FE_OFN21730_sa03_3),
	.B(FE_OFN28689_sa03_5),
	.C(FE_OCPN27405_sa03_4));
   NAND2xp5_ASAP7_75t_L U15549 (.Y(n16560),
	.A(n16559),
	.B(n16558));
   NAND2xp5_ASAP7_75t_L U15550 (.Y(n16561),
	.A(n16557),
	.B(n16558));
   NAND3xp33_ASAP7_75t_SL U15551 (.Y(n21900),
	.A(n23121),
	.B(n19674),
	.C(n19673));
   NAND2xp33_ASAP7_75t_R U15552 (.Y(n19674),
	.A(FE_OFN26161_sa10_4),
	.B(FE_OCPN27900_n23949));
   NOR3xp33_ASAP7_75t_R U15553 (.Y(n19673),
	.A(n19672),
	.B(n19671),
	.C(n19670));
   NOR3x1_ASAP7_75t_R U15554 (.Y(n21894),
	.A(n16556),
	.B(FE_OFN28751_n),
	.C(n16610));
   INVx1_ASAP7_75t_SL U15555 (.Y(n19771),
	.A(n23137));
   NOR3x1_ASAP7_75t_L U15556 (.Y(n19661),
	.A(n23036),
	.B(FE_OFN27196_n),
	.C(FE_OCPN27636_sa10_4));
   NOR2x1p5_ASAP7_75t_L U15557 (.Y(n24944),
	.A(FE_OFN28751_n),
	.B(n16556));
   OAI21xp5_ASAP7_75t_L U15559 (.Y(n24943),
	.A1(n23012),
	.A2(n16533),
	.B(n16642));
   NAND3xp33_ASAP7_75t_SL U15560 (.Y(n19573),
	.A(FE_OFN28744_FE_OCPN27908),
	.B(FE_OFN28514_sa00_1),
	.C(FE_OCPN27818_n17267));
   NOR2x1_ASAP7_75t_SL U15561 (.Y(n21479),
	.A(FE_OCPN29463_n),
	.B(n17262));
   NOR3x1_ASAP7_75t_SL U15562 (.Y(n21166),
	.A(FE_OFN28514_sa00_1),
	.B(FE_OCPN27818_n17267),
	.C(FE_OFN28744_FE_OCPN27908));
   NAND2xp5_ASAP7_75t_SL U15564 (.Y(n18387),
	.A(n17610),
	.B(n18360));
   NOR2xp67_ASAP7_75t_L U15566 (.Y(n22640),
	.A(n18364),
	.B(FE_OFN25901_n22133));
   NAND2xp33_ASAP7_75t_L U15567 (.Y(n22132),
	.A(n17602),
	.B(FE_OCPN8207_n18497));
   NOR2x1_ASAP7_75t_L U15568 (.Y(n21823),
	.A(FE_OCPN27313_n21845),
	.B(FE_OCPN28447_n23392));
   NOR3xp33_ASAP7_75t_SL U15569 (.Y(n19824),
	.A(n17298),
	.B(FE_OFN29249_n),
	.C(n18651));
   NAND2x1_ASAP7_75t_L U15570 (.Y(n19166),
	.A(n19206),
	.B(FE_OCPN27228_sa11_2));
   NAND3xp33_ASAP7_75t_SL U15571 (.Y(n17475),
	.A(FE_OCPN27625_sa11_5),
	.B(FE_OCPN29504_sa11_4),
	.C(n19170));
   NAND2xp5_ASAP7_75t_SL U15572 (.Y(n21385),
	.A(n17512),
	.B(n17511));
   NOR3x1_ASAP7_75t_L U15573 (.Y(n21373),
	.A(n19214),
	.B(FE_OFN29137_FE_OCPN27228_sa11_2),
	.C(FE_OCPN27592_n17501));
   NOR3xp33_ASAP7_75t_SL U15574 (.Y(n25793),
	.A(n21399),
	.B(n24551),
	.C(n23373));
   NAND2xp5_ASAP7_75t_L U15575 (.Y(n22495),
	.A(n17444),
	.B(FE_OFN29054_n17453));
   NOR2x1_ASAP7_75t_L U15576 (.Y(n21428),
	.A(n19192),
	.B(n21823));
   NAND2xp5_ASAP7_75t_R U15577 (.Y(n19194),
	.A(n21851),
	.B(FE_OFN16391_n22490));
   NAND3xp33_ASAP7_75t_SL U15578 (.Y(n22142),
	.A(n25108),
	.B(n17646),
	.C(FE_OFN16247_sa30_1));
   NAND2x1p5_ASAP7_75t_L U15579 (.Y(n19072),
	.A(FE_OCPN8207_n18497),
	.B(FE_OFN27176_n));
   NAND3xp33_ASAP7_75t_SL U15580 (.Y(n23721),
	.A(FE_OFN29139_n18527),
	.B(n18529),
	.C(FE_OFN29131_FE_OCPN27371_sa20_2));
   NOR2x1_ASAP7_75t_L U15581 (.Y(n23791),
	.A(FE_OFN28815_n18523),
	.B(FE_OCPN27891_n18561));
   NOR2xp33_ASAP7_75t_SL U15582 (.Y(n20646),
	.A(n25632),
	.B(n23797));
   NAND2x1p5_ASAP7_75t_SL U15583 (.Y(n18561),
	.A(FE_OFN29251_n18536),
	.B(n18524));
   NAND3xp33_ASAP7_75t_SL U15584 (.Y(n23302),
	.A(FE_OFN26136_sa22_3),
	.B(FE_OFN55_sa22_5),
	.C(FE_OFN16135_sa22_4));
   NAND3xp33_ASAP7_75t_L U15585 (.Y(n22312),
	.A(FE_OCPN29269_sa22_1),
	.B(sa22_0_),
	.C(FE_OFN28688_sa22_2));
   NAND2x2_ASAP7_75t_SL U15587 (.Y(n21123),
	.A(FE_OFN26136_sa22_3),
	.B(FE_OFN55_sa22_5));
   NOR2x1_ASAP7_75t_SL U15588 (.Y(n21787),
	.A(FE_OFN29238_n22811),
	.B(n21804));
   NAND2xp5_ASAP7_75t_SL U15589 (.Y(n23162),
	.A(n22802),
	.B(n22317));
   NOR3x1_ASAP7_75t_SL U15590 (.Y(n23792),
	.A(FE_OFN28815_n18523),
	.B(FE_OCPN27580_n),
	.C(n18602));
   NOR2x1_ASAP7_75t_L U15592 (.Y(n23864),
	.A(FE_OCPN27371_sa20_2),
	.B(n18547));
   NOR2x1_ASAP7_75t_R U15593 (.Y(n18431),
	.A(FE_OCPN27604_n16421),
	.B(n16947));
   NOR3xp33_ASAP7_75t_SL U15594 (.Y(n18141),
	.A(FE_OCPN27460_n16913),
	.B(FE_OFN26055_n),
	.C(n16676));
   NAND2xp5_ASAP7_75t_SL U15595 (.Y(n18405),
	.A(FE_OFN26055_n),
	.B(n16960));
   OAI21xp33_ASAP7_75t_L U15596 (.Y(n18104),
	.A1(FE_OFN26545_n16447),
	.A2(FE_OFN25960_n),
	.B(n16922));
   NOR2x1_ASAP7_75t_R U15597 (.Y(n18433),
	.A(FE_OCPN27604_n16421),
	.B(n16473));
   OAI21xp33_ASAP7_75t_R U15598 (.Y(n18135),
	.A1(n16925),
	.A2(FE_OFN29208_n16436),
	.B(n16924));
   NOR2x1_ASAP7_75t_L U15599 (.Y(n18143),
	.A(n16925),
	.B(FE_OFN29208_n16436));
   NAND2xp5_ASAP7_75t_R U15600 (.Y(n16416),
	.A(FE_OFN28727_sa33_1),
	.B(FE_OFN28643_sa33_0));
   NAND2x1p5_ASAP7_75t_L U15601 (.Y(n16847),
	.A(n16873),
	.B(FE_OCPN29438_sa33_2));
   NOR2xp67_ASAP7_75t_R U15602 (.Y(n23553),
	.A(n16847),
	.B(FE_OCPN27604_n16421));
   NOR3xp33_ASAP7_75t_SL U15603 (.Y(n18425),
	.A(n16473),
	.B(FE_OFN25938_sa33_3),
	.C(FE_OCPN28354_n16677));
   NOR2xp33_ASAP7_75t_L U15604 (.Y(n20942),
	.A(FE_OCPN28071_n25092),
	.B(FE_OFN29187_FE_OCPN27571_n20235));
   NOR3x1_ASAP7_75t_SL U15605 (.Y(n22925),
	.A(n22980),
	.B(FE_OCPN29374_FE_OFN29191_sa23_2),
	.C(FE_OCPN28107_n23504));
   NAND2xp5_ASAP7_75t_L U15606 (.Y(n20930),
	.A(n19313),
	.B(FE_OFN29026_n20911));
   NAND3xp33_ASAP7_75t_SL U15607 (.Y(n20270),
	.A(n23476),
	.B(n19328),
	.C(n22020));
   NAND3x1_ASAP7_75t_SL U15609 (.Y(n22046),
	.A(FE_OCPN28112_n26664),
	.B(FE_OCPN27727_n22964),
	.C(FE_OCPN29551_n));
   NOR2xp33_ASAP7_75t_L U15610 (.Y(n18668),
	.A(n17318),
	.B(n23107));
   NOR3xp33_ASAP7_75t_SL U15611 (.Y(n21571),
	.A(n18667),
	.B(FE_OFN28736_FE_OCPN28216_sa01_5),
	.C(n18684));
   NOR2xp33_ASAP7_75t_L U15612 (.Y(n21568),
	.A(n21560),
	.B(n23060));
   NAND3xp33_ASAP7_75t_SL U15613 (.Y(n21566),
	.A(n24396),
	.B(n21565),
	.C(n21564));
   NOR3xp33_ASAP7_75t_SL U15614 (.Y(n22601),
	.A(FE_OCPN29406_n18710),
	.B(FE_OFN28736_FE_OCPN28216_sa01_5),
	.C(n18684));
   NOR2xp33_ASAP7_75t_R U15615 (.Y(n17378),
	.A(n22436),
	.B(n23075));
   OAI21xp33_ASAP7_75t_R U15616 (.Y(n17376),
	.A1(FE_OFN27152_n17315),
	.A2(FE_OFN60_n27007),
	.B(n18677));
   OAI21xp33_ASAP7_75t_R U15617 (.Y(n17383),
	.A1(n18693),
	.A2(n17318),
	.B(n17372));
   NAND2xp5_ASAP7_75t_L U15618 (.Y(n23079),
	.A(FE_OFN29254_n),
	.B(n20371));
   NAND2x1p5_ASAP7_75t_L U15619 (.Y(n17389),
	.A(FE_OCPN28217_sa01_5),
	.B(n17326));
   NOR3x1_ASAP7_75t_SL U15620 (.Y(n23093),
	.A(FE_OCPN29406_n18710),
	.B(FE_OCPN29429_FE_OFN16141_sa01_3),
	.C(n17389));
   NAND3xp33_ASAP7_75t_SL U15621 (.Y(n23101),
	.A(FE_OFN28672_sa01_2),
	.B(FE_OFN28718_sa01_1),
	.C(FE_OCPN27423_sa01_0));
   NAND3x2_ASAP7_75t_SL U15622 (.Y(n22223),
	.A(FE_OCPN29484_sa12_3),
	.B(FE_OCPN29476_sa12_5),
	.C(FE_OCPN29453_sa12_4));
   NAND2x2_ASAP7_75t_SL U15623 (.Y(n17949),
	.A(FE_OCPN29485_sa12_3),
	.B(FE_OFN73_sa12_5));
   NAND2xp5_ASAP7_75t_L U15624 (.Y(n20549),
	.A(n20548),
	.B(n20547));
   NAND2xp5_ASAP7_75t_R U15626 (.Y(n20812),
	.A(FE_OCPN29485_sa12_3),
	.B(n17954));
   NOR2x1_ASAP7_75t_L U15627 (.Y(n17675),
	.A(FE_OCPN27230_sa32_3),
	.B(n17712));
   NOR2x1_ASAP7_75t_R U15628 (.Y(n19713),
	.A(FE_OFN28893_n),
	.B(FE_OFN26035_n));
   NOR2x1_ASAP7_75t_SL U15629 (.Y(n17693),
	.A(FE_OCPN29298_n25028),
	.B(n18836));
   NOR3xp33_ASAP7_75t_SRAM U15630 (.Y(n19726),
	.A(n18842),
	.B(n22369),
	.C(n17587));
   NOR3x1_ASAP7_75t_SL U15631 (.Y(n18813),
	.A(n17583),
	.B(n22384),
	.C(n18307));
   NAND2x1p5_ASAP7_75t_L U15632 (.Y(n18827),
	.A(n17565),
	.B(n17564));
   NAND2xp5_ASAP7_75t_L U15633 (.Y(n18800),
	.A(n18298),
	.B(n17560));
   NAND2x1p5_ASAP7_75t_SL U15634 (.Y(n18818),
	.A(FE_OCPN29405_FE_OFN27148_sa32_3),
	.B(n17553));
   NOR2xp33_ASAP7_75t_L U15635 (.Y(n18833),
	.A(n19710),
	.B(n19739));
   NOR2x1p5_ASAP7_75t_L U15636 (.Y(n20095),
	.A(FE_OCPN29323_n19721),
	.B(n18828));
   NAND3x1_ASAP7_75t_SL U15637 (.Y(n19889),
	.A(FE_OFN29023_n16750),
	.B(FE_OFN16153_n16747),
	.C(FE_OCPN5126_sa21_2));
   NAND3xp33_ASAP7_75t_L U15638 (.Y(n19972),
	.A(FE_OFN28836_FE_OCPN27631_n16774),
	.B(FE_OCPN27616_n16760),
	.C(FE_OCPN29265_FE_OFN28698_sa21_1));
   NAND2xp5_ASAP7_75t_L U15639 (.Y(n17878),
	.A(n17877),
	.B(n17874));
   NAND2xp33_ASAP7_75t_SL U15640 (.Y(n17879),
	.A(n17875),
	.B(n17874));
   NOR3x1_ASAP7_75t_SL U15642 (.Y(n22676),
	.A(n23633),
	.B(FE_OCPN29293_FE_OFN28678_sa21_3),
	.C(n16806));
   NOR2xp33_ASAP7_75t_L U15643 (.Y(n21924),
	.A(n18081),
	.B(n18080));
   NAND2xp33_ASAP7_75t_SRAM U15644 (.Y(n18080),
	.A(n18079),
	.B(n20066));
   NOR2x1_ASAP7_75t_L U15645 (.Y(n21935),
	.A(FE_OFN26570_n20866),
	.B(n18091));
   NAND2xp5_ASAP7_75t_SL U15646 (.Y(n16350),
	.A(n20868),
	.B(n16300));
   NAND3x1_ASAP7_75t_L U15647 (.Y(n21932),
	.A(n16348),
	.B(FE_OCPN27444_n20064),
	.C(FE_OCPN29483_FE_OFN26014_sa31_3));
   NOR2x1p5_ASAP7_75t_SL U15648 (.Y(n26290),
	.A(FE_OCPN28314_n20842),
	.B(n16408));
   NOR3xp33_ASAP7_75t_SL U15650 (.Y(n17031),
	.A(n17030),
	.B(n17045),
	.C(n19379));
   NAND3xp33_ASAP7_75t_SL U15651 (.Y(n17030),
	.A(n17162),
	.B(n20510),
	.C(n17029));
   NAND2xp5_ASAP7_75t_SL U15652 (.Y(n20312),
	.A(FE_OFN29023_n16750),
	.B(FE_OCPN27642_n16758));
   NAND2xp5_ASAP7_75t_SL U15653 (.Y(n22667),
	.A(n16771),
	.B(FE_OFN28779_n24257));
   NOR3xp33_ASAP7_75t_L U15654 (.Y(n16887),
	.A(n24617),
	.B(n16838),
	.C(n23530));
   NOR2xp33_ASAP7_75t_L U15655 (.Y(n23538),
	.A(FE_OCPN27604_n16421),
	.B(FE_OCPN27460_n16913));
   NAND2xp5_ASAP7_75t_R U15657 (.Y(n24385),
	.A(n24382),
	.B(FE_OFN28904_n25733));
   NAND2xp33_ASAP7_75t_R U15659 (.Y(n24410),
	.A(n24403),
	.B(n24402));
   NAND2xp33_ASAP7_75t_SRAM U15660 (.Y(n24402),
	.A(n24401),
	.B(n24400));
   NAND2xp33_ASAP7_75t_R U15661 (.Y(n24403),
	.A(n24398),
	.B(n24400));
   NOR3xp33_ASAP7_75t_L U15663 (.Y(n24728),
	.A(n24727),
	.B(n24726),
	.C(n24725));
   NOR3x1_ASAP7_75t_L U15664 (.Y(n26995),
	.A(n24763),
	.B(n24762),
	.C(n24761));
   NOR2xp33_ASAP7_75t_SL U15665 (.Y(n26311),
	.A(n26309),
	.B(n26308));
   OAI222xp33_ASAP7_75t_R U15666 (.Y(n26309),
	.A1(n26302),
	.A2(n27075),
	.B1(n26301),
	.B2(n27075),
	.C1(n26300),
	.C2(n27075));
   A2O1A1Ixp33_ASAP7_75t_L U15667 (.Y(n26308),
	.A1(n26307),
	.A2(n26306),
	.B(n27168),
	.C(n26305));
   NAND2xp5_ASAP7_75t_SL U15668 (.Y(n24269),
	.A(n19971),
	.B(n19970));
   NAND2xp33_ASAP7_75t_SL U15669 (.Y(n19970),
	.A(n19969),
	.B(FE_OCPN5167_n22336));
   NOR3xp33_ASAP7_75t_L U15670 (.Y(n25163),
	.A(n20592),
	.B(n20591),
	.C(n25438));
   NAND3xp33_ASAP7_75t_R U15671 (.Y(n20592),
	.A(n25399),
	.B(n25398),
	.C(n23234));
   NAND2xp5_ASAP7_75t_SL U15672 (.Y(n23265),
	.A(n21831),
	.B(n21830));
   NAND2xp33_ASAP7_75t_L U15673 (.Y(n21830),
	.A(n21829),
	.B(n21828));
   NAND2xp33_ASAP7_75t_L U15674 (.Y(n21831),
	.A(n21826),
	.B(n21828));
   NOR2xp33_ASAP7_75t_SRAM U15675 (.Y(n21829),
	.A(FE_OFN29034_FE_OCPN27414_n23359),
	.B(n21827));
   NOR2xp33_ASAP7_75t_R U15676 (.Y(n16890),
	.A(n16937),
	.B(n16446));
   NAND2xp33_ASAP7_75t_SRAM U15677 (.Y(n16446),
	.A(n16893),
	.B(n18446));
   NAND2xp33_ASAP7_75t_L U15678 (.Y(n23763),
	.A(n23752),
	.B(FE_OFN29096_n25188));
   NOR3x1_ASAP7_75t_R U15679 (.Y(n23787),
	.A(n21673),
	.B(n23835),
	.C(n23791));
   NOR3xp33_ASAP7_75t_L U15680 (.Y(n23771),
	.A(n23758),
	.B(n23812),
	.C(n23757));
   NAND3xp33_ASAP7_75t_L U15681 (.Y(n23758),
	.A(n23752),
	.B(n23751),
	.C(n23750));
   NAND3x2_ASAP7_75t_L U15682 (.Y(n25029),
	.A(FE_OFN28686_FE_OCPN27812),
	.B(FE_OFN26035_n),
	.C(FE_OFN28892_n));
   NAND3xp33_ASAP7_75t_SL U15683 (.Y(n18794),
	.A(FE_OFN28696_sa32_4),
	.B(FE_OCPN27499_FE_OFN16151_sa32_5),
	.C(FE_OFN27148_sa32_3));
   NAND2xp33_ASAP7_75t_SRAM U15684 (.Y(n19282),
	.A(n19280),
	.B(n19279));
   NAND3xp33_ASAP7_75t_L U15685 (.Y(n25208),
	.A(n19278),
	.B(n20127),
	.C(n19277));
   NAND2xp33_ASAP7_75t_SRAM U15686 (.Y(n19276),
	.A(n22534),
	.B(n22554));
   NAND3x1_ASAP7_75t_L U15687 (.Y(n25217),
	.A(n22573),
	.B(n22067),
	.C(n22906));
   NAND3xp33_ASAP7_75t_L U15689 (.Y(n25210),
	.A(n20204),
	.B(n22891),
	.C(n25301));
   NOR2xp33_ASAP7_75t_L U15690 (.Y(n20202),
	.A(n20186),
	.B(FE_OFN28897_n20132));
   NOR2xp67_ASAP7_75t_L U15691 (.Y(n22573),
	.A(n26972),
	.B(n22873));
   NAND3x2_ASAP7_75t_SL U15693 (.Y(n21441),
	.A(n12998),
	.B(FE_OFN28835_n),
	.C(FE_OCPN29370_FE_OFN28744));
   NAND3xp33_ASAP7_75t_SL U15694 (.Y(n27039),
	.A(FE_OFN16392_n24102),
	.B(n18621),
	.C(n18620));
   NOR3xp33_ASAP7_75t_SRAM U15695 (.Y(n18621),
	.A(n19121),
	.B(n19839),
	.C(n19813));
   NOR3x1_ASAP7_75t_L U15696 (.Y(n25635),
	.A(n18566),
	.B(n23775),
	.C(n18546));
   NOR3xp33_ASAP7_75t_SRAM U15697 (.Y(n18546),
	.A(n20670),
	.B(FE_OFN29251_n18536),
	.C(FE_OFN27045_n));
   NAND2xp33_ASAP7_75t_SL U15698 (.Y(n20683),
	.A(n20679),
	.B(n20680));
   NOR2xp33_ASAP7_75t_L U15699 (.Y(n20591),
	.A(FE_OFN27145_n23216),
	.B(FE_OFN26158_n22224));
   NOR3x1_ASAP7_75t_SL U15700 (.Y(n23214),
	.A(n20554),
	.B(FE_OCPN29494_sa12_4),
	.C(FE_OCPN28232_n17949));
   OAI22xp33_ASAP7_75t_SRAM U15701 (.Y(n19472),
	.A1(FE_OFN28589_n21048),
	.A2(FE_OCPN27918_n21042),
	.B1(FE_OCPN27617_n18016),
	.B2(FE_OCPN27918_n21042));
   NAND2xp5_ASAP7_75t_L U15702 (.Y(n19468),
	.A(n19467),
	.B(n19466));
   NAND2xp5_ASAP7_75t_L U15704 (.Y(n23476),
	.A(FE_OCPN28112_n26664),
	.B(FE_OFN16272_n24767));
   NAND2xp33_ASAP7_75t_R U15706 (.Y(n17669),
	.A(n17668),
	.B(n17667));
   NOR3xp33_ASAP7_75t_SRAM U15707 (.Y(n17670),
	.A(n25107),
	.B(n20481),
	.C(n22161));
   NAND2xp33_ASAP7_75t_SRAM U15708 (.Y(n17667),
	.A(n17666),
	.B(n17665));
   NAND3xp33_ASAP7_75t_SRAM U15709 (.Y(n18943),
	.A(n25994),
	.B(n27090),
	.C(n18939));
   NAND2xp5_ASAP7_75t_L U15710 (.Y(n18942),
	.A(n18941),
	.B(n18940));
   NOR3xp33_ASAP7_75t_SRAM U15711 (.Y(n17140),
	.A(FE_OCPN27684_n17139),
	.B(n18919),
	.C(n17144));
   NOR2xp33_ASAP7_75t_L U15712 (.Y(n17156),
	.A(FE_OFN29234_n16996),
	.B(n17154));
   NOR2xp33_ASAP7_75t_SRAM U15716 (.Y(n17176),
	.A(n16996),
	.B(n17174));
   NAND2xp5_ASAP7_75t_R U15717 (.Y(n24853),
	.A(FE_OCPN27230_sa32_3),
	.B(n17559));
   NOR2xp33_ASAP7_75t_R U15718 (.Y(n17559),
	.A(FE_OFN69_sa32_4),
	.B(n19920));
   NOR2xp33_ASAP7_75t_L U15719 (.Y(n21721),
	.A(FE_OCPN27628_n23455),
	.B(n23450));
   NAND3xp33_ASAP7_75t_SL U15720 (.Y(n17986),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2),
	.B(FE_OFN141_sa03_1),
	.C(FE_OCPN27726_n));
   NOR2xp33_ASAP7_75t_SL U15721 (.Y(n21272),
	.A(n21504),
	.B(n21505));
   NOR3xp33_ASAP7_75t_SL U15722 (.Y(n21277),
	.A(n19490),
	.B(n21296),
	.C(n18899));
   NAND2xp5_ASAP7_75t_SL U15723 (.Y(n18864),
	.A(n21069),
	.B(n18047));
   NOR3xp33_ASAP7_75t_L U15724 (.Y(n21282),
	.A(n19448),
	.B(n18859),
	.C(n18858));
   NAND3x1_ASAP7_75t_SL U15725 (.Y(n23441),
	.A(n18037),
	.B(n21047),
	.C(n21724));
   NOR3x1_ASAP7_75t_L U15726 (.Y(n18037),
	.A(n18036),
	.B(n21746),
	.C(n23449));
   NOR3xp33_ASAP7_75t_L U15728 (.Y(n25502),
	.A(n22540),
	.B(n22539),
	.C(FE_OCPN27424_n22560));
   NAND3xp33_ASAP7_75t_SL U15729 (.Y(n18734),
	.A(n17253),
	.B(n19094),
	.C(n18642));
   NOR3xp33_ASAP7_75t_SL U15730 (.Y(n24625),
	.A(n24094),
	.B(n24089),
	.C(FE_OFN28569_n18755));
   NOR3xp33_ASAP7_75t_L U15731 (.Y(n24626),
	.A(n17259),
	.B(FE_OFN28593_n18627),
	.C(n24093));
   NOR3xp33_ASAP7_75t_SL U15733 (.Y(n17085),
	.A(n17081),
	.B(n17171),
	.C(n17114));
   INVxp33_ASAP7_75t_SRAM U15734 (.Y(n17083),
	.A(n19431));
   NOR3x1_ASAP7_75t_L U15735 (.Y(n25307),
	.A(n17773),
	.B(n25211),
	.C(n20205));
   NOR2xp33_ASAP7_75t_R U15736 (.Y(n19269),
	.A(n25523),
	.B(FE_OCPN27424_n22560));
   NAND2xp33_ASAP7_75t_L U15737 (.Y(n19267),
	.A(n19266),
	.B(n19265));
   NOR3xp33_ASAP7_75t_SL U15738 (.Y(n19694),
	.A(n16626),
	.B(n23044),
	.C(n16625));
   NAND2xp33_ASAP7_75t_SL U15739 (.Y(n16626),
	.A(n19784),
	.B(n16624));
   NAND2xp5_ASAP7_75t_SRAM U15740 (.Y(n16624),
	.A(FE_OFN26161_sa10_4),
	.B(n16623));
   NAND2xp5_ASAP7_75t_R U15741 (.Y(n16651),
	.A(n23950),
	.B(n19771));
   NOR2x1_ASAP7_75t_L U15742 (.Y(n18490),
	.A(n17656),
	.B(n25082));
   NAND3xp33_ASAP7_75t_L U15743 (.Y(n18363),
	.A(n22639),
	.B(FE_PSN8333_n18478),
	.C(n18452));
   NOR2x1_ASAP7_75t_R U15745 (.Y(n20434),
	.A(n22636),
	.B(n17652));
   NAND2xp5_ASAP7_75t_SRAM U15746 (.Y(n17652),
	.A(n22626),
	.B(n20467));
   NAND3x1_ASAP7_75t_L U15748 (.Y(n26076),
	.A(n17472),
	.B(n17471),
	.C(n17512));
   NOR3xp33_ASAP7_75t_SL U15749 (.Y(n17472),
	.A(n21403),
	.B(FE_PSN8309_n21372),
	.C(n21422));
   NOR3xp33_ASAP7_75t_L U15750 (.Y(n17471),
	.A(n17469),
	.B(n21838),
	.C(n21368));
   NOR2x1p5_ASAP7_75t_L U15751 (.Y(n25082),
	.A(FE_OCPN27966_n18473),
	.B(FE_OFN25901_n22133));
   NOR3xp33_ASAP7_75t_L U15752 (.Y(n21599),
	.A(n17607),
	.B(FE_OFN28563_n20480),
	.C(n20438));
   NAND2xp33_ASAP7_75t_SRAM U15753 (.Y(n17607),
	.A(n22633),
	.B(n25104));
   NOR2xp33_ASAP7_75t_R U15755 (.Y(n20710),
	.A(n22828),
	.B(n21764));
   NOR2xp33_ASAP7_75t_L U15756 (.Y(n22276),
	.A(n21778),
	.B(n21789));
   NOR2xp33_ASAP7_75t_SRAM U15757 (.Y(n21778),
	.A(n21770),
	.B(FE_OFN25987_n23322));
   NAND2xp5_ASAP7_75t_SL U15758 (.Y(n25899),
	.A(n21206),
	.B(n21205));
   NAND2xp33_ASAP7_75t_L U15759 (.Y(n21205),
	.A(n23839),
	.B(n21204));
   AND3x1_ASAP7_75t_SL U15760 (.Y(n23862),
	.A(n20645),
	.B(n23766),
	.C(n20644));
   OAI222xp33_ASAP7_75t_SL U15761 (.Y(n24609),
	.A1(n18437),
	.A2(n24331),
	.B1(n18435),
	.B2(n24331),
	.C1(n18438),
	.C2(n24331));
   NOR2xp33_ASAP7_75t_L U15762 (.Y(n18435),
	.A(FE_OCPN29577_n24298),
	.B(FE_RN_193_0));
   OAI22xp33_ASAP7_75t_L U15764 (.Y(n18138),
	.A1(n16417),
	.A2(FE_OFN16241_n23552),
	.B1(n16418),
	.B2(FE_OFN16241_n23552));
   NAND2xp5_ASAP7_75t_L U15765 (.Y(n16696),
	.A(n16695),
	.B(n16694));
   NAND2xp5_ASAP7_75t_L U15766 (.Y(n16697),
	.A(n16693),
	.B(n16694));
   NOR3xp33_ASAP7_75t_SL U15767 (.Y(n18107),
	.A(n16436),
	.B(FE_OFN25938_sa33_3),
	.C(FE_OCPN28354_n16677));
   NAND3xp33_ASAP7_75t_SRAM U15768 (.Y(n25100),
	.A(n26557),
	.B(n26556),
	.C(n26553));
   NAND2xp33_ASAP7_75t_R U15769 (.Y(n26573),
	.A(n18984),
	.B(n18983));
   NAND2xp33_ASAP7_75t_R U15770 (.Y(n18984),
	.A(n18980),
	.B(n18981));
   NAND2xp5_ASAP7_75t_L U15771 (.Y(n26160),
	.A(FE_OFN29026_n20911),
	.B(n19000));
   NAND3xp33_ASAP7_75t_SL U15772 (.Y(n24767),
	.A(FE_OCPN27803_sa23_4),
	.B(FE_OFN27078_sa23_5),
	.C(FE_OFN27126_sa23_3));
   NAND3xp33_ASAP7_75t_L U15773 (.Y(n26551),
	.A(n22987),
	.B(n19012),
	.C(n20249));
   NAND2xp33_ASAP7_75t_R U15775 (.Y(n17367),
	.A(n17366),
	.B(n17365));
   NOR3xp33_ASAP7_75t_L U15776 (.Y(n24219),
	.A(n17328),
	.B(FE_OCPN28365_n21549),
	.C(n17356));
   NAND2xp5_ASAP7_75t_L U15777 (.Y(n17327),
	.A(n17325),
	.B(n17324));
   NAND2xp33_ASAP7_75t_L U15778 (.Y(n17324),
	.A(n17323),
	.B(n17322));
   NAND3xp33_ASAP7_75t_SL U15780 (.Y(n17962),
	.A(n23612),
	.B(n20795),
	.C(n17961));
   NAND2xp5_ASAP7_75t_L U15781 (.Y(n17959),
	.A(n17958),
	.B(n22735));
   NOR2xp33_ASAP7_75t_L U15784 (.Y(n22266),
	.A(n22730),
	.B(n17968));
   NAND3xp33_ASAP7_75t_L U15785 (.Y(n17968),
	.A(n20558),
	.B(n23236),
	.C(n23584));
   NAND2xp5_ASAP7_75t_L U15786 (.Y(n20112),
	.A(n17589),
	.B(n17588));
   NOR2xp33_ASAP7_75t_R U15787 (.Y(n17588),
	.A(n17675),
	.B(n17587));
   NOR2xp33_ASAP7_75t_L U15788 (.Y(n17589),
	.A(n17586),
	.B(n17585));
   OAI21xp33_ASAP7_75t_SRAM U15789 (.Y(n17586),
	.A1(n25029),
	.A2(FE_OCPN29298_n25028),
	.B(n18335));
   OAI21xp5_ASAP7_75t_SL U15790 (.Y(n18343),
	.A1(n22380),
	.A2(n18342),
	.B(n25367));
   NOR3xp33_ASAP7_75t_SL U15791 (.Y(n18344),
	.A(n18328),
	.B(n22369),
	.C(n18327));
   NAND3xp33_ASAP7_75t_SL U15792 (.Y(n18342),
	.A(n22395),
	.B(n18341),
	.C(n18340));
   NOR2x1_ASAP7_75t_R U15793 (.Y(n19908),
	.A(FE_OCPN27882_n18829),
	.B(n18818));
   NOR2x1_ASAP7_75t_SL U15794 (.Y(n25024),
	.A(n22383),
	.B(n18314));
   NAND2xp33_ASAP7_75t_L U15795 (.Y(n18311),
	.A(FE_OFN16231_n17691),
	.B(n18336));
   A2O1A1Ixp33_ASAP7_75t_SL U15797 (.Y(n23961),
	.A1(n26829),
	.A2(n25005),
	.B(n25002),
	.C(n23960));
   NAND2xp5_ASAP7_75t_L U15798 (.Y(n23962),
	.A(n25000),
	.B(n23959));
   NAND2xp33_ASAP7_75t_L U15801 (.Y(n16351),
	.A(n16349),
	.B(n20054));
   NOR3xp33_ASAP7_75t_SRAM U15802 (.Y(n25234),
	.A(n25220),
	.B(FE_OFN16220_n25219),
	.C(FE_OFN29228_n25218));
   NOR3xp33_ASAP7_75t_SRAM U15803 (.Y(n25233),
	.A(n25226),
	.B(n25225),
	.C(n25224));
   NAND2xp5_ASAP7_75t_L U15805 (.Y(n24276),
	.A(n24826),
	.B(n24449));
   O2A1O1Ixp33_ASAP7_75t_L U15806 (.Y(n26016),
	.A1(n26315),
	.A2(n26015),
	.B(n26014),
	.C(n26013));
   A2O1A1Ixp33_ASAP7_75t_SL U15807 (.Y(n25972),
	.A1(n27117),
	.A2(FE_PSN8300_n26482),
	.B(FE_OCPN27494_n26479),
	.C(n25971));
   A2O1A1Ixp33_ASAP7_75t_SL U15809 (.Y(n25661),
	.A1(n26829),
	.A2(n25959),
	.B(n25655),
	.C(n25654));
   O2A1O1Ixp33_ASAP7_75t_L U15810 (.Y(n25660),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25659),
	.C(n25658));
   A2O1A1Ixp33_ASAP7_75t_L U15811 (.Y(n25654),
	.A1(n25959),
	.A2(n26829),
	.B(FE_OFN16249_n25956),
	.C(FE_OFN25896_w3_4));
   NAND3xp33_ASAP7_75t_L U15812 (.Y(n24355),
	.A(n24356),
	.B(FE_OCPN28235_n26631),
	.C(n24502));
   NOR3xp33_ASAP7_75t_SL U15813 (.Y(n24352),
	.A(FE_OCPN27357_n26369),
	.B(n24353),
	.C(n24354));
   A2O1A1Ixp33_ASAP7_75t_SL U15814 (.Y(n25126),
	.A1(FE_OFN16164_n25081),
	.A2(n25080),
	.B(n25079),
	.C(n25078));
   A2O1A1Ixp33_ASAP7_75t_L U15815 (.Y(n25078),
	.A1(FE_OFN16164_n25081),
	.A2(n25080),
	.B(n25077),
	.C(w1_12_));
   NAND2xp5_ASAP7_75t_L U15816 (.Y(n25079),
	.A(n25076),
	.B(n25128));
   NAND2xp33_ASAP7_75t_L U15817 (.Y(n24448),
	.A(n24446),
	.B(n24445));
   NAND2xp33_ASAP7_75t_SRAM U15818 (.Y(n24446),
	.A(n24439),
	.B(FE_OFN118_sa03_7));
   A2O1A1Ixp33_ASAP7_75t_L U15819 (.Y(n24558),
	.A1(n27127),
	.A2(n24543),
	.B(n24542),
	.C(n24541));
   O2A1O1Ixp5_ASAP7_75t_SL U15820 (.Y(n24557),
	.A1(n17463),
	.A2(n24556),
	.B(n24555),
	.C(n24554));
   A2O1A1Ixp33_ASAP7_75t_SL U15821 (.Y(n25388),
	.A1(n25575),
	.A2(n25382),
	.B(n25381),
	.C(n25380));
   A2O1A1Ixp33_ASAP7_75t_SL U15822 (.Y(n25387),
	.A1(FE_OCPN29586_n26857),
	.A2(n26793),
	.B(n25386),
	.C(n25385));
   A2O1A1Ixp33_ASAP7_75t_SL U15823 (.Y(n25917),
	.A1(n26915),
	.A2(n26753),
	.B(n26750),
	.C(FE_OFN27142_n25934));
   A2O1A1Ixp33_ASAP7_75t_SL U15824 (.Y(n24982),
	.A1(n24974),
	.A2(n24939),
	.B(n24938),
	.C(n24937));
   NAND2xp33_ASAP7_75t_SL U15825 (.Y(n24938),
	.A(n24935),
	.B(FE_OFN28571_w3_28));
   NOR2xp33_ASAP7_75t_L U15827 (.Y(n26323),
	.A(sa20_6_),
	.B(sa20_7_));
   NAND2xp5_ASAP7_75t_L U15828 (.Y(n14578),
	.A(n14575),
	.B(n14574));
   NAND2xp33_ASAP7_75t_R U15829 (.Y(n14575),
	.A(n14571),
	.B(n14572));
   INVxp33_ASAP7_75t_L U15830 (.Y(n14580),
	.A(n14576));
   OR2x2_ASAP7_75t_L U15831 (.Y(n14160),
	.A(n14607),
	.B(n15975));
   NAND2xp33_ASAP7_75t_R U15833 (.Y(n14124),
	.A(n14116),
	.B(n14938));
   NOR2xp33_ASAP7_75t_R U15834 (.Y(n14138),
	.A(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(n15380));
   INVxp67_ASAP7_75t_L U15835 (.Y(n13980),
	.A(n13978));
   NOR2xp33_ASAP7_75t_SL U15836 (.Y(n13985),
	.A(FE_OFN26007_n16010),
	.B(n15956));
   NOR2xp33_ASAP7_75t_L U15837 (.Y(n14858),
	.A(n15835),
	.B(n15045));
   NOR3x1_ASAP7_75t_L U15840 (.Y(n14498),
	.A(FE_OCPN27655_w3_25),
	.B(FE_OCPN8232_FE_OFN27206_w3_30),
	.C(FE_OFN28891_n));
   NAND3xp33_ASAP7_75t_SL U15841 (.Y(n15253),
	.A(FE_OFN28530_n14593),
	.B(FE_OFN16159_w3_24),
	.C(FE_OFN16412_w3_26));
   NAND3xp33_ASAP7_75t_SRAM U15842 (.Y(n15822),
	.A(FE_OFN27124_w3_1),
	.B(FE_OFN26645_n),
	.C(FE_OCPN27978_w3_3));
   NAND2xp33_ASAP7_75t_R U15843 (.Y(n13976),
	.A(n13975),
	.B(n14112));
   INVxp67_ASAP7_75t_L U15844 (.Y(n13975),
	.A(n15959));
   NAND2x1p5_ASAP7_75t_L U15846 (.Y(n13870),
	.A(FE_OFN16426_w3_20),
	.B(w3_21_));
   OAI21x1_ASAP7_75t_R U15847 (.Y(n14795),
	.A1(FE_OFN27096_n),
	.A2(FE_OFN27214_w3_17),
	.B(FE_OFN27151_n));
   NOR2xp33_ASAP7_75t_L U15852 (.Y(n18946),
	.A(FE_OFN16162_n25869),
	.B(n19410));
   NAND2xp5_ASAP7_75t_SL U15853 (.Y(n20137),
	.A(FE_OFN28812_FE_OCPN27261_sa02_0),
	.B(n20982));
   NOR2x1p5_ASAP7_75t_L U15855 (.Y(n18776),
	.A(FE_OFN26651_n19573),
	.B(FE_OCPN28270_n17237));
   NAND2xp5_ASAP7_75t_R U15857 (.Y(n19489),
	.A(FE_OCPN28214_n21500),
	.B(FE_OCPN27285_n18011));
   NAND2xp5_ASAP7_75t_SL U15858 (.Y(n18040),
	.A(sa03_2_),
	.B(sa03_1_));
   INVxp33_ASAP7_75t_L U15859 (.Y(n17622),
	.A(FE_OCPN27428_n26027));
   NOR2x1_ASAP7_75t_SL U15860 (.Y(n21824),
	.A(n21406),
	.B(n21400));
   NAND2xp67_ASAP7_75t_SL U15861 (.Y(n21400),
	.A(n23370),
	.B(n22486));
   NAND3xp33_ASAP7_75t_SL U15862 (.Y(n21655),
	.A(FE_OFN28776_n18532),
	.B(FE_OFN29140_n18527),
	.C(FE_OCPN7660_FE_OFN28720_sa20_1));
   NAND3xp33_ASAP7_75t_L U15864 (.Y(n23688),
	.A(FE_OFN29251_n18536),
	.B(n18532),
	.C(FE_OCPN29380_sa20_1));
   NAND2x1_ASAP7_75t_L U15868 (.Y(n18989),
	.A(FE_OCPN27803_sa23_4),
	.B(FE_OFN28850_FE_OCPN27840));
   NOR3xp33_ASAP7_75t_SRAM U15870 (.Y(n20371),
	.A(n22450),
	.B(FE_OCPN27423_sa01_0),
	.C(FE_OFN28718_sa01_1));
   NOR3xp33_ASAP7_75t_SL U15872 (.Y(n20339),
	.A(n22663),
	.B(FE_OFN28903_sa21_0),
	.C(n17881));
   NAND2xp33_ASAP7_75t_SRAM U15873 (.Y(n16814),
	.A(FE_OCPN27328_sa21_2),
	.B(n19967));
   NAND2xp5_ASAP7_75t_L U15875 (.Y(n17591),
	.A(n17563),
	.B(n17564));
   NOR2xp33_ASAP7_75t_L U15876 (.Y(n23037),
	.A(n23035),
	.B(n23038));
   NOR3xp33_ASAP7_75t_SL U15878 (.Y(n17747),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(n17760),
	.C(n17763));
   NAND2xp33_ASAP7_75t_SRAM U15879 (.Y(n14018),
	.A(n15338),
	.B(n12994));
   NOR2xp33_ASAP7_75t_SRAM U15880 (.Y(n14493),
	.A(FE_OCPN28096_w3_31),
	.B(FE_OFN27129_w3_28));
   INVx1_ASAP7_75t_L U15881 (.Y(n14439),
	.A(n15601));
   INVxp67_ASAP7_75t_R U15882 (.Y(n15434),
	.A(n15999));
   NAND3xp33_ASAP7_75t_SL U15883 (.Y(n13876),
	.A(FE_OFN28908_w3_23),
	.B(w3_21_),
	.C(FE_OFN16426_w3_20));
   NAND2x1p5_ASAP7_75t_SL U15884 (.Y(n15339),
	.A(FE_OFN26538_w3_19),
	.B(FE_OCPN27929_FE_OFN4_w3_22));
   NOR2x1_ASAP7_75t_L U15885 (.Y(n15636),
	.A(FE_OCPN28072_w3_3),
	.B(FE_OFN28695_n));
   NOR2xp33_ASAP7_75t_R U15886 (.Y(n15792),
	.A(n15080),
	.B(n13725));
   NOR2x1p5_ASAP7_75t_L U15887 (.Y(n15438),
	.A(FE_OCPN29535_FE_OFN8_w3_14),
	.B(n15963));
   NAND2xp5_ASAP7_75t_L U15888 (.Y(n15936),
	.A(FE_OFN26633_w3_14),
	.B(FE_OFN27115_n));
   NOR2xp33_ASAP7_75t_R U15889 (.Y(n15275),
	.A(FE_PSN8280_n15660),
	.B(n13869));
   INVxp33_ASAP7_75t_L U15890 (.Y(n13577),
	.A(n13575));
   NAND3xp33_ASAP7_75t_SRAM U15891 (.Y(n13574),
	.A(FE_OFN25895_n13662),
	.B(n15156),
	.C(FE_OFN16193_n15200));
   NOR2xp33_ASAP7_75t_L U15892 (.Y(n13776),
	.A(FE_OCPN28072_w3_3),
	.B(FE_OFN28889_n15845));
   NAND2xp5_ASAP7_75t_SL U15893 (.Y(n15825),
	.A(FE_OFN28671_FE_OCPN28076),
	.B(FE_OFN25912_n15848));
   OR3x1_ASAP7_75t_SRAM U15894 (.Y(n14845),
	.A(n13726),
	.B(FE_OFN28662_w3_7),
	.C(n14996));
   NOR2xp33_ASAP7_75t_L U15895 (.Y(n14449),
	.A(n15061),
	.B(n13725));
   NAND3xp33_ASAP7_75t_SRAM U15896 (.Y(n14931),
	.A(FE_PSN8271_n15924),
	.B(n13804),
	.C(FE_OFN27200_n));
   OAI21xp5_ASAP7_75t_L U15897 (.Y(n15539),
	.A1(FE_OFN27096_n),
	.A2(FE_PSN8292_FE_OFN26041_w3_17),
	.B(FE_OFN26114_n));
   OA21x2_ASAP7_75t_R U15898 (.Y(n15308),
	.A1(n15478),
	.A2(n13890),
	.B(n15304));
   NAND2xp33_ASAP7_75t_SL U15899 (.Y(n15304),
	.A(n15303),
	.B(n15302));
   NAND2xp33_ASAP7_75t_L U15900 (.Y(n15302),
	.A(n15301),
	.B(n15300));
   NAND2xp33_ASAP7_75t_L U15901 (.Y(n15303),
	.A(n15299),
	.B(n15300));
   NAND2xp33_ASAP7_75t_L U15902 (.Y(n13502),
	.A(n14573),
	.B(n14593));
   NAND3xp33_ASAP7_75t_L U15903 (.Y(n15870),
	.A(FE_OFN25897_w3_4),
	.B(n14430),
	.C(n15857));
   NAND2xp5_ASAP7_75t_L U15904 (.Y(n15601),
	.A(FE_OCPN27978_w3_3),
	.B(FE_OFN26057_w3_1));
   NAND3xp33_ASAP7_75t_L U15905 (.Y(n15626),
	.A(n25140),
	.B(FE_OFN28732_n),
	.C(FE_OCPN29537_FE_OFN28699_w3_6));
   NOR2xp33_ASAP7_75t_SRAM U15906 (.Y(n14980),
	.A(n14976),
	.B(n13725));
   NAND3xp33_ASAP7_75t_SL U15907 (.Y(n14985),
	.A(FE_OFN28829_n),
	.B(FE_OFN28732_n),
	.C(FE_OFN29209_FE_OCPN27978_w3_3));
   NAND2xp5_ASAP7_75t_R U15908 (.Y(n15446),
	.A(FE_OFN26642_w3_14),
	.B(FE_OCPN29506_FE_OFN16184_w3_9));
   NOR3xp33_ASAP7_75t_SL U15909 (.Y(n15953),
	.A(n15969),
	.B(FE_OCPN29521_n24755),
	.C(n14913));
   INVxp33_ASAP7_75t_L U15910 (.Y(n15403),
	.A(n15399));
   NAND3xp33_ASAP7_75t_SRAM U15911 (.Y(n15397),
	.A(n15948),
	.B(n15956),
	.C(FE_OFN28758_n15422));
   NOR2x1p5_ASAP7_75t_SL U15912 (.Y(n15528),
	.A(FE_OFN28_w3_23),
	.B(n13870));
   NAND3xp33_ASAP7_75t_L U15914 (.Y(n14254),
	.A(n15514),
	.B(n14795),
	.C(n12994));
   NAND3x1_ASAP7_75t_SL U15915 (.Y(n14276),
	.A(FE_OFN26045_n25377),
	.B(FE_OFN5_w3_22),
	.C(FE_OFN26539_w3_19));
   NAND3xp33_ASAP7_75t_SRAM U15916 (.Y(n13462),
	.A(n13713),
	.B(n15156),
	.C(n13691));
   NOR3x1_ASAP7_75t_R U15917 (.Y(n14986),
	.A(FE_OFN28695_n),
	.B(FE_OCPN27978_w3_3),
	.C(FE_OFN26057_w3_1));
   NAND2xp5_ASAP7_75t_L U15918 (.Y(n14442),
	.A(FE_OFN27124_w3_1),
	.B(FE_OFN26645_n));
   OAI21xp33_ASAP7_75t_SRAM U15919 (.Y(n14914),
	.A1(FE_OCPN29535_FE_OFN8_w3_14),
	.A2(FE_OFN28856_n15450),
	.B(n14938));
   OAI21xp5_ASAP7_75t_SL U15920 (.Y(n15477),
	.A1(FE_OFN27151_n),
	.A2(n14778),
	.B(n15339));
   NAND2x1p5_ASAP7_75t_R U15921 (.Y(n15484),
	.A(FE_OFN26045_n25377),
	.B(FE_OFN26053_n25415));
   NAND2xp5_ASAP7_75t_L U15923 (.Y(n15861),
	.A(FE_OFN25912_n15848),
	.B(n15842));
   OAI21xp5_ASAP7_75t_L U15924 (.Y(n15983),
	.A1(FE_OFN27115_n),
	.A2(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(FE_OCPN29534_FE_OFN8_w3_14));
   NAND3xp33_ASAP7_75t_L U15925 (.Y(n15949),
	.A(n25051),
	.B(FE_OFN25961_w3_8),
	.C(n15934));
   NAND2xp5_ASAP7_75t_R U15926 (.Y(n15668),
	.A(n13873),
	.B(n15743));
   NAND2xp33_ASAP7_75t_L U15927 (.Y(n13873),
	.A(n13872),
	.B(FE_OFN28600_n14289));
   NAND3xp33_ASAP7_75t_SRAM U15928 (.Y(n15710),
	.A(n13867),
	.B(FE_OFN28712_n),
	.C(n15667));
   NAND2xp33_ASAP7_75t_L U15929 (.Y(n15743),
	.A(n15487),
	.B(FE_OFN28600_n14289));
   NOR2x1_ASAP7_75t_L U15930 (.Y(n14573),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN26049_w3_27));
   OAI21xp5_ASAP7_75t_SL U15931 (.Y(n15158),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OCPN27659_w3_25),
	.B(FE_OFN27206_w3_30));
   INVxp67_ASAP7_75t_L U15932 (.Y(n13692),
	.A(n15171));
   NAND3xp33_ASAP7_75t_SL U15933 (.Y(n13636),
	.A(FE_OCPN29571_n26355),
	.B(n13530),
	.C(n15167));
   NOR2xp33_ASAP7_75t_L U15935 (.Y(n15171),
	.A(FE_OFN26051_w3_27),
	.B(FE_OFN27211_w3_30));
   NAND3xp33_ASAP7_75t_SL U15936 (.Y(n15233),
	.A(FE_OCPN28096_w3_31),
	.B(FE_OFN27130_w3_28),
	.C(FE_OFN28452_w3_29));
   NAND3xp33_ASAP7_75t_L U15937 (.Y(n15205),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN27207_w3_30),
	.C(FE_OFN26049_w3_27));
   NAND2xp5_ASAP7_75t_SL U15938 (.Y(n14410),
	.A(n13752),
	.B(n13751));
   INVxp67_ASAP7_75t_L U15940 (.Y(n13752),
	.A(n14996));
   NOR3xp33_ASAP7_75t_L U15941 (.Y(n15845),
	.A(FE_OFN25896_w3_4),
	.B(FE_OFN29052_w3_5),
	.C(FE_OFN28661_w3_7));
   NOR2xp33_ASAP7_75t_SRAM U15942 (.Y(n23905),
	.A(n26819),
	.B(n23906));
   NAND2xp5_ASAP7_75t_L U15944 (.Y(n25027),
	.A(n18298),
	.B(FE_OCPN28434_n17546));
   O2A1O1Ixp33_ASAP7_75t_SL U15945 (.Y(n24707),
	.A1(n26880),
	.A2(n26879),
	.B(n26878),
	.C(n24706));
   NOR3xp33_ASAP7_75t_L U15947 (.Y(n24704),
	.A(n24703),
	.B(n26870),
	.C(n26876));
   NOR2x1_ASAP7_75t_SL U15948 (.Y(n21351),
	.A(n19222),
	.B(FE_OCPN27496_n21820));
   NAND2xp5_ASAP7_75t_L U15949 (.Y(n22771),
	.A(n19532),
	.B(n19531));
   NAND2xp33_ASAP7_75t_L U15950 (.Y(n19531),
	.A(n19530),
	.B(FE_OCPN27252_n22753));
   NAND2xp33_ASAP7_75t_L U15951 (.Y(n19532),
	.A(n19528),
	.B(FE_OCPN27252_n22753));
   NAND2xp33_ASAP7_75t_L U15952 (.Y(n22122),
	.A(n18505),
	.B(n18504));
   NAND2xp33_ASAP7_75t_L U15955 (.Y(n19036),
	.A(n18463),
	.B(FE_PSN8308_n22624));
   NAND2xp5_ASAP7_75t_SL U15956 (.Y(n18390),
	.A(n18389),
	.B(n19047));
   NOR2xp33_ASAP7_75t_R U15957 (.Y(n22631),
	.A(n22642),
	.B(n19061));
   OAI21xp33_ASAP7_75t_SRAM U15958 (.Y(n19061),
	.A1(FE_OFN28896_sa30_2),
	.A2(n25105),
	.B(n21584));
   NAND2x1p5_ASAP7_75t_SL U15960 (.Y(n18306),
	.A(FE_OCPN29449_n17521),
	.B(n17525));
   NOR2xp33_ASAP7_75t_L U15961 (.Y(n18843),
	.A(n19739),
	.B(n17714));
   OAI21xp33_ASAP7_75t_L U15962 (.Y(n17714),
	.A1(n18818),
	.A2(FE_OCPN28423_n18836),
	.B(n17713));
   NOR3x1_ASAP7_75t_L U15964 (.Y(n24869),
	.A(n18827),
	.B(FE_OCPN29459_n),
	.C(n17592));
   NAND2x1p5_ASAP7_75t_L U15965 (.Y(n24867),
	.A(n18847),
	.B(n19940));
   INVx1_ASAP7_75t_L U15966 (.Y(n18324),
	.A(FE_OCPN27267_n18794));
   NOR3x1_ASAP7_75t_SL U15968 (.Y(n25711),
	.A(n20235),
	.B(FE_OCPN29441_sa23_4),
	.C(n22971));
   NAND2x1_ASAP7_75t_SL U15970 (.Y(n22272),
	.A(n22795),
	.B(FE_OCPN27947_n18177));
   INVx1_ASAP7_75t_R U15971 (.Y(n21118),
	.A(n22277));
   NAND2xp5_ASAP7_75t_L U15972 (.Y(n23951),
	.A(n19641),
	.B(n16643));
   AND3x1_ASAP7_75t_SRAM U15973 (.Y(n20693),
	.A(n23699),
	.B(n21637),
	.C(n25189));
   NOR2xp33_ASAP7_75t_L U15974 (.Y(n20678),
	.A(n20636),
	.B(n23688));
   NAND2x1_ASAP7_75t_SL U15976 (.Y(n21544),
	.A(n20367),
	.B(n22470));
   NOR2xp67_ASAP7_75t_L U15978 (.Y(n23138),
	.A(n17191),
	.B(n16576));
   NOR3xp33_ASAP7_75t_SL U15980 (.Y(n21733),
	.A(n17993),
	.B(FE_OCPN29451_n),
	.C(n18040));
   NAND3xp33_ASAP7_75t_R U15981 (.Y(n22194),
	.A(n22458),
	.B(n20386),
	.C(n21535));
   NAND2xp5_ASAP7_75t_L U15982 (.Y(n20081),
	.A(n24181),
	.B(FE_OCPN27516_n26292));
   NAND3xp33_ASAP7_75t_L U15983 (.Y(n25359),
	.A(n20296),
	.B(n20295),
	.C(n20324));
   NAND2xp33_ASAP7_75t_SRAM U15984 (.Y(n20295),
	.A(n20294),
	.B(n20293));
   NAND2xp33_ASAP7_75t_SRAM U15985 (.Y(n20293),
	.A(n20292),
	.B(n20291));
   NAND2xp33_ASAP7_75t_SRAM U15986 (.Y(n20294),
	.A(n20290),
	.B(n20291));
   NAND2x1_ASAP7_75t_SL U15987 (.Y(n16953),
	.A(FE_OCPN8256_n16873),
	.B(n16430));
   OAI22xp33_ASAP7_75t_SRAM U15988 (.Y(n17643),
	.A1(FE_OCPN8207_n18497),
	.A2(n22156),
	.B1(n17603),
	.B2(n22156));
   NOR2x1_ASAP7_75t_SL U15989 (.Y(n18373),
	.A(n20429),
	.B(n18473));
   NAND2xp33_ASAP7_75t_L U15990 (.Y(n19364),
	.A(n17146),
	.B(n17145));
   NAND3xp33_ASAP7_75t_L U15991 (.Y(n17117),
	.A(FE_OCPN27761_n16977),
	.B(FE_OCPN28137_n17170),
	.C(FE_OFN29173_n));
   NAND2xp5_ASAP7_75t_SL U15992 (.Y(n19698),
	.A(n22378),
	.B(n25027));
   NAND2x1_ASAP7_75t_SL U15993 (.Y(n20103),
	.A(n18321),
	.B(n19741));
   NAND3xp33_ASAP7_75t_L U15994 (.Y(n20105),
	.A(n19943),
	.B(n19942),
	.C(n19941));
   NAND2xp5_ASAP7_75t_L U15995 (.Y(n17765),
	.A(n20993),
	.B(FE_OCPN27273_sa02_3));
   NAND2x1_ASAP7_75t_SL U15996 (.Y(n17771),
	.A(n17760),
	.B(n17763));
   NAND2xp5_ASAP7_75t_R U15997 (.Y(n21069),
	.A(FE_OCPN27393_sa03_0),
	.B(n18046));
   NOR2x1_ASAP7_75t_SL U15998 (.Y(n18859),
	.A(n23457),
	.B(FE_OCPN27599_n18875));
   NAND3xp33_ASAP7_75t_SL U15999 (.Y(n21719),
	.A(n21295),
	.B(FE_OCPN28214_n21500),
	.C(FE_OFN29109_n));
   NOR2x1_ASAP7_75t_L U16000 (.Y(n18904),
	.A(FE_OFN26581_n21317),
	.B(FE_OFN28951_n18011));
   NOR3xp33_ASAP7_75t_SL U16003 (.Y(n21475),
	.A(n21454),
	.B(n21453),
	.C(n21452));
   NAND2xp33_ASAP7_75t_SL U16004 (.Y(n21454),
	.A(n21451),
	.B(n21450));
   NAND3xp33_ASAP7_75t_SL U16005 (.Y(n18755),
	.A(n19572),
	.B(n18635),
	.C(n18620));
   NAND2xp33_ASAP7_75t_SL U16007 (.Y(n17280),
	.A(n17279),
	.B(n17278));
   NAND2xp33_ASAP7_75t_SL U16008 (.Y(n17281),
	.A(n17277),
	.B(n17278));
   NOR2x1_ASAP7_75t_L U16009 (.Y(n17102),
	.A(FE_OCPN27589_n25987),
	.B(n17043));
   NAND2xp33_ASAP7_75t_R U16010 (.Y(n17095),
	.A(FE_OFN28801_n16978),
	.B(n16983));
   NOR2x1p5_ASAP7_75t_L U16012 (.Y(n20170),
	.A(FE_OFN28665_FE_OCPN27566),
	.B(n17771));
   NAND3xp33_ASAP7_75t_L U16013 (.Y(n19257),
	.A(FE_OCPN28357_n22882),
	.B(FE_OCPN29469_n17747),
	.C(FE_OFN28812_FE_OCPN27261_sa02_0));
   NAND3xp33_ASAP7_75t_L U16014 (.Y(n22554),
	.A(FE_OCPN28357_n22882),
	.B(n22089),
	.C(FE_OCPN27261_sa02_0));
   NOR2x1_ASAP7_75t_L U16015 (.Y(n22539),
	.A(FE_OFN28800_n22526),
	.B(n22529));
   NOR2xp67_ASAP7_75t_L U16016 (.Y(n20174),
	.A(n22095),
	.B(n17798));
   NAND2x1_ASAP7_75t_L U16017 (.Y(n22065),
	.A(FE_OFN28703_FE_OCPN27740_sa02_4),
	.B(n20189));
   NAND3xp33_ASAP7_75t_L U16018 (.Y(n20204),
	.A(FE_OCPN27634_n20169),
	.B(FE_OCPN29469_n17747),
	.C(FE_OFN16234_sa02_2));
   NOR2x1_ASAP7_75t_L U16019 (.Y(n22561),
	.A(FE_OFN28941_sa02_2),
	.B(n22076));
   NOR3xp33_ASAP7_75t_SL U16020 (.Y(n25912),
	.A(FE_OFN29148_n),
	.B(FE_OFN29102_FE_OCPN27261_sa02_0),
	.C(n20196));
   NOR3x1_ASAP7_75t_SL U16022 (.Y(n17776),
	.A(n22873),
	.B(n20194),
	.C(FE_OCPN27972_n20988));
   NAND2x1p5_ASAP7_75t_SL U16023 (.Y(n17033),
	.A(n17060),
	.B(FE_OCPN28121_n16975));
   NAND2x1_ASAP7_75t_L U16024 (.Y(n25221),
	.A(FE_OCPN27859_n25868),
	.B(n19376));
   NAND2x1_ASAP7_75t_SL U16025 (.Y(n18272),
	.A(FE_OCPN27859_n25868),
	.B(FE_OCPN28212_n16980));
   NAND3xp33_ASAP7_75t_L U16026 (.Y(n19414),
	.A(FE_OFN16162_n25869),
	.B(FE_OCPN28121_n16975),
	.C(FE_OFN28491_sa13_3));
   NOR2xp33_ASAP7_75t_L U16027 (.Y(n19475),
	.A(FE_OCPN28184_n18020),
	.B(FE_OFN28950_n18011));
   NOR2x1_ASAP7_75t_R U16030 (.Y(n21058),
	.A(FE_OFN27189_n),
	.B(n21292));
   NAND2xp5_ASAP7_75t_L U16031 (.Y(n21047),
	.A(FE_OFN29124_n),
	.B(n21733));
   NAND2xp5_ASAP7_75t_R U16032 (.Y(n21060),
	.A(n21295),
	.B(FE_OFN28589_n21048));
   NAND3xp33_ASAP7_75t_SL U16033 (.Y(n21755),
	.A(n21272),
	.B(n17999),
	.C(FE_OCPN28297_n23417));
   NOR2xp33_ASAP7_75t_L U16034 (.Y(n17999),
	.A(n23430),
	.B(n23412));
   NOR3xp33_ASAP7_75t_SL U16035 (.Y(n21525),
	.A(n21067),
	.B(FE_OCPN29451_n),
	.C(n18040));
   NOR2x1_ASAP7_75t_SL U16036 (.Y(n21529),
	.A(n18891),
	.B(n18890));
   OAI21xp5_ASAP7_75t_SL U16037 (.Y(n18890),
	.A1(FE_OCPN28184_n18020),
	.A2(FE_OCPN27733_n17996),
	.B(n18889));
   NOR3x1_ASAP7_75t_L U16038 (.Y(n21524),
	.A(n18015),
	.B(FE_OCPN27483_FE_OFN16132_sa03_5),
	.C(FE_OFN28997_sa03_4));
   NOR3x1_ASAP7_75t_L U16039 (.Y(n21297),
	.A(FE_OFN26581_n21317),
	.B(FE_OCPN7619_FE_OFN28689_sa03_5),
	.C(n18029));
   OAI21xp5_ASAP7_75t_L U16040 (.Y(n21518),
	.A1(FE_OCPN27998_n18019),
	.A2(FE_OFN28588_n21048),
	.B(n18878));
   NAND2xp33_ASAP7_75t_L U16041 (.Y(n18878),
	.A(n21295),
	.B(n21738));
   NAND2xp5_ASAP7_75t_L U16042 (.Y(n17186),
	.A(n17222),
	.B(n23135));
   NOR2x1p5_ASAP7_75t_SL U16043 (.Y(n23995),
	.A(n16648),
	.B(n21902));
   NOR2xp33_ASAP7_75t_L U16044 (.Y(n19660),
	.A(n17190),
	.B(n21888));
   NOR2xp33_ASAP7_75t_L U16045 (.Y(n19635),
	.A(n17221),
	.B(n17220));
   NAND2xp5_ASAP7_75t_R U16046 (.Y(n17220),
	.A(n17219),
	.B(n23128));
   NAND2xp5_ASAP7_75t_SL U16047 (.Y(n17222),
	.A(FE_OCPN28157_n16534),
	.B(n19787));
   NOR2xp33_ASAP7_75t_L U16048 (.Y(n21896),
	.A(n24734),
	.B(n19772));
   OAI21xp5_ASAP7_75t_L U16049 (.Y(n21890),
	.A1(FE_OFN25956_n16575),
	.A2(n19677),
	.B(n16655));
   NOR3xp33_ASAP7_75t_L U16050 (.Y(n16655),
	.A(n19774),
	.B(n19791),
	.C(n21872));
   NOR2xp33_ASAP7_75t_L U16051 (.Y(n19625),
	.A(FE_OFN130_sa10_5),
	.B(n23951));
   NAND2xp5_ASAP7_75t_SL U16052 (.Y(n21901),
	.A(n17194),
	.B(n17193));
   NAND2xp5_ASAP7_75t_SL U16053 (.Y(n16637),
	.A(n23148),
	.B(n19787));
   NAND2x1p5_ASAP7_75t_L U16054 (.Y(n19644),
	.A(n23980),
	.B(FE_OCPN28157_n16534));
   NAND3x2_ASAP7_75t_SL U16056 (.Y(n21902),
	.A(FE_OFN26161_sa10_4),
	.B(FE_OFN130_sa10_5),
	.C(FE_OFN27196_n));
   NAND2xp5_ASAP7_75t_L U16057 (.Y(n19646),
	.A(FE_OCPN27636_sa10_4),
	.B(n23996));
   NOR2x1_ASAP7_75t_L U16058 (.Y(n23948),
	.A(n16610),
	.B(n16648));
   NOR2x1_ASAP7_75t_L U16059 (.Y(n21453),
	.A(n18651),
	.B(n17237));
   OAI21xp33_ASAP7_75t_SRAM U16060 (.Y(n18768),
	.A1(FE_PSN8288_n17275),
	.A2(FE_OFN26651_n19573),
	.B(n18766));
   NAND2x1_ASAP7_75t_SL U16061 (.Y(n24085),
	.A(FE_OFN28796_n17301),
	.B(n17245));
   INVxp67_ASAP7_75t_L U16062 (.Y(n19116),
	.A(n17247));
   NAND2x1p5_ASAP7_75t_L U16064 (.Y(n21473),
	.A(FE_OFN26146_n18774),
	.B(n19116));
   NOR3x1_ASAP7_75t_SL U16065 (.Y(n21177),
	.A(n19101),
	.B(n19588),
	.C(n19102));
   NOR2x1_ASAP7_75t_R U16066 (.Y(n19117),
	.A(n17275),
	.B(FE_OCPN27649_n17236));
   NOR2x1_ASAP7_75t_L U16067 (.Y(n22167),
	.A(n22124),
	.B(n19073));
   NOR2xp67_ASAP7_75t_L U16068 (.Y(n20450),
	.A(FE_OFN28790_n),
	.B(FE_OFN25901_n22133));
   NAND2xp33_ASAP7_75t_L U16069 (.Y(n19063),
	.A(FE_OFN28610_n22125),
	.B(n17622));
   NOR2xp33_ASAP7_75t_L U16070 (.Y(n20431),
	.A(FE_OFN28563_n20480),
	.B(n18500));
   NAND2xp33_ASAP7_75t_L U16071 (.Y(n18500),
	.A(n18499),
	.B(n18498));
   NOR2xp67_ASAP7_75t_L U16072 (.Y(n20421),
	.A(n21626),
	.B(FE_OFN29121_n26026));
   NOR2x1_ASAP7_75t_L U16073 (.Y(n19139),
	.A(FE_OCPN27908_FE_OFN16156_sa00_2),
	.B(n21473));
   NOR2x1_ASAP7_75t_L U16074 (.Y(n21444),
	.A(FE_OCPN28250_n19573),
	.B(n19817));
   NAND2x2_ASAP7_75t_SL U16075 (.Y(n17298),
	.A(FE_OCPN29302_sa00_4),
	.B(FE_OCPN27227_sa00_5));
   NOR2x1_ASAP7_75t_L U16077 (.Y(n19106),
	.A(n19097),
	.B(n17300));
   NAND3x1_ASAP7_75t_L U16079 (.Y(n21383),
	.A(FE_OCPN27730_n17464),
	.B(FE_OCPN27903_n19223),
	.C(n17473));
   NOR3xp33_ASAP7_75t_SL U16080 (.Y(n21372),
	.A(FE_OCPN27313_n21845),
	.B(FE_OFN138_sa11_0),
	.C(n17489));
   NAND2xp5_ASAP7_75t_SL U16081 (.Y(n21362),
	.A(n17464),
	.B(n17453));
   NAND2xp33_ASAP7_75t_L U16082 (.Y(n22502),
	.A(n26064),
	.B(n23380));
   NOR2x1_ASAP7_75t_L U16083 (.Y(n23282),
	.A(n23366),
	.B(n21414));
   NAND2xp5_ASAP7_75t_L U16084 (.Y(n21414),
	.A(n21413),
	.B(n23378));
   NAND2xp5_ASAP7_75t_SL U16085 (.Y(n21419),
	.A(n21418),
	.B(FE_OFN16351_n26084));
   NAND2xp5_ASAP7_75t_L U16086 (.Y(n23381),
	.A(n17464),
	.B(FE_OCPN28038_n23252));
   NOR3x1_ASAP7_75t_L U16087 (.Y(n21820),
	.A(FE_OCPN27601_n17475),
	.B(FE_OFN138_sa11_0),
	.C(n17489));
   NOR2xp33_ASAP7_75t_SRAM U16088 (.Y(n23273),
	.A(FE_OCPN27757_n21819),
	.B(n21374));
   NAND3xp33_ASAP7_75t_SL U16090 (.Y(n21396),
	.A(FE_OCPN28038_n23252),
	.B(n17447),
	.C(FE_OFN28915_FE_OCPN27241_sa11_1));
   NOR3x1_ASAP7_75t_SL U16091 (.Y(n17616),
	.A(FE_OFN25901_n22133),
	.B(n17618),
	.C(n18381));
   NOR2xp33_ASAP7_75t_SL U16092 (.Y(n18492),
	.A(n21619),
	.B(n22169));
   NOR3xp33_ASAP7_75t_SL U16093 (.Y(n18506),
	.A(n21625),
	.B(FE_OCPN29400_sa30_3),
	.C(FE_OCPN27971_n21627));
   NOR2x1_ASAP7_75t_L U16094 (.Y(n18483),
	.A(FE_OFN28901_sa30_4),
	.B(FE_OCPN29398_sa30_3));
   NOR3xp33_ASAP7_75t_SL U16095 (.Y(n22162),
	.A(n21625),
	.B(FE_OCPN29413_sa30_5),
	.C(n18381));
   NAND3xp33_ASAP7_75t_R U16096 (.Y(n18489),
	.A(FE_OCPN7643_n17646),
	.B(FE_OFN25917_n21591),
	.C(FE_OCPN29368_FE_OFN16247_sa30_1));
   NAND3xp33_ASAP7_75t_SL U16097 (.Y(n22643),
	.A(FE_OCPN8207_n18497),
	.B(FE_OCPN7643_n17646),
	.C(FE_OCPN29368_FE_OFN16247_sa30_1));
   NOR2xp67_ASAP7_75t_L U16098 (.Y(n21608),
	.A(n20428),
	.B(FE_OFN25901_n22133));
   NOR3xp33_ASAP7_75t_L U16099 (.Y(n20439),
	.A(FE_OCPN27829_n25102),
	.B(FE_OCPN29432_sa30_3),
	.C(FE_OCPN27971_n21627));
   OAI21xp5_ASAP7_75t_SL U16100 (.Y(n21587),
	.A1(n19054),
	.A2(FE_OFN16200_sa30_2),
	.B(n18478));
   NAND3xp33_ASAP7_75t_L U16101 (.Y(n20467),
	.A(FE_OCPN28057_n17603),
	.B(FE_OFN25917_n21591),
	.C(FE_OFN28896_sa30_2));
   NAND2xp5_ASAP7_75t_SL U16102 (.Y(n20466),
	.A(n17650),
	.B(n17649));
   NAND2xp33_ASAP7_75t_SL U16103 (.Y(n17649),
	.A(n18376),
	.B(n17648));
   NAND2xp33_ASAP7_75t_R U16104 (.Y(n17650),
	.A(n18374),
	.B(n17648));
   AND2x2_ASAP7_75t_L U16105 (.Y(n17648),
	.A(n17653),
	.B(n19046));
   NOR2xp33_ASAP7_75t_SL U16107 (.Y(n18481),
	.A(n26023),
	.B(n17651));
   NOR2xp33_ASAP7_75t_SRAM U16108 (.Y(n17651),
	.A(n21604),
	.B(FE_OFN25901_n22133));
   OAI21xp5_ASAP7_75t_SL U16110 (.Y(n18531),
	.A1(n18530),
	.A2(n23711),
	.B(n23752));
   INVx1_ASAP7_75t_SL U16111 (.Y(n18599),
	.A(FE_OCPN27606_n23869));
   NAND2x1p5_ASAP7_75t_SL U16112 (.Y(n23192),
	.A(n24691),
	.B(n18162));
   NAND2xp33_ASAP7_75t_SRAM U16113 (.Y(n23191),
	.A(FE_OFN25952_n22312),
	.B(n21084));
   NOR2x1_ASAP7_75t_SL U16114 (.Y(n22321),
	.A(FE_OFN25987_n23322),
	.B(n18178));
   NOR2xp33_ASAP7_75t_SRAM U16115 (.Y(n20760),
	.A(n23315),
	.B(n21122));
   NOR2x1_ASAP7_75t_L U16116 (.Y(n22862),
	.A(n22278),
	.B(n20722));
   NOR2x1_ASAP7_75t_L U16117 (.Y(n20721),
	.A(n24694),
	.B(n21798));
   NAND2xp5_ASAP7_75t_SL U16118 (.Y(n23195),
	.A(n22842),
	.B(n22841));
   NAND2xp33_ASAP7_75t_L U16119 (.Y(n22842),
	.A(n22837),
	.B(n22839));
   NAND2xp33_ASAP7_75t_R U16120 (.Y(n22841),
	.A(n22840),
	.B(n22839));
   NOR2xp33_ASAP7_75t_SL U16121 (.Y(n22807),
	.A(n18166),
	.B(n18186));
   NOR2x1_ASAP7_75t_SL U16122 (.Y(n22828),
	.A(n21803),
	.B(n20729));
   NAND2xp5_ASAP7_75t_SL U16123 (.Y(n22292),
	.A(n21120),
	.B(n21119));
   NAND2x1_ASAP7_75t_L U16124 (.Y(n22825),
	.A(n23172),
	.B(n22272));
   NAND2xp33_ASAP7_75t_SL U16125 (.Y(n22271),
	.A(FE_OCPN29557_n18161),
	.B(n18159));
   NAND2xp5_ASAP7_75t_SL U16127 (.Y(n21126),
	.A(n18159),
	.B(n23336));
   A2O1A1Ixp33_ASAP7_75t_L U16128 (.Y(n18197),
	.A1(FE_OFN26133_sa22_3),
	.A2(n18159),
	.B(n22305),
	.C(FE_OFN16135_sa22_4));
   NAND2xp5_ASAP7_75t_R U16129 (.Y(n22319),
	.A(n20723),
	.B(n18192));
   NAND2xp33_ASAP7_75t_SRAM U16130 (.Y(n18192),
	.A(FE_OCPN27750_n22293),
	.B(n23336));
   NOR3xp33_ASAP7_75t_SL U16131 (.Y(n21111),
	.A(n21774),
	.B(n21764),
	.C(n18190));
   OAI21xp5_ASAP7_75t_SL U16132 (.Y(n21802),
	.A1(n20729),
	.A2(n23160),
	.B(n18197));
   NAND2xp5_ASAP7_75t_SL U16134 (.Y(n18222),
	.A(n18221),
	.B(FE_OFN29237_n22811));
   NAND2xp5_ASAP7_75t_SL U16135 (.Y(n18223),
	.A(n18219),
	.B(FE_OFN29237_n22811));
   NOR2x1_ASAP7_75t_R U16136 (.Y(n22848),
	.A(FE_OCPN29585_n22281),
	.B(n21779));
   NAND3xp33_ASAP7_75t_SL U16137 (.Y(n21789),
	.A(n21777),
	.B(n21776),
	.C(n21775));
   NOR2xp33_ASAP7_75t_L U16138 (.Y(n21776),
	.A(n21774),
	.B(n21773));
   OAI21xp5_ASAP7_75t_L U16139 (.Y(n21773),
	.A1(n18186),
	.A2(n21772),
	.B(n22801));
   NOR3xp33_ASAP7_75t_R U16141 (.Y(n21258),
	.A(n18606),
	.B(n23719),
	.C(n23739));
   NAND2xp33_ASAP7_75t_R U16142 (.Y(n18606),
	.A(n20674),
	.B(n21667));
   NAND3xp33_ASAP7_75t_SL U16143 (.Y(n23799),
	.A(n21655),
	.B(n25189),
	.C(n21255));
   NOR2xp33_ASAP7_75t_SRAM U16144 (.Y(n21255),
	.A(n23698),
	.B(FE_OCPN28432_n23829));
   NAND2xp5_ASAP7_75t_L U16145 (.Y(n21220),
	.A(n21219),
	.B(n21218));
   NAND2xp33_ASAP7_75t_SL U16146 (.Y(n21221),
	.A(n21216),
	.B(n21218));
   AND2x2_ASAP7_75t_SL U16148 (.Y(n23832),
	.A(n21209),
	.B(n25188));
   NOR3xp33_ASAP7_75t_SL U16149 (.Y(n21209),
	.A(n21208),
	.B(n21648),
	.C(n18548));
   NAND2xp67_ASAP7_75t_L U16150 (.Y(n23726),
	.A(n21655),
	.B(FE_OFN29096_n25188));
   NOR2x1p5_ASAP7_75t_L U16151 (.Y(n21682),
	.A(n23838),
	.B(FE_OCPN28353_n18534));
   NOR3x2_ASAP7_75t_L U16152 (.Y(n21642),
	.A(n20670),
	.B(FE_OCPN27580_n),
	.C(FE_OCPN29563_n18602));
   OAI21xp33_ASAP7_75t_L U16153 (.Y(n23810),
	.A1(n23855),
	.A2(n23840),
	.B(FE_OCPN27580_n));
   NOR2xp33_ASAP7_75t_L U16154 (.Y(n23731),
	.A(n23740),
	.B(n21682));
   OAI222xp33_ASAP7_75t_L U16155 (.Y(n23714),
	.A1(FE_OFN29091_n),
	.A2(n23814),
	.B1(n18532),
	.B2(n23814),
	.C1(FE_OFN29076_n18540),
	.C2(n23814));
   NAND2xp33_ASAP7_75t_L U16156 (.Y(n23709),
	.A(FE_OFN29251_n18536),
	.B(n23855));
   NAND3xp33_ASAP7_75t_SL U16157 (.Y(n23774),
	.A(FE_OCPN29380_sa20_1),
	.B(n18522),
	.C(FE_RN_168_0));
   NAND2xp5_ASAP7_75t_R U16158 (.Y(n23680),
	.A(n25328),
	.B(n21692));
   NOR3xp33_ASAP7_75t_SRAM U16159 (.Y(n23866),
	.A(FE_OFN28815_n18523),
	.B(FE_OFN28791_n),
	.C(n18571));
   NAND3xp33_ASAP7_75t_L U16160 (.Y(n23880),
	.A(n21194),
	.B(FE_OFN28477_n23853),
	.C(n21690));
   NOR2xp33_ASAP7_75t_SL U16163 (.Y(n18424),
	.A(n18430),
	.B(n16936));
   OAI21xp33_ASAP7_75t_R U16164 (.Y(n17425),
	.A1(n16874),
	.A2(n16473),
	.B(n16918));
   NOR3xp33_ASAP7_75t_L U16165 (.Y(n16949),
	.A(FE_OCPN28127_n16872),
	.B(FE_OFN25938_sa33_3),
	.C(FE_OCPN28354_n16677));
   NOR3xp33_ASAP7_75t_SL U16166 (.Y(n18125),
	.A(n16723),
	.B(n23553),
	.C(FE_OFN28918_n16949));
   NAND2xp5_ASAP7_75t_SL U16167 (.Y(n16871),
	.A(n16919),
	.B(n16726));
   NOR3xp33_ASAP7_75t_SRAM U16168 (.Y(n16474),
	.A(FE_OCPN27539_n16875),
	.B(FE_OCPN29391_FE_OFN29162_sa33_2),
	.C(n23556));
   NOR3xp33_ASAP7_75t_SL U16169 (.Y(n23562),
	.A(n16451),
	.B(n16450),
	.C(n18136));
   NAND2xp33_ASAP7_75t_R U16170 (.Y(n16450),
	.A(n16888),
	.B(n16448));
   NOR2xp33_ASAP7_75t_SL U16171 (.Y(n18426),
	.A(n23556),
	.B(n16473));
   NAND2x1_ASAP7_75t_L U16173 (.Y(n16924),
	.A(n16479),
	.B(FE_OFN28998_n16923));
   NAND2x1p5_ASAP7_75t_L U16174 (.Y(n23504),
	.A(FE_OFN29189_sa23_0),
	.B(FE_OCPN27627_sa23_1));
   NOR3xp33_ASAP7_75t_SL U16177 (.Y(n22928),
	.A(n20921),
	.B(n22048),
	.C(n23496));
   OAI21xp33_ASAP7_75t_L U16178 (.Y(n20921),
	.A1(FE_OCPN28363_n22979),
	.A2(FE_OCPN28266_n20920),
	.B(n20919));
   NOR2x1_ASAP7_75t_L U16179 (.Y(n22926),
	.A(n22980),
	.B(FE_OCPN28289_n20235));
   NOR3xp33_ASAP7_75t_SL U16180 (.Y(n20268),
	.A(n20228),
	.B(FE_OFN25890_n23497),
	.C(n20227));
   NAND3xp33_ASAP7_75t_SL U16181 (.Y(n20228),
	.A(n20238),
	.B(n22046),
	.C(n26146));
   NOR2x1_ASAP7_75t_L U16183 (.Y(n20928),
	.A(FE_OCPN28266_n20920),
	.B(FE_OCPN28289_n20235));
   NAND3xp33_ASAP7_75t_R U16184 (.Y(n20941),
	.A(FE_OFN29189_sa23_0),
	.B(n19000),
	.C(FE_OCPN29373_FE_OFN29191_sa23_2));
   NOR2xp33_ASAP7_75t_L U16185 (.Y(n26152),
	.A(n22935),
	.B(n20928));
   NOR3xp33_ASAP7_75t_L U16186 (.Y(n19332),
	.A(n23499),
	.B(n22997),
	.C(n22930));
   NOR2x1_ASAP7_75t_SL U16187 (.Y(n22048),
	.A(FE_OCPN27954_n22945),
	.B(n22952));
   NOR3xp33_ASAP7_75t_L U16188 (.Y(n22043),
	.A(n19330),
	.B(n20270),
	.C(n22003));
   NOR2x1_ASAP7_75t_L U16189 (.Y(n22930),
	.A(n22952),
	.B(FE_OFN25889_n20913));
   NOR3x1_ASAP7_75t_L U16190 (.Y(n23499),
	.A(FE_OCPN27710_n19011),
	.B(FE_OCPN27881_FE_OFN27126_sa23_3),
	.C(FE_OCPN27954_n22945));
   NOR2xp33_ASAP7_75t_L U16191 (.Y(n22039),
	.A(n22926),
	.B(n20265));
   NAND3x1_ASAP7_75t_SL U16193 (.Y(n26556),
	.A(FE_OCPN27986_n18970),
	.B(n19000),
	.C(FE_OFN29191_sa23_2));
   NAND2xp5_ASAP7_75t_SL U16194 (.Y(n20238),
	.A(n19019),
	.B(n19000));
   NAND2xp5_ASAP7_75t_SL U16196 (.Y(n22996),
	.A(n23480),
	.B(FE_OCPN28098_n20907));
   NOR2x1_ASAP7_75t_SL U16197 (.Y(n26660),
	.A(FE_OFN27127_sa23_3),
	.B(n18989));
   NAND2x2_ASAP7_75t_SL U16198 (.Y(n22980),
	.A(FE_OCPN27482_sa23_5),
	.B(n20933));
   NOR2x1_ASAP7_75t_SL U16199 (.Y(n23517),
	.A(n22993),
	.B(n22992));
   NAND2x1p5_ASAP7_75t_SL U16200 (.Y(n22971),
	.A(FE_OCPN29489_sa23_3),
	.B(FE_OFN27078_sa23_5));
   NAND2xp5_ASAP7_75t_L U16201 (.Y(n22973),
	.A(n23513),
	.B(n22030));
   NAND2xp5_ASAP7_75t_L U16202 (.Y(n18716),
	.A(n17331),
	.B(n23059));
   NAND2xp5_ASAP7_75t_L U16203 (.Y(n22435),
	.A(n18716),
	.B(FE_OFN27150_n22175));
   NOR2xp67_ASAP7_75t_R U16204 (.Y(n21560),
	.A(FE_OFN26648_n22197),
	.B(n17330));
   NOR2xp67_ASAP7_75t_SL U16207 (.Y(n23075),
	.A(n23107),
	.B(FE_OFN27052_n21551));
   NAND2xp33_ASAP7_75t_R U16208 (.Y(n18723),
	.A(n22191),
	.B(n22183));
   NAND2xp5_ASAP7_75t_L U16209 (.Y(n23074),
	.A(n20394),
	.B(n20393));
   NAND2xp5_ASAP7_75t_L U16210 (.Y(n20393),
	.A(n20392),
	.B(FE_OCPN27433_n21571));
   NAND2xp33_ASAP7_75t_L U16211 (.Y(n20394),
	.A(n20390),
	.B(FE_OCPN27433_n21571));
   NAND2xp5_ASAP7_75t_R U16212 (.Y(n23094),
	.A(n22422),
	.B(n22421));
   OAI21x1_ASAP7_75t_SL U16213 (.Y(n20365),
	.A1(n23107),
	.A2(n17318),
	.B(n17375));
   NOR2xp33_ASAP7_75t_SL U16214 (.Y(n20401),
	.A(FE_OCPN27423_sa01_0),
	.B(n18709));
   NAND2xp33_ASAP7_75t_R U16215 (.Y(n18709),
	.A(FE_OFN29135_n21551),
	.B(n18708));
   NAND3x1_ASAP7_75t_L U16217 (.Y(n22451),
	.A(n18721),
	.B(n17369),
	.C(n22415));
   NAND2xp5_ASAP7_75t_L U16218 (.Y(n22583),
	.A(n20368),
	.B(n18727));
   NOR2xp33_ASAP7_75t_L U16220 (.Y(n22467),
	.A(n22177),
	.B(FE_OCPN8236_n22438));
   NAND2xp33_ASAP7_75t_L U16221 (.Y(n23083),
	.A(n23103),
	.B(n22468));
   NOR3xp33_ASAP7_75t_SRAM U16222 (.Y(n22753),
	.A(n19527),
	.B(FE_OCPN29493_sa12_4),
	.C(n19526));
   NAND3xp33_ASAP7_75t_SRAM U16224 (.Y(n23613),
	.A(FE_OCPN28198_n22776),
	.B(FE_OCPN8265_n24362),
	.C(FE_OFN25907_sa12_2));
   NOR2x1_ASAP7_75t_L U16225 (.Y(n23602),
	.A(n23217),
	.B(FE_OFN26158_n22224));
   NAND2xp5_ASAP7_75t_SL U16226 (.Y(n19540),
	.A(n17973),
	.B(n17972));
   NOR2xp33_ASAP7_75t_L U16228 (.Y(n17973),
	.A(n17970),
	.B(FE_OCPN27888_sa12_2));
   NOR2xp33_ASAP7_75t_L U16229 (.Y(n23242),
	.A(n22724),
	.B(n22723));
   OAI21xp33_ASAP7_75t_SRAM U16230 (.Y(n22723),
	.A1(n22722),
	.A2(FE_OFN27070_n),
	.B(n23612));
   NOR3xp33_ASAP7_75t_L U16231 (.Y(n22261),
	.A(n20559),
	.B(n25439),
	.C(n22718));
   NOR3xp33_ASAP7_75t_L U16232 (.Y(n22764),
	.A(n22240),
	.B(n22239),
	.C(n22238));
   OAI21xp33_ASAP7_75t_SRAM U16233 (.Y(n22240),
	.A1(FE_OCPN29492_sa12_4),
	.A2(n22237),
	.B(n22236));
   OAI222xp33_ASAP7_75t_R U16234 (.Y(n22762),
	.A1(FE_OFN25907_sa12_2),
	.A2(n22235),
	.B1(FE_OFN28882_FE_OCPN27356_sa12_0),
	.B2(n22235),
	.C1(FE_OFN28739_n17898),
	.C2(n22235));
   NAND3xp33_ASAP7_75t_SL U16235 (.Y(n19512),
	.A(FE_OFN28882_FE_OCPN27356_sa12_0),
	.B(n23600),
	.C(FE_OFN28764_n17928));
   NAND3xp33_ASAP7_75t_SL U16236 (.Y(n22226),
	.A(n17906),
	.B(FE_OCPN28386_n17899),
	.C(FE_OCPN27429_sa12_3));
   NOR3x1_ASAP7_75t_R U16237 (.Y(n20596),
	.A(n19527),
	.B(FE_OCPN29494_sa12_4),
	.C(n17949));
   NAND2xp5_ASAP7_75t_L U16238 (.Y(n23596),
	.A(FE_OFN28834_FE_OCPN28371_n17900),
	.B(n20796));
   NAND3x1_ASAP7_75t_L U16239 (.Y(n23609),
	.A(FE_OCPN5137_n23600),
	.B(FE_OCPN28386_n17899),
	.C(FE_OFN28764_n17928));
   NOR3xp33_ASAP7_75t_SL U16240 (.Y(n22225),
	.A(n20784),
	.B(n22750),
	.C(n23602));
   NAND2xp5_ASAP7_75t_SL U16241 (.Y(n22228),
	.A(n25741),
	.B(n20796));
   NAND3xp33_ASAP7_75t_R U16242 (.Y(n27091),
	.A(n19425),
	.B(n19424),
	.C(n19423));
   NAND2xp5_ASAP7_75t_SL U16243 (.Y(n27088),
	.A(n17169),
	.B(n17168));
   NAND2xp33_ASAP7_75t_SL U16244 (.Y(n17168),
	.A(n17167),
	.B(n17166));
   NAND2xp33_ASAP7_75t_L U16245 (.Y(n17169),
	.A(n17164),
	.B(n17166));
   NAND3x1_ASAP7_75t_SL U16247 (.Y(n18335),
	.A(n19911),
	.B(n19940),
	.C(FE_OCPN29404_FE_OFN27148_sa32_3));
   NAND2xp5_ASAP7_75t_L U16249 (.Y(n18307),
	.A(n19934),
	.B(n24988));
   NOR2xp67_ASAP7_75t_R U16250 (.Y(n20106),
	.A(FE_OCPN27267_n18794),
	.B(FE_OFN26577_n));
   NOR2xp67_ASAP7_75t_L U16251 (.Y(n18799),
	.A(n17564),
	.B(n18832));
   NOR3x1_ASAP7_75t_L U16253 (.Y(n19712),
	.A(n17591),
	.B(FE_OCPN29405_FE_OFN27148_sa32_3),
	.C(FE_OCPN29459_n));
   NAND2xp5_ASAP7_75t_L U16254 (.Y(n18329),
	.A(n17525),
	.B(FE_OCPN29524_n25029));
   NAND2xp5_ASAP7_75t_L U16255 (.Y(n17704),
	.A(n24861),
	.B(n25025));
   NOR3x1_ASAP7_75t_L U16256 (.Y(n22395),
	.A(n18334),
	.B(FE_OCPN27792_n18333),
	.C(n18332));
   NAND2xp5_ASAP7_75t_R U16257 (.Y(n18334),
	.A(n18330),
	.B(n18329));
   OAI21xp33_ASAP7_75t_L U16258 (.Y(n18332),
	.A1(FE_OCPN27267_n18794),
	.A2(n18836),
	.B(n18331));
   NAND2xp33_ASAP7_75t_SRAM U16259 (.Y(n18331),
	.A(FE_OCPN28229_n17529),
	.B(n22392));
   NAND2xp5_ASAP7_75t_L U16260 (.Y(n17697),
	.A(FE_OCPN28229_n17529),
	.B(n17560));
   NAND2xp5_ASAP7_75t_L U16261 (.Y(n18309),
	.A(n18298),
	.B(n22392));
   NOR2xp33_ASAP7_75t_L U16262 (.Y(n17711),
	.A(n19710),
	.B(n22399));
   NAND2xp5_ASAP7_75t_R U16263 (.Y(n20117),
	.A(n17560),
	.B(n17690));
   OAI21xp33_ASAP7_75t_SRAM U16264 (.Y(n17690),
	.A1(FE_OFN28686_FE_OCPN27812),
	.A2(FE_OFN26035_n),
	.B(FE_OCPN27882_n18829));
   NAND2x1_ASAP7_75t_L U16265 (.Y(n18839),
	.A(n17560),
	.B(n18799));
   NOR2x1_ASAP7_75t_SL U16266 (.Y(n19728),
	.A(FE_OCPN29420_FE_OFN16128_sa32_2),
	.B(n18826));
   NAND2xp5_ASAP7_75t_L U16267 (.Y(n18299),
	.A(n22392),
	.B(n19940));
   OAI22xp5_ASAP7_75t_L U16268 (.Y(n20303),
	.A1(FE_OCPN28298_n),
	.A2(FE_OCPN27454_n16789),
	.B1(FE_OCPN27642_n16758),
	.B2(FE_OCPN27454_n16789));
   NAND2xp5_ASAP7_75t_SL U16269 (.Y(n20009),
	.A(FE_OCPN29265_FE_OFN28698_sa21_1),
	.B(n22694));
   NAND3xp33_ASAP7_75t_L U16270 (.Y(n20332),
	.A(FE_OFN28779_n24257),
	.B(FE_OFN16153_n16747),
	.C(FE_OCPN5126_sa21_2));
   NOR2x1_ASAP7_75t_L U16271 (.Y(n19890),
	.A(n16762),
	.B(n23633));
   NAND2xp5_ASAP7_75t_L U16272 (.Y(n17856),
	.A(n22353),
	.B(n19974));
   NAND3xp33_ASAP7_75t_L U16273 (.Y(n20299),
	.A(FE_OCPN27616_n16760),
	.B(FE_OFN16447_n16749),
	.C(FE_OCPN29265_FE_OFN28698_sa21_1));
   NOR3x1_ASAP7_75t_L U16275 (.Y(n23643),
	.A(n17860),
	.B(FE_OFN28903_sa21_0),
	.C(n17881));
   NAND3x1_ASAP7_75t_L U16276 (.Y(n23628),
	.A(FE_OCPN29293_FE_OFN28678_sa21_3),
	.B(n16760),
	.C(FE_OCPN29265_FE_OFN28698_sa21_1));
   NOR3x1_ASAP7_75t_SL U16277 (.Y(n25353),
	.A(n19982),
	.B(FE_OCPN29293_FE_OFN28678_sa21_3),
	.C(FE_OCPN28187_n16806));
   NOR2x1_ASAP7_75t_SL U16278 (.Y(n21989),
	.A(FE_OCPN29482_FE_OFN26014_sa31_3),
	.B(n16340));
   NOR3x1_ASAP7_75t_SL U16279 (.Y(n21984),
	.A(n20024),
	.B(n20023),
	.C(FE_OFN26550_n16331));
   NAND3xp33_ASAP7_75t_L U16280 (.Y(n16519),
	.A(n16300),
	.B(n16512),
	.C(FE_OFN26060_sa31_4));
   NOR3xp33_ASAP7_75t_L U16281 (.Y(n21975),
	.A(n20057),
	.B(n20056),
	.C(n20055));
   NAND2xp33_ASAP7_75t_SRAM U16282 (.Y(n20055),
	.A(n20856),
	.B(n20054));
   NOR3xp33_ASAP7_75t_L U16283 (.Y(n20837),
	.A(n20854),
	.B(FE_OCPN29482_FE_OFN26014_sa31_3),
	.C(n16340));
   OAI21xp33_ASAP7_75t_L U16284 (.Y(n21944),
	.A1(FE_OCPN28008_n16290),
	.A2(n20074),
	.B(n20065));
   NOR2xp33_ASAP7_75t_L U16285 (.Y(n21946),
	.A(FE_OFN26629_sa31_4),
	.B(FE_OFN26015_sa31_3));
   NAND2x1_ASAP7_75t_L U16288 (.Y(n16407),
	.A(FE_OCPN27516_n26292),
	.B(n20050));
   NOR2x1_ASAP7_75t_SL U16289 (.Y(n20840),
	.A(FE_OFN26095_n16293),
	.B(n18093));
   NAND3x1_ASAP7_75t_L U16290 (.Y(n20832),
	.A(n16295),
	.B(n20050),
	.C(FE_OFN16415_sa31_2));
   OAI22xp33_ASAP7_75t_L U16292 (.Y(n20070),
	.A1(FE_OCPN28008_n16290),
	.A2(FE_OFN29117_n),
	.B1(n16408),
	.B2(FE_OFN29117_n));
   NAND2xp5_ASAP7_75t_L U16293 (.Y(n16335),
	.A(FE_OFN28669_sa31_5),
	.B(n18073));
   NAND2xp5_ASAP7_75t_L U16294 (.Y(n20874),
	.A(FE_OCPN29483_FE_OFN26014_sa31_3),
	.B(n16507));
   NAND3xp33_ASAP7_75t_L U16295 (.Y(n20034),
	.A(n20050),
	.B(n20060),
	.C(FE_OFN26095_n16293));
   NAND2xp5_ASAP7_75t_L U16296 (.Y(n20052),
	.A(FE_OFN29016_n16512),
	.B(n16299));
   NAND2xp33_ASAP7_75t_SRAM U16297 (.Y(n21940),
	.A(n24181),
	.B(FE_OFN26015_sa31_3));
   OAI22xp33_ASAP7_75t_R U16298 (.Y(n19919),
	.A1(FE_OCPN27882_n18829),
	.A2(n18828),
	.B1(n18827),
	.B2(n18828));
   NAND2x1_ASAP7_75t_SL U16299 (.Y(n20093),
	.A(n18324),
	.B(n17527));
   NOR2x1p5_ASAP7_75t_SL U16300 (.Y(n19907),
	.A(FE_OCPN29421_FE_OFN16128_sa32_2),
	.B(n18306));
   NOR2x1_ASAP7_75t_L U16301 (.Y(n22399),
	.A(FE_OCPN27420_n18794),
	.B(n17591));
   NAND2xp5_ASAP7_75t_R U16302 (.Y(n25196),
	.A(n17039),
	.B(n17038));
   NAND2xp33_ASAP7_75t_L U16303 (.Y(n17038),
	.A(n17037),
	.B(n17036));
   NAND2xp33_ASAP7_75t_L U16304 (.Y(n17039),
	.A(n17035),
	.B(n17036));
   NOR2x1_ASAP7_75t_L U16306 (.Y(n21986),
	.A(n18096),
	.B(n20837));
   NAND2xp5_ASAP7_75t_R U16307 (.Y(n18063),
	.A(FE_OCPN27877_n21980),
	.B(FE_OFN29016_n16512));
   NAND2xp33_ASAP7_75t_L U16308 (.Y(n18065),
	.A(n20838),
	.B(n20052));
   NOR2x1_ASAP7_75t_SL U16310 (.Y(n26154),
	.A(FE_OCPN27916_n),
	.B(n22969));
   NOR3xp33_ASAP7_75t_L U16311 (.Y(n25601),
	.A(n24476),
	.B(n24475),
	.C(n24474));
   NOR2xp33_ASAP7_75t_SRAM U16313 (.Y(n15986),
	.A(FE_OFN28715_w3_15),
	.B(FE_OCPN29520_n24755));
   NAND2xp5_ASAP7_75t_L U16315 (.Y(n14915),
	.A(n16000),
	.B(n15959));
   NAND2xp33_ASAP7_75t_SRAM U16316 (.Y(n14907),
	.A(n15434),
	.B(n14919));
   NAND2x1_ASAP7_75t_L U16317 (.Y(n15876),
	.A(FE_OFN28747_n),
	.B(FE_OFN16195_n13771));
   NOR3xp33_ASAP7_75t_SRAM U16318 (.Y(n15449),
	.A(n15987),
	.B(FE_OFN26642_w3_14),
	.C(FE_OCPN29570_n15423));
   OA222x2_ASAP7_75t_R U16319 (.Y(n14875),
	.A1(n14862),
	.A2(FE_OFN28682_n15888),
	.B1(n14861),
	.B2(FE_OFN28682_n15888),
	.C1(n14880),
	.C2(FE_OFN28682_n15888));
   NAND3xp33_ASAP7_75t_SRAM U16320 (.Y(n14861),
	.A(FE_OFN26073_n),
	.B(n15610),
	.C(n15857));
   NAND2xp33_ASAP7_75t_L U16321 (.Y(n14862),
	.A(n14854),
	.B(n14853));
   NAND2xp33_ASAP7_75t_L U16322 (.Y(n14853),
	.A(n15802),
	.B(n14890));
   O2A1O1Ixp5_ASAP7_75t_SRAM U16323 (.Y(n14890),
	.A1(FE_OFN28747_n),
	.A2(FE_OFN26532_n13766),
	.B(n15859),
	.C(n14852));
   NOR2xp33_ASAP7_75t_L U16324 (.Y(n14852),
	.A(FE_OFN16195_n13771),
	.B(n15825));
   NAND2xp5_ASAP7_75t_L U16325 (.Y(n14844),
	.A(n14449),
	.B(n14985));
   NOR2xp33_ASAP7_75t_R U16326 (.Y(n15298),
	.A(n14778),
	.B(n15480));
   OAI21xp33_ASAP7_75t_R U16327 (.Y(n13670),
	.A1(FE_OFN27208_w3_30),
	.A2(FE_OCPN27655_w3_25),
	.B(n25675));
   NAND2xp5_ASAP7_75t_SL U16328 (.Y(n15959),
	.A(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(FE_OFN26635_w3_14));
   NAND3xp33_ASAP7_75t_SRAM U16329 (.Y(n14896),
	.A(FE_OFN27115_n),
	.B(n15986),
	.C(FE_OFN26633_w3_14));
   NOR2xp33_ASAP7_75t_SL U16330 (.Y(n14897),
	.A(FE_OFN27115_n),
	.B(FE_OFN26635_w3_14));
   NAND3xp33_ASAP7_75t_SL U16331 (.Y(n15376),
	.A(FE_OCPN29427_w3_15),
	.B(n24755),
	.C(FE_OFN26162_w3_13));
   NAND3xp33_ASAP7_75t_L U16332 (.Y(n15180),
	.A(FE_OCPN29428_FE_OFN27131_w3_29),
	.B(FE_OFN28571_w3_28),
	.C(FE_OCPN28096_w3_31));
   NOR2x1p5_ASAP7_75t_L U16333 (.Y(n15859),
	.A(FE_OFN28662_w3_7),
	.B(n13726));
   NOR3xp33_ASAP7_75t_R U16334 (.Y(n15577),
	.A(n13730),
	.B(FE_OFN28662_w3_7),
	.C(n15061));
   NAND3xp33_ASAP7_75t_SL U16335 (.Y(n16010),
	.A(n24755),
	.B(n25782),
	.C(FE_OFN27200_n));
   NOR3x1_ASAP7_75t_L U16336 (.Y(n15422),
	.A(n24755),
	.B(FE_OFN26162_w3_13),
	.C(FE_OCPN29427_w3_15));
   OAI21xp33_ASAP7_75t_L U16337 (.Y(n13713),
	.A1(n25675),
	.A2(w3_25_),
	.B(FE_OFN27206_w3_30));
   NOR3x1_ASAP7_75t_SL U16339 (.Y(n14996),
	.A(FE_OFN25886_w3_3),
	.B(FE_OCPN27985_n24831),
	.C(FE_OFN26531_n));
   NAND3xp33_ASAP7_75t_R U16341 (.Y(n24550),
	.A(n24549),
	.B(n24548),
	.C(n24547));
   NOR3xp33_ASAP7_75t_L U16342 (.Y(n24549),
	.A(n24546),
	.B(n24545),
	.C(n24544));
   NAND2xp33_ASAP7_75t_L U16343 (.Y(n24224),
	.A(n24220),
	.B(n24219));
   NAND3xp33_ASAP7_75t_SRAM U16344 (.Y(n25796),
	.A(n25795),
	.B(n25794),
	.C(n25793));
   NAND2xp33_ASAP7_75t_R U16345 (.Y(n25791),
	.A(n25790),
	.B(n25789));
   NOR3xp33_ASAP7_75t_SL U16347 (.Y(n24020),
	.A(FE_OCPN27226_n25357),
	.B(n24021),
	.C(n24659));
   NAND3xp33_ASAP7_75t_SRAM U16348 (.Y(n24922),
	.A(n24921),
	.B(n23630),
	.C(n24920));
   NAND2xp5_ASAP7_75t_L U16349 (.Y(n25709),
	.A(n26679),
	.B(n25694));
   NOR2xp33_ASAP7_75t_SL U16350 (.Y(n25700),
	.A(FE_OCPN29532_n25697),
	.B(FE_OCPN27507_n25695));
   O2A1O1Ixp33_ASAP7_75t_SL U16351 (.Y(n25699),
	.A1(n27027),
	.A2(n25701),
	.B(n25698),
	.C(n25697));
   NOR3xp33_ASAP7_75t_L U16352 (.Y(n19209),
	.A(FE_OFN28630_n23385),
	.B(n21385),
	.C(n19208));
   NOR3xp33_ASAP7_75t_L U16353 (.Y(n24570),
	.A(n19169),
	.B(n19168),
	.C(n19167));
   OAI21xp33_ASAP7_75t_SRAM U16354 (.Y(n19169),
	.A1(FE_OFN28874_FE_OCPN27551_sa11_4),
	.A2(FE_OFN29033_FE_OCPN27414_n23359),
	.B(n22495));
   OAI21xp33_ASAP7_75t_SRAM U16355 (.Y(n19167),
	.A1(n19166),
	.A2(FE_OCPN27757_n21819),
	.B(n23372));
   NAND2xp33_ASAP7_75t_L U16356 (.Y(n19168),
	.A(n23387),
	.B(n19165));
   OAI222xp33_ASAP7_75t_R U16357 (.Y(n25818),
	.A1(FE_OFN28669_sa31_5),
	.A2(n18070),
	.B1(FE_OCPN27516_n26292),
	.B2(n18070),
	.C1(FE_OCPN29483_FE_OFN26014_sa31_3),
	.C2(n18070));
   NAND3xp33_ASAP7_75t_L U16358 (.Y(n18070),
	.A(n18069),
	.B(n21979),
	.C(n18068));
   NOR3xp33_ASAP7_75t_R U16359 (.Y(n25817),
	.A(n18091),
	.B(n18076),
	.C(n18084));
   NOR3xp33_ASAP7_75t_L U16361 (.Y(n18092),
	.A(n18090),
	.B(n18089),
	.C(n18088));
   NAND3xp33_ASAP7_75t_L U16362 (.Y(n18089),
	.A(n18087),
	.B(n24182),
	.C(n18086));
   NOR3xp33_ASAP7_75t_L U16363 (.Y(n18099),
	.A(n18097),
	.B(n18096),
	.C(n18095));
   NOR2x1_ASAP7_75t_L U16364 (.Y(n19056),
	.A(n18373),
	.B(n17616));
   NOR3xp33_ASAP7_75t_SL U16366 (.Y(n22625),
	.A(n17612),
	.B(n18387),
	.C(n17611));
   NAND2xp33_ASAP7_75t_SRAM U16367 (.Y(n17611),
	.A(FE_OCPN28241_n22142),
	.B(n17619));
   NOR2x1_ASAP7_75t_L U16368 (.Y(n22628),
	.A(FE_OFN26597_n),
	.B(FE_OFN28790_n));
   NAND2xp5_ASAP7_75t_L U16369 (.Y(n23352),
	.A(n23319),
	.B(n23318));
   NAND2xp33_ASAP7_75t_R U16370 (.Y(n23318),
	.A(n23317),
	.B(n23316));
   NAND2xp33_ASAP7_75t_R U16371 (.Y(n23319),
	.A(n23313),
	.B(n23316));
   NOR3xp33_ASAP7_75t_R U16372 (.Y(n24483),
	.A(n16426),
	.B(n23553),
	.C(n16912));
   NOR3x1_ASAP7_75t_L U16373 (.Y(n24489),
	.A(FE_OFN29005_n23558),
	.B(n24297),
	.C(n17424));
   NOR2xp33_ASAP7_75t_SL U16374 (.Y(n18418),
	.A(n16442),
	.B(n16441));
   OAI22xp33_ASAP7_75t_SL U16375 (.Y(n16437),
	.A1(FE_OFN28999_n16923),
	.A2(n16937),
	.B1(FE_OFN29101_n16418),
	.B2(n16937));
   NAND3x1_ASAP7_75t_SL U16376 (.Y(n22378),
	.A(FE_OCPN28268_n19911),
	.B(n17527),
	.C(FE_OCPN27230_sa32_3));
   NAND2xp5_ASAP7_75t_SL U16378 (.Y(n17716),
	.A(n18335),
	.B(n22386));
   NAND2xp33_ASAP7_75t_L U16379 (.Y(n17722),
	.A(n18306),
	.B(n19951));
   NAND3xp33_ASAP7_75t_SRAM U16380 (.Y(n17727),
	.A(n18843),
	.B(n18825),
	.C(n18813));
   NAND2xp33_ASAP7_75t_SL U16381 (.Y(n17047),
	.A(n18268),
	.B(n18242));
   NOR3x2_ASAP7_75t_SL U16382 (.Y(n19379),
	.A(FE_OFN28738_n16989),
	.B(FE_OCPN29543_FE_OFN28862_n),
	.C(FE_OCPN28149_n17121));
   NAND2xp33_ASAP7_75t_SL U16383 (.Y(n19950),
	.A(n19700),
	.B(n19699));
   NOR3xp33_ASAP7_75t_SL U16384 (.Y(n19699),
	.A(n19698),
	.B(n22399),
	.C(n19908));
   NAND2xp5_ASAP7_75t_R U16385 (.Y(n19697),
	.A(n18298),
	.B(n18324));
   OAI22xp33_ASAP7_75t_SRAM U16386 (.Y(n22393),
	.A1(FE_OCPN28229_n17529),
	.A2(n20095),
	.B1(FE_OCPN28268_n19911),
	.B2(n20095));
   NAND2xp5_ASAP7_75t_SL U16387 (.Y(n24872),
	.A(n19940),
	.B(FE_OCPN28434_n17546));
   NAND2xp33_ASAP7_75t_L U16388 (.Y(n24854),
	.A(n19708),
	.B(n19707));
   NAND2xp33_ASAP7_75t_R U16389 (.Y(n19707),
	.A(n19706),
	.B(FE_OFN16402_n19704));
   NOR3xp33_ASAP7_75t_SL U16390 (.Y(n24216),
	.A(n20902),
	.B(n20901),
	.C(n20900));
   NAND2xp33_ASAP7_75t_SRAM U16391 (.Y(n20900),
	.A(n20899),
	.B(n26162));
   NOR3xp33_ASAP7_75t_R U16392 (.Y(n24040),
	.A(n19295),
	.B(n19294),
	.C(n20942));
   NAND2xp33_ASAP7_75t_L U16393 (.Y(n19295),
	.A(n19293),
	.B(n22986));
   NAND2xp33_ASAP7_75t_L U16394 (.Y(n19293),
	.A(n19292),
	.B(n19291));
   NOR3xp33_ASAP7_75t_SL U16395 (.Y(n22024),
	.A(n22979),
	.B(FE_OCPN29441_sa23_4),
	.C(n22971));
   NOR2xp33_ASAP7_75t_L U16396 (.Y(n22269),
	.A(n21786),
	.B(n23164));
   NOR2xp33_ASAP7_75t_SRAM U16397 (.Y(n21786),
	.A(n18186),
	.B(n21785));
   NAND2xp33_ASAP7_75t_L U16398 (.Y(n22273),
	.A(n22311),
	.B(n21118));
   NOR2xp33_ASAP7_75t_SL U16399 (.Y(n19754),
	.A(n21902),
	.B(n16564));
   AND3x1_ASAP7_75t_L U16400 (.Y(n20649),
	.A(n20647),
	.B(n23793),
	.C(n20646));
   NAND2xp33_ASAP7_75t_SRAM U16401 (.Y(n20632),
	.A(n21692),
	.B(n21684));
   NOR3xp33_ASAP7_75t_SL U16402 (.Y(n22182),
	.A(n22205),
	.B(n23076),
	.C(n17383));
   NAND2xp5_ASAP7_75t_SL U16403 (.Y(n20377),
	.A(n22428),
	.B(n20376));
   NOR3xp33_ASAP7_75t_R U16404 (.Y(n20376),
	.A(n22438),
	.B(n22447),
	.C(n20387));
   NAND2xp33_ASAP7_75t_L U16405 (.Y(n21538),
	.A(n21535),
	.B(n21534));
   NOR2x1p5_ASAP7_75t_L U16406 (.Y(n21147),
	.A(FE_OFN29079_FE_OCPN27518_n17251),
	.B(FE_OCPN28270_n17237));
   NAND2xp5_ASAP7_75t_R U16407 (.Y(n27037),
	.A(n18619),
	.B(n18618));
   NAND2xp33_ASAP7_75t_SRAM U16408 (.Y(n18618),
	.A(n18617),
	.B(n18616));
   NAND2xp33_ASAP7_75t_SRAM U16409 (.Y(n18619),
	.A(n18615),
	.B(n18616));
   NOR3xp33_ASAP7_75t_L U16411 (.Y(n25637),
	.A(FE_PSN8305_n21217),
	.B(n23866),
	.C(n23719));
   NOR3xp33_ASAP7_75t_R U16412 (.Y(n20603),
	.A(n20813),
	.B(n22730),
	.C(n22242));
   NOR3x1_ASAP7_75t_L U16413 (.Y(n21750),
	.A(n23432),
	.B(FE_OFN28614_n21715),
	.C(n21297));
   NAND3xp33_ASAP7_75t_L U16415 (.Y(n23474),
	.A(n25090),
	.B(n20904),
	.C(n23501));
   NOR2xp33_ASAP7_75t_L U16416 (.Y(n23475),
	.A(n20928),
	.B(n20927));
   NAND3xp33_ASAP7_75t_L U16417 (.Y(n20927),
	.A(n22941),
	.B(n26146),
	.C(n20926));
   NOR2xp67_ASAP7_75t_L U16418 (.Y(n26402),
	.A(FE_OFN29117_n),
	.B(FE_OCPN7597_n21981));
   NOR2xp33_ASAP7_75t_SRAM U16419 (.Y(n20040),
	.A(n26292),
	.B(n21968));
   NAND3xp33_ASAP7_75t_R U16420 (.Y(n19373),
	.A(n19372),
	.B(n25994),
	.C(n25880));
   NAND2xp5_ASAP7_75t_L U16421 (.Y(n18924),
	.A(FE_OFN29173_n),
	.B(n24156));
   NOR3xp33_ASAP7_75t_L U16422 (.Y(n20116),
	.A(FE_OFN28552_n20105),
	.B(n20104),
	.C(n20103));
   NOR3xp33_ASAP7_75t_L U16423 (.Y(n26001),
	.A(FE_OCPN8231_n20522),
	.B(n19380),
	.C(n19379));
   NAND2xp5_ASAP7_75t_L U16424 (.Y(n18944),
	.A(n18938),
	.B(n18937));
   NAND2xp33_ASAP7_75t_L U16425 (.Y(n18938),
	.A(n18934),
	.B(FE_OFN25999_n25875));
   NAND2x1_ASAP7_75t_SL U16426 (.Y(n22075),
	.A(FE_OCPN27570_n17791),
	.B(n17741));
   NOR2xp33_ASAP7_75t_R U16427 (.Y(n17741),
	.A(FE_OCPN27273_sa02_3),
	.B(n17740));
   NOR2xp33_ASAP7_75t_SRAM U16428 (.Y(n18862),
	.A(FE_OCPN29327_n21017),
	.B(n21715));
   NOR2x1_ASAP7_75t_SL U16429 (.Y(n21521),
	.A(n18873),
	.B(n18872));
   NAND2xp5_ASAP7_75t_L U16430 (.Y(n18872),
	.A(n21711),
	.B(n18051));
   NAND3xp33_ASAP7_75t_L U16431 (.Y(n18873),
	.A(n21719),
	.B(FE_OFN16294_n19461),
	.C(n21071));
   NOR3xp33_ASAP7_75t_SL U16432 (.Y(n23946),
	.A(n18027),
	.B(FE_OCPN5140_n21049),
	.C(n21503));
   NOR3xp33_ASAP7_75t_SRAM U16435 (.Y(n25503),
	.A(n22873),
	.B(n22872),
	.C(n22871));
   INVxp67_ASAP7_75t_SL U16436 (.Y(n22883),
	.A(n22879));
   OAI21xp33_ASAP7_75t_SRAM U16437 (.Y(n21880),
	.A1(n16542),
	.A2(n23132),
	.B(n24944));
   NOR3xp33_ASAP7_75t_SRAM U16440 (.Y(n24345),
	.A(n21148),
	.B(n21147),
	.C(n17297));
   NOR3xp33_ASAP7_75t_L U16441 (.Y(n21495),
	.A(n19576),
	.B(n19575),
	.C(n21452));
   NOR3xp33_ASAP7_75t_SRAM U16442 (.Y(n17296),
	.A(n19836),
	.B(n19090),
	.C(n19813));
   NAND2xp5_ASAP7_75t_L U16443 (.Y(n19089),
	.A(n19811),
	.B(n24085));
   NOR3x1_ASAP7_75t_L U16444 (.Y(n19122),
	.A(n17298),
	.B(FE_OCPN29396_n19149),
	.C(FE_OCPN29370_FE_OFN28744));
   NOR2xp33_ASAP7_75t_SRAM U16445 (.Y(n17104),
	.A(n17103),
	.B(FE_OCPN28202_n16991));
   NAND2xp33_ASAP7_75t_L U16446 (.Y(n20953),
	.A(n20170),
	.B(FE_OCPN27634_n20169));
   NAND3xp33_ASAP7_75t_L U16447 (.Y(n22874),
	.A(n20188),
	.B(n20187),
	.C(n25274));
   OAI21xp5_ASAP7_75t_SL U16448 (.Y(n25298),
	.A1(FE_OFN26159_n22080),
	.A2(n22103),
	.B(n22106));
   NOR2xp33_ASAP7_75t_SL U16449 (.Y(n17764),
	.A(n25202),
	.B(n17762));
   NAND3x1_ASAP7_75t_SL U16450 (.Y(n22114),
	.A(n22104),
	.B(n22103),
	.C(n22102));
   NOR2x1_ASAP7_75t_L U16451 (.Y(n20502),
	.A(n17042),
	.B(FE_OCPN29446_n17115));
   NOR2x1_ASAP7_75t_SL U16453 (.Y(n21888),
	.A(n21902),
	.B(n23036));
   NOR3xp33_ASAP7_75t_SL U16454 (.Y(n21877),
	.A(n21901),
	.B(n19625),
	.C(n19758));
   NAND2xp5_ASAP7_75t_L U16455 (.Y(n24956),
	.A(n19788),
	.B(n16618));
   NOR3xp33_ASAP7_75t_L U16456 (.Y(n24979),
	.A(n16562),
	.B(n24901),
	.C(n23143));
   O2A1O1Ixp5_ASAP7_75t_L U16458 (.Y(n25599),
	.A1(n19116),
	.A2(n19609),
	.B(FE_OCPN29346_n12998),
	.C(n19115));
   NAND3xp33_ASAP7_75t_L U16459 (.Y(n19115),
	.A(n19114),
	.B(n19113),
	.C(n19598));
   NAND3x1_ASAP7_75t_SL U16460 (.Y(n19132),
	.A(FE_OFN28835_n),
	.B(n21479),
	.C(FE_OCPN27908_FE_OFN16156_sa00_2));
   INVxp33_ASAP7_75t_SRAM U16461 (.Y(n19107),
	.A(n19106));
   NOR2x1_ASAP7_75t_L U16462 (.Y(n22169),
	.A(FE_OCPN27428_n26027),
	.B(FE_OFN29121_n26026));
   NOR2xp33_ASAP7_75t_L U16463 (.Y(n22153),
	.A(FE_OCPN27764_n22152),
	.B(n24792));
   NAND3xp33_ASAP7_75t_SL U16464 (.Y(n22149),
	.A(n22147),
	.B(n22146),
	.C(n22145));
   OAI222xp33_ASAP7_75t_SL U16465 (.Y(n26036),
	.A1(n24131),
	.A2(n24800),
	.B1(n22165),
	.B2(n24800),
	.C1(n22164),
	.C2(n24800));
   NOR3xp33_ASAP7_75t_SRAM U16466 (.Y(n22164),
	.A(n22163),
	.B(FE_OCPN29289_n22162),
	.C(n22161));
   NOR3xp33_ASAP7_75t_SL U16467 (.Y(n22165),
	.A(n22160),
	.B(n22159),
	.C(n25088));
   NAND2xp33_ASAP7_75t_L U16468 (.Y(n22160),
	.A(n22158),
	.B(n22622));
   NOR3x1_ASAP7_75t_L U16469 (.Y(n26023),
	.A(n21605),
	.B(n17618),
	.C(n18381));
   NAND2x1_ASAP7_75t_SL U16470 (.Y(n22130),
	.A(n17637),
	.B(n22628));
   NOR3xp33_ASAP7_75t_L U16471 (.Y(n22654),
	.A(n20459),
	.B(n20458),
	.C(n20457));
   NAND2xp33_ASAP7_75t_L U16472 (.Y(n20458),
	.A(n20455),
	.B(n22151));
   OAI21xp33_ASAP7_75t_R U16473 (.Y(n20457),
	.A1(FE_OFN28896_sa30_2),
	.A2(n25105),
	.B(n20456));
   NAND2xp33_ASAP7_75t_L U16474 (.Y(n20459),
	.A(n20454),
	.B(n20453));
   NOR2xp33_ASAP7_75t_L U16475 (.Y(n20473),
	.A(n25087),
	.B(n20482));
   NAND3xp33_ASAP7_75t_SL U16476 (.Y(n22486),
	.A(FE_OCPN28321_n21341),
	.B(n17445),
	.C(FE_OFN94_sa11_5));
   NAND3x1_ASAP7_75t_SL U16477 (.Y(n23255),
	.A(FE_OCPN28321_n21341),
	.B(FE_OCPN27903_n19223),
	.C(FE_OFN94_sa11_5));
   NOR3xp33_ASAP7_75t_L U16478 (.Y(n19860),
	.A(FE_OCPN28111_n19091),
	.B(n19090),
	.C(n19139));
   NOR3xp33_ASAP7_75t_SL U16479 (.Y(n26104),
	.A(n21153),
	.B(n19813),
	.C(n21444));
   NOR3x1_ASAP7_75t_L U16480 (.Y(n26099),
	.A(FE_OCPN27518_n17251),
	.B(FE_OCPN29396_n19149),
	.C(n17298));
   OAI21xp33_ASAP7_75t_L U16481 (.Y(n24081),
	.A1(n21373),
	.A2(n21372),
	.B(FE_OFN94_sa11_5));
   OAI22xp33_ASAP7_75t_SRAM U16482 (.Y(n24083),
	.A1(n17444),
	.A2(n21817),
	.B1(FE_OFN29034_FE_OCPN27414_n23359),
	.B2(n21817));
   NAND3xp33_ASAP7_75t_L U16483 (.Y(n21864),
	.A(n25793),
	.B(n23282),
	.C(n23369));
   NAND2xp5_ASAP7_75t_SL U16484 (.Y(n21839),
	.A(n21836),
	.B(n21835));
   NAND2xp5_ASAP7_75t_SL U16485 (.Y(n22498),
	.A(n21850),
	.B(n21849));
   NOR3xp33_ASAP7_75t_SL U16486 (.Y(n22497),
	.A(n21819),
	.B(FE_OFN29137_FE_OCPN27228_sa11_2),
	.C(FE_OCPN27592_n17501));
   NOR2x1_ASAP7_75t_SL U16487 (.Y(n24559),
	.A(n19194),
	.B(n19193));
   NAND2xp5_ASAP7_75t_SL U16488 (.Y(n19199),
	.A(n21393),
	.B(n21396));
   NOR3x1_ASAP7_75t_SL U16489 (.Y(n22629),
	.A(n20428),
	.B(FE_OFN28895_sa30_2),
	.C(n19051));
   NOR3x1_ASAP7_75t_SL U16490 (.Y(n18368),
	.A(FE_OFN25901_n22133),
	.B(FE_OCPN29431_sa30_3),
	.C(n21627));
   NAND2xp5_ASAP7_75t_L U16491 (.Y(n22151),
	.A(n17621),
	.B(n21591));
   NOR2xp33_ASAP7_75t_R U16492 (.Y(n17621),
	.A(FE_OFN16200_sa30_2),
	.B(n18352));
   NAND2x1_ASAP7_75t_L U16494 (.Y(n21626),
	.A(n17630),
	.B(FE_OCPN29398_sa30_3));
   NAND3xp33_ASAP7_75t_L U16495 (.Y(n21628),
	.A(n19056),
	.B(n24787),
	.C(n18481));
   NOR3x1_ASAP7_75t_SL U16496 (.Y(n23831),
	.A(n18561),
	.B(FE_OCPN29430_FE_OFN31_sa20_0),
	.C(n18582));
   NOR2x1_ASAP7_75t_L U16497 (.Y(n23884),
	.A(FE_OCPN27891_n18561),
	.B(n18599));
   NAND2x1_ASAP7_75t_SL U16498 (.Y(n21658),
	.A(n18588),
	.B(n21239));
   NOR2x1_ASAP7_75t_L U16499 (.Y(n22305),
	.A(n20753),
	.B(FE_OCPN29305_n23302));
   NOR2x1_ASAP7_75t_L U16500 (.Y(n23165),
	.A(n21093),
	.B(n21092));
   NAND2xp33_ASAP7_75t_L U16501 (.Y(n21093),
	.A(FE_OFN28966_n23329),
	.B(n21782));
   OAI222xp33_ASAP7_75t_L U16502 (.Y(n21091),
	.A1(FE_OCPN27979_FE_OFN16147_sa22_1),
	.A2(n23297),
	.B1(FE_PSN8320_n18176),
	.B2(n23297),
	.C1(FE_OCPN27722_n23336),
	.C2(n23297));
   NAND2xp5_ASAP7_75t_SL U16503 (.Y(n18209),
	.A(n21126),
	.B(n23325));
   NOR2xp33_ASAP7_75t_SL U16504 (.Y(n22808),
	.A(FE_OFN26548_n18206),
	.B(n21772));
   NAND2xp5_ASAP7_75t_R U16505 (.Y(n22308),
	.A(n22269),
	.B(n24702));
   NAND2x1_ASAP7_75t_SL U16506 (.Y(n22309),
	.A(n18227),
	.B(n18226));
   NAND2xp33_ASAP7_75t_SRAM U16507 (.Y(n18226),
	.A(FE_OFN26141_n23307),
	.B(n18162));
   NOR3xp33_ASAP7_75t_SL U16508 (.Y(n18227),
	.A(n23162),
	.B(n23297),
	.C(n22796));
   NAND2xp33_ASAP7_75t_L U16509 (.Y(n21766),
	.A(n21787),
	.B(n20704));
   NAND2x1_ASAP7_75t_SL U16510 (.Y(n23745),
	.A(n23714),
	.B(n21233));
   NOR2xp67_ASAP7_75t_SL U16511 (.Y(n21233),
	.A(n21232),
	.B(n21231));
   NAND2xp33_ASAP7_75t_L U16512 (.Y(n21231),
	.A(n21230),
	.B(n21229));
   NAND2xp33_ASAP7_75t_SL U16513 (.Y(n21229),
	.A(n21228),
	.B(n21227));
   NOR3x1_ASAP7_75t_L U16514 (.Y(n25902),
	.A(n23726),
	.B(FE_OCPN29567_n23806),
	.C(n23880));
   NOR2xp33_ASAP7_75t_R U16515 (.Y(n23704),
	.A(FE_OFN29081_n18526),
	.B(n23792));
   NAND3xp33_ASAP7_75t_R U16516 (.Y(n18559),
	.A(n23803),
	.B(n23833),
	.C(n18595));
   NOR2x1_ASAP7_75t_L U16517 (.Y(n23685),
	.A(n21654),
	.B(n21653));
   NOR3xp33_ASAP7_75t_R U16518 (.Y(n18438),
	.A(n18434),
	.B(n18433),
	.C(n23530));
   NOR2x1_ASAP7_75t_L U16519 (.Y(n18437),
	.A(n16935),
	.B(n16920));
   NOR2x1_ASAP7_75t_SL U16520 (.Y(n18445),
	.A(n16867),
	.B(n16929));
   NOR3xp33_ASAP7_75t_L U16521 (.Y(n18441),
	.A(n18143),
	.B(n18142),
	.C(FE_OCPN28322_n18141));
   NAND2xp5_ASAP7_75t_L U16522 (.Y(n23557),
	.A(n16887),
	.B(n16454));
   NOR2xp33_ASAP7_75t_SL U16523 (.Y(n16719),
	.A(n18425),
	.B(n18143));
   NOR3x1_ASAP7_75t_L U16525 (.Y(n23539),
	.A(n16925),
	.B(FE_OFN29164_sa33_2),
	.C(FE_OCPN29299_FE_OFN29232_n16875));
   OR3x1_ASAP7_75t_L U16526 (.Y(n23535),
	.A(n16692),
	.B(n23553),
	.C(n16859));
   NAND3xp33_ASAP7_75t_L U16527 (.Y(n16692),
	.A(n17429),
	.B(n16724),
	.C(n16691));
   NOR3x1_ASAP7_75t_L U16530 (.Y(n16867),
	.A(n16429),
	.B(FE_OFN29164_sa33_2),
	.C(FE_OCPN29299_FE_OFN29232_n16875));
   NOR2x1_ASAP7_75t_L U16531 (.Y(n24300),
	.A(n16473),
	.B(n16429));
   NOR2xp67_ASAP7_75t_L U16532 (.Y(n18145),
	.A(n16847),
	.B(n16925));
   NOR3xp33_ASAP7_75t_SL U16533 (.Y(n16927),
	.A(n16844),
	.B(n16843),
	.C(n16842));
   NAND2xp33_ASAP7_75t_SRAM U16534 (.Y(n16842),
	.A(n16841),
	.B(n16840));
   NAND2xp33_ASAP7_75t_SRAM U16535 (.Y(n16843),
	.A(n23529),
	.B(n16945));
   NAND2xp33_ASAP7_75t_L U16536 (.Y(n18144),
	.A(n16924),
	.B(n18121));
   NOR3xp33_ASAP7_75t_SRAM U16538 (.Y(n26161),
	.A(n22926),
	.B(FE_OFN26127_n22925),
	.C(n25095));
   NAND3xp33_ASAP7_75t_R U16540 (.Y(n26162),
	.A(FE_OCPN29331_n20933),
	.B(FE_OCPN27986_n18970),
	.C(FE_OFN27078_sa23_5));
   NAND2xp5_ASAP7_75t_L U16541 (.Y(n24769),
	.A(FE_OCPN5191_n20272),
	.B(n20268));
   NAND2xp5_ASAP7_75t_L U16542 (.Y(n22984),
	.A(n20231),
	.B(n20233));
   NAND2xp33_ASAP7_75t_L U16543 (.Y(n20233),
	.A(n20232),
	.B(n20919));
   NOR2xp33_ASAP7_75t_L U16544 (.Y(n19346),
	.A(FE_PSN8328_n20260),
	.B(n25093));
   NAND2xp5_ASAP7_75t_SL U16545 (.Y(n22969),
	.A(FE_OCPN27743_n22009),
	.B(n19000));
   NAND2xp33_ASAP7_75t_SRAM U16546 (.Y(n22968),
	.A(FE_OCPN27727_n22964),
	.B(FE_OCPN29480_n20913));
   NOR3xp33_ASAP7_75t_SL U16547 (.Y(n18675),
	.A(n20369),
	.B(n21560),
	.C(n23060));
   NAND2x1_ASAP7_75t_SL U16548 (.Y(n22470),
	.A(n17321),
	.B(FE_OCPN29454_n18671));
   NOR2x1_ASAP7_75t_L U16549 (.Y(n23076),
	.A(FE_OFN27152_n17315),
	.B(n18716));
   NAND2xp5_ASAP7_75t_L U16550 (.Y(n24396),
	.A(FE_OCPN29388_n22461),
	.B(n23059));
   NAND3xp33_ASAP7_75t_SL U16551 (.Y(n24392),
	.A(n20395),
	.B(FE_OFN25954_n18719),
	.C(n21539));
   NOR3xp33_ASAP7_75t_L U16552 (.Y(n23097),
	.A(n22464),
	.B(n22463),
	.C(n22462));
   OAI21xp33_ASAP7_75t_L U16553 (.Y(n22462),
	.A1(FE_OCPN29320_n22461),
	.A2(FE_OCPN29334_n17330),
	.B(n22460));
   NOR3x1_ASAP7_75t_SL U16554 (.Y(n27007),
	.A(n21561),
	.B(FE_OCPN29429_FE_OFN16141_sa01_3),
	.C(n17389));
   NAND3xp33_ASAP7_75t_SRAM U16555 (.Y(n22609),
	.A(n22590),
	.B(n22589),
	.C(n22588));
   NOR3xp33_ASAP7_75t_L U16556 (.Y(n27017),
	.A(n22434),
	.B(n22584),
	.C(FE_OCPN28380_n22433));
   OR2x2_ASAP7_75t_SRAM U16557 (.Y(n27015),
	.A(sa01_6_),
	.B(n17392));
   NAND3xp33_ASAP7_75t_SL U16558 (.Y(n25750),
	.A(n17921),
	.B(n22256),
	.C(n17918));
   NAND2xp5_ASAP7_75t_L U16559 (.Y(n22779),
	.A(FE_OCPN5137_n23600),
	.B(n25741));
   NOR2x1_ASAP7_75t_SL U16561 (.Y(n20824),
	.A(n23574),
	.B(n17951));
   NAND3xp33_ASAP7_75t_SL U16562 (.Y(n17951),
	.A(n22725),
	.B(n17950),
	.C(n22254));
   NAND2xp33_ASAP7_75t_SL U16563 (.Y(n20803),
	.A(n20798),
	.B(n20800));
   NAND2xp33_ASAP7_75t_SL U16564 (.Y(n17969),
	.A(n17967),
	.B(n17966));
   NAND2xp33_ASAP7_75t_R U16565 (.Y(n17966),
	.A(n17965),
	.B(n17964));
   NAND2xp33_ASAP7_75t_R U16566 (.Y(n17967),
	.A(n17963),
	.B(n17964));
   NOR3xp33_ASAP7_75t_L U16567 (.Y(n26594),
	.A(n20794),
	.B(n20793),
	.C(n20792));
   NAND2xp5_ASAP7_75t_L U16568 (.Y(n20589),
	.A(n20585),
	.B(FE_OFN16380_n20584));
   NOR3xp33_ASAP7_75t_SL U16570 (.Y(n18841),
	.A(FE_OCPN29348_n17592),
	.B(FE_OCPN29459_n),
	.C(n25029));
   NOR3xp33_ASAP7_75t_L U16571 (.Y(n18798),
	.A(n18818),
	.B(FE_OFN28892_n),
	.C(n17566));
   NAND3x1_ASAP7_75t_SL U16572 (.Y(n25025),
	.A(n17560),
	.B(n19713),
	.C(FE_OCPN8259_FE_OFN28686_FE_OCPN27812));
   NOR2x1_ASAP7_75t_SL U16573 (.Y(n25022),
	.A(FE_OCPN7586_n17693),
	.B(n17692));
   NAND3xp33_ASAP7_75t_SL U16574 (.Y(n17692),
	.A(n20094),
	.B(FE_OFN28965_n24869),
	.C(n19924));
   NAND2xp5_ASAP7_75t_L U16575 (.Y(n24988),
	.A(n17525),
	.B(n18799));
   NAND3xp33_ASAP7_75t_SL U16576 (.Y(n24998),
	.A(n17545),
	.B(n18321),
	.C(n18815));
   NOR3xp33_ASAP7_75t_L U16577 (.Y(n17545),
	.A(n22381),
	.B(n19728),
	.C(n19732));
   NAND2xp33_ASAP7_75t_L U16578 (.Y(n24012),
	.A(n19726),
	.B(n17543));
   NAND2xp5_ASAP7_75t_L U16579 (.Y(n24991),
	.A(n18800),
	.B(n17547));
   NOR2x1_ASAP7_75t_L U16580 (.Y(n22370),
	.A(n18818),
	.B(n19920));
   NOR2xp33_ASAP7_75t_SL U16582 (.Y(n23639),
	.A(n23926),
	.B(n16764));
   NOR2x1_ASAP7_75t_L U16583 (.Y(n17880),
	.A(n17872),
	.B(n23926));
   NAND3xp33_ASAP7_75t_L U16584 (.Y(n25588),
	.A(n19888),
	.B(n19887),
	.C(n19886));
   NOR3xp33_ASAP7_75t_L U16585 (.Y(n19899),
	.A(n19978),
	.B(FE_OCPN29294_n23925),
	.C(n22694));
   AND3x1_ASAP7_75t_SL U16586 (.Y(n23645),
	.A(n23641),
	.B(n23640),
	.C(n23639));
   OAI22xp33_ASAP7_75t_SRAM U16587 (.Y(n23641),
	.A1(FE_OFN28836_FE_OCPN27631_n16774),
	.A2(n23638),
	.B1(n16771),
	.B2(n23638));
   NAND2xp5_ASAP7_75t_L U16588 (.Y(n21972),
	.A(n21933),
	.B(n21932));
   NAND2xp5_ASAP7_75t_L U16590 (.Y(n25318),
	.A(n18063),
	.B(n16326));
   NOR2xp33_ASAP7_75t_SL U16591 (.Y(n25315),
	.A(n21977),
	.B(n20077));
   OAI21xp5_ASAP7_75t_L U16592 (.Y(n20077),
	.A1(FE_OCPN28061_n20076),
	.A2(n20853),
	.B(n20075));
   NAND2xp5_ASAP7_75t_L U16593 (.Y(n25314),
	.A(n16318),
	.B(n16317));
   NAND2xp33_ASAP7_75t_SL U16594 (.Y(n16317),
	.A(n16316),
	.B(n16315));
   NAND2xp33_ASAP7_75t_SL U16595 (.Y(n16318),
	.A(n16314),
	.B(n16315));
   OAI21xp5_ASAP7_75t_SL U16596 (.Y(n20850),
	.A1(FE_OFN26060_sa31_4),
	.A2(n16350),
	.B(n16327));
   NAND2xp5_ASAP7_75t_L U16597 (.Y(n16382),
	.A(n16381),
	.B(n16380));
   OAI222xp33_ASAP7_75t_L U16598 (.Y(n25856),
	.A1(n16393),
	.A2(n27168),
	.B1(n25846),
	.B2(n27168),
	.C1(n25847),
	.C2(n27168));
   NOR2x1_ASAP7_75t_L U16599 (.Y(n25815),
	.A(n21977),
	.B(n26290));
   NOR2x1_ASAP7_75t_L U16600 (.Y(n26347),
	.A(n19919),
	.B(n19918));
   NAND3xp33_ASAP7_75t_L U16601 (.Y(n19918),
	.A(n19917),
	.B(n20093),
	.C(n19916));
   NAND2xp5_ASAP7_75t_L U16602 (.Y(n26345),
	.A(n19915),
	.B(n19914));
   NAND2xp33_ASAP7_75t_L U16603 (.Y(n19915),
	.A(n19909),
	.B(FE_OFN28927_n22374));
   NAND2xp33_ASAP7_75t_L U16604 (.Y(n19914),
	.A(n19913),
	.B(FE_OFN28927_n22374));
   NOR3xp33_ASAP7_75t_SRAM U16605 (.Y(n26344),
	.A(n19908),
	.B(n19907),
	.C(n22399));
   OAI222xp33_ASAP7_75t_R U16606 (.Y(n27186),
	.A1(n17040),
	.A2(n27102),
	.B1(n25196),
	.B2(n27102),
	.C1(n25197),
	.C2(n27102));
   NAND3xp33_ASAP7_75t_L U16608 (.Y(n24147),
	.A(sa23_7_),
	.B(n24045),
	.C(FE_OFN45_sa23_6));
   NAND2xp33_ASAP7_75t_SRAM U16611 (.Y(n22672),
	.A(n22669),
	.B(FE_OFN25968_n22668));
   NOR3xp33_ASAP7_75t_SRAM U16613 (.Y(n24888),
	.A(n22660),
	.B(n22659),
	.C(n22658));
   NAND2xp5_ASAP7_75t_L U16615 (.Y(n26822),
	.A(n24682),
	.B(n24681));
   NAND2xp33_ASAP7_75t_R U16616 (.Y(n24681),
	.A(n24680),
	.B(n24679));
   NAND2xp33_ASAP7_75t_L U16618 (.Y(n24417),
	.A(FE_OFN16164_n25081),
	.B(n24422));
   NAND3xp33_ASAP7_75t_SL U16620 (.Y(n23050),
	.A(n23034),
	.B(n23033),
	.C(n23994));
   NOR3xp33_ASAP7_75t_SRAM U16621 (.Y(n23046),
	.A(FE_OFN27048_n23045),
	.B(n23044),
	.C(n23043));
   NOR3xp33_ASAP7_75t_SL U16623 (.Y(n25831),
	.A(n24154),
	.B(sa20_7_),
	.C(n24153));
   NAND3xp33_ASAP7_75t_L U16624 (.Y(n24169),
	.A(n24163),
	.B(n24162),
	.C(n25197));
   NOR3xp33_ASAP7_75t_L U16626 (.Y(n17151),
	.A(n17150),
	.B(n19378),
	.C(FE_OCPN8253_n17149));
   NAND2xp5_ASAP7_75t_L U16627 (.Y(n17150),
	.A(n17143),
	.B(n17142));
   NOR3xp33_ASAP7_75t_SRAM U16628 (.Y(n16891),
	.A(n16889),
	.B(n24328),
	.C(n23538));
   NOR2xp33_ASAP7_75t_SRAM U16630 (.Y(n16898),
	.A(n17405),
	.B(n17424));
   NOR3xp33_ASAP7_75t_SL U16631 (.Y(n16899),
	.A(n16897),
	.B(n16896),
	.C(n24299));
   NOR2xp33_ASAP7_75t_L U16632 (.Y(n13634),
	.A(w3_26_),
	.B(w3_24_));
   NOR2xp33_ASAP7_75t_L U16633 (.Y(n15884),
	.A(w3_0_),
	.B(w3_2_));
   O2A1O1Ixp33_ASAP7_75t_SL U16634 (.Y(n26589),
	.A1(n26710),
	.A2(n26709),
	.B(n26577),
	.C(n26576));
   NOR2xp33_ASAP7_75t_SRAM U16635 (.Y(n26577),
	.A(FE_OCPN28083_n26574),
	.B(n26703));
   NAND2xp33_ASAP7_75t_L U16636 (.Y(n24528),
	.A(n26110),
	.B(n24521));
   NAND2xp33_ASAP7_75t_SRAM U16637 (.Y(n24521),
	.A(n24520),
	.B(FE_OFN163_sa00_7));
   A2O1A1Ixp33_ASAP7_75t_SL U16638 (.Y(n26383),
	.A1(n27117),
	.A2(n27116),
	.B(n25608),
	.C(n25607));
   NAND2xp33_ASAP7_75t_L U16639 (.Y(n25608),
	.A(FE_OFN29011_n27113),
	.B(n26630));
   O2A1O1Ixp5_ASAP7_75t_L U16640 (.Y(n26890),
	.A1(n26889),
	.A2(n26888),
	.B(n26887),
	.C(n26886));
   A2O1A1Ixp33_ASAP7_75t_SL U16641 (.Y(n26891),
	.A1(n27127),
	.A2(n27126),
	.B(n26869),
	.C(n26868));
   NOR2xp33_ASAP7_75t_R U16642 (.Y(n26887),
	.A(w0_20_),
	.B(n26883));
   NAND2xp33_ASAP7_75t_SRAM U16643 (.Y(n27125),
	.A(w0_5_),
	.B(FE_OFN29024_n));
   O2A1O1Ixp5_ASAP7_75t_SL U16644 (.Y(n26259),
	.A1(FE_OFN16413_n26687),
	.A2(n26258),
	.B(n26257),
	.C(n26256));
   O2A1O1Ixp33_ASAP7_75t_SL U16645 (.Y(n25560),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(n25559),
	.C(n25558));
   NOR2xp33_ASAP7_75t_SL U16646 (.Y(n25559),
	.A(w2_27_),
	.B(n26954));
   NOR2xp33_ASAP7_75t_R U16647 (.Y(n24716),
	.A(w0_27_),
	.B(n24713));
   NOR2xp33_ASAP7_75t_SRAM U16648 (.Y(n25429),
	.A(FE_OCPN28407_FE_OFN16433_w3_11),
	.B(n25667));
   NOR2xp33_ASAP7_75t_SRAM U16649 (.Y(n26126),
	.A(FE_OFN46_w0_12),
	.B(FE_OCPN27641_n27121));
   NOR2xp33_ASAP7_75t_SRAM U16650 (.Y(n25671),
	.A(FE_OFN27100_n25675),
	.B(n25667));
   NAND2xp33_ASAP7_75t_L U16651 (.Y(n25046),
	.A(n25037),
	.B(n25036));
   OAI21xp33_ASAP7_75t_R U16652 (.Y(n25047),
	.A1(n25149),
	.A2(n26346),
	.B(n25021));
   O2A1O1Ixp33_ASAP7_75t_L U16653 (.Y(n26092),
	.A1(FE_OFN16180_n26542),
	.A2(n18158),
	.B(n26090),
	.C(n26089));
   NOR2xp33_ASAP7_75t_SRAM U16654 (.Y(n26090),
	.A(w0_11_),
	.B(FE_OFN25973_n26087));
   NOR3xp33_ASAP7_75t_SL U16655 (.Y(n24110),
	.A(FE_OFN28934_n24552),
	.B(n24111),
	.C(n24112));
   NAND2xp33_ASAP7_75t_R U16656 (.Y(n24116),
	.A(FE_OFN106_n24511),
	.B(n26764));
   A2O1A1Ixp33_ASAP7_75t_L U16657 (.Y(n24753),
	.A1(n22405),
	.A2(n24930),
	.B(n24748),
	.C(n24747));
   NAND2xp33_ASAP7_75t_SL U16658 (.Y(n24746),
	.A(FE_OCPN7599_n26721),
	.B(n24743));
   O2A1O1Ixp33_ASAP7_75t_L U16660 (.Y(n25687),
	.A1(FE_OFN16413_n26687),
	.A2(n26258),
	.B(n25686),
	.C(n25685));
   NOR2xp33_ASAP7_75t_SL U16661 (.Y(n25686),
	.A(w1_11_),
	.B(FE_OFN16311_n26252));
   NAND2xp5_ASAP7_75t_L U16662 (.Y(n26225),
	.A(FE_OCPN27394_n26223),
	.B(n26221));
   NAND2xp33_ASAP7_75t_SRAM U16663 (.Y(n26182),
	.A(FE_OFN47_w1_2),
	.B(n26179));
   NAND2xp5_ASAP7_75t_L U16664 (.Y(n24814),
	.A(n26179),
	.B(n24821));
   NAND3xp33_ASAP7_75t_L U16665 (.Y(n24408),
	.A(n24409),
	.B(n24410),
	.C(n24405));
   A2O1A1Ixp33_ASAP7_75t_L U16666 (.Y(n24409),
	.A1(FE_OFN16169_n26567),
	.A2(FE_OFN28506_n26996),
	.B(n24407),
	.C(n24406));
   NAND2xp33_ASAP7_75t_R U16667 (.Y(n24125),
	.A(n24122),
	.B(n26467));
   NAND2xp5_ASAP7_75t_SRAM U16669 (.Y(n25181),
	.A(n25179),
	.B(n25184));
   A2O1A1Ixp33_ASAP7_75t_SL U16670 (.Y(n25268),
	.A1(n27117),
	.A2(FE_OFN28690_n25979),
	.B(n25267),
	.C(n25266));
   A2O1A1Ixp33_ASAP7_75t_SL U16671 (.Y(n25266),
	.A1(FE_OFN28690_n25979),
	.A2(n27117),
	.B(n25974),
	.C(n25265));
   NAND2xp5_ASAP7_75t_L U16672 (.Y(n25267),
	.A(w0_1_),
	.B(FE_OFN16263_n25976));
   O2A1O1Ixp5_ASAP7_75t_SL U16673 (.Y(n24314),
	.A1(FE_OFN16180_n26542),
	.A2(n26431),
	.B(n24308),
	.C(n24307));
   O2A1O1Ixp33_ASAP7_75t_L U16674 (.Y(n26924),
	.A1(n26926),
	.A2(n26995),
	.B(n26992),
	.C(FE_OFN25926_n26922));
   A2O1A1Ixp33_ASAP7_75t_SL U16675 (.Y(n25980),
	.A1(n27117),
	.A2(FE_OFN28690_n25979),
	.B(n25978),
	.C(n25977));
   A2O1A1Ixp33_ASAP7_75t_L U16676 (.Y(n25977),
	.A1(FE_OFN28690_n25979),
	.A2(n27117),
	.B(n25974),
	.C(n25975));
   NAND2xp5_ASAP7_75t_L U16677 (.Y(n25978),
	.A(FE_OFN38_w0_17),
	.B(FE_OFN16263_n25976));
   NAND2xp33_ASAP7_75t_SL U16678 (.Y(n24452),
	.A(n26850),
	.B(n24449));
   NAND2xp33_ASAP7_75t_SRAM U16679 (.Y(n25335),
	.A(w2_9_),
	.B(n26936));
   A2O1A1Ixp33_ASAP7_75t_R U16681 (.Y(n25456),
	.A1(n26139),
	.A2(n25455),
	.B(n25454),
	.C(n25453));
   NAND2xp33_ASAP7_75t_L U16682 (.Y(n25454),
	.A(w1_25_),
	.B(n25451));
   A2O1A1Ixp33_ASAP7_75t_L U16683 (.Y(n24468),
	.A1(n26857),
	.A2(n19640),
	.B(n24251),
	.C(n24250));
   NAND2xp33_ASAP7_75t_SRAM U16684 (.Y(n24251),
	.A(n25010),
	.B(n25384));
   NAND2xp33_ASAP7_75t_L U16685 (.Y(n25920),
	.A(n25910),
	.B(n25909));
   NAND2xp33_ASAP7_75t_R U16686 (.Y(n25910),
	.A(n25900),
	.B(n25907));
   NOR2xp33_ASAP7_75t_SRAM U16687 (.Y(n27138),
	.A(w2_17_),
	.B(FE_OCPN29514_n27136));
   A2O1A1Ixp33_ASAP7_75t_SL U16688 (.Y(n26140),
	.A1(n26139),
	.A2(n26138),
	.B(n26137),
	.C(n26136));
   NAND2xp5_ASAP7_75t_L U16689 (.Y(n26137),
	.A(w1_28_),
	.B(n26134));
   A2O1A1Ixp33_ASAP7_75t_L U16690 (.Y(n26373),
	.A1(n27062),
	.A2(n26372),
	.B(n26371),
	.C(n26370));
   NAND2xp33_ASAP7_75t_R U16691 (.Y(n26371),
	.A(w0_28_),
	.B(n26368));
   O2A1O1Ixp33_ASAP7_75t_SL U16692 (.Y(n26518),
	.A1(n26517),
	.A2(n26516),
	.B(n26515),
	.C(n26514));
   O2A1O1Ixp33_ASAP7_75t_L U16693 (.Y(n26514),
	.A1(n26517),
	.A2(n26516),
	.B(n26513),
	.C(n26512));
   O2A1O1Ixp33_ASAP7_75t_SL U16694 (.Y(n25150),
	.A1(n26346),
	.A2(n25149),
	.B(n25148),
	.C(n25147));
   O2A1O1Ixp33_ASAP7_75t_L U16695 (.Y(n25151),
	.A1(n25420),
	.A2(FE_OFN28561_n25419),
	.B(n25142),
	.C(n25141));
   O2A1O1Ixp33_ASAP7_75t_SL U16696 (.Y(n25147),
	.A1(n26346),
	.A2(n25149),
	.B(FE_OFN29020_n25146),
	.C(n25145));
   O2A1O1Ixp33_ASAP7_75t_SL U16697 (.Y(n26960),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(n26957),
	.C(n26956));
   NOR2xp33_ASAP7_75t_SRAM U16698 (.Y(n26957),
	.A(w2_11_),
	.B(n26954));
   O2A1O1Ixp33_ASAP7_75t_SL U16699 (.Y(n27029),
	.A1(n26926),
	.A2(n26995),
	.B(n26994),
	.C(n26993));
   NOR2xp33_ASAP7_75t_SL U16700 (.Y(n26994),
	.A(w1_1_),
	.B(FE_OFN28451_n26990));
   O2A1O1Ixp33_ASAP7_75t_R U16701 (.Y(n26312),
	.A1(n26315),
	.A2(n26314),
	.B(n26311),
	.C(n26310));
   NOR2xp33_ASAP7_75t_L U16702 (.Y(n26498),
	.A(n26495),
	.B(n26954));
   NAND2xp5_ASAP7_75t_R U16704 (.Y(n25804),
	.A(n26364),
	.B(n25802));
   O2A1O1Ixp33_ASAP7_75t_SL U16705 (.Y(n26712),
	.A1(n27004),
	.A2(n26702),
	.B(n26701),
	.C(n26700));
   NOR2xp33_ASAP7_75t_R U16706 (.Y(n26708),
	.A(n26704),
	.B(n26703));
   A2O1A1Ixp33_ASAP7_75t_L U16707 (.Y(n26727),
	.A1(n26819),
	.A2(n26725),
	.B(n26724),
	.C(n26723));
   NAND2xp5_ASAP7_75t_L U16708 (.Y(n26724),
	.A(FE_OCPN7599_n26721),
	.B(FE_OFN28713_n));
   OAI21xp33_ASAP7_75t_R U16709 (.Y(n25472),
	.A1(n20019),
	.A2(n24263),
	.B(n20018));
   NOR3xp33_ASAP7_75t_SRAM U16710 (.Y(n20019),
	.A(n24252),
	.B(n24253),
	.C(n19995));
   NAND3xp33_ASAP7_75t_SRAM U16712 (.Y(n25475),
	.A(n24269),
	.B(n19991),
	.C(n24921));
   A2O1A1Ixp33_ASAP7_75t_SL U16717 (.Y(n27058),
	.A1(n23293),
	.A2(n23292),
	.B(n17463),
	.C(n23291));
   NOR3xp33_ASAP7_75t_SRAM U16718 (.Y(n23293),
	.A(n24564),
	.B(n23267),
	.C(n23277));
   NOR3xp33_ASAP7_75t_SRAM U16719 (.Y(n23292),
	.A(n23271),
	.B(n26076),
	.C(n23270));
   NAND2x1_ASAP7_75t_SL U16720 (.Y(n27061),
	.A(n23265),
	.B(n23264));
   NOR3xp33_ASAP7_75t_L U16721 (.Y(n23264),
	.A(n23263),
	.B(n23262),
	.C(n23261));
   NAND3x1_ASAP7_75t_L U16722 (.Y(n27052),
	.A(n23321),
	.B(n23320),
	.C(n23352));
   NOR3xp33_ASAP7_75t_R U16723 (.Y(n23321),
	.A(n23298),
	.B(n23297),
	.C(FE_OFN28505_n23296));
   NOR3xp33_ASAP7_75t_SL U16724 (.Y(n23320),
	.A(n23305),
	.B(n23304),
	.C(n26876));
   A2O1A1Ixp33_ASAP7_75t_SL U16726 (.Y(n26825),
	.A1(n22715),
	.A2(n22714),
	.B(n24263),
	.C(n22713));
   NAND3xp33_ASAP7_75t_SRAM U16727 (.Y(n22711),
	.A(n22707),
	.B(n22710),
	.C(n24268));
   NOR3xp33_ASAP7_75t_SL U16728 (.Y(n23788),
	.A(n23763),
	.B(n23762),
	.C(n23761));
   NAND3xp33_ASAP7_75t_SL U16729 (.Y(n23784),
	.A(n23783),
	.B(n23782),
	.C(FE_PSN8316_n23781));
   NAND3x1_ASAP7_75t_L U16730 (.Y(n27192),
	.A(n23760),
	.B(n23759),
	.C(n23771));
   NOR3xp33_ASAP7_75t_SRAM U16731 (.Y(n23760),
	.A(n23741),
	.B(n23740),
	.C(n23739));
   NAND2xp33_ASAP7_75t_L U16732 (.Y(n23759),
	.A(n23749),
	.B(n23748));
   NAND2xp33_ASAP7_75t_L U16733 (.Y(n23749),
	.A(n23744),
	.B(n23746));
   OAI21xp5_ASAP7_75t_L U16734 (.Y(n25834),
	.A1(n19285),
	.A2(n26976),
	.B(n19284));
   NOR3xp33_ASAP7_75t_SRAM U16735 (.Y(n19285),
	.A(n19260),
	.B(n25202),
	.C(n25201));
   NAND2xp5_ASAP7_75t_SRAM U16736 (.Y(n25837),
	.A(n19247),
	.B(n19254));
   NOR3xp33_ASAP7_75t_SL U16737 (.Y(n19750),
	.A(n19724),
	.B(n19723),
	.C(n19722));
   OAI21xp33_ASAP7_75t_SRAM U16738 (.Y(n19722),
	.A1(FE_OCPN29323_n19721),
	.A2(FE_OCPN29298_n25028),
	.B(n19720));
   NOR2xp33_ASAP7_75t_L U16739 (.Y(n22572),
	.A(n22904),
	.B(n22546));
   NAND3xp33_ASAP7_75t_R U16740 (.Y(n22546),
	.A(n22545),
	.B(n22544),
	.C(n25307));
   NOR2xp33_ASAP7_75t_SRAM U16741 (.Y(n22537),
	.A(n22536),
	.B(n22541));
   NOR3xp33_ASAP7_75t_SRAM U16742 (.Y(n22538),
	.A(n22532),
	.B(n22531),
	.C(n22530));
   NOR3xp33_ASAP7_75t_L U16744 (.Y(n18663),
	.A(n18637),
	.B(n27039),
	.C(n26106));
   NAND3xp33_ASAP7_75t_R U16745 (.Y(n18637),
	.A(n24084),
	.B(n18630),
	.C(n18629));
   NAND3xp33_ASAP7_75t_L U16747 (.Y(n25465),
	.A(n23429),
	.B(n23428),
	.C(n23427));
   NOR3xp33_ASAP7_75t_L U16748 (.Y(n23428),
	.A(n23424),
	.B(n23423),
	.C(n23442));
   NOR3xp33_ASAP7_75t_SL U16749 (.Y(n19962),
	.A(n19937),
	.B(n19936),
	.C(n19935));
   NAND3x1_ASAP7_75t_L U16750 (.Y(n24830),
	.A(n26344),
	.B(n26345),
	.C(n26347));
   NAND3xp33_ASAP7_75t_L U16753 (.Y(n25950),
	.A(n21277),
	.B(n21276),
	.C(n21275));
   NOR3xp33_ASAP7_75t_L U16754 (.Y(n21276),
	.A(n21274),
	.B(n17989),
	.C(n21273));
   OAI21xp33_ASAP7_75t_SRAM U16755 (.Y(n21273),
	.A1(FE_OFN28886_FE_OCPN27675_n17986),
	.A2(FE_OFN27133_n21725),
	.B(n21272));
   INVxp67_ASAP7_75t_L U16757 (.Y(n25961),
	.A(w3_21_));
   NOR3xp33_ASAP7_75t_L U16758 (.Y(n21188),
	.A(n21161),
	.B(n21160),
	.C(n21159));
   NOR2xp33_ASAP7_75t_R U16759 (.Y(n21189),
	.A(n21464),
	.B(n21153));
   NOR2xp33_ASAP7_75t_L U16760 (.Y(n26637),
	.A(sa00_7_),
	.B(n17305));
   NOR3x1_ASAP7_75t_SL U16761 (.Y(n25258),
	.A(n17256),
	.B(n18734),
	.C(n21465));
   OAI22xp33_ASAP7_75t_L U16762 (.Y(n25549),
	.A1(n16983),
	.A2(n19411),
	.B1(n16975),
	.B2(n19411));
   NAND3xp33_ASAP7_75t_SL U16763 (.Y(n24844),
	.A(n24247),
	.B(n21508),
	.C(n24245));
   NAND2xp33_ASAP7_75t_SRAM U16764 (.Y(n21507),
	.A(n24241),
	.B(n21506));
   NAND2xp5_ASAP7_75t_SL U16765 (.Y(n25044),
	.A(n17189),
	.B(n17188));
   NOR2xp33_ASAP7_75t_R U16766 (.Y(n17188),
	.A(n24901),
	.B(n24459));
   NOR3xp33_ASAP7_75t_R U16767 (.Y(n17189),
	.A(n17185),
	.B(n24458),
	.C(n24460));
   NAND2xp33_ASAP7_75t_SRAM U16768 (.Y(n17185),
	.A(n24461),
	.B(n24964));
   NOR3xp33_ASAP7_75t_SL U16769 (.Y(n23157),
	.A(n23130),
	.B(n24726),
	.C(n24727));
   NOR2xp67_ASAP7_75t_L U16771 (.Y(n24974),
	.A(sa10_7_),
	.B(sa10_6_));
   NOR3xp33_ASAP7_75t_SL U16772 (.Y(n24581),
	.A(n17658),
	.B(n20460),
	.C(n17657));
   OAI21xp33_ASAP7_75t_SRAM U16773 (.Y(n17657),
	.A1(n20471),
	.A2(FE_OCPN27428_n26027),
	.B(n18490));
   NAND2xp33_ASAP7_75t_L U16775 (.Y(n24580),
	.A(n18357),
	.B(n18356));
   NAND2xp33_ASAP7_75t_SRAM U16776 (.Y(n18356),
	.A(n18355),
	.B(n18354));
   NAND2xp33_ASAP7_75t_R U16777 (.Y(n18357),
	.A(n18353),
	.B(n18354));
   NOR3xp33_ASAP7_75t_L U16778 (.Y(n18399),
	.A(n18367),
	.B(n24128),
	.C(n22148));
   NOR2xp33_ASAP7_75t_SRAM U16779 (.Y(n23400),
	.A(sa11_6_),
	.B(n19161));
   NOR2xp67_ASAP7_75t_L U16781 (.Y(n27062),
	.A(FE_OFN150_sa11_7),
	.B(n21340));
   NOR3xp33_ASAP7_75t_L U16782 (.Y(n24153),
	.A(n25191),
	.B(FE_OFN16301_n25905),
	.C(n21646));
   NAND2xp33_ASAP7_75t_SRAM U16783 (.Y(n21646),
	.A(n25189),
	.B(FE_OFN29096_n25188));
   NAND2xp33_ASAP7_75t_L U16784 (.Y(n21700),
	.A(n21662),
	.B(n21661));
   INVxp33_ASAP7_75t_SRAM U16785 (.Y(n21701),
	.A(FE_OCPN8233_n21647));
   NAND2xp5_ASAP7_75t_L U16786 (.Y(n23861),
	.A(n23860),
	.B(n23859));
   NAND2xp33_ASAP7_75t_SRAM U16787 (.Y(n23859),
	.A(n23858),
	.B(n23857));
   NAND2xp33_ASAP7_75t_SL U16788 (.Y(n23860),
	.A(n23854),
	.B(n23857));
   NOR2x1_ASAP7_75t_L U16789 (.Y(n26770),
	.A(FE_OFN173_sa33_6),
	.B(FE_OFN90_sa33_7));
   INVxp67_ASAP7_75t_L U16790 (.Y(n26124),
	.A(FE_OCPN27641_n27121));
   INVxp67_ASAP7_75t_L U16793 (.Y(n25698),
	.A(FE_OCPN27507_n25695));
   INVxp33_ASAP7_75t_SRAM U16794 (.Y(n25179),
	.A(n25681));
   NOR2x1_ASAP7_75t_L U16795 (.Y(n25682),
	.A(FE_OFN175_sa12_6),
	.B(FE_OFN165_sa12_7));
   NAND3xp33_ASAP7_75t_SL U16796 (.Y(n24214),
	.A(n24586),
	.B(n22232),
	.C(n24585));
   NOR2xp33_ASAP7_75t_SRAM U16797 (.Y(n22232),
	.A(FE_OCPN8235_n24589),
	.B(n22231));
   NOR2xp33_ASAP7_75t_SRAM U16798 (.Y(n27100),
	.A(w2_25_),
	.B(n27097));
   NOR2x1_ASAP7_75t_L U16800 (.Y(n18855),
	.A(n18817),
	.B(n18816));
   NAND3xp33_ASAP7_75t_SL U16801 (.Y(n26842),
	.A(n18804),
	.B(n18803),
	.C(n25024));
   NAND2xp33_ASAP7_75t_L U16802 (.Y(n18804),
	.A(n18792),
	.B(n18791));
   NAND2xp33_ASAP7_75t_SRAM U16803 (.Y(n18791),
	.A(n24858),
	.B(n18790));
   NOR2x1_ASAP7_75t_R U16804 (.Y(n25367),
	.A(FE_OFN25946_sa32_6),
	.B(FE_OFN25997_n));
   NOR2xp67_ASAP7_75t_L U16806 (.Y(n25575),
	.A(sa21_6_),
	.B(sa21_7_));
   NAND3xp33_ASAP7_75t_L U16807 (.Y(n25005),
	.A(n22338),
	.B(n22337),
	.C(n24920));
   NAND2xp33_ASAP7_75t_R U16808 (.Y(n13332),
	.A(n13329),
	.B(n27129));
   OAI21xp5_ASAP7_75t_L U16809 (.Y(n13333),
	.A1(n14491),
	.A2(n14504),
	.B(n13285));
   OAI21xp5_ASAP7_75t_SL U16810 (.Y(n16201),
	.A1(n16179),
	.A2(n26018),
	.B(n16178));
   NAND2xp33_ASAP7_75t_R U16811 (.Y(n15655),
	.A(n15652),
	.B(n26744));
   NAND2xp33_ASAP7_75t_R U16812 (.Y(n15656),
	.A(n15584),
	.B(n15583));
   NAND2xp5_ASAP7_75t_L U16813 (.Y(n13454),
	.A(n13450),
	.B(n13449));
   NAND2xp33_ASAP7_75t_L U16814 (.Y(n13449),
	.A(n13448),
	.B(FE_OFN28455_n13348));
   NOR2xp33_ASAP7_75t_R U16815 (.Y(n13448),
	.A(FE_OFN28603_n14534),
	.B(n14479));
   NAND2xp33_ASAP7_75t_L U16816 (.Y(n14547),
	.A(n14546),
	.B(n15224));
   NOR2xp33_ASAP7_75t_L U16817 (.Y(n14546),
	.A(FE_OFN26051_w3_27),
	.B(FE_OFN26552_n14545));
   OA21x2_ASAP7_75t_L U16818 (.Y(n13584),
	.A1(n14515),
	.A2(FE_OFN27085_n),
	.B(n13647));
   NOR2xp67_ASAP7_75t_L U16819 (.Y(n14500),
	.A(FE_OFN27209_w3_30),
	.B(n15183));
   NOR2xp33_ASAP7_75t_R U16820 (.Y(n13456),
	.A(FE_OFN25895_n13662),
	.B(n13454));
   NOR2xp33_ASAP7_75t_SRAM U16821 (.Y(n13453),
	.A(n15170),
	.B(n13454));
   NOR3xp33_ASAP7_75t_SRAM U16822 (.Y(n15985),
	.A(n15983),
	.B(FE_OFN26129_w3_15),
	.C(FE_OCPN29520_n24755));
   NAND2xp5_ASAP7_75t_R U16825 (.Y(n16459),
	.A(FE_OFN26055_n),
	.B(n16456));
   NAND2xp33_ASAP7_75t_SRAM U16826 (.Y(n14542),
	.A(n14541),
	.B(n14540));
   NOR2xp33_ASAP7_75t_R U16827 (.Y(n14541),
	.A(FE_OFN16145_n15214),
	.B(n14539));
   NAND2xp33_ASAP7_75t_SRAM U16828 (.Y(n14543),
	.A(n14538),
	.B(n14540));
   NOR2xp33_ASAP7_75t_R U16829 (.Y(n14538),
	.A(n15234),
	.B(n14539));
   NAND2xp33_ASAP7_75t_L U16830 (.Y(n14584),
	.A(n14583),
	.B(n14582));
   NAND2xp33_ASAP7_75t_R U16831 (.Y(n14582),
	.A(n14581),
	.B(n14580));
   INVxp67_ASAP7_75t_L U16832 (.Y(n13847),
	.A(n13845));
   NOR2xp33_ASAP7_75t_L U16833 (.Y(n15680),
	.A(FE_OFN28977_n),
	.B(FE_OFN27151_n));
   NAND2xp33_ASAP7_75t_L U16834 (.Y(n15243),
	.A(n15237),
	.B(FE_OFN16206_n15240));
   NAND2xp33_ASAP7_75t_L U16835 (.Y(n15242),
	.A(n15241),
	.B(FE_OFN16206_n15240));
   NOR2xp33_ASAP7_75t_SRAM U16836 (.Y(n15237),
	.A(n13596),
	.B(n15238));
   INVxp33_ASAP7_75t_L U16837 (.Y(n15210),
	.A(n15206));
   NOR2xp33_ASAP7_75t_SRAM U16838 (.Y(n15191),
	.A(n15189),
	.B(n15188));
   NOR3xp33_ASAP7_75t_R U16839 (.Y(n15154),
	.A(n15200),
	.B(FE_OFN27212_w3_30),
	.C(FE_OFN28859_FE_OCPN27664_w3_25));
   NOR2xp33_ASAP7_75t_SRAM U16840 (.Y(n15170),
	.A(n15155),
	.B(FE_OFN26104_n13659));
   NAND2xp33_ASAP7_75t_SL U16841 (.Y(n13314),
	.A(n13311),
	.B(n13358));
   NOR2xp33_ASAP7_75t_SRAM U16842 (.Y(n13311),
	.A(n14479),
	.B(n13312));
   NOR2xp33_ASAP7_75t_SL U16843 (.Y(n13604),
	.A(FE_OFN25893_n15214),
	.B(n15158));
   NOR2xp33_ASAP7_75t_L U16844 (.Y(n13778),
	.A(n14439),
	.B(n15825));
   NOR2xp33_ASAP7_75t_R U16845 (.Y(n14140),
	.A(FE_OCPN28407_FE_OFN16433_w3_11),
	.B(n15380));
   OA21x2_ASAP7_75t_SL U16846 (.Y(n13920),
	.A1(n15735),
	.A2(FE_OFN27074_n13868),
	.B(n13918));
   NAND3xp33_ASAP7_75t_SL U16848 (.Y(n13904),
	.A(FE_OFN26091_n24663),
	.B(FE_OFN28624_n13874),
	.C(n15729));
   NAND2xp33_ASAP7_75t_L U16849 (.Y(n13586),
	.A(n13585),
	.B(n13584));
   NOR2xp33_ASAP7_75t_L U16850 (.Y(n13585),
	.A(FE_OFN28455_n13348),
	.B(n15168));
   NAND2xp33_ASAP7_75t_SL U16851 (.Y(n13587),
	.A(n13583),
	.B(n13584));
   NOR2xp33_ASAP7_75t_L U16852 (.Y(n13583),
	.A(n14557),
	.B(n15168));
   NAND2xp5_ASAP7_75t_L U16853 (.Y(n13590),
	.A(n13589),
	.B(n13588));
   NAND2xp33_ASAP7_75t_SRAM U16854 (.Y(n13589),
	.A(n15209),
	.B(FE_OFN25966_n13646));
   OAI21xp33_ASAP7_75t_R U16855 (.Y(n15235),
	.A1(FE_OFN27211_w3_30),
	.A2(n14498),
	.B(FE_OFN28604_n14534));
   NOR2xp33_ASAP7_75t_SRAM U16856 (.Y(n13611),
	.A(n15254),
	.B(n13612));
   NOR2xp33_ASAP7_75t_R U16857 (.Y(n13615),
	.A(n13613),
	.B(n13612));
   NAND2xp5_ASAP7_75t_R U16858 (.Y(n15199),
	.A(FE_OFN27211_w3_30),
	.B(n15224));
   OR3x1_ASAP7_75t_SRAM U16859 (.Y(n14868),
	.A(n15808),
	.B(FE_OFN16195_n13771),
	.C(n13741));
   INVx1_ASAP7_75t_L U16860 (.Y(n15333),
	.A(n15280));
   NAND3xp33_ASAP7_75t_SL U16861 (.Y(n15280),
	.A(FE_OFN28683_w3_21),
	.B(n15338),
	.C(FE_OFN16426_w3_20));
   OA21x2_ASAP7_75t_R U16862 (.Y(n13358),
	.A1(n13421),
	.A2(FE_OFN16451_n),
	.B(n13310));
   NAND3xp33_ASAP7_75t_L U16864 (.Y(n13682),
	.A(FE_OFN27209_w3_30),
	.B(n15145),
	.C(n13659));
   NAND2xp5_ASAP7_75t_R U16865 (.Y(n14221),
	.A(n15787),
	.B(n15814));
   NOR2xp33_ASAP7_75t_R U16866 (.Y(n14291),
	.A(n14804),
	.B(n14292));
   NOR2xp33_ASAP7_75t_L U16867 (.Y(n14294),
	.A(n14766),
	.B(n14292));
   NOR3xp33_ASAP7_75t_R U16868 (.Y(n14310),
	.A(FE_OFN29192_n13870),
	.B(FE_OFN27214_w3_17),
	.C(FE_OFN4_w3_22));
   NOR2xp33_ASAP7_75t_L U16869 (.Y(n14315),
	.A(n15694),
	.B(FE_OFN29192_n13870));
   NOR3xp33_ASAP7_75t_R U16870 (.Y(n15615),
	.A(n15888),
	.B(FE_OCPN8252_FE_OFN28661_w3_7),
	.C(n13730));
   OAI21xp33_ASAP7_75t_SRAM U16871 (.Y(n14942),
	.A1(n14941),
	.A2(n14940),
	.B(n25782));
   NOR2xp33_ASAP7_75t_L U16872 (.Y(n15541),
	.A(FE_OFN37_w3_23),
	.B(n14795));
   OA21x2_ASAP7_75t_R U16873 (.Y(n15497),
	.A1(n15494),
	.A2(n13875),
	.B(n15493));
   OAI22xp33_ASAP7_75t_SRAM U16874 (.Y(n15494),
	.A1(FE_PSN8298_FE_OFN27151_n),
	.A2(FE_OFN26535_w3_19),
	.B1(FE_OFN27082_n25377),
	.B2(FE_OFN26535_w3_19));
   INVxp67_ASAP7_75t_R U16875 (.Y(n13484),
	.A(n13713));
   NAND2xp33_ASAP7_75t_SRAM U16876 (.Y(n13527),
	.A(n15240),
	.B(n15183));
   NAND2xp5_ASAP7_75t_SL U16878 (.Y(n13534),
	.A(n13384),
	.B(n13383));
   NAND2xp5_ASAP7_75t_L U16879 (.Y(n13383),
	.A(n13382),
	.B(FE_OFN26567_n));
   NOR2xp33_ASAP7_75t_SL U16880 (.Y(n13382),
	.A(FE_OFN28929_n15182),
	.B(n13551));
   NAND3xp33_ASAP7_75t_R U16881 (.Y(n15099),
	.A(FE_OFN26073_n),
	.B(FE_OFN16276_w3_5),
	.C(n14846));
   NAND2xp5_ASAP7_75t_SL U16882 (.Y(n15864),
	.A(n15109),
	.B(n15108));
   NAND2xp5_ASAP7_75t_L U16883 (.Y(n15109),
	.A(n15107),
	.B(FE_OFN25918_n15813));
   O2A1O1Ixp33_ASAP7_75t_SRAM U16884 (.Y(n14719),
	.A1(n16016),
	.A2(n14714),
	.B(n15921),
	.C(n14713));
   OAI22xp33_ASAP7_75t_SRAM U16885 (.Y(n14713),
	.A1(FE_OFN26642_w3_14),
	.A2(FE_OCPN28408_FE_OFN16433_w3_11),
	.B1(FE_OCPN29509_FE_OFN16184_w3_9),
	.B2(FE_OCPN28408_FE_OFN16433_w3_11));
   NOR2xp33_ASAP7_75t_SL U16886 (.Y(n14718),
	.A(n14715),
	.B(n14719));
   NOR2xp33_ASAP7_75t_SRAM U16887 (.Y(n14715),
	.A(n13804),
	.B(FE_OFN26007_n16010));
   NOR2xp33_ASAP7_75t_L U16888 (.Y(n14696),
	.A(FE_OFN28848_n14912),
	.B(n13804));
   NAND2xp5_ASAP7_75t_R U16889 (.Y(n14697),
	.A(n15927),
	.B(n14919));
   OR2x2_ASAP7_75t_SL U16890 (.Y(n15343),
	.A(FE_OFN28_w3_23),
	.B(n15658));
   NOR2xp33_ASAP7_75t_R U16892 (.Y(n13683),
	.A(FE_OFN16193_n15200),
	.B(n15162));
   NAND2xp33_ASAP7_75t_R U16893 (.Y(n14430),
	.A(FE_OFN26531_n),
	.B(FE_OFN26058_w3_1));
   NOR2xp33_ASAP7_75t_R U16894 (.Y(n15128),
	.A(n25140),
	.B(n15639));
   NOR2xp33_ASAP7_75t_R U16896 (.Y(n24946),
	.A(FE_OFN28807_n24944),
	.B(n24943));
   NAND2xp33_ASAP7_75t_L U16897 (.Y(n24948),
	.A(n24942),
	.B(n24945));
   NOR2xp33_ASAP7_75t_SL U16898 (.Y(n19232),
	.A(FE_OFN29054_n17453),
	.B(n23402));
   NAND3xp33_ASAP7_75t_R U16902 (.Y(n23754),
	.A(n21195),
	.B(n18529),
	.C(FE_OCPN27633_sa20_5));
   NOR2xp33_ASAP7_75t_L U16903 (.Y(n20405),
	.A(n20404),
	.B(n22438));
   NOR3x1_ASAP7_75t_SL U16904 (.Y(n20406),
	.A(n22463),
	.B(n22584),
	.C(FE_OFN16252_n27003));
   NAND2xp33_ASAP7_75t_L U16906 (.Y(n21323),
	.A(n21319),
	.B(n21320));
   NOR2xp33_ASAP7_75t_SL U16907 (.Y(n21319),
	.A(n21318),
	.B(n21502));
   NOR2xp33_ASAP7_75t_SL U16908 (.Y(n19249),
	.A(n25297),
	.B(n22063));
   NOR2x1_ASAP7_75t_L U16911 (.Y(n20208),
	.A(FE_OCPN29436_n22080),
	.B(n22076));
   NOR3x1_ASAP7_75t_L U16912 (.Y(n20971),
	.A(n20208),
	.B(n22533),
	.C(n22871));
   NAND2xp5_ASAP7_75t_R U16914 (.Y(n22892),
	.A(FE_OCPN27771_n19275),
	.B(n22089));
   NOR2x1_ASAP7_75t_SL U16915 (.Y(n16988),
	.A(FE_OFN16444_sa13_1),
	.B(FE_OFN26600_sa13_0));
   NAND2xp67_ASAP7_75t_SL U16917 (.Y(n17006),
	.A(n17005),
	.B(n17004));
   NOR2xp33_ASAP7_75t_L U16920 (.Y(n21019),
	.A(FE_OFN25986_n21012),
	.B(n21017));
   O2A1O1Ixp33_ASAP7_75t_SRAM U16921 (.Y(n18014),
	.A1(FE_OCPN27483_FE_OFN16132_sa03_5),
	.A2(FE_OFN21730_sa03_3),
	.B(FE_OCPN29349_FE_OCPN27405_sa03_4),
	.C(n17998));
   NOR2x1_ASAP7_75t_SL U16922 (.Y(n21318),
	.A(FE_OFN21730_sa03_3),
	.B(n17992));
   NOR3xp33_ASAP7_75t_SL U16925 (.Y(n23137),
	.A(n23036),
	.B(FE_OFN26161_sa10_4),
	.C(n16581));
   NOR3xp33_ASAP7_75t_SL U16926 (.Y(n16534),
	.A(FE_OFN26585_n23011),
	.B(FE_OFN28722_sa10_3),
	.C(FE_OCPN27635_sa10_4));
   NOR3xp33_ASAP7_75t_SL U16927 (.Y(n17194),
	.A(FE_OCPN5015_n23031),
	.B(n21894),
	.C(n19663));
   NAND3xp33_ASAP7_75t_R U16928 (.Y(n18764),
	.A(n17245),
	.B(FE_OFN28835_n),
	.C(FE_OCPN29370_FE_OFN28744));
   NOR2x1p5_ASAP7_75t_SL U16929 (.Y(n19578),
	.A(FE_OCPN28270_n17237),
	.B(FE_OFN26172_n19609));
   NAND2x1_ASAP7_75t_SL U16930 (.Y(n19101),
	.A(n18614),
	.B(n18652));
   NOR3xp33_ASAP7_75t_SL U16931 (.Y(n18614),
	.A(n21438),
	.B(n21439),
	.C(n18746));
   NOR2xp33_ASAP7_75t_L U16932 (.Y(n18392),
	.A(n22614),
	.B(n21586));
   NOR3x1_ASAP7_75t_L U16933 (.Y(n19044),
	.A(FE_OFN29121_n26026),
	.B(FE_OCPN29399_sa30_3),
	.C(FE_OCPN27971_n21627));
   NAND2xp5_ASAP7_75t_SL U16936 (.Y(n18757),
	.A(n18742),
	.B(FE_OCPN29376_n24099));
   NAND2x1p5_ASAP7_75t_L U16937 (.Y(n17247),
	.A(FE_OCPN27818_n17267),
	.B(FE_OFN148_sa00_1));
   NAND2xp5_ASAP7_75t_SL U16938 (.Y(n17300),
	.A(n17271),
	.B(FE_OCPN29464_n));
   NAND2xp5_ASAP7_75t_L U16939 (.Y(n18756),
	.A(FE_OCPN28021_n21445),
	.B(n17245));
   NAND2xp5_ASAP7_75t_L U16941 (.Y(n23393),
	.A(FE_OCPN27625_sa11_5),
	.B(FE_OFN26554_n19170));
   NAND2xp5_ASAP7_75t_L U16943 (.Y(n23356),
	.A(FE_OCPN27730_n17464),
	.B(n17445));
   NAND3xp33_ASAP7_75t_SL U16944 (.Y(n19046),
	.A(FE_OFN29094_n21607),
	.B(FE_OCPN28057_n17603),
	.C(FE_OFN28896_sa30_2));
   NAND2xp5_ASAP7_75t_SL U16945 (.Y(n20654),
	.A(FE_OCPN27591_n23742),
	.B(n23721));
   NAND2xp5_ASAP7_75t_L U16946 (.Y(n22282),
	.A(n23312),
	.B(n21105));
   INVx1_ASAP7_75t_L U16947 (.Y(n20772),
	.A(n21114));
   NAND2x1_ASAP7_75t_SL U16948 (.Y(n18174),
	.A(FE_OFN28688_sa22_2),
	.B(n23183));
   NOR3x1_ASAP7_75t_L U16949 (.Y(n22277),
	.A(n23160),
	.B(FE_OFN16135_sa22_4),
	.C(n21123));
   NAND2xp33_ASAP7_75t_SL U16950 (.Y(n21774),
	.A(n21094),
	.B(n23325));
   NAND3xp33_ASAP7_75t_L U16951 (.Y(n21129),
	.A(n18176),
	.B(n18177),
	.C(FE_OCPN29269_sa22_1));
   NAND2xp5_ASAP7_75t_L U16952 (.Y(n22317),
	.A(n23315),
	.B(n18162));
   NAND2xp5_ASAP7_75t_SL U16954 (.Y(n18544),
	.A(n18524),
	.B(FE_OFN29021_sa20_3));
   NAND3x2_ASAP7_75t_SL U16955 (.Y(n21637),
	.A(FE_OFN28987_n18597),
	.B(FE_OFN29200_n18521),
	.C(FE_OCPN27542_sa20_3));
   NAND2xp33_ASAP7_75t_SL U16956 (.Y(n23697),
	.A(n23692),
	.B(n23694));
   NAND2xp33_ASAP7_75t_SL U16957 (.Y(n23696),
	.A(n23695),
	.B(n23694));
   NOR3x1_ASAP7_75t_SL U16958 (.Y(n23693),
	.A(n18571),
	.B(FE_OFN28791_n),
	.C(n23838));
   NAND2xp5_ASAP7_75t_L U16959 (.Y(n23753),
	.A(n18540),
	.B(n23869));
   NOR3xp33_ASAP7_75t_L U16961 (.Y(n18603),
	.A(n23838),
	.B(n18536),
	.C(n18602));
   NOR2xp67_ASAP7_75t_L U16962 (.Y(n21690),
	.A(n21193),
	.B(n23693));
   NAND2x1p5_ASAP7_75t_SL U16963 (.Y(n18551),
	.A(n18522),
	.B(FE_OCPN29379_sa20_1));
   NAND2x1p5_ASAP7_75t_SL U16965 (.Y(n23689),
	.A(FE_OCPN27558_sa20_4),
	.B(FE_OFN16368_n18545));
   NAND3xp33_ASAP7_75t_SRAM U16966 (.Y(n16717),
	.A(FE_OFN29164_sa33_2),
	.B(FE_OCPN27782_n16873),
	.C(n16427));
   NOR2xp33_ASAP7_75t_L U16967 (.Y(n16910),
	.A(n26122),
	.B(n18141));
   NOR3xp33_ASAP7_75t_L U16968 (.Y(n19303),
	.A(n22008),
	.B(n20931),
	.C(n26154));
   NOR2xp67_ASAP7_75t_SL U16969 (.Y(n22020),
	.A(n22004),
	.B(n19327));
   NOR2xp33_ASAP7_75t_R U16971 (.Y(n17347),
	.A(FE_OFN29135_n21551),
	.B(FE_OFN16252_n27003));
   NAND2x1p5_ASAP7_75t_SL U16973 (.Y(n25054),
	.A(FE_OCPN28217_sa01_5),
	.B(FE_OCPN27712_sa01_4));
   NOR2xp33_ASAP7_75t_SL U16975 (.Y(n18694),
	.A(n22438),
	.B(n20388));
   NOR3xp33_ASAP7_75t_L U16976 (.Y(n17381),
	.A(n17330),
	.B(FE_OCPN27423_sa01_0),
	.C(n17345));
   NAND2xp5_ASAP7_75t_SL U16977 (.Y(n17375),
	.A(FE_OCPN29409_n22461),
	.B(FE_OFN29135_n21551));
   NOR2x1_ASAP7_75t_SL U16978 (.Y(n20404),
	.A(FE_OCPN29475_n25054),
	.B(n18693));
   NOR2x1_ASAP7_75t_L U16979 (.Y(n22177),
	.A(FE_OFN27152_n17315),
	.B(FE_OFN60_n27007));
   NAND3xp33_ASAP7_75t_R U16980 (.Y(n22468),
	.A(FE_OCPN29409_n22461),
	.B(n21553),
	.C(n17326));
   NAND2xp33_ASAP7_75t_SRAM U16981 (.Y(n23103),
	.A(n23059),
	.B(FE_OFN28594_n26454));
   NAND2x1_ASAP7_75t_R U16982 (.Y(n17916),
	.A(FE_OCPN29493_sa12_4),
	.B(FE_OCPN29485_sa12_3));
   NOR2xp33_ASAP7_75t_SL U16983 (.Y(n23605),
	.A(n23603),
	.B(n23602));
   NAND2xp33_ASAP7_75t_L U16984 (.Y(n23607),
	.A(n23601),
	.B(n23604));
   NOR2xp33_ASAP7_75t_R U16985 (.Y(n23601),
	.A(FE_OCPN5137_n23600),
	.B(n23602));
   NAND2xp5_ASAP7_75t_R U16987 (.Y(n20797),
	.A(FE_OFN28739_n17898),
	.B(FE_OCPN28386_n17899));
   NOR3x1_ASAP7_75t_SL U16990 (.Y(n23590),
	.A(FE_OFN27145_n23216),
	.B(FE_OFN25908_sa12_2),
	.C(FE_OCPN28248_n17971));
   NAND2xp5_ASAP7_75t_L U16991 (.Y(n19941),
	.A(n18847),
	.B(n17527));
   OAI21xp5_ASAP7_75t_L U16992 (.Y(n17557),
	.A1(FE_OCPN29348_n17592),
	.A2(n17700),
	.B(n18299));
   NAND3xp33_ASAP7_75t_SL U16993 (.Y(n18795),
	.A(n24867),
	.B(n24872),
	.C(n18839));
   NAND3xp33_ASAP7_75t_SL U16994 (.Y(n17873),
	.A(n16760),
	.B(FE_OCPN28298_n),
	.C(FE_OCPN29265_FE_OFN28698_sa21_1));
   NAND3xp33_ASAP7_75t_R U16995 (.Y(n20008),
	.A(n16771),
	.B(n19979),
	.C(FE_OCPN27289_sa21_5));
   NAND2xp5_ASAP7_75t_SL U16996 (.Y(n20289),
	.A(FE_OFN28678_sa21_3),
	.B(FE_OCPN27388_FE_OFN25990_sa21_4));
   NOR3xp33_ASAP7_75t_L U16997 (.Y(n17833),
	.A(FE_OFN27140_n20007),
	.B(FE_OCPN5083_sa21_2),
	.C(n17860));
   NAND2xp5_ASAP7_75t_SL U16999 (.Y(n20866),
	.A(n16399),
	.B(n16398));
   INVx1_ASAP7_75t_L U17000 (.Y(n16399),
	.A(n16490));
   NAND2xp33_ASAP7_75t_SL U17001 (.Y(n16334),
	.A(n24181),
	.B(n16303));
   NAND2xp5_ASAP7_75t_L U17002 (.Y(n25875),
	.A(n19425),
	.B(n19424));
   NAND2xp5_ASAP7_75t_L U17003 (.Y(n20559),
	.A(n24592),
	.B(n20812));
   NAND2xp33_ASAP7_75t_SL U17004 (.Y(n19651),
	.A(n19650),
	.B(n19649));
   NAND2xp33_ASAP7_75t_SL U17005 (.Y(n19652),
	.A(n19648),
	.B(n19649));
   NAND2x1_ASAP7_75t_SL U17008 (.Y(n19429),
	.A(n19425),
	.B(n20532));
   NOR2x1_ASAP7_75t_L U17009 (.Y(n16479),
	.A(FE_OCPN29438_sa33_2),
	.B(n17418));
   NOR3xp33_ASAP7_75t_SL U17010 (.Y(n16434),
	.A(FE_OCPN27568_sa33_3),
	.B(FE_OFN28694_sa33_4),
	.C(FE_OFN28679_sa33_5));
   NOR2x1_ASAP7_75t_L U17011 (.Y(n16854),
	.A(FE_OFN26055_n),
	.B(n16676));
   OAI21xp33_ASAP7_75t_L U17012 (.Y(n16449),
	.A1(FE_OCPN28127_n16872),
	.A2(n16925),
	.B(n16707));
   NOR2xp33_ASAP7_75t_L U17015 (.Y(n14036),
	.A(n15349),
	.B(FE_OFN16210_n13876));
   OA21x2_ASAP7_75t_L U17016 (.Y(n14037),
	.A1(n15319),
	.A2(n13875),
	.B(n14034));
   O2A1O1Ixp33_ASAP7_75t_L U17017 (.Y(n14034),
	.A1(n15729),
	.A2(n12994),
	.B(n14303),
	.C(n14033));
   NAND2xp33_ASAP7_75t_L U17018 (.Y(n14033),
	.A(n14032),
	.B(n14031));
   NAND2xp33_ASAP7_75t_L U17019 (.Y(n14031),
	.A(n14030),
	.B(FE_OFN28600_n14289));
   INVxp33_ASAP7_75t_L U17020 (.Y(n14205),
	.A(n14202));
   OA21x2_ASAP7_75t_L U17021 (.Y(n14198),
	.A1(FE_OFN16195_n13771),
	.A2(n15797),
	.B(n14195));
   NOR2xp33_ASAP7_75t_R U17022 (.Y(n13837),
	.A(FE_OFN28856_n15450),
	.B(FE_OFN26007_n16010));
   NAND3xp33_ASAP7_75t_SRAM U17023 (.Y(n13834),
	.A(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(n15934),
	.C(FE_OFN28883_n));
   NAND2xp5_ASAP7_75t_SL U17024 (.Y(n15679),
	.A(n14804),
	.B(n15339));
   NAND2xp5_ASAP7_75t_L U17026 (.Y(n14351),
	.A(FE_OFN28909_w3_23),
	.B(n14310));
   NOR2xp33_ASAP7_75t_R U17027 (.Y(n14352),
	.A(FE_OFN27066_n13869),
	.B(n14350));
   NAND2xp33_ASAP7_75t_R U17028 (.Y(n14350),
	.A(n14349),
	.B(n14348));
   NAND2xp33_ASAP7_75t_SRAM U17029 (.Y(n14348),
	.A(n14371),
	.B(FE_OFN28600_n14289));
   NAND2xp33_ASAP7_75t_SRAM U17030 (.Y(n14349),
	.A(n14377),
	.B(FE_OFN28600_n14289));
   NOR2xp33_ASAP7_75t_R U17031 (.Y(n15850),
	.A(n15841),
	.B(n15840));
   NOR3xp33_ASAP7_75t_SRAM U17032 (.Y(n15844),
	.A(n15842),
	.B(FE_OCPN8252_FE_OFN28661_w3_7),
	.C(FE_OFN25900_w3_4));
   INVxp33_ASAP7_75t_SRAM U17033 (.Y(n15852),
	.A(n15851));
   NAND2xp5_ASAP7_75t_R U17034 (.Y(n14114),
	.A(n15414),
	.B(n14112));
   NOR2xp33_ASAP7_75t_SRAM U17035 (.Y(n14125),
	.A(FE_OFN29017_n15921),
	.B(n14126));
   NOR2xp33_ASAP7_75t_R U17036 (.Y(n14128),
	.A(n15375),
	.B(n14126));
   NAND2xp33_ASAP7_75t_SRAM U17037 (.Y(n14131),
	.A(n15438),
	.B(n15954));
   NOR3xp33_ASAP7_75t_SRAM U17038 (.Y(n14137),
	.A(n15423),
	.B(FE_OCPN29535_FE_OFN8_w3_14),
	.C(n14912));
   NOR2xp33_ASAP7_75t_SRAM U17039 (.Y(n14165),
	.A(w3_8_),
	.B(n25051));
   NOR2xp33_ASAP7_75t_R U17040 (.Y(n14154),
	.A(FE_OCPN28296_n15386),
	.B(n14152));
   OAI22xp33_ASAP7_75t_SRAM U17041 (.Y(n14932),
	.A1(FE_OFN27115_n),
	.A2(FE_OCPN29508_FE_OFN16184_w3_9),
	.B1(FE_OCPN29535_FE_OFN8_w3_14),
	.B2(FE_OCPN29508_FE_OFN16184_w3_9));
   NOR2x1_ASAP7_75t_L U17042 (.Y(n14804),
	.A(n15338),
	.B(n14289));
   NOR3xp33_ASAP7_75t_SRAM U17043 (.Y(n14790),
	.A(FE_OFN29192_n13870),
	.B(FE_OFN26114_n),
	.C(n15484));
   NAND2xp5_ASAP7_75t_L U17044 (.Y(n14784),
	.A(n14771),
	.B(n14770));
   NAND2xp33_ASAP7_75t_SRAM U17045 (.Y(n14770),
	.A(FE_OCPN28278_n15512),
	.B(FE_OFN27066_n13869));
   NAND2xp33_ASAP7_75t_R U17046 (.Y(n14771),
	.A(n14769),
	.B(FE_OFN27066_n13869));
   NOR2xp33_ASAP7_75t_SRAM U17047 (.Y(n14769),
	.A(FE_OFN25915_n15514),
	.B(n15713));
   OA21x2_ASAP7_75t_L U17048 (.Y(n14785),
	.A1(FE_OFN28683_w3_21),
	.A2(n15551),
	.B(n14782));
   NAND2xp5_ASAP7_75t_SL U17049 (.Y(n14782),
	.A(n14781),
	.B(n14780));
   NAND2xp33_ASAP7_75t_SL U17050 (.Y(n14781),
	.A(n14777),
	.B(n14776));
   NAND2xp5_ASAP7_75t_L U17051 (.Y(n14766),
	.A(FE_OFN4_w3_22),
	.B(FE_OFN28706_n));
   NAND2xp33_ASAP7_75t_L U17052 (.Y(n15255),
	.A(FE_OFN27212_w3_30),
	.B(FE_OFN28929_n15182));
   NOR2xp33_ASAP7_75t_L U17053 (.Y(n13290),
	.A(n15185),
	.B(n14535));
   OAI21xp33_ASAP7_75t_L U17055 (.Y(n14214),
	.A1(n25140),
	.A2(FE_OFN28732_n),
	.B(FE_OCPN29537_FE_OFN28699_w3_6));
   AND2x2_ASAP7_75t_R U17056 (.Y(n13762),
	.A(n13755),
	.B(n13754));
   NAND2xp33_ASAP7_75t_SRAM U17057 (.Y(n13755),
	.A(n14410),
	.B(n15615));
   NAND2xp33_ASAP7_75t_R U17058 (.Y(n13754),
	.A(n13753),
	.B(n15615));
   NOR2xp33_ASAP7_75t_R U17059 (.Y(n13753),
	.A(FE_OFN26057_w3_1),
	.B(n15592));
   NOR2xp33_ASAP7_75t_SL U17060 (.Y(n15841),
	.A(n13741),
	.B(n15813));
   NOR2xp33_ASAP7_75t_SL U17062 (.Y(n13981),
	.A(n14941),
	.B(n14951));
   NOR2xp33_ASAP7_75t_L U17064 (.Y(n13987),
	.A(FE_OFN25985_n15997),
	.B(n13985));
   NAND3xp33_ASAP7_75t_L U17065 (.Y(n13966),
	.A(n15936),
	.B(n15956),
	.C(n15934));
   NAND2xp33_ASAP7_75t_L U17066 (.Y(n13922),
	.A(n13921),
	.B(n13920));
   NOR2xp33_ASAP7_75t_R U17067 (.Y(n13921),
	.A(FE_OFN27066_n13869),
	.B(n15281));
   NAND2xp33_ASAP7_75t_SL U17068 (.Y(n13923),
	.A(n13919),
	.B(n13920));
   NOR2xp33_ASAP7_75t_R U17069 (.Y(n13919),
	.A(n13915),
	.B(n15281));
   OAI22xp33_ASAP7_75t_SRAM U17070 (.Y(n13915),
	.A1(FE_OFN4_w3_22),
	.A2(n15341),
	.B1(FE_OFN26538_w3_19),
	.B2(n15341));
   NOR3xp33_ASAP7_75t_L U17071 (.Y(n15184),
	.A(FE_OFN27222_n14593),
	.B(FE_OFN27210_w3_30),
	.C(FE_OFN26049_w3_27));
   A2O1A1Ixp33_ASAP7_75t_L U17072 (.Y(n14864),
	.A1(n13736),
	.A2(n15835),
	.B(n14837),
	.C(FE_OFN26645_n));
   NAND2xp33_ASAP7_75t_SRAM U17073 (.Y(n14870),
	.A(n14869),
	.B(n14868));
   NOR2xp33_ASAP7_75t_SRAM U17074 (.Y(n14869),
	.A(n15079),
	.B(n14867));
   NAND2xp33_ASAP7_75t_R U17075 (.Y(n14871),
	.A(n14866),
	.B(n14868));
   NOR2xp33_ASAP7_75t_SRAM U17076 (.Y(n14866),
	.A(FE_OFN28831_n15838),
	.B(n14867));
   NOR2xp33_ASAP7_75t_R U17078 (.Y(n13851),
	.A(n15975),
	.B(n15983));
   NOR2xp33_ASAP7_75t_L U17079 (.Y(n15451),
	.A(n15414),
	.B(n13805));
   NAND2xp5_ASAP7_75t_SL U17080 (.Y(n15431),
	.A(FE_OFN29017_n15921),
	.B(n14622));
   OAI22xp5_ASAP7_75t_L U17081 (.Y(n14623),
	.A1(n15455),
	.A2(n14100),
	.B1(FE_OFN28574_n16016),
	.B2(n14100));
   NAND3xp33_ASAP7_75t_R U17082 (.Y(n14143),
	.A(FE_OFN26635_w3_14),
	.B(FE_OCPN29520_n24755),
	.C(n15922));
   NOR2xp33_ASAP7_75t_L U17083 (.Y(n15286),
	.A(FE_OFN37_w3_23),
	.B(n15280));
   NOR2x1p5_ASAP7_75t_L U17084 (.Y(n15536),
	.A(FE_OFN26539_w3_19),
	.B(FE_OFN28706_n));
   INVxp67_ASAP7_75t_L U17085 (.Y(n13398),
	.A(n13395));
   NAND2xp33_ASAP7_75t_SRAM U17086 (.Y(n13394),
	.A(FE_OFN16412_w3_26),
	.B(FE_OFN16193_n15200));
   INVxp33_ASAP7_75t_L U17087 (.Y(n13365),
	.A(n13361));
   OAI21xp33_ASAP7_75t_SRAM U17088 (.Y(n13338),
	.A1(FE_OFN25893_n15214),
	.A2(n13335),
	.B(n14503));
   INVxp33_ASAP7_75t_SRAM U17089 (.Y(n14997),
	.A(n15822));
   NOR2xp33_ASAP7_75t_SL U17090 (.Y(n15596),
	.A(n13729),
	.B(n15813));
   NOR2xp33_ASAP7_75t_L U17092 (.Y(n15032),
	.A(n14439),
	.B(n14221));
   NAND2xp33_ASAP7_75t_L U17093 (.Y(n15036),
	.A(n15035),
	.B(FE_OFN25918_n15813));
   NOR2xp33_ASAP7_75t_R U17094 (.Y(n15872),
	.A(n13736),
	.B(FE_OFN25928_n15779));
   NOR3xp33_ASAP7_75t_R U17095 (.Y(n15871),
	.A(n13730),
	.B(FE_OFN28661_w3_7),
	.C(n15080));
   NOR2xp33_ASAP7_75t_SL U17096 (.Y(n15382),
	.A(n15993),
	.B(n14645));
   OAI21xp33_ASAP7_75t_L U17097 (.Y(n15385),
	.A1(FE_OCPN29535_FE_OFN8_w3_14),
	.A2(n16012),
	.B(n14924));
   NOR3xp33_ASAP7_75t_SRAM U17099 (.Y(n14645),
	.A(FE_OFN26639_w3_14),
	.B(FE_OCPN28407_FE_OFN16433_w3_11),
	.C(FE_OCPN29506_FE_OFN16184_w3_9));
   NAND3xp33_ASAP7_75t_SL U17100 (.Y(n15958),
	.A(FE_OCPN29583_n15422),
	.B(FE_OFN25961_w3_8),
	.C(w3_10_));
   INVxp67_ASAP7_75t_R U17101 (.Y(n15418),
	.A(n15415));
   NAND3xp33_ASAP7_75t_R U17102 (.Y(n14316),
	.A(FE_OFN28628_n15667),
	.B(n15349),
	.C(FE_OFN16426_w3_20));
   OAI21xp33_ASAP7_75t_L U17103 (.Y(n14270),
	.A1(n14061),
	.A2(n15491),
	.B(n14265));
   NOR3xp33_ASAP7_75t_SRAM U17104 (.Y(n14264),
	.A(n13890),
	.B(FE_OFN28701_w3_16),
	.C(FE_OFN50_w3_18));
   OA21x2_ASAP7_75t_L U17105 (.Y(n14272),
	.A1(n14268),
	.A2(n15710),
	.B(n14267));
   OAI22xp33_ASAP7_75t_SRAM U17106 (.Y(n14268),
	.A1(FE_OFN5_w3_22),
	.A2(n15487),
	.B1(FE_OCPN29578_FE_OFN27214_w3_17),
	.B2(n15487));
   NOR3xp33_ASAP7_75t_SRAM U17107 (.Y(n14266),
	.A(FE_OFN16211_n13876),
	.B(FE_OFN28701_w3_16),
	.C(FE_OFN50_w3_18));
   NAND2xp33_ASAP7_75t_L U17108 (.Y(n15236),
	.A(FE_OFN27206_w3_30),
	.B(FE_OFN26049_w3_27));
   OAI21xp5_ASAP7_75t_L U17109 (.Y(n15196),
	.A1(FE_OFN27210_w3_30),
	.A2(FE_OFN26049_w3_27),
	.B(n13556));
   NAND2xp33_ASAP7_75t_L U17110 (.Y(n13444),
	.A(n13443),
	.B(n13442));
   NOR2xp33_ASAP7_75t_SRAM U17111 (.Y(n15569),
	.A(FE_OFN29052_w3_5),
	.B(FE_OCPN8252_FE_OFN28661_w3_7));
   OAI21xp33_ASAP7_75t_SRAM U17112 (.Y(n15575),
	.A1(n24831),
	.A2(FE_OCPN29537_FE_OFN28699_w3_6),
	.B(n15787));
   OAI22xp5_ASAP7_75t_L U17113 (.Y(n14957),
	.A1(FE_OFN29125_n),
	.A2(FE_OCPN29535_FE_OFN8_w3_14),
	.B1(FE_OCPN29508_FE_OFN16184_w3_9),
	.B2(FE_OCPN29535_FE_OFN8_w3_14));
   NAND2xp33_ASAP7_75t_SL U17114 (.Y(n14922),
	.A(n14920),
	.B(n14919));
   NOR2xp33_ASAP7_75t_L U17115 (.Y(n14920),
	.A(FE_OCPN28296_n15386),
	.B(n15963));
   OAI22xp33_ASAP7_75t_L U17116 (.Y(n14930),
	.A1(FE_PSN8271_n15924),
	.A2(FE_OFN28758_n15422),
	.B1(FE_OFN27200_n),
	.B2(FE_OFN28758_n15422));
   NOR2xp33_ASAP7_75t_L U17117 (.Y(n14928),
	.A(FE_OCPN28402_w3_13),
	.B(n24755));
   NAND2xp5_ASAP7_75t_L U17118 (.Y(n14933),
	.A(FE_OFN26641_w3_14),
	.B(n13844));
   NOR2xp33_ASAP7_75t_SL U17119 (.Y(n15978),
	.A(FE_OFN28898_n13805),
	.B(n16000));
   NOR3x1_ASAP7_75t_SL U17120 (.Y(n15739),
	.A(FE_OFN28706_n),
	.B(FE_OFN26539_w3_19),
	.C(FE_OFN26091_n24663));
   NAND2xp5_ASAP7_75t_SL U17121 (.Y(n15551),
	.A(n14774),
	.B(n14773));
   NOR2x1_ASAP7_75t_SL U17122 (.Y(n15501),
	.A(FE_OFN26535_w3_19),
	.B(FE_OFN28977_n));
   NOR3xp33_ASAP7_75t_SRAM U17123 (.Y(n15471),
	.A(FE_OCPN4685_n15658),
	.B(FE_OFN28909_w3_23),
	.C(n15739));
   NAND3x2_ASAP7_75t_L U17124 (.Y(n15197),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN26051_w3_27),
	.C(FE_OFN27211_w3_30));
   NOR2xp67_ASAP7_75t_L U17127 (.Y(n15814),
	.A(FE_OCPN28076_FE_OFN9_w3_6),
	.B(n15862));
   NOR2xp33_ASAP7_75t_SRAM U17128 (.Y(n15117),
	.A(n15859),
	.B(n15118));
   NOR2xp33_ASAP7_75t_SRAM U17129 (.Y(n15125),
	.A(n15838),
	.B(n15124));
   NAND3xp33_ASAP7_75t_SRAM U17130 (.Y(n15127),
	.A(n15567),
	.B(FE_OFN25900_w3_4),
	.C(n15857));
   NAND2xp33_ASAP7_75t_SRAM U17131 (.Y(n15115),
	.A(n24831),
	.B(n15787));
   NOR2xp33_ASAP7_75t_SRAM U17132 (.Y(n15110),
	.A(n15787),
	.B(n15864));
   NOR2xp33_ASAP7_75t_SRAM U17133 (.Y(n15112),
	.A(n15610),
	.B(n15864));
   NOR3xp33_ASAP7_75t_R U17134 (.Y(n15064),
	.A(n13771),
	.B(FE_OFN28695_n),
	.C(n13726));
   INVxp67_ASAP7_75t_R U17135 (.Y(n15065),
	.A(n15062));
   NOR3xp33_ASAP7_75t_SL U17136 (.Y(n15061),
	.A(FE_OFN26058_w3_1),
	.B(FE_OFN26591_w3_3),
	.C(FE_OFN26531_n));
   NOR2x1_ASAP7_75t_L U17137 (.Y(n16009),
	.A(FE_OCPN29534_FE_OFN8_w3_14),
	.B(FE_OFN27115_n));
   NOR3x1_ASAP7_75t_SL U17138 (.Y(n15660),
	.A(FE_OFN4_w3_22),
	.B(FE_OFN26538_w3_19),
	.C(FE_OFN27214_w3_17));
   OAI21xp5_ASAP7_75t_L U17139 (.Y(n15674),
	.A1(FE_OFN26053_n25415),
	.A2(FE_OFN28706_n),
	.B(FE_OFN5_w3_22));
   NOR3xp33_ASAP7_75t_L U17140 (.Y(n15666),
	.A(n13870),
	.B(FE_OFN28_w3_23),
	.C(n15665));
   NAND2x1p5_ASAP7_75t_L U17143 (.Y(n15257),
	.A(FE_OFN27211_w3_30),
	.B(FE_OCPN27656_w3_25));
   NOR2xp33_ASAP7_75t_L U17144 (.Y(n13665),
	.A(FE_OFN27210_w3_30),
	.B(n13551));
   OAI22xp33_ASAP7_75t_SRAM U17145 (.Y(n13669),
	.A1(n14557),
	.A2(n14514),
	.B1(FE_OFN27211_w3_30),
	.B2(n14514));
   INVxp67_ASAP7_75t_R U17146 (.Y(n14557),
	.A(FE_OCPN29547_n15183));
   NOR2xp33_ASAP7_75t_R U17147 (.Y(n14571),
	.A(FE_OFN27211_w3_30),
	.B(FE_OFN26049_w3_27));
   NAND2xp5_ASAP7_75t_L U17148 (.Y(n13648),
	.A(n15240),
	.B(n14579));
   NAND3xp33_ASAP7_75t_SRAM U17150 (.Y(n14441),
	.A(FE_OFN28721_n),
	.B(n15787),
	.C(n24831));
   NAND3xp33_ASAP7_75t_L U17151 (.Y(n14440),
	.A(FE_OCPN8252_FE_OFN28661_w3_7),
	.B(n14439),
	.C(FE_OFN28721_n));
   NAND3xp33_ASAP7_75t_L U17152 (.Y(n15848),
	.A(FE_OFN29052_w3_5),
	.B(FE_OFN28661_w3_7),
	.C(w3_4_));
   INVxp67_ASAP7_75t_L U17153 (.Y(n14431),
	.A(n14427));
   NOR2xp33_ASAP7_75t_L U17154 (.Y(n14846),
	.A(FE_OCPN29537_FE_OFN28699_w3_6),
	.B(n25140));
   NOR2xp33_ASAP7_75t_L U17155 (.Y(n15939),
	.A(n15455),
	.B(FE_OFN112_n15994));
   NAND2x1p5_ASAP7_75t_SL U17156 (.Y(n25328),
	.A(n18540),
	.B(FE_OFN28986_n18597));
   NAND3xp33_ASAP7_75t_L U17157 (.Y(n26879),
	.A(n24701),
	.B(n24700),
	.C(n24699));
   NAND2xp33_ASAP7_75t_R U17158 (.Y(n24700),
	.A(n24698),
	.B(n24697));
   NAND2xp33_ASAP7_75t_R U17159 (.Y(n24697),
	.A(n24696),
	.B(n24695));
   NAND2xp33_ASAP7_75t_SRAM U17160 (.Y(n24698),
	.A(n24693),
	.B(n24695));
   NAND3xp33_ASAP7_75t_R U17161 (.Y(n18892),
	.A(n21304),
	.B(n21295),
	.C(FE_OCPN29451_n));
   NAND2xp33_ASAP7_75t_SL U17162 (.Y(n18055),
	.A(n21024),
	.B(n18052));
   NAND3xp33_ASAP7_75t_SL U17164 (.Y(n26971),
	.A(n17763),
	.B(FE_OCPN27566_FE_OFN16138_sa02_5),
	.C(n17760));
   NAND2xp33_ASAP7_75t_R U17165 (.Y(n25790),
	.A(n25785),
	.B(n25787));
   NAND2xp33_ASAP7_75t_SRAM U17166 (.Y(n25789),
	.A(n25788),
	.B(n25787));
   NAND2xp5_ASAP7_75t_L U17167 (.Y(n25031),
	.A(n17685),
	.B(n18329));
   NAND2xp33_ASAP7_75t_SRAM U17168 (.Y(n18990),
	.A(FE_OCPN27743_n22009),
	.B(n26660));
   NAND2xp5_ASAP7_75t_L U17169 (.Y(n20565),
	.A(n23603),
	.B(n23587));
   NAND2xp5_ASAP7_75t_L U17170 (.Y(n20563),
	.A(n22222),
	.B(n20542));
   NOR2xp33_ASAP7_75t_SRAM U17171 (.Y(n24398),
	.A(n26282),
	.B(n24399));
   NAND2xp5_ASAP7_75t_SL U17172 (.Y(n25111),
	.A(n25110),
	.B(n25109));
   NOR2xp33_ASAP7_75t_SL U17173 (.Y(n25110),
	.A(n25108),
	.B(n25107));
   NAND2xp5_ASAP7_75t_SL U17174 (.Y(n25112),
	.A(n25106),
	.B(n25109));
   NOR2xp33_ASAP7_75t_SL U17175 (.Y(n25106),
	.A(FE_OCPN29467_n25102),
	.B(n25107));
   NAND2xp33_ASAP7_75t_L U17176 (.Y(n24259),
	.A(n24258),
	.B(n24883));
   NOR2xp33_ASAP7_75t_R U17177 (.Y(n24258),
	.A(FE_OFN28779_n24257),
	.B(n24256));
   NAND3xp33_ASAP7_75t_L U17178 (.Y(n24271),
	.A(n24269),
	.B(n24268),
	.C(n24921));
   NAND2xp5_ASAP7_75t_SL U17179 (.Y(n24786),
	.A(n24784),
	.B(n24783));
   NAND2xp33_ASAP7_75t_L U17180 (.Y(n24784),
	.A(n24778),
	.B(FE_OFN16326_n19058));
   NOR3xp33_ASAP7_75t_SRAM U17182 (.Y(n24793),
	.A(n24792),
	.B(n24791),
	.C(n24790));
   NOR2x1p5_ASAP7_75t_L U17183 (.Y(n24087),
	.A(n19817),
	.B(n17236));
   NAND2xp33_ASAP7_75t_SRAM U17186 (.Y(n22141),
	.A(FE_OFN25917_n21591),
	.B(FE_OFN27176_n));
   NAND2xp33_ASAP7_75t_SRAM U17187 (.Y(n19066),
	.A(FE_OFN28901_sa30_4),
	.B(FE_OCPN29398_sa30_3));
   NAND2xp33_ASAP7_75t_L U17188 (.Y(n19067),
	.A(n25103),
	.B(n22621));
   INVxp33_ASAP7_75t_L U17189 (.Y(n23278),
	.A(n23277));
   NOR2xp33_ASAP7_75t_SRAM U17190 (.Y(n23286),
	.A(FE_OFN28877_FE_OCPN27730_n17464),
	.B(n23281));
   AND3x1_ASAP7_75t_L U17191 (.Y(n23285),
	.A(n23284),
	.B(n23283),
	.C(n23282));
   NOR2xp33_ASAP7_75t_L U17192 (.Y(n23288),
	.A(n21854),
	.B(n24565));
   NOR3x1_ASAP7_75t_L U17193 (.Y(n22287),
	.A(n23303),
	.B(FE_OFN16135_sa22_4),
	.C(n21123));
   NAND2xp5_ASAP7_75t_SL U17194 (.Y(n23335),
	.A(n22295),
	.B(n22294));
   NOR3x1_ASAP7_75t_L U17196 (.Y(n23300),
	.A(n22310),
	.B(FE_OCPN27673_n18163),
	.C(n21123));
   NAND3xp33_ASAP7_75t_SRAM U17198 (.Y(n22693),
	.A(FE_OFN29215_n24262),
	.B(n22690),
	.C(n22689));
   NAND2xp33_ASAP7_75t_R U17199 (.Y(n22700),
	.A(n22695),
	.B(n22697));
   NOR2xp67_ASAP7_75t_L U17201 (.Y(n23765),
	.A(n21193),
	.B(n18535));
   NOR2xp33_ASAP7_75t_R U17202 (.Y(n18535),
	.A(n18534),
	.B(n20670));
   INVxp67_ASAP7_75t_R U17203 (.Y(n23767),
	.A(n23725));
   NOR2xp67_ASAP7_75t_SL U17204 (.Y(n23769),
	.A(FE_OCPN27606_n23869),
	.B(n23798));
   NAND2xp33_ASAP7_75t_L U17205 (.Y(n23812),
	.A(n23754),
	.B(n23753));
   NAND2xp5_ASAP7_75t_SRAM U17207 (.Y(n20510),
	.A(FE_OFN28801_n16978),
	.B(FE_OCPN27761_n16977));
   NOR3xp33_ASAP7_75t_SL U17208 (.Y(n20144),
	.A(FE_OCPN27838_n17747),
	.B(FE_OFN29210_FE_OCPN27261_sa02_0),
	.C(n17799));
   NAND2xp33_ASAP7_75t_L U17209 (.Y(n19272),
	.A(n22076),
	.B(n19255));
   NOR3xp33_ASAP7_75t_SL U17210 (.Y(n23031),
	.A(FE_OFN28832_n19789),
	.B(FE_OFN26160_sa10_4),
	.C(FE_OCPN29498_n16581));
   NAND3xp33_ASAP7_75t_SL U17211 (.Y(n23699),
	.A(n18583),
	.B(n18529),
	.C(FE_OFN29131_FE_OCPN27371_sa20_2));
   NOR2x1_ASAP7_75t_L U17213 (.Y(n23840),
	.A(n23677),
	.B(n20670));
   NAND2xp5_ASAP7_75t_SL U17214 (.Y(n21246),
	.A(n23753),
	.B(n25188));
   NOR2xp33_ASAP7_75t_SRAM U17216 (.Y(n26999),
	.A(n18698),
	.B(n22177));
   NOR2xp33_ASAP7_75t_L U17217 (.Y(n21558),
	.A(n18678),
	.B(n18714));
   NAND3xp33_ASAP7_75t_L U17220 (.Y(n22258),
	.A(n20600),
	.B(n20599),
	.C(n20598));
   NOR2xp33_ASAP7_75t_SRAM U17221 (.Y(n20600),
	.A(n24055),
	.B(n20596));
   NOR3xp33_ASAP7_75t_L U17222 (.Y(n20599),
	.A(n22248),
	.B(n23590),
	.C(n24363));
   NOR2x1_ASAP7_75t_SL U17223 (.Y(n20784),
	.A(n20554),
	.B(n22223));
   NAND2xp33_ASAP7_75t_R U17224 (.Y(n20578),
	.A(n20574),
	.B(n20575));
   NAND2xp33_ASAP7_75t_R U17225 (.Y(n20577),
	.A(n20576),
	.B(n20575));
   NAND2xp33_ASAP7_75t_SL U17226 (.Y(n16660),
	.A(n16656),
	.B(FE_OFN29153_n19753));
   NAND2xp33_ASAP7_75t_SL U17227 (.Y(n16659),
	.A(n16658),
	.B(FE_OFN29153_n19753));
   NOR2x1_ASAP7_75t_L U17231 (.Y(n23413),
	.A(FE_OFN29182_n21708),
	.B(FE_OFN27133_n21725));
   NOR3xp33_ASAP7_75t_SL U17232 (.Y(n21042),
	.A(n21725),
	.B(FE_OCPN27393_sa03_0),
	.C(n18040));
   NOR3xp33_ASAP7_75t_SRAM U17233 (.Y(n21070),
	.A(n23430),
	.B(n23447),
	.C(n21068));
   NAND2xp5_ASAP7_75t_L U17234 (.Y(n23432),
	.A(n18028),
	.B(n19449));
   NOR2xp33_ASAP7_75t_L U17235 (.Y(n18028),
	.A(n21023),
	.B(n21301));
   NOR2x1_ASAP7_75t_SL U17236 (.Y(n21751),
	.A(FE_OFN29182_n21708),
	.B(FE_OFN28955_n18011));
   NOR3xp33_ASAP7_75t_R U17237 (.Y(n23519),
	.A(FE_OFN28562_n19342),
	.B(FE_OFN25890_n23497),
	.C(n20265));
   NAND2xp33_ASAP7_75t_SL U17238 (.Y(n23513),
	.A(n19313),
	.B(FE_OCPN27953_n22945));
   NAND2xp5_ASAP7_75t_L U17239 (.Y(n25090),
	.A(n19019),
	.B(FE_OFN28752_n));
   OAI21xp5_ASAP7_75t_L U17241 (.Y(n26460),
	.A1(n23107),
	.A2(FE_OCPN28000_n22450),
	.B(n23104));
   NOR2xp33_ASAP7_75t_L U17243 (.Y(n16400),
	.A(FE_OCPN27516_n26292),
	.B(n18076));
   NOR2xp67_ASAP7_75t_R U17244 (.Y(n20060),
	.A(FE_OFN28719_n20025),
	.B(FE_OFN29147_sa31_1));
   NOR2xp33_ASAP7_75t_SL U17245 (.Y(n20325),
	.A(FE_OCPN27246_n22663),
	.B(FE_OFN28820_n));
   NOR2xp33_ASAP7_75t_SL U17246 (.Y(n22352),
	.A(n23643),
	.B(n20329));
   NAND2xp5_ASAP7_75t_SL U17247 (.Y(n20327),
	.A(n16771),
	.B(n16808));
   NAND3xp33_ASAP7_75t_L U17248 (.Y(n20288),
	.A(n22667),
	.B(n20002),
	.C(n19976));
   NOR2xp33_ASAP7_75t_SL U17249 (.Y(n16729),
	.A(n16937),
	.B(n23537));
   NAND2xp5_ASAP7_75t_L U17250 (.Y(n16725),
	.A(n16427),
	.B(n16946));
   NOR2x1_ASAP7_75t_L U17252 (.Y(n18939),
	.A(FE_OCPN27589_n25987),
	.B(n17087));
   NAND2xp5_ASAP7_75t_L U17253 (.Y(n17087),
	.A(n19372),
	.B(n18272));
   NOR2xp67_ASAP7_75t_R U17254 (.Y(n24156),
	.A(n19360),
	.B(n17115));
   NOR2x1_ASAP7_75t_SL U17255 (.Y(n18286),
	.A(n20527),
	.B(FE_OFN28738_n16989));
   NOR2x1_ASAP7_75t_SL U17256 (.Y(n20100),
	.A(n18789),
	.B(n17573));
   NAND2xp5_ASAP7_75t_SL U17257 (.Y(n17573),
	.A(n17581),
	.B(n19720));
   NAND2xp5_ASAP7_75t_L U17258 (.Y(n17542),
	.A(n17553),
	.B(FE_OCPN28245_n));
   NOR2xp33_ASAP7_75t_SRAM U17259 (.Y(n19380),
	.A(n16992),
	.B(n18932));
   NOR2xp33_ASAP7_75t_SL U17260 (.Y(n17172),
	.A(n20502),
	.B(n18276));
   NAND2xp5_ASAP7_75t_R U17262 (.Y(n17796),
	.A(n17795),
	.B(n17794));
   NAND2xp33_ASAP7_75t_L U17263 (.Y(n17795),
	.A(n17793),
	.B(n17792));
   NAND3xp33_ASAP7_75t_SL U17265 (.Y(n17713),
	.A(n19725),
	.B(n17527),
	.C(FE_OFN69_sa32_4));
   NAND2xp5_ASAP7_75t_SL U17266 (.Y(n21290),
	.A(n18897),
	.B(n18896));
   NAND2xp33_ASAP7_75t_SL U17267 (.Y(n18897),
	.A(n18894),
	.B(n18895));
   NAND2xp33_ASAP7_75t_R U17268 (.Y(n18896),
	.A(FE_OFN27125_n21057),
	.B(n18895));
   NAND2x1_ASAP7_75t_L U17272 (.Y(n21735),
	.A(n18039),
	.B(n23419));
   NOR3xp33_ASAP7_75t_L U17273 (.Y(n18039),
	.A(n23430),
	.B(n18038),
	.C(n21747));
   NOR3xp33_ASAP7_75t_L U17274 (.Y(n18038),
	.A(FE_OFN28949_n18011),
	.B(FE_OCPN27393_sa03_0),
	.C(FE_OFN141_sa03_1));
   NAND2xp5_ASAP7_75t_SL U17275 (.Y(n18869),
	.A(n18031),
	.B(n18892));
   NOR2xp33_ASAP7_75t_SL U17276 (.Y(n18031),
	.A(n21524),
	.B(n18008));
   NAND2xp5_ASAP7_75t_L U17277 (.Y(n23462),
	.A(n18007),
	.B(n18006));
   NAND2xp33_ASAP7_75t_SL U17278 (.Y(n18006),
	.A(n18005),
	.B(n18004));
   NAND2xp33_ASAP7_75t_L U17279 (.Y(n18007),
	.A(n18003),
	.B(n18004));
   NOR2x1_ASAP7_75t_SL U17281 (.Y(n18889),
	.A(n18879),
	.B(n21740));
   OAI21xp33_ASAP7_75t_R U17282 (.Y(n22893),
	.A1(n22083),
	.A2(n20962),
	.B(n22069));
   NAND2xp5_ASAP7_75t_L U17283 (.Y(n16576),
	.A(FE_OFN27196_n),
	.B(FE_OFN26161_sa10_4));
   INVxp67_ASAP7_75t_R U17284 (.Y(n16552),
	.A(n16597));
   NAND2x1p5_ASAP7_75t_L U17285 (.Y(n18652),
	.A(n19609),
	.B(FE_OCPN28389_n21479));
   NAND2xp5_ASAP7_75t_SL U17286 (.Y(n19835),
	.A(FE_OFN28835_n),
	.B(n19122));
   NOR3x1_ASAP7_75t_SL U17287 (.Y(n18746),
	.A(n19817),
	.B(FE_OCPN29385_n),
	.C(FE_OCPN29292_n18640));
   NAND2xp33_ASAP7_75t_L U17288 (.Y(n21452),
	.A(n21175),
	.B(n19574));
   NOR2xp33_ASAP7_75t_L U17290 (.Y(n19812),
	.A(n17297),
	.B(n18760));
   NAND2x1p5_ASAP7_75t_SL U17292 (.Y(n21442),
	.A(FE_OCPN29411_n),
	.B(n17274));
   NOR2x1_ASAP7_75t_L U17293 (.Y(n18752),
	.A(n19839),
	.B(n18776));
   NOR3x1_ASAP7_75t_SL U17294 (.Y(n18750),
	.A(FE_OCPN29291_n17282),
	.B(FE_OCPN29411_n),
	.C(FE_OFN26651_n19573));
   NOR3x1_ASAP7_75t_SL U17295 (.Y(n19818),
	.A(FE_OCPN27518_n17251),
	.B(FE_OCPN29411_n),
	.C(FE_OCPN29291_n17282));
   NAND2x1p5_ASAP7_75t_L U17296 (.Y(n21468),
	.A(FE_OFN16216_n19573),
	.B(FE_OCPN27819_n17245));
   NOR2xp67_ASAP7_75t_L U17298 (.Y(n18632),
	.A(FE_PSN8273_n24087),
	.B(n24086));
   NAND3xp33_ASAP7_75t_L U17299 (.Y(n18247),
	.A(FE_OCPN27902_n20514),
	.B(n25868),
	.C(FE_OCPN29351_FE_OFN26116_sa13_1));
   NOR2x1_ASAP7_75t_L U17300 (.Y(n20981),
	.A(FE_OCPN27919_n20155),
	.B(FE_OCPN27503_n20195));
   NAND3xp33_ASAP7_75t_SL U17301 (.Y(n26970),
	.A(n17763),
	.B(FE_OCPN27771_n19275),
	.C(FE_OFN28703_FE_OCPN27740_sa02_4));
   NAND2xp33_ASAP7_75t_R U17302 (.Y(n18925),
	.A(FE_OFN26170_n19361),
	.B(n19399));
   NOR2x1_ASAP7_75t_SL U17304 (.Y(n19438),
	.A(n17021),
	.B(n20529));
   NOR2xp33_ASAP7_75t_L U17305 (.Y(n20509),
	.A(n18276),
	.B(FE_OFN132_n18247));
   NOR2xp33_ASAP7_75t_L U17307 (.Y(n20500),
	.A(n19430),
	.B(n19429));
   NAND2xp5_ASAP7_75t_R U17308 (.Y(n25222),
	.A(FE_OFN28801_n16978),
	.B(n17060));
   NAND2x1_ASAP7_75t_SL U17309 (.Y(n20522),
	.A(n18272),
	.B(FE_OCPN29568_n18257));
   NOR3xp33_ASAP7_75t_R U17310 (.Y(n20525),
	.A(n17066),
	.B(n25990),
	.C(n19408));
   OAI21xp33_ASAP7_75t_SRAM U17311 (.Y(n17066),
	.A1(FE_OCPN29446_n17115),
	.A2(FE_OFN29243_n17065),
	.B(n25988));
   OAI21xp33_ASAP7_75t_L U17312 (.Y(n19462),
	.A1(FE_OCPN27733_n17996),
	.A2(FE_OCPN28184_n18020),
	.B(n23418));
   NOR2xp33_ASAP7_75t_SL U17313 (.Y(n19464),
	.A(n21752),
	.B(n18010));
   NAND2xp5_ASAP7_75t_L U17314 (.Y(n19480),
	.A(n18880),
	.B(FE_OFN16294_n19461));
   NOR2x1_ASAP7_75t_L U17315 (.Y(n21043),
	.A(FE_OCPN27675_n17986),
	.B(FE_OFN28952_n18011));
   NOR2xp33_ASAP7_75t_SL U17316 (.Y(n21068),
	.A(FE_OFN28677_n17998),
	.B(FE_OCPN27998_n18019));
   NAND2xp5_ASAP7_75t_L U17317 (.Y(n18048),
	.A(n21724),
	.B(n21271));
   NAND3xp33_ASAP7_75t_SL U17318 (.Y(n18041),
	.A(n21327),
	.B(n21708),
	.C(FE_OFN29124_n));
   NOR2x1_ASAP7_75t_SL U17320 (.Y(n19487),
	.A(n18904),
	.B(n21747));
   NOR2x1_ASAP7_75t_R U17321 (.Y(n21504),
	.A(FE_OCPN27675_n17986),
	.B(FE_OCPN27733_n17996));
   OAI21xp33_ASAP7_75t_L U17322 (.Y(n21280),
	.A1(n23431),
	.A2(n23430),
	.B(FE_OCPN29314_n));
   NAND3x1_ASAP7_75t_L U17323 (.Y(n23038),
	.A(n19685),
	.B(n19684),
	.C(n19683));
   NAND2xp5_ASAP7_75t_SL U17324 (.Y(n19684),
	.A(n19682),
	.B(FE_OFN28916_sa10_4));
   NAND2xp33_ASAP7_75t_SL U17325 (.Y(n19682),
	.A(n19681),
	.B(n19680));
   NOR2xp33_ASAP7_75t_SL U17327 (.Y(n17190),
	.A(n16648),
	.B(n19677));
   NOR2x1_ASAP7_75t_L U17328 (.Y(n16663),
	.A(n16565),
	.B(n19686));
   NOR2xp33_ASAP7_75t_L U17329 (.Y(n16580),
	.A(n21894),
	.B(n23132));
   NAND2xp5_ASAP7_75t_L U17330 (.Y(n16620),
	.A(n19788),
	.B(n19775));
   NOR2xp33_ASAP7_75t_L U17331 (.Y(n19671),
	.A(n16533),
	.B(n23982));
   NAND2xp5_ASAP7_75t_L U17332 (.Y(n17197),
	.A(FE_OFN130_sa10_5),
	.B(n23138));
   NOR2xp33_ASAP7_75t_L U17333 (.Y(n19781),
	.A(n23141),
	.B(n17196));
   NAND2xp33_ASAP7_75t_L U17334 (.Y(n17196),
	.A(n17195),
	.B(n21885));
   NOR3xp33_ASAP7_75t_SL U17335 (.Y(n19784),
	.A(n16619),
	.B(n23133),
	.C(n16640));
   NAND2xp5_ASAP7_75t_SL U17336 (.Y(n16619),
	.A(n19802),
	.B(n16618));
   OAI21xp33_ASAP7_75t_R U17337 (.Y(n23129),
	.A1(n17216),
	.A2(n19791),
	.B(FE_OCPN28157_n16534));
   NOR2xp33_ASAP7_75t_SL U17338 (.Y(n16632),
	.A(FE_OCPN5015_n23031),
	.B(n16548));
   NAND2xp33_ASAP7_75t_L U17339 (.Y(n16548),
	.A(n16637),
	.B(n17201));
   NAND2xp33_ASAP7_75t_SL U17340 (.Y(n16586),
	.A(n16585),
	.B(n16584));
   NAND2xp33_ASAP7_75t_SRAM U17341 (.Y(n16644),
	.A(n19788),
	.B(n23951));
   NOR2xp33_ASAP7_75t_SL U17342 (.Y(n16641),
	.A(FE_OCPN28358_n21899),
	.B(n19672));
   NOR2x1_ASAP7_75t_R U17343 (.Y(n23132),
	.A(FE_OFN29204_sa10_2),
	.B(n16616));
   NOR2x1_ASAP7_75t_L U17344 (.Y(n23131),
	.A(n16610),
	.B(n17191));
   NOR2x1_ASAP7_75t_SL U17345 (.Y(n23141),
	.A(n21902),
	.B(FE_OFN28832_n19789));
   OAI21xp5_ASAP7_75t_L U17346 (.Y(n19772),
	.A1(FE_OCPN27636_sa10_4),
	.A2(n16646),
	.B(n17219));
   NAND2xp5_ASAP7_75t_L U17347 (.Y(n19770),
	.A(n17216),
	.B(n16542));
   NAND3xp33_ASAP7_75t_SL U17348 (.Y(n19769),
	.A(FE_OCPN28040_n19766),
	.B(n23980),
	.C(FE_OFN27196_n));
   NAND3xp33_ASAP7_75t_SL U17349 (.Y(n23135),
	.A(n19766),
	.B(n24944),
	.C(FE_OFN27196_n));
   INVx1_ASAP7_75t_SL U17350 (.Y(n16650),
	.A(n16543));
   NAND3xp33_ASAP7_75t_SL U17351 (.Y(n19121),
	.A(n21468),
	.B(n21441),
	.C(n18639));
   NOR2xp33_ASAP7_75t_SRAM U17352 (.Y(n19143),
	.A(FE_OCPN28021_n21445),
	.B(n19144));
   OAI222xp33_ASAP7_75t_SL U17353 (.Y(n19131),
	.A1(FE_OCPN29463_n),
	.A2(FE_OCPN27588_n19824),
	.B1(n19609),
	.B2(FE_OCPN27588_n19824),
	.C1(FE_OCPN29542_n21151),
	.C2(FE_OCPN27588_n19824));
   NOR2xp33_ASAP7_75t_SL U17354 (.Y(n19113),
	.A(n19578),
	.B(n19106));
   NOR2x1p5_ASAP7_75t_SL U17356 (.Y(n17301),
	.A(FE_OCPN29284_n19821),
	.B(n17247));
   NOR2xp33_ASAP7_75t_L U17357 (.Y(n19087),
	.A(FE_OCPN27518_n17251),
	.B(n17300));
   NOR2x1_ASAP7_75t_L U17358 (.Y(n19150),
	.A(FE_OCPN27951_n19098),
	.B(FE_OCPN27518_n17251));
   NOR2xp33_ASAP7_75t_SL U17359 (.Y(n22147),
	.A(FE_OFN26037_n22144),
	.B(n22143));
   NAND2xp5_ASAP7_75t_L U17360 (.Y(n22124),
	.A(FE_OFN28513_n20470),
	.B(n19072));
   NOR2x1_ASAP7_75t_L U17362 (.Y(n22641),
	.A(FE_OCPN28027_n22125),
	.B(FE_OCPN27428_n26027));
   NOR2xp33_ASAP7_75t_L U17363 (.Y(n18499),
	.A(FE_OCPN29289_n22162),
	.B(n20440));
   NAND2x1p5_ASAP7_75t_L U17364 (.Y(n20470),
	.A(FE_OCPN29467_n25102),
	.B(FE_OFN25917_n21591));
   NAND2xp5_ASAP7_75t_L U17365 (.Y(n22636),
	.A(n18481),
	.B(n18489));
   NOR3x1_ASAP7_75t_R U17366 (.Y(n19222),
	.A(FE_OCPN29378_n23266),
	.B(n21844),
	.C(n17489));
   NOR2x1_ASAP7_75t_R U17367 (.Y(n19088),
	.A(n19817),
	.B(FE_OFN29079_FE_OCPN27518_n17251));
   NOR3xp33_ASAP7_75t_SL U17370 (.Y(n24097),
	.A(n17300),
	.B(FE_OCPN27818_n17267),
	.C(FE_PSN8289_FE_OFN28514_sa00_1));
   NAND3xp33_ASAP7_75t_SL U17371 (.Y(n19846),
	.A(n21468),
	.B(n19835),
	.C(n19828));
   AND3x1_ASAP7_75t_L U17372 (.Y(n19854),
	.A(n19095),
	.B(n18751),
	.C(n19595));
   NOR3xp33_ASAP7_75t_R U17373 (.Y(n18751),
	.A(n19836),
	.B(FE_PSN8290_n21439),
	.C(FE_PSN8284_n21438));
   NOR2x1_ASAP7_75t_L U17374 (.Y(n21150),
	.A(n19817),
	.B(n19097));
   NOR3xp33_ASAP7_75t_SL U17375 (.Y(n19847),
	.A(n17247),
	.B(FE_OFN29249_n),
	.C(n17298));
   NOR3xp33_ASAP7_75t_SL U17376 (.Y(n19828),
	.A(n17294),
	.B(n26100),
	.C(n26099));
   NAND3xp33_ASAP7_75t_SL U17377 (.Y(n17294),
	.A(n18752),
	.B(n21178),
	.C(n19592));
   NOR3x2_ASAP7_75t_L U17378 (.Y(n21834),
	.A(FE_OCPN29378_n23266),
	.B(FE_OFN28915_FE_OCPN27241_sa11_1),
	.C(n21844));
   NAND2x1_ASAP7_75t_L U17379 (.Y(n23250),
	.A(n17446),
	.B(n17453));
   NOR2x1_ASAP7_75t_SL U17380 (.Y(n23247),
	.A(FE_OCPN28175_n21818),
	.B(FE_OCPN27601_n17475));
   INVx1_ASAP7_75t_L U17381 (.Y(n21344),
	.A(n22486));
   NOR2xp33_ASAP7_75t_SL U17382 (.Y(n17512),
	.A(n22500),
	.B(n17470));
   NAND2xp5_ASAP7_75t_R U17383 (.Y(n17470),
	.A(n22487),
	.B(n23390));
   NOR2x1_ASAP7_75t_R U17384 (.Y(n21422),
	.A(FE_OCPN27313_n21845),
	.B(n21374));
   NAND2xp5_ASAP7_75t_L U17386 (.Y(n22504),
	.A(n23356),
	.B(FE_OCPN28417_n21396));
   NOR3x1_ASAP7_75t_SL U17387 (.Y(n22500),
	.A(FE_OCPN27313_n21845),
	.B(FE_OFN29137_FE_OCPN27228_sa11_2),
	.C(FE_OCPN27592_n17501));
   NAND3xp33_ASAP7_75t_L U17388 (.Y(n22490),
	.A(FE_OCPN28038_n23252),
	.B(n17446),
	.C(FE_OFN28915_FE_OCPN27241_sa11_1));
   NAND2xp5_ASAP7_75t_SL U17390 (.Y(n23378),
	.A(n21365),
	.B(n17447));
   NAND2xp5_ASAP7_75t_L U17391 (.Y(n23388),
	.A(n23387),
	.B(n23386));
   NAND3xp33_ASAP7_75t_SL U17393 (.Y(n23357),
	.A(n17473),
	.B(FE_OCPN27903_n19223),
	.C(n21366));
   NAND2x1p5_ASAP7_75t_L U17394 (.Y(n21851),
	.A(FE_OCPN27730_n17464),
	.B(n21365));
   NAND2xp5_ASAP7_75t_L U17395 (.Y(n18467),
	.A(n21596),
	.B(n22166));
   NOR3x1_ASAP7_75t_SL U17396 (.Y(n24759),
	.A(n18474),
	.B(FE_PSN8308_n22624),
	.C(n21597));
   NAND3xp33_ASAP7_75t_L U17397 (.Y(n18474),
	.A(n21596),
	.B(n22621),
	.C(n18472));
   NOR3xp33_ASAP7_75t_SRAM U17398 (.Y(n24760),
	.A(n22641),
	.B(n21586),
	.C(n26029));
   NAND2xp5_ASAP7_75t_SL U17399 (.Y(n24762),
	.A(n19082),
	.B(n18509));
   NOR2xp33_ASAP7_75t_R U17400 (.Y(n18509),
	.A(n18508),
	.B(FE_OCPN27764_n22152));
   NAND3xp33_ASAP7_75t_L U17401 (.Y(n24761),
	.A(n22138),
	.B(n18501),
	.C(n20431));
   NOR2x1_ASAP7_75t_L U17402 (.Y(n22156),
	.A(n18503),
	.B(FE_OFN29121_n26026));
   NOR3xp33_ASAP7_75t_SRAM U17403 (.Y(n20440),
	.A(FE_PSN8270_n26027),
	.B(FE_OFN28895_sa30_2),
	.C(n19051));
   NAND2xp5_ASAP7_75t_SL U17404 (.Y(n20438),
	.A(n22621),
	.B(n18475));
   NOR2xp33_ASAP7_75t_R U17405 (.Y(n20480),
	.A(n20471),
	.B(FE_OCPN27428_n26027));
   NAND2xp5_ASAP7_75t_R U17406 (.Y(n22633),
	.A(n22125),
	.B(n25108));
   NAND3xp33_ASAP7_75t_L U17407 (.Y(n19047),
	.A(n17603),
	.B(n25108),
	.C(FE_OFN28895_sa30_2));
   NAND2x1_ASAP7_75t_SL U17410 (.Y(n21604),
	.A(n18483),
	.B(FE_OCPN29412_sa30_5));
   NAND2xp5_ASAP7_75t_SL U17411 (.Y(n23694),
	.A(FE_OFN28791_n),
	.B(n23725));
   NAND2xp5_ASAP7_75t_L U17412 (.Y(n23764),
	.A(n18549),
	.B(n21655));
   NOR2xp33_ASAP7_75t_SL U17413 (.Y(n18549),
	.A(n23864),
	.B(FE_OCPN28017_n18548));
   NOR2xp33_ASAP7_75t_L U17414 (.Y(n22307),
	.A(FE_OFN25941_n22857),
	.B(n21122));
   NAND3xp33_ASAP7_75t_SL U17415 (.Y(n20773),
	.A(FE_OCPN27750_n22293),
	.B(n18161),
	.C(FE_OFN28688_sa22_2));
   NAND3xp33_ASAP7_75t_L U17417 (.Y(n21135),
	.A(FE_OCPN27750_n22293),
	.B(n23336),
	.C(FE_OFN28688_sa22_2));
   NAND3xp33_ASAP7_75t_SL U17418 (.Y(n21134),
	.A(n23341),
	.B(n20733),
	.C(n22307));
   NOR3x1_ASAP7_75t_L U17419 (.Y(n21114),
	.A(n21772),
	.B(FE_OCPN27521_n18163),
	.C(FE_OFN29080_n22310));
   NAND2xp5_ASAP7_75t_SL U17422 (.Y(n21121),
	.A(n21104),
	.B(n21103));
   NAND2xp5_ASAP7_75t_L U17423 (.Y(n21104),
	.A(n21102),
	.B(n21101));
   NAND2xp33_ASAP7_75t_SL U17424 (.Y(n21102),
	.A(n21098),
	.B(n21099));
   NAND2xp33_ASAP7_75t_L U17425 (.Y(n21101),
	.A(n21100),
	.B(n21099));
   NAND2xp5_ASAP7_75t_SL U17426 (.Y(n22821),
	.A(n20774),
	.B(n23192));
   NAND2xp5_ASAP7_75t_L U17427 (.Y(n22854),
	.A(n22828),
	.B(n18159));
   NAND2xp5_ASAP7_75t_L U17429 (.Y(n22815),
	.A(n22810),
	.B(n22812));
   NAND2xp5_ASAP7_75t_L U17430 (.Y(n22814),
	.A(n22813),
	.B(n22812));
   NOR2x1_ASAP7_75t_L U17431 (.Y(n22295),
	.A(n22321),
	.B(n21107));
   NOR3xp33_ASAP7_75t_L U17432 (.Y(n21117),
	.A(FE_OFN29080_n22310),
	.B(FE_OCPN27521_n18163),
	.C(n18166));
   NOR2x1_ASAP7_75t_L U17433 (.Y(n18190),
	.A(FE_OCPN27979_FE_OFN16147_sa22_1),
	.B(n23192));
   NAND2xp5_ASAP7_75t_R U17434 (.Y(n20723),
	.A(n23322),
	.B(n23336));
   NOR2x1_ASAP7_75t_R U17436 (.Y(n21107),
	.A(n23160),
	.B(FE_OCPN29478_n23306));
   NOR2x1_ASAP7_75t_L U17437 (.Y(n21669),
	.A(FE_OFN28537_sa20_2),
	.B(n18551));
   NOR2xp33_ASAP7_75t_SL U17439 (.Y(n20626),
	.A(FE_OFN28988_n18597),
	.B(n21193));
   NOR2xp33_ASAP7_75t_SRAM U17440 (.Y(n20618),
	.A(FE_OCPN27715_n23875),
	.B(FE_OCPN29567_n23806));
   NOR2xp33_ASAP7_75t_SRAM U17441 (.Y(n20620),
	.A(n20617),
	.B(FE_OCPN29567_n23806));
   AND3x1_ASAP7_75t_L U17442 (.Y(n21659),
	.A(n21656),
	.B(n21655),
	.C(n23685));
   NOR2xp33_ASAP7_75t_R U17443 (.Y(n23728),
	.A(n23725),
	.B(n23724));
   NAND3xp33_ASAP7_75t_R U17445 (.Y(n23723),
	.A(n23722),
	.B(FE_OCPN5110_n23721),
	.C(n23720));
   NAND3xp33_ASAP7_75t_SRAM U17446 (.Y(n21663),
	.A(n23869),
	.B(n18521),
	.C(FE_OFN29251_n18536));
   NAND3xp33_ASAP7_75t_SL U17447 (.Y(n23865),
	.A(n23753),
	.B(n25188),
	.C(n21681));
   NAND2xp33_ASAP7_75t_SL U17448 (.Y(n21681),
	.A(n21680),
	.B(n21679));
   NAND2xp33_ASAP7_75t_SL U17449 (.Y(n21679),
	.A(n21678),
	.B(n21677));
   NAND2xp33_ASAP7_75t_L U17450 (.Y(n21680),
	.A(n21675),
	.B(n21677));
   NOR2x1_ASAP7_75t_L U17451 (.Y(n23863),
	.A(FE_OFN29131_FE_OCPN27371_sa20_2),
	.B(n21240));
   NAND2xp5_ASAP7_75t_L U17452 (.Y(n20691),
	.A(n20689),
	.B(n20688));
   NAND2xp33_ASAP7_75t_SL U17453 (.Y(n20688),
	.A(n20687),
	.B(n18570));
   NOR3x1_ASAP7_75t_L U17454 (.Y(n23855),
	.A(n20670),
	.B(FE_OFN28791_n),
	.C(FE_OCPN28163_FE_OFN99_sa20_5));
   NAND2xp5_ASAP7_75t_L U17455 (.Y(n16918),
	.A(FE_OFN28999_n16923),
	.B(n16705));
   NOR2x1_ASAP7_75t_L U17456 (.Y(n16852),
	.A(n16923),
	.B(FE_OFN29208_n16436));
   INVxp67_ASAP7_75t_R U17457 (.Y(n18408),
	.A(n24617));
   NOR2x1_ASAP7_75t_R U17459 (.Y(n16928),
	.A(FE_OFN29134_sa33_0),
	.B(n16423));
   NAND2xp33_ASAP7_75t_L U17460 (.Y(n16943),
	.A(n16939),
	.B(n16940));
   NAND2xp33_ASAP7_75t_L U17461 (.Y(n16942),
	.A(n16941),
	.B(n16940));
   NOR2x1_ASAP7_75t_L U17462 (.Y(n16960),
	.A(FE_OFN26545_n16447),
	.B(n16673));
   NAND3xp33_ASAP7_75t_SL U17463 (.Y(n23550),
	.A(n16854),
	.B(FE_OCPN27555_n16422),
	.C(FE_OCPN29391_FE_OFN29162_sa33_2));
   NAND3xp33_ASAP7_75t_L U17465 (.Y(n18136),
	.A(n16698),
	.B(n24614),
	.C(n16895));
   NAND2xp5_ASAP7_75t_L U17466 (.Y(n18134),
	.A(n16854),
	.B(FE_OCPN27555_n16422));
   NOR2xp33_ASAP7_75t_L U17468 (.Y(n23542),
	.A(n18107),
	.B(n16929));
   NAND2xp33_ASAP7_75t_L U17469 (.Y(n23554),
	.A(n23551),
	.B(n23550));
   NAND3xp33_ASAP7_75t_L U17470 (.Y(n16724),
	.A(n16424),
	.B(n16909),
	.C(FE_OCPN29487_FE_OFN28694_sa33_4));
   INVxp67_ASAP7_75t_R U17471 (.Y(n18420),
	.A(n16855));
   NOR2xp33_ASAP7_75t_SRAM U17472 (.Y(n16861),
	.A(FE_OFN29101_n16418),
	.B(n16859));
   OAI21xp33_ASAP7_75t_SL U17473 (.Y(n19458),
	.A1(FE_OFN29122_n),
	.A2(n19450),
	.B(n19449));
   NAND2x1p5_ASAP7_75t_SL U17474 (.Y(n20241),
	.A(n20256),
	.B(FE_OFN27127_sa23_3));
   OAI21xp5_ASAP7_75t_L U17475 (.Y(n20227),
	.A1(FE_OFN29187_FE_OCPN27571_n20235),
	.A2(FE_OCPN28266_n20920),
	.B(n22019));
   OAI21xp33_ASAP7_75t_R U17476 (.Y(n23483),
	.A1(FE_OCPN27955_n22945),
	.A2(n18970),
	.B(FE_OFN28752_n));
   NAND3xp33_ASAP7_75t_L U17477 (.Y(n22990),
	.A(FE_OCPN27627_sa23_1),
	.B(n18971),
	.C(FE_OCPN29551_n));
   NAND2xp33_ASAP7_75t_L U17478 (.Y(n20277),
	.A(n20273),
	.B(n20274));
   NAND2xp33_ASAP7_75t_R U17479 (.Y(n20276),
	.A(n20275),
	.B(n20274));
   NOR3xp33_ASAP7_75t_SL U17482 (.Y(n19342),
	.A(n20913),
	.B(FE_OCPN29441_sa23_4),
	.C(n22971));
   NOR2xp67_ASAP7_75t_SL U17483 (.Y(n22033),
	.A(FE_OCPN27627_sa23_1),
	.B(n18987));
   NAND2xp5_ASAP7_75t_R U17484 (.Y(n18987),
	.A(n18971),
	.B(FE_OFN16272_n24767));
   NOR2xp67_ASAP7_75t_L U17485 (.Y(n20255),
	.A(n18989),
	.B(n20911));
   NOR2xp33_ASAP7_75t_SL U17486 (.Y(n20262),
	.A(FE_OFN28580_n23491),
	.B(n20260));
   NAND2xp5_ASAP7_75t_L U17487 (.Y(n20264),
	.A(n20259),
	.B(n20261));
   NOR2xp33_ASAP7_75t_L U17488 (.Y(n20259),
	.A(FE_OFN29026_n20911),
	.B(n20260));
   NOR2x1_ASAP7_75t_SL U17489 (.Y(n22998),
	.A(FE_OCPN28266_n20920),
	.B(FE_OFN25889_n20913));
   NOR2x1p5_ASAP7_75t_SL U17490 (.Y(n20260),
	.A(FE_OCPN29488_FE_OFN25883_n22945),
	.B(n22010));
   NAND2xp5_ASAP7_75t_L U17491 (.Y(n22986),
	.A(FE_OCPN27881_FE_OFN27126_sa23_3),
	.B(n20255));
   OAI21xp33_ASAP7_75t_SL U17492 (.Y(n22988),
	.A1(FE_OCPN27916_n),
	.A2(n22969),
	.B(n20272));
   NOR2xp33_ASAP7_75t_SL U17493 (.Y(n18678),
	.A(FE_OCPN29320_n22461),
	.B(FE_OCPN27399_n22598));
   NAND2xp5_ASAP7_75t_SL U17494 (.Y(n22596),
	.A(n18681),
	.B(n18680));
   NAND2xp5_ASAP7_75t_R U17495 (.Y(n18680),
	.A(FE_OCPN29320_n22461),
	.B(FE_OCPN5188_n22414));
   NAND2xp33_ASAP7_75t_SL U17496 (.Y(n18681),
	.A(n18679),
	.B(FE_OCPN5188_n22414));
   NOR2xp33_ASAP7_75t_R U17497 (.Y(n23105),
	.A(FE_OCPN27871_n17317),
	.B(n23106));
   NAND3x1_ASAP7_75t_L U17498 (.Y(n22457),
	.A(FE_OCPN27871_n17317),
	.B(n17386),
	.C(FE_OFN26054_sa01_3));
   NOR2xp33_ASAP7_75t_SRAM U17499 (.Y(n23086),
	.A(FE_OCPN27988_n26454),
	.B(n23087));
   INVxp33_ASAP7_75t_SRAM U17500 (.Y(n23064),
	.A(n23060));
   AND2x2_ASAP7_75t_L U17501 (.Y(n23088),
	.A(n21558),
	.B(n17357));
   NOR3xp33_ASAP7_75t_SL U17502 (.Y(n17357),
	.A(n17356),
	.B(n22177),
	.C(n17355));
   INVxp67_ASAP7_75t_L U17504 (.Y(n17322),
	.A(n20365));
   NAND2xp5_ASAP7_75t_SL U17505 (.Y(n23104),
	.A(FE_OCPN27423_sa01_0),
	.B(n20360));
   NOR3xp33_ASAP7_75t_SL U17507 (.Y(n23102),
	.A(n22193),
	.B(n22602),
	.C(n22603));
   NOR2x1_ASAP7_75t_SL U17508 (.Y(n22588),
	.A(n21546),
	.B(n17381));
   NOR2xp33_ASAP7_75t_SRAM U17509 (.Y(n22591),
	.A(FE_OFN26648_n22197),
	.B(FE_OFN27052_n21551));
   OAI22xp33_ASAP7_75t_L U17510 (.Y(n22432),
	.A1(n23059),
	.A2(n18668),
	.B1(FE_OCPN29409_n22461),
	.B2(n18668));
   NOR2xp33_ASAP7_75t_SL U17511 (.Y(n18706),
	.A(n18678),
	.B(n17381));
   NOR2xp33_ASAP7_75t_SL U17512 (.Y(n18699),
	.A(n17331),
	.B(n21544));
   NOR3xp33_ASAP7_75t_SL U17513 (.Y(n22448),
	.A(n23101),
	.B(FE_OFN28736_FE_OCPN28216_sa01_5),
	.C(n18684));
   NAND2xp5_ASAP7_75t_R U17516 (.Y(n22235),
	.A(n19552),
	.B(n22227));
   NOR2x1_ASAP7_75t_SL U17517 (.Y(n24055),
	.A(n23215),
	.B(n23217));
   NOR2x1_ASAP7_75t_SL U17518 (.Y(n17953),
	.A(FE_OCPN29499_FE_OFN16131_sa12_1),
	.B(FE_OFN28931_n17897));
   NOR3xp33_ASAP7_75t_SL U17520 (.Y(n17954),
	.A(n19527),
	.B(FE_OCPN29493_sa12_4),
	.C(FE_OFN73_sa12_5));
   INVx1_ASAP7_75t_L U17521 (.Y(n19546),
	.A(n22223));
   NOR2x1_ASAP7_75t_L U17524 (.Y(n22734),
	.A(FE_OFN25907_sa12_2),
	.B(n19512));
   NAND3xp33_ASAP7_75t_SL U17525 (.Y(n22760),
	.A(n19533),
	.B(n23235),
	.C(n22771));
   NAND2xp33_ASAP7_75t_R U17526 (.Y(n19524),
	.A(n19523),
	.B(FE_OFN122_n22751));
   NAND2xp33_ASAP7_75t_R U17527 (.Y(n19525),
	.A(n19521),
	.B(FE_OFN122_n22751));
   NOR3xp33_ASAP7_75t_SL U17528 (.Y(n23611),
	.A(FE_OFN28520_n22753),
	.B(n22752),
	.C(FE_OFN28654_n22751));
   NOR3x1_ASAP7_75t_SL U17529 (.Y(n22781),
	.A(n17952),
	.B(FE_OFN28882_FE_OCPN27356_sa12_0),
	.C(n23217));
   NAND2xp5_ASAP7_75t_SL U17530 (.Y(n23236),
	.A(FE_OFN26125_n22742),
	.B(n25741));
   NOR2xp33_ASAP7_75t_SL U17531 (.Y(n22724),
	.A(n19527),
	.B(n17916));
   NAND3xp33_ASAP7_75t_SL U17532 (.Y(n20814),
	.A(n17906),
	.B(n24364),
	.C(FE_OCPN29485_sa12_3));
   NAND2xp5_ASAP7_75t_R U17533 (.Y(n22227),
	.A(FE_OCPN28198_n22776),
	.B(n23587));
   NAND2x1_ASAP7_75t_L U17534 (.Y(n27089),
	.A(n25869),
	.B(FE_OFN29234_n16996));
   NOR2xp33_ASAP7_75t_SL U17535 (.Y(n18842),
	.A(FE_OCPN29298_n25028),
	.B(n19920));
   NAND2xp5_ASAP7_75t_SL U17536 (.Y(n19954),
	.A(n19934),
	.B(n18800));
   NOR3xp33_ASAP7_75t_SL U17537 (.Y(n17579),
	.A(n18830),
	.B(n22375),
	.C(n24864));
   NOR3xp33_ASAP7_75t_L U17538 (.Y(n17691),
	.A(FE_OCPN29579_n18837),
	.B(FE_OCPN27230_sa32_3),
	.C(FE_OCPN27882_n18829));
   NAND3x1_ASAP7_75t_SL U17539 (.Y(n18321),
	.A(FE_OCPN28268_n19911),
	.B(n17529),
	.C(FE_OCPN27230_sa32_3));
   NAND2x1p5_ASAP7_75t_L U17540 (.Y(n19718),
	.A(n17540),
	.B(n17539));
   NAND2xp5_ASAP7_75t_SL U17541 (.Y(n17539),
	.A(n17538),
	.B(n17537));
   NAND2xp5_ASAP7_75t_SL U17542 (.Y(n17540),
	.A(n17536),
	.B(n17537));
   NOR2x1_ASAP7_75t_L U17543 (.Y(n24855),
	.A(FE_OFN28991_n19938),
	.B(FE_OCPN27267_n18794));
   NOR2x1_ASAP7_75t_L U17544 (.Y(n18820),
	.A(n22367),
	.B(n17593));
   NAND2xp5_ASAP7_75t_L U17545 (.Y(n17593),
	.A(n19941),
	.B(n19943));
   NAND3xp33_ASAP7_75t_SL U17546 (.Y(n18826),
	.A(FE_OFN26035_n),
	.B(n17525),
	.C(FE_OFN16463_sa32_0));
   NAND2x1_ASAP7_75t_L U17547 (.Y(n18830),
	.A(n22378),
	.B(n24866));
   NOR2xp33_ASAP7_75t_L U17549 (.Y(n18815),
	.A(n17557),
	.B(n17544));
   NAND2xp33_ASAP7_75t_L U17550 (.Y(n17544),
	.A(n17551),
	.B(n20093));
   NOR2x1_ASAP7_75t_R U17552 (.Y(n18325),
	.A(n20096),
	.B(n19703));
   NOR2x1_ASAP7_75t_L U17553 (.Y(n22396),
	.A(n19926),
	.B(n22370));
   NAND3xp33_ASAP7_75t_L U17554 (.Y(n22398),
	.A(n18844),
	.B(n24872),
	.C(n18843));
   NOR3xp33_ASAP7_75t_L U17555 (.Y(n18844),
	.A(n18842),
	.B(FE_OCPN27937_n18841),
	.C(n22369));
   NAND2xp33_ASAP7_75t_L U17556 (.Y(n22387),
	.A(n18840),
	.B(n18839));
   NAND2x1_ASAP7_75t_L U17557 (.Y(n22386),
	.A(n17522),
	.B(n17560));
   NAND2xp5_ASAP7_75t_SL U17558 (.Y(n22397),
	.A(n17525),
	.B(n19940));
   NOR3xp33_ASAP7_75t_L U17559 (.Y(n16768),
	.A(FE_OFN28820_n),
	.B(FE_OCPN29293_FE_OFN28678_sa21_3),
	.C(n16806));
   NOR3xp33_ASAP7_75t_L U17560 (.Y(n23661),
	.A(n22662),
	.B(FE_OCPN29414_n),
	.C(n16801));
   NAND2xp33_ASAP7_75t_R U17561 (.Y(n17850),
	.A(n17846),
	.B(n17847));
   NAND2xp5_ASAP7_75t_L U17562 (.Y(n20305),
	.A(FE_OFN29215_n24262),
	.B(n22690));
   NAND2xp33_ASAP7_75t_SL U17563 (.Y(n20329),
	.A(n19993),
	.B(n17873));
   NAND2xp5_ASAP7_75t_L U17564 (.Y(n19881),
	.A(n16776),
	.B(n16780));
   NAND2xp5_ASAP7_75t_L U17565 (.Y(n16780),
	.A(n16779),
	.B(FE_OFN28969_n19890));
   NAND3xp33_ASAP7_75t_L U17567 (.Y(n19885),
	.A(n19867),
	.B(n19889),
	.C(n22690));
   NAND3xp33_ASAP7_75t_L U17568 (.Y(n19978),
	.A(n20312),
	.B(n24918),
	.C(n20315));
   NAND3x1_ASAP7_75t_SL U17569 (.Y(n22354),
	.A(FE_OFN16153_n16747),
	.B(FE_OCPN28298_n),
	.C(FE_OCPN5126_sa21_2));
   NOR3xp33_ASAP7_75t_L U17570 (.Y(n20287),
	.A(n19982),
	.B(FE_OCPN29414_n),
	.C(n16801));
   NAND2x1_ASAP7_75t_L U17571 (.Y(n22349),
	.A(n19992),
	.B(n16775));
   NAND2xp5_ASAP7_75t_L U17572 (.Y(n16775),
	.A(FE_OCPN5126_sa21_2),
	.B(n22675));
   NAND3x1_ASAP7_75t_L U17573 (.Y(n22343),
	.A(FE_OFN16153_n16747),
	.B(FE_OFN16447_n16749),
	.C(FE_OCPN5126_sa21_2));
   NAND3xp33_ASAP7_75t_L U17574 (.Y(n17871),
	.A(n22665),
	.B(n19872),
	.C(n17862));
   NOR3xp33_ASAP7_75t_L U17575 (.Y(n17862),
	.A(n22696),
	.B(n17861),
	.C(n22676));
   NOR2x1_ASAP7_75t_R U17576 (.Y(n22356),
	.A(FE_OCPN29279_n25353),
	.B(FE_OFN28970_n19890));
   NAND2xp5_ASAP7_75t_L U17577 (.Y(n23651),
	.A(n16802),
	.B(n16814));
   NAND3xp33_ASAP7_75t_SL U17578 (.Y(n23652),
	.A(n22354),
	.B(n22353),
	.C(n22352));
   NAND3xp33_ASAP7_75t_SL U17579 (.Y(n22678),
	.A(n22343),
	.B(n20332),
	.C(FE_OFN29215_n24262));
   NAND2xp33_ASAP7_75t_R U17580 (.Y(n22683),
	.A(n22682),
	.B(n24917));
   NAND2xp33_ASAP7_75t_SRAM U17581 (.Y(n22684),
	.A(n22681),
	.B(n24917));
   NOR2xp67_ASAP7_75t_L U17584 (.Y(n21988),
	.A(FE_OCPN29483_FE_OFN26014_sa31_3),
	.B(FE_OFN27168_n16334));
   NOR3xp33_ASAP7_75t_SL U17585 (.Y(n20080),
	.A(n20079),
	.B(n20078),
	.C(n21968));
   NAND3xp33_ASAP7_75t_L U17586 (.Y(n20079),
	.A(n20882),
	.B(n20856),
	.C(n25315));
   NAND2xp5_ASAP7_75t_R U17587 (.Y(n21979),
	.A(FE_OFN29032_FE_OCPN27728_n21981),
	.B(n21946));
   NAND2xp5_ASAP7_75t_L U17588 (.Y(n16296),
	.A(FE_OCPN29526_sa31_4),
	.B(n16512));
   NAND2xp5_ASAP7_75t_L U17589 (.Y(n18085),
	.A(n25323),
	.B(FE_OFN26584_n20059));
   NAND2xp5_ASAP7_75t_L U17591 (.Y(n20833),
	.A(n25316),
	.B(n24182));
   NOR2x1_ASAP7_75t_SL U17592 (.Y(n16496),
	.A(FE_OCPN28314_n20842),
	.B(FE_OCPN28334_n16497));
   NOR2xp33_ASAP7_75t_L U17593 (.Y(n25848),
	.A(FE_OFN26095_n16293),
	.B(n16308));
   NAND2xp33_ASAP7_75t_SRAM U17594 (.Y(n16308),
	.A(n20050),
	.B(n16307));
   NAND2xp33_ASAP7_75t_R U17595 (.Y(n16307),
	.A(FE_OFN29147_sa31_1),
	.B(FE_OFN29136_n));
   NOR2xp33_ASAP7_75t_SL U17596 (.Y(n18078),
	.A(n26290),
	.B(n21988));
   NOR3x1_ASAP7_75t_SL U17597 (.Y(n16338),
	.A(n16305),
	.B(n16362),
	.C(n16304));
   NAND2xp5_ASAP7_75t_SL U17598 (.Y(n16305),
	.A(n24182),
	.B(n18079));
   NOR3xp33_ASAP7_75t_SL U17599 (.Y(n18094),
	.A(n16312),
	.B(n26402),
	.C(n16495));
   NAND2xp33_ASAP7_75t_SL U17600 (.Y(n16312),
	.A(n18068),
	.B(n21948));
   NOR2x1p5_ASAP7_75t_SL U17602 (.Y(n18096),
	.A(FE_OCPN29483_FE_OFN26014_sa31_3),
	.B(n16289));
   OAI21xp33_ASAP7_75t_L U17605 (.Y(n25225),
	.A1(FE_OCPN28204_n20526),
	.A2(n20527),
	.B(n16984));
   NAND3xp33_ASAP7_75t_SL U17606 (.Y(n25820),
	.A(n25818),
	.B(n25817),
	.C(n26302));
   NAND3xp33_ASAP7_75t_L U17608 (.Y(n22668),
	.A(n19979),
	.B(FE_OFN16153_n16747),
	.C(FE_OCPN27289_sa21_5));
   NAND2xp33_ASAP7_75t_R U17609 (.Y(n24674),
	.A(n24673),
	.B(FE_OFN131_sa10_6));
   NOR2xp33_ASAP7_75t_SRAM U17610 (.Y(n24673),
	.A(n24671),
	.B(FE_OFN59_sa10_7));
   NOR2xp33_ASAP7_75t_SRAM U17612 (.Y(n24645),
	.A(n17561),
	.B(n20095));
   NOR2xp33_ASAP7_75t_SRAM U17613 (.Y(n17561),
	.A(FE_OFN26553_n24644),
	.B(n19920));
   NAND2xp33_ASAP7_75t_R U17615 (.Y(n24860),
	.A(n24856),
	.B(FE_OFN26166_n24855));
   NAND2xp33_ASAP7_75t_SRAM U17616 (.Y(n24859),
	.A(n24858),
	.B(FE_OFN26166_n24855));
   NOR3xp33_ASAP7_75t_SRAM U17617 (.Y(n24871),
	.A(n24870),
	.B(n24869),
	.C(n24868));
   NAND3xp33_ASAP7_75t_SRAM U17618 (.Y(n24900),
	.A(n24898),
	.B(n24897),
	.C(n24896));
   INVxp33_ASAP7_75t_SRAM U17619 (.Y(n24898),
	.A(n24892));
   NAND2xp33_ASAP7_75t_L U17620 (.Y(n27041),
	.A(n21158),
	.B(n18625));
   NOR2xp33_ASAP7_75t_L U17621 (.Y(n25240),
	.A(FE_OCPN8234_n25199),
	.B(n25198));
   NAND2xp33_ASAP7_75t_SRAM U17622 (.Y(n25198),
	.A(n25197),
	.B(n25196));
   NOR3xp33_ASAP7_75t_SL U17623 (.Y(n25987),
	.A(FE_OCPN28202_n16991),
	.B(FE_OFN28862_n),
	.C(n17121));
   NOR2xp33_ASAP7_75t_L U17624 (.Y(n19408),
	.A(FE_OCPN28202_n16991),
	.B(FE_OCPN27836_n16976));
   NOR3x1_ASAP7_75t_SL U17625 (.Y(n16507),
	.A(n21981),
	.B(FE_OCPN29526_sa31_4),
	.C(FE_OFN28669_sa31_5));
   NOR3xp33_ASAP7_75t_L U17626 (.Y(n21934),
	.A(n16329),
	.B(FE_OCPN29482_FE_OFN26014_sa31_3),
	.C(n16340));
   NAND2xp5_ASAP7_75t_SL U17627 (.Y(n25399),
	.A(FE_OCPN29477_sa12_5),
	.B(n22724));
   NAND3xp33_ASAP7_75t_L U17628 (.Y(n16888),
	.A(n16417),
	.B(n16946),
	.C(FE_OFN25938_sa33_3));
   INVxp33_ASAP7_75t_SRAM U17629 (.Y(n26665),
	.A(n26661));
   NAND2xp33_ASAP7_75t_R U17630 (.Y(n14024),
	.A(n14020),
	.B(n14019));
   NAND2xp33_ASAP7_75t_L U17631 (.Y(n14023),
	.A(n14022),
	.B(n14019));
   OAI21xp33_ASAP7_75t_SRAM U17632 (.Y(n14021),
	.A1(FE_OFN5_w3_22),
	.A2(FE_OFN28712_n),
	.B(n14276));
   NOR2xp33_ASAP7_75t_R U17633 (.Y(n14025),
	.A(n15739),
	.B(n13875));
   NOR3xp33_ASAP7_75t_L U17634 (.Y(n14369),
	.A(FE_OFN26053_n25415),
	.B(FE_OFN5_w3_22),
	.C(FE_OFN28706_n));
   NAND3xp33_ASAP7_75t_SRAM U17635 (.Y(n14013),
	.A(FE_OFN5_w3_22),
	.B(n14774),
	.C(FE_OFN26539_w3_19));
   NOR2xp33_ASAP7_75t_R U17636 (.Y(n14015),
	.A(FE_OFN27096_n),
	.B(FE_OFN16211_n13876));
   NAND2xp5_ASAP7_75t_L U17637 (.Y(n14605),
	.A(n14497),
	.B(n14496));
   NAND2xp33_ASAP7_75t_L U17638 (.Y(n14496),
	.A(n14495),
	.B(n14494));
   OAI222xp33_ASAP7_75t_L U17639 (.Y(n14238),
	.A1(n14864),
	.A2(n15881),
	.B1(n14237),
	.B2(n15881),
	.C1(n14236),
	.C2(n15881));
   NAND2xp5_ASAP7_75t_L U17640 (.Y(n14237),
	.A(n14227),
	.B(n14226));
   NAND2xp5_ASAP7_75t_L U17641 (.Y(n14236),
	.A(n14235),
	.B(n14234));
   NAND2xp33_ASAP7_75t_L U17642 (.Y(n14226),
	.A(n14225),
	.B(n14224));
   NAND2xp33_ASAP7_75t_SRAM U17643 (.Y(n14209),
	.A(n15034),
	.B(n15609));
   NAND2xp33_ASAP7_75t_L U17644 (.Y(n14208),
	.A(n14203),
	.B(n14205));
   NOR2xp33_ASAP7_75t_SRAM U17645 (.Y(n14203),
	.A(n15810),
	.B(n14204));
   NAND2xp33_ASAP7_75t_L U17646 (.Y(n14207),
	.A(n14206),
	.B(n14205));
   NOR2xp33_ASAP7_75t_SRAM U17647 (.Y(n14206),
	.A(n15859),
	.B(n14204));
   NAND2xp33_ASAP7_75t_R U17648 (.Y(n14200),
	.A(n14199),
	.B(n14198));
   NOR2xp33_ASAP7_75t_SRAM U17649 (.Y(n14199),
	.A(n15838),
	.B(n14197));
   NAND2xp33_ASAP7_75t_R U17650 (.Y(n14201),
	.A(n14196),
	.B(n14198));
   NOR2xp33_ASAP7_75t_SRAM U17651 (.Y(n14196),
	.A(n14210),
	.B(n14197));
   NOR2xp33_ASAP7_75t_SRAM U17652 (.Y(n13806),
	.A(FE_OFN26131_n15376),
	.B(n14611));
   NOR2xp33_ASAP7_75t_SRAM U17653 (.Y(n13808),
	.A(n16004),
	.B(n14611));
   NOR2x1_ASAP7_75t_SL U17654 (.Y(n15992),
	.A(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(FE_OFN26635_w3_14));
   NAND2xp33_ASAP7_75t_R U17655 (.Y(n15407),
	.A(FE_OFN26635_w3_14),
	.B(FE_OCPN29520_n24755));
   NAND2xp33_ASAP7_75t_SRAM U17656 (.Y(n13801),
	.A(n15934),
	.B(FE_OFN16459_n));
   NOR2x1_ASAP7_75t_L U17657 (.Y(n15534),
	.A(FE_OFN26538_w3_19),
	.B(FE_OFN6_w3_22));
   NOR2xp33_ASAP7_75t_R U17658 (.Y(n14093),
	.A(n15434),
	.B(n15939));
   NOR2xp33_ASAP7_75t_R U17659 (.Y(n14095),
	.A(n14928),
	.B(n15939));
   NOR3xp33_ASAP7_75t_L U17660 (.Y(n15682),
	.A(FE_OFN16210_n13876),
	.B(FE_OFN6_w3_22),
	.C(FE_OFN26053_n25415));
   NOR2xp67_ASAP7_75t_L U17661 (.Y(n15281),
	.A(n15536),
	.B(n15738));
   NOR2xp33_ASAP7_75t_R U17662 (.Y(n14751),
	.A(n15528),
	.B(n15315));
   NAND2xp33_ASAP7_75t_L U17663 (.Y(n14759),
	.A(n14758),
	.B(n14757));
   NAND2xp33_ASAP7_75t_SRAM U17664 (.Y(n14757),
	.A(n14756),
	.B(n14755));
   NAND2xp33_ASAP7_75t_L U17665 (.Y(n14758),
	.A(n14754),
	.B(n14755));
   INVxp33_ASAP7_75t_SRAM U17666 (.Y(n14756),
	.A(FE_PSN8334_n15539));
   NAND3xp33_ASAP7_75t_SRAM U17667 (.Y(n14760),
	.A(FE_OFN28628_n15667),
	.B(n15536),
	.C(FE_OFN6_w3_22));
   OAI222xp33_ASAP7_75t_R U17668 (.Y(n13774),
	.A1(n15865),
	.A2(n13770),
	.B1(FE_OFN26073_n),
	.B2(n13770),
	.C1(n15857),
	.C2(n13770));
   NOR2xp33_ASAP7_75t_SRAM U17669 (.Y(n13770),
	.A(n14214),
	.B(FE_OFN28792_n15787));
   OAI22xp33_ASAP7_75t_L U17671 (.Y(n13788),
	.A1(n15841),
	.A2(n13775),
	.B1(n15876),
	.B2(n13775));
   O2A1O1Ixp33_ASAP7_75t_SRAM U17672 (.Y(n13786),
	.A1(n15835),
	.A2(n13785),
	.B(n14442),
	.C(n13784));
   NAND2xp5_ASAP7_75t_R U17673 (.Y(n13787),
	.A(n13782),
	.B(n13781));
   OAI21xp33_ASAP7_75t_SRAM U17674 (.Y(n13791),
	.A1(n13769),
	.A2(FE_OFN26084_n15106),
	.B(n13768));
   NAND2xp33_ASAP7_75t_SRAM U17675 (.Y(n13768),
	.A(FE_OFN25897_w3_4),
	.B(n13767));
   INVxp33_ASAP7_75t_SRAM U17676 (.Y(n13769),
	.A(n15810));
   NOR2x1p5_ASAP7_75t_L U17677 (.Y(n15341),
	.A(FE_OFN26041_w3_17),
	.B(FE_OFN5_w3_22));
   AND3x1_ASAP7_75t_L U17678 (.Y(n13883),
	.A(n13879),
	.B(n14254),
	.C(n13878));
   OAI222xp33_ASAP7_75t_SRAM U17679 (.Y(n13879),
	.A1(n15528),
	.A2(n13871),
	.B1(n15484),
	.B2(n13871),
	.C1(FE_OFN26091_n24663),
	.C2(n13871));
   NOR2xp33_ASAP7_75t_L U17680 (.Y(n13871),
	.A(n15484),
	.B(n13875));
   NOR2xp33_ASAP7_75t_L U17681 (.Y(n13413),
	.A(n13556),
	.B(FE_OFN16225_n15195));
   NOR2xp33_ASAP7_75t_L U17682 (.Y(n14614),
	.A(FE_OCPN28407_FE_OFN16433_w3_11),
	.B(n14143));
   NOR2xp33_ASAP7_75t_SRAM U17683 (.Y(n14617),
	.A(n14615),
	.B(n14614));
   NOR2xp33_ASAP7_75t_L U17684 (.Y(n14607),
	.A(n15972),
	.B(n15455));
   NOR2xp33_ASAP7_75t_L U17685 (.Y(n14611),
	.A(n13804),
	.B(FE_OFN28898_n13805));
   OAI21xp33_ASAP7_75t_SRAM U17686 (.Y(n14633),
	.A1(n15963),
	.A2(n15998),
	.B(n14629));
   INVxp33_ASAP7_75t_SRAM U17687 (.Y(n14651),
	.A(n15953));
   NAND2xp5_ASAP7_75t_SL U17688 (.Y(n14716),
	.A(n14628),
	.B(n14627));
   NAND3xp33_ASAP7_75t_R U17689 (.Y(n14628),
	.A(n15451),
	.B(n16012),
	.C(FE_OFN26642_w3_14));
   NAND2xp33_ASAP7_75t_SL U17690 (.Y(n14627),
	.A(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(n14927));
   NOR2xp33_ASAP7_75t_SL U17691 (.Y(n14940),
	.A(n15992),
	.B(n16010));
   INVxp67_ASAP7_75t_R U17692 (.Y(n14626),
	.A(n14143));
   NAND2xp33_ASAP7_75t_L U17693 (.Y(n15353),
	.A(n15337),
	.B(n15336));
   NAND2xp5_ASAP7_75t_L U17694 (.Y(n15354),
	.A(n15327),
	.B(n15326));
   NAND2xp33_ASAP7_75t_L U17695 (.Y(n15311),
	.A(n15305),
	.B(n15308));
   NOR2xp33_ASAP7_75t_R U17696 (.Y(n15305),
	.A(n12994),
	.B(n15306));
   NAND2xp33_ASAP7_75t_R U17697 (.Y(n15310),
	.A(n15309),
	.B(n15308));
   NOR2xp33_ASAP7_75t_R U17698 (.Y(n15309),
	.A(n15307),
	.B(n15306));
   NAND2xp33_ASAP7_75t_SRAM U17699 (.Y(n15317),
	.A(n15316),
	.B(n15313));
   NOR2xp33_ASAP7_75t_R U17700 (.Y(n15316),
	.A(FE_OCPN27987_FE_OFN4_w3_22),
	.B(n15315));
   NAND2xp33_ASAP7_75t_SRAM U17701 (.Y(n15318),
	.A(n15314),
	.B(n15313));
   NOR2xp33_ASAP7_75t_SRAM U17702 (.Y(n15314),
	.A(n15479),
	.B(n15315));
   NAND2xp5_ASAP7_75t_R U17703 (.Y(n15744),
	.A(FE_OFN5_w3_22),
	.B(FE_OFN26053_n25415));
   NAND2xp5_ASAP7_75t_L U17704 (.Y(n13401),
	.A(n13396),
	.B(n13398));
   NOR2xp33_ASAP7_75t_SL U17705 (.Y(n13396),
	.A(n13691),
	.B(n13397));
   NAND2xp33_ASAP7_75t_SL U17706 (.Y(n13400),
	.A(n13399),
	.B(n13398));
   NOR2xp33_ASAP7_75t_L U17707 (.Y(n13399),
	.A(n15181),
	.B(n13397));
   NAND2xp5_ASAP7_75t_L U17709 (.Y(n13378),
	.A(n13377),
	.B(n13376));
   NAND2xp33_ASAP7_75t_SL U17710 (.Y(n13376),
	.A(n13375),
	.B(n13374));
   NOR2xp33_ASAP7_75t_SRAM U17711 (.Y(n14979),
	.A(FE_OFN25912_n15848),
	.B(n14980));
   NOR2xp33_ASAP7_75t_SRAM U17712 (.Y(n14982),
	.A(n15856),
	.B(n14980));
   NAND2xp33_ASAP7_75t_SRAM U17713 (.Y(n14989),
	.A(FE_OFN27156_n),
	.B(n13766));
   NOR2xp33_ASAP7_75t_SRAM U17714 (.Y(n14988),
	.A(n14985),
	.B(n15813));
   OR3x1_ASAP7_75t_SRAM U17715 (.Y(n14990),
	.A(n13726),
	.B(FE_OFN28661_w3_7),
	.C(n15788));
   NOR2xp33_ASAP7_75t_SRAM U17716 (.Y(n15389),
	.A(n13805),
	.B(n15955));
   OAI21x1_ASAP7_75t_SL U17717 (.Y(n15375),
	.A1(FE_OFN26642_w3_14),
	.A2(n16012),
	.B(FE_OFN27135_n15992));
   NAND2xp5_ASAP7_75t_L U17719 (.Y(n15441),
	.A(n15440),
	.B(n15439));
   A2O1A1Ixp33_ASAP7_75t_SL U17720 (.Y(n15459),
	.A1(n15458),
	.A2(n15457),
	.B(n15969),
	.C(n15456));
   NOR2xp33_ASAP7_75t_SRAM U17721 (.Y(n15458),
	.A(n15449),
	.B(n15448));
   NOR2x1_ASAP7_75t_R U17722 (.Y(n15460),
	.A(n13957),
	.B(n15958));
   NAND2xp33_ASAP7_75t_L U17723 (.Y(n15406),
	.A(n15400),
	.B(n15403));
   NAND2xp33_ASAP7_75t_L U17724 (.Y(n15405),
	.A(n15404),
	.B(n15403));
   NAND2xp33_ASAP7_75t_R U17725 (.Y(n15420),
	.A(n15419),
	.B(n15418));
   NOR2xp33_ASAP7_75t_SRAM U17726 (.Y(n15419),
	.A(n16012),
	.B(n15417));
   NAND2xp33_ASAP7_75t_R U17727 (.Y(n15421),
	.A(n15416),
	.B(n15418));
   NOR2xp33_ASAP7_75t_SRAM U17728 (.Y(n15416),
	.A(n15412),
	.B(n15417));
   NAND2xp33_ASAP7_75t_SRAM U17729 (.Y(n15412),
	.A(n15410),
	.B(FE_OFN28658_n15934));
   NAND2xp33_ASAP7_75t_SRAM U17730 (.Y(n15410),
	.A(n15408),
	.B(FE_OFN28715_w3_15));
   NAND3xp33_ASAP7_75t_L U17731 (.Y(n14361),
	.A(FE_OFN26053_n25415),
	.B(FE_OFN27082_n25377),
	.C(FE_OFN6_w3_22));
   NAND2xp33_ASAP7_75t_L U17732 (.Y(n14253),
	.A(n14252),
	.B(n14251));
   NOR2xp33_ASAP7_75t_R U17734 (.Y(n14252),
	.A(FE_OFN28827_n15683),
	.B(n14250));
   NAND2xp5_ASAP7_75t_L U17735 (.Y(n14260),
	.A(n14259),
	.B(n14258));
   NAND2xp33_ASAP7_75t_SL U17736 (.Y(n14258),
	.A(n14257),
	.B(n14256));
   NAND2xp33_ASAP7_75t_L U17737 (.Y(n14259),
	.A(n14255),
	.B(n14256));
   OA21x2_ASAP7_75t_SRAM U17738 (.Y(n14256),
	.A1(n15760),
	.A2(n13875),
	.B(n14254));
   NAND3xp33_ASAP7_75t_SL U17739 (.Y(n13421),
	.A(FE_OFN27210_w3_30),
	.B(FE_OCPN27655_w3_25),
	.C(FE_OFN26049_w3_27));
   NOR3xp33_ASAP7_75t_SL U17740 (.Y(n13659),
	.A(FE_OFN27130_w3_28),
	.B(FE_OFN28663_n),
	.C(FE_OCPN28096_w3_31));
   A2O1A1Ixp33_ASAP7_75t_SL U17741 (.Y(n15623),
	.A1(n15622),
	.A2(n15621),
	.B(n15881),
	.C(n15620));
   NAND2xp5_ASAP7_75t_L U17742 (.Y(n15621),
	.A(n15614),
	.B(n15613));
   NAND2xp5_ASAP7_75t_L U17743 (.Y(n15622),
	.A(n15605),
	.B(n15604));
   NAND2xp33_ASAP7_75t_SRAM U17744 (.Y(n15566),
	.A(n15835),
	.B(n15814));
   NOR2xp33_ASAP7_75t_SL U17745 (.Y(n15571),
	.A(FE_OFN28695_n),
	.B(n13729));
   OAI22xp33_ASAP7_75t_SRAM U17746 (.Y(n15570),
	.A1(n15569),
	.A2(FE_OFN25912_n15848),
	.B1(n13771),
	.B2(FE_OFN25912_n15848));
   NAND2xp5_ASAP7_75t_L U17747 (.Y(n15578),
	.A(FE_OCPN28072_w3_3),
	.B(n14442));
   NOR2xp33_ASAP7_75t_SRAM U17748 (.Y(n15576),
	.A(n15859),
	.B(n15577));
   NAND2xp5_ASAP7_75t_R U17749 (.Y(n14901),
	.A(n15948),
	.B(n15959));
   NAND2xp33_ASAP7_75t_L U17750 (.Y(n15476),
	.A(n15475),
	.B(n15474));
   NAND2xp33_ASAP7_75t_SRAM U17751 (.Y(n15475),
	.A(n15472),
	.B(n15473));
   NAND2xp33_ASAP7_75t_R U17752 (.Y(n15474),
	.A(n14354),
	.B(n15473));
   OAI22xp33_ASAP7_75t_SRAM U17753 (.Y(n15486),
	.A1(n15485),
	.A2(n15683),
	.B1(n15484),
	.B2(n15683));
   NOR2x1_ASAP7_75t_R U17754 (.Y(n15188),
	.A(FE_OFN27210_w3_30),
	.B(FE_OFN25893_n15214));
   NAND3xp33_ASAP7_75t_L U17755 (.Y(n14503),
	.A(n14593),
	.B(FE_OFN26111_n13288),
	.C(FE_OCPN8232_FE_OFN27206_w3_30));
   NOR2xp33_ASAP7_75t_L U17756 (.Y(n15167),
	.A(FE_OFN28452_w3_29),
	.B(FE_OFN27130_w3_28));
   NOR2xp33_ASAP7_75t_SRAM U17758 (.Y(n14731),
	.A(n15455),
	.B(FE_OFN16348_n15949));
   NAND2xp5_ASAP7_75t_L U17761 (.Y(n14734),
	.A(n14706),
	.B(n14705));
   NAND2xp33_ASAP7_75t_L U17762 (.Y(n14705),
	.A(n14704),
	.B(n14703));
   NAND2xp5_ASAP7_75t_L U17763 (.Y(n14706),
	.A(n14701),
	.B(n14703));
   NAND2xp33_ASAP7_75t_L U17764 (.Y(n14733),
	.A(n14711),
	.B(n14710));
   NAND2xp33_ASAP7_75t_SL U17765 (.Y(n14711),
	.A(n14708),
	.B(n14709));
   NAND2xp33_ASAP7_75t_R U17766 (.Y(n14710),
	.A(FE_OFN28848_n14912),
	.B(n14709));
   NOR2xp33_ASAP7_75t_SRAM U17767 (.Y(n14708),
	.A(n15934),
	.B(n14707));
   NAND2xp33_ASAP7_75t_L U17768 (.Y(n14691),
	.A(n14690),
	.B(n14689));
   NAND2xp33_ASAP7_75t_L U17769 (.Y(n14689),
	.A(n14688),
	.B(n14687));
   NAND2xp33_ASAP7_75t_L U17770 (.Y(n14690),
	.A(n14684),
	.B(n14687));
   NAND2xp33_ASAP7_75t_SRAM U17771 (.Y(n14692),
	.A(FE_OFN26131_n15376),
	.B(n16009));
   OAI21xp33_ASAP7_75t_SL U17772 (.Y(n15450),
	.A1(FE_OFN29063_n25433),
	.A2(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(n16012));
   NAND3xp33_ASAP7_75t_L U17773 (.Y(n15995),
	.A(FE_OFN29063_n25433),
	.B(FE_OCPN29509_FE_OFN16184_w3_9),
	.C(FE_OFN26642_w3_14));
   NAND2xp33_ASAP7_75t_SRAM U17774 (.Y(n14670),
	.A(n14927),
	.B(FE_OFN29063_n25433));
   NAND2xp33_ASAP7_75t_R U17775 (.Y(n14669),
	.A(n14668),
	.B(FE_OFN29063_n25433));
   NOR2xp33_ASAP7_75t_R U17776 (.Y(n14671),
	.A(n15934),
	.B(n14672));
   NOR2xp33_ASAP7_75t_SRAM U17777 (.Y(n14674),
	.A(n15923),
	.B(n14672));
   NAND2xp5_ASAP7_75t_L U17778 (.Y(n15738),
	.A(FE_PSN8298_FE_OFN27151_n),
	.B(n15683));
   NAND2xp5_ASAP7_75t_L U17779 (.Y(n15758),
	.A(n15756),
	.B(n15755));
   OAI22xp33_ASAP7_75t_L U17780 (.Y(n15756),
	.A1(n15746),
	.A2(n15745),
	.B1(n15744),
	.B2(n15745));
   NAND2xp33_ASAP7_75t_SL U17781 (.Y(n15755),
	.A(n15754),
	.B(n15753));
   NAND2xp33_ASAP7_75t_L U17782 (.Y(n15745),
	.A(n15743),
	.B(n15742));
   NAND3xp33_ASAP7_75t_SRAM U17783 (.Y(n15760),
	.A(FE_OFN27151_n),
	.B(FE_OFN28706_n),
	.C(FE_OFN27096_n));
   NOR2xp33_ASAP7_75t_SL U17784 (.Y(n14534),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN26051_w3_27));
   NOR3x1_ASAP7_75t_L U17785 (.Y(n14479),
	.A(FE_OCPN27655_w3_25),
	.B(FE_OFN27206_w3_30),
	.C(n25675));
   NAND2xp5_ASAP7_75t_SL U17787 (.Y(n13668),
	.A(n13667),
	.B(n13666));
   NAND2xp5_ASAP7_75t_R U17788 (.Y(n13666),
	.A(n13665),
	.B(n13664));
   NAND2xp5_ASAP7_75t_L U17789 (.Y(n13667),
	.A(n13663),
	.B(n13664));
   NOR2xp33_ASAP7_75t_L U17790 (.Y(n15246),
	.A(n15200),
	.B(n15238));
   NOR2xp33_ASAP7_75t_L U17791 (.Y(n13702),
	.A(n13700),
	.B(n13699));
   NOR2xp33_ASAP7_75t_SRAM U17792 (.Y(n13700),
	.A(FE_OFN27211_w3_30),
	.B(FE_OFN26112_n13288));
   INVx1_ASAP7_75t_SL U17793 (.Y(n13701),
	.A(n13697));
   A2O1A1Ixp33_ASAP7_75t_SL U17794 (.Y(n13697),
	.A1(n14579),
	.A2(n13696),
	.B(n13695),
	.C(n13694));
   NOR2xp33_ASAP7_75t_SRAM U17796 (.Y(n13642),
	.A(n14557),
	.B(n13636));
   INVxp33_ASAP7_75t_R U17797 (.Y(n13640),
	.A(n13639));
   OAI21xp33_ASAP7_75t_SRAM U17798 (.Y(n13638),
	.A1(n13637),
	.A2(n15171),
	.B(FE_OFN25875_n15227));
   NOR2xp33_ASAP7_75t_L U17799 (.Y(n13649),
	.A(FE_OFN25893_n15214),
	.B(n13643));
   NOR2xp33_ASAP7_75t_R U17800 (.Y(n13709),
	.A(FE_OFN25966_n13646),
	.B(n13649));
   INVxp33_ASAP7_75t_SRAM U17801 (.Y(n23903),
	.A(n23902));
   NOR3xp33_ASAP7_75t_L U17802 (.Y(n26015),
	.A(n26010),
	.B(FE_OCPN7617_n26009),
	.C(n26008));
   NAND2xp33_ASAP7_75t_SRAM U17803 (.Y(n26010),
	.A(FE_OFN28521_n26007),
	.B(FE_OFN25996_n26006));
   NAND2xp5_ASAP7_75t_R U17804 (.Y(n25749),
	.A(n25747),
	.B(n25746));
   NAND2xp33_ASAP7_75t_L U17806 (.Y(n25746),
	.A(n25745),
	.B(n25744));
   NAND3xp33_ASAP7_75t_L U17808 (.Y(n24741),
	.A(n24739),
	.B(n24738),
	.C(n24737));
   NOR3xp33_ASAP7_75t_SL U17810 (.Y(n24738),
	.A(n24735),
	.B(n24734),
	.C(n24733));
   NOR3xp33_ASAP7_75t_R U17811 (.Y(n25853),
	.A(n26008),
	.B(n24180),
	.C(FE_OCPN7617_n26009));
   A2O1A1Ixp33_ASAP7_75t_SL U17812 (.Y(n25982),
	.A1(n27117),
	.A2(n26531),
	.B(n25969),
	.C(n25968));
   A2O1A1Ixp33_ASAP7_75t_SL U17814 (.Y(n25644),
	.A1(n25643),
	.A2(n25642),
	.B(n25641),
	.C(n25640));
   NOR3xp33_ASAP7_75t_SL U17815 (.Y(n26516),
	.A(n25633),
	.B(n25632),
	.C(n25631));
   NOR2xp33_ASAP7_75t_L U17817 (.Y(n27025),
	.A(FE_OFN28972_n27021),
	.B(FE_OFN28512_n27020));
   A2O1A1Ixp33_ASAP7_75t_SL U17818 (.Y(n25855),
	.A1(FE_OFN28521_n26007),
	.A2(n25853),
	.B(n26315),
	.C(n25851));
   NOR2x1_ASAP7_75t_L U17819 (.Y(n26958),
	.A(FE_OFN28548_n27092),
	.B(n25542));
   O2A1O1Ixp33_ASAP7_75t_L U17821 (.Y(n26570),
	.A1(n26569),
	.A2(n26568),
	.B(n26567),
	.C(n26566));
   NAND2xp33_ASAP7_75t_SL U17822 (.Y(n26566),
	.A(n26565),
	.B(n26564));
   NAND2xp5_ASAP7_75t_L U17823 (.Y(n26565),
	.A(n26554),
	.B(n26562));
   NOR3xp33_ASAP7_75t_SL U17824 (.Y(n26709),
	.A(n26552),
	.B(FE_OCPN5109_n26551),
	.C(n26550));
   NAND2xp33_ASAP7_75t_SRAM U17825 (.Y(n26552),
	.A(n26549),
	.B(n19010));
   NOR2xp33_ASAP7_75t_R U17826 (.Y(n24566),
	.A(FE_PSN8304_n24565),
	.B(n24564));
   NAND3xp33_ASAP7_75t_SL U17827 (.Y(n24262),
	.A(n19979),
	.B(FE_OCPN27642_n16758),
	.C(FE_OCPN27289_sa21_5));
   NAND2xp33_ASAP7_75t_L U17828 (.Y(n25397),
	.A(n23212),
	.B(n23211));
   NAND2xp33_ASAP7_75t_R U17829 (.Y(n23211),
	.A(n23210),
	.B(n23209));
   NAND2xp5_ASAP7_75t_L U17830 (.Y(n22772),
	.A(n22770),
	.B(n22769));
   NAND2xp33_ASAP7_75t_SRAM U17831 (.Y(n22769),
	.A(n22768),
	.B(n22767));
   NOR3xp33_ASAP7_75t_R U17832 (.Y(n24031),
	.A(n19041),
	.B(n22640),
	.C(n19040));
   NAND2xp33_ASAP7_75t_R U17833 (.Y(n19040),
	.A(n19039),
	.B(n19054));
   NAND2xp33_ASAP7_75t_SRAM U17834 (.Y(n19039),
	.A(n24780),
	.B(n19038));
   NOR2xp33_ASAP7_75t_SRAM U17835 (.Y(n24032),
	.A(n24791),
	.B(n19034));
   NAND2xp5_ASAP7_75t_SL U17836 (.Y(n23325),
	.A(n23308),
	.B(n23170));
   NOR2xp33_ASAP7_75t_SL U17837 (.Y(n23296),
	.A(n23160),
	.B(n21772));
   NOR2x1_ASAP7_75t_SL U17838 (.Y(n23297),
	.A(FE_OCPN29305_n23302),
	.B(FE_OCPN28037_n22855));
   NAND2xp5_ASAP7_75t_R U17839 (.Y(n23739),
	.A(n18605),
	.B(n18604));
   NAND2xp33_ASAP7_75t_L U17840 (.Y(n18604),
	.A(FE_OFN29112_FE_OCPN27870_n18527),
	.B(FE_OFN29081_n18526));
   NAND2xp5_ASAP7_75t_SL U17841 (.Y(n17703),
	.A(FE_OFN69_sa32_4),
	.B(n17534));
   NAND2xp33_ASAP7_75t_L U17842 (.Y(n19729),
	.A(n17708),
	.B(n17707));
   NAND2x1p5_ASAP7_75t_SL U17843 (.Y(n18336),
	.A(n17560),
	.B(FE_OCPN29524_n25029));
   NAND3xp33_ASAP7_75t_SL U17844 (.Y(n20102),
	.A(n17706),
	.B(n17705),
	.C(n22389));
   NAND2xp33_ASAP7_75t_R U17846 (.Y(n17023),
	.A(n17022),
	.B(FE_OFN25977_n18922));
   NOR2x1_ASAP7_75t_L U17847 (.Y(n19430),
	.A(FE_OCPN28202_n16991),
	.B(FE_OCPN29446_n17115));
   NAND2xp33_ASAP7_75t_L U17848 (.Y(n25231),
	.A(n16994),
	.B(n16993));
   NOR2xp33_ASAP7_75t_SRAM U17849 (.Y(n16994),
	.A(FE_OCPN29510_n16996),
	.B(n19411));
   NAND2xp33_ASAP7_75t_L U17851 (.Y(n19723),
	.A(n17570),
	.B(n17569));
   NOR3xp33_ASAP7_75t_L U17852 (.Y(n24217),
	.A(n20910),
	.B(n20909),
	.C(n20908));
   NOR2xp33_ASAP7_75t_L U17853 (.Y(n17782),
	.A(n22881),
	.B(n22539));
   NOR2xp33_ASAP7_75t_SRAM U17855 (.Y(n19664),
	.A(n19663),
	.B(n23015));
   NAND2xp33_ASAP7_75t_R U17857 (.Y(n19804),
	.A(n19795),
	.B(n19794));
   NOR3x1_ASAP7_75t_SL U17858 (.Y(n19803),
	.A(n24893),
	.B(n23958),
	.C(n24941));
   NAND2xp33_ASAP7_75t_SRAM U17859 (.Y(n19794),
	.A(n19793),
	.B(n19792));
   NOR3xp33_ASAP7_75t_SL U17860 (.Y(n24667),
	.A(n19779),
	.B(n24733),
	.C(n19778));
   NAND3xp33_ASAP7_75t_SRAM U17861 (.Y(n19779),
	.A(n23994),
	.B(n19768),
	.C(n19767));
   OAI22xp33_ASAP7_75t_R U17862 (.Y(n24729),
	.A1(FE_OCPN28040_n19766),
	.A2(n19765),
	.B1(n19787),
	.B2(n19765));
   NAND2xp33_ASAP7_75t_L U17863 (.Y(n20641),
	.A(n20637),
	.B(n20638));
   NOR3x1_ASAP7_75t_L U17864 (.Y(n23802),
	.A(n18600),
	.B(n23691),
	.C(n21246));
   OAI21xp5_ASAP7_75t_SL U17865 (.Y(n18600),
	.A1(n23711),
	.A2(n18599),
	.B(n23766));
   NOR3xp33_ASAP7_75t_L U17866 (.Y(n24206),
	.A(n21543),
	.B(n22187),
	.C(n21542));
   NAND2xp33_ASAP7_75t_SRAM U17867 (.Y(n21542),
	.A(n21541),
	.B(n21540));
   NAND2xp5_ASAP7_75t_SRAM U17869 (.Y(n27040),
	.A(n19591),
	.B(n21152));
   NOR3x1_ASAP7_75t_SL U17870 (.Y(n20556),
	.A(n22223),
	.B(FE_OFN28476_sa12_0),
	.C(n17952));
   OAI21xp33_ASAP7_75t_L U17871 (.Y(n27073),
	.A1(FE_OFN26095_n16293),
	.A2(n18093),
	.B(n16504));
   OAI21x1_ASAP7_75t_SL U17872 (.Y(n19683),
	.A1(n23138),
	.A2(n24734),
	.B(FE_OFN130_sa10_5));
   NOR2xp33_ASAP7_75t_L U17873 (.Y(n16596),
	.A(FE_OFN28916_sa10_4),
	.B(n16594));
   NAND3x1_ASAP7_75t_SL U17874 (.Y(n21064),
	.A(n21304),
	.B(FE_OFN28655_FE_OFN25986_n21012),
	.C(FE_OCPN27393_sa03_0));
   OAI22xp33_ASAP7_75t_R U17875 (.Y(n21039),
	.A1(FE_OFN29122_n),
	.A2(n21038),
	.B1(FE_OFN28614_n21715),
	.B2(n21038));
   NAND3x1_ASAP7_75t_SL U17876 (.Y(n21726),
	.A(FE_OFN21730_sa03_3),
	.B(n21708),
	.C(FE_OCPN27405_sa03_4));
   NOR2xp33_ASAP7_75t_SL U17877 (.Y(n23429),
	.A(n21068),
	.B(n21043));
   NOR3xp33_ASAP7_75t_L U17878 (.Y(n21737),
	.A(n21732),
	.B(n21756),
	.C(n21731));
   NAND2xp67_ASAP7_75t_L U17879 (.Y(n23507),
	.A(n23503),
	.B(n23502));
   NAND2xp33_ASAP7_75t_L U17880 (.Y(n23495),
	.A(n23489),
	.B(n23492));
   NAND2xp33_ASAP7_75t_L U17881 (.Y(n23494),
	.A(n23493),
	.B(n23492));
   NAND2xp33_ASAP7_75t_SRAM U17882 (.Y(n23484),
	.A(n20930),
	.B(n22046));
   NAND2xp33_ASAP7_75t_L U17884 (.Y(n20938),
	.A(FE_OCPN27627_sa23_1),
	.B(n20937));
   NAND2xp33_ASAP7_75t_SRAM U17885 (.Y(n20399),
	.A(n20389),
	.B(n24396));
   NOR2x1_ASAP7_75t_L U17886 (.Y(n25071),
	.A(n26465),
	.B(n26464));
   AND3x1_ASAP7_75t_SL U17887 (.Y(n20319),
	.A(n20316),
	.B(n20315),
	.C(n22363));
   NOR3xp33_ASAP7_75t_L U17888 (.Y(n24014),
	.A(n25359),
	.B(n25353),
	.C(n20297));
   NOR3xp33_ASAP7_75t_L U17889 (.Y(n25354),
	.A(n20288),
	.B(n24881),
	.C(FE_OCPN5079_n20287));
   NOR2xp33_ASAP7_75t_L U17890 (.Y(n16742),
	.A(n16859),
	.B(n16708));
   NAND3xp33_ASAP7_75t_SRAM U17891 (.Y(n16708),
	.A(n24489),
	.B(n16707),
	.C(n18424));
   OAI22xp33_ASAP7_75t_L U17892 (.Y(n16737),
	.A1(n16946),
	.A2(n16929),
	.B1(n16427),
	.B2(n16929));
   NAND2xp33_ASAP7_75t_SRAM U17893 (.Y(n16736),
	.A(n16417),
	.B(n16705));
   NAND3xp33_ASAP7_75t_SL U17894 (.Y(n24133),
	.A(n19070),
	.B(n20466),
	.C(n20434));
   NAND2xp5_ASAP7_75t_L U17895 (.Y(n24134),
	.A(n18455),
	.B(n17636));
   NAND2xp33_ASAP7_75t_L U17896 (.Y(n17636),
	.A(n17635),
	.B(n17634));
   NAND2xp33_ASAP7_75t_R U17897 (.Y(n17634),
	.A(n17633),
	.B(n17632));
   NAND2xp33_ASAP7_75t_R U17898 (.Y(n17635),
	.A(n17631),
	.B(n17632));
   NAND2xp33_ASAP7_75t_L U17899 (.Y(n17626),
	.A(n18352),
	.B(n17623));
   NAND2xp33_ASAP7_75t_SL U17900 (.Y(n17625),
	.A(n17624),
	.B(n17623));
   NOR3xp33_ASAP7_75t_SL U17901 (.Y(n24137),
	.A(n17604),
	.B(n18373),
	.C(n18393));
   NOR3xp33_ASAP7_75t_L U17903 (.Y(n24136),
	.A(n17614),
	.B(n22148),
	.C(n20433));
   NOR3xp33_ASAP7_75t_SRAM U17904 (.Y(n19391),
	.A(n19378),
	.B(n20502),
	.C(n19377));
   OAI21xp5_ASAP7_75t_SL U17905 (.Y(n19389),
	.A1(n19388),
	.A2(n19387),
	.B(n26915));
   NOR3xp33_ASAP7_75t_R U17906 (.Y(n25561),
	.A(n19364),
	.B(n19363),
	.C(n19362));
   NOR2xp33_ASAP7_75t_SRAM U17907 (.Y(n19362),
	.A(FE_OCPN5143_n19361),
	.B(n19360));
   NOR2x1_ASAP7_75t_SL U17908 (.Y(n22403),
	.A(n19698),
	.B(n18337));
   NOR3xp33_ASAP7_75t_SRAM U17909 (.Y(n20109),
	.A(n22384),
	.B(n20107),
	.C(n20106));
   NAND2xp5_ASAP7_75t_SL U17914 (.Y(n18918),
	.A(n25221),
	.B(n18256));
   NAND3xp33_ASAP7_75t_SL U17915 (.Y(n18916),
	.A(n18915),
	.B(n27090),
	.C(n25290));
   NAND2xp33_ASAP7_75t_SRAM U17916 (.Y(n18915),
	.A(FE_OCPN27859_n25868),
	.B(FE_OFN16396_n25869));
   NAND3xp33_ASAP7_75t_SL U17917 (.Y(n23419),
	.A(n21327),
	.B(FE_OFN28589_n21048),
	.C(FE_OFN29124_n));
   NOR3x1_ASAP7_75t_L U17918 (.Y(n19670),
	.A(n16576),
	.B(FE_OFN130_sa10_5),
	.C(n17191));
   NOR2x1_ASAP7_75t_SL U17920 (.Y(n21182),
	.A(n21180),
	.B(n21179));
   NAND3xp33_ASAP7_75t_SL U17921 (.Y(n21179),
	.A(n21467),
	.B(n21178),
	.C(n21177));
   NOR2xp33_ASAP7_75t_SL U17922 (.Y(n21463),
	.A(n21147),
	.B(n24517));
   NAND2xp33_ASAP7_75t_R U17923 (.Y(n18778),
	.A(n18777),
	.B(n19123));
   NAND2xp33_ASAP7_75t_SRAM U17924 (.Y(n18753),
	.A(n24084),
	.B(n19811));
   NAND3xp33_ASAP7_75t_SL U17925 (.Y(n24516),
	.A(FE_OFN28767_n26103),
	.B(n17249),
	.C(n24473));
   NAND2xp5_ASAP7_75t_R U17926 (.Y(n17249),
	.A(FE_OFN16216_n19573),
	.B(FE_OCPN28389_n21479));
   NOR2x1_ASAP7_75t_L U17928 (.Y(n18276),
	.A(FE_OCPN5143_n19361),
	.B(FE_OCPN28204_n20526));
   INVx1_ASAP7_75t_L U17929 (.Y(n17100),
	.A(n19414));
   NOR3xp33_ASAP7_75t_SL U17930 (.Y(n17028),
	.A(n17027),
	.B(n17144),
	.C(n19409));
   NAND3xp33_ASAP7_75t_SL U17931 (.Y(n25870),
	.A(n17061),
	.B(n20492),
	.C(n17152));
   NOR2xp67_ASAP7_75t_L U17932 (.Y(n25306),
	.A(n22901),
	.B(n20201));
   NOR3xp33_ASAP7_75t_SRAM U17934 (.Y(n20216),
	.A(n25276),
	.B(n25277),
	.C(FE_OCPN29387_n25273));
   NAND2xp33_ASAP7_75t_SRAM U17935 (.Y(n25911),
	.A(FE_OCPN27773_n22070),
	.B(n22069));
   NAND2x1p5_ASAP7_75t_L U17936 (.Y(n18254),
	.A(FE_OCPN28212_n16980),
	.B(FE_OFN29234_n16996));
   NAND3xp33_ASAP7_75t_SL U17938 (.Y(n25281),
	.A(n19414),
	.B(n19413),
	.C(n19412));
   NAND2xp33_ASAP7_75t_SRAM U17939 (.Y(n19413),
	.A(n19376),
	.B(FE_OCPN29510_n16996));
   NOR3xp33_ASAP7_75t_SL U17940 (.Y(n20491),
	.A(FE_OCPN5143_n19361),
	.B(FE_OFN28478_sa13_2),
	.C(FE_OCPN29340_n17079));
   NOR2x1_ASAP7_75t_L U17941 (.Y(n19405),
	.A(FE_OCPN5143_n19361),
	.B(n17042));
   NOR2x1p5_ASAP7_75t_L U17942 (.Y(n25990),
	.A(n16992),
	.B(FE_OCPN5143_n19361));
   NAND2x1_ASAP7_75t_SL U17944 (.Y(n24164),
	.A(n17126),
	.B(n17125));
   NAND2xp5_ASAP7_75t_L U17945 (.Y(n17125),
	.A(n17124),
	.B(n17122));
   NAND2xp5_ASAP7_75t_L U17946 (.Y(n17126),
	.A(n17123),
	.B(n17122));
   OAI21xp33_ASAP7_75t_L U17947 (.Y(n19447),
	.A1(FE_OFN27133_n21725),
	.A2(FE_OCPN27675_n17986),
	.B(n18041));
   NAND3xp33_ASAP7_75t_SRAM U17948 (.Y(n24839),
	.A(n21047),
	.B(n21060),
	.C(n19487));
   OAI21xp33_ASAP7_75t_L U17952 (.Y(n21528),
	.A1(n23457),
	.A2(FE_OCPN27675_n17986),
	.B(n21526));
   NOR3xp33_ASAP7_75t_L U17953 (.Y(n21526),
	.A(n21525),
	.B(n21524),
	.C(FE_OCPN27628_n23455));
   NAND2xp5_ASAP7_75t_R U17954 (.Y(n23027),
	.A(FE_OFN28946_n23135),
	.B(n23120));
   NAND3xp33_ASAP7_75t_L U17955 (.Y(n24976),
	.A(n16544),
	.B(n19646),
	.C(n16650));
   NOR3xp33_ASAP7_75t_SL U17957 (.Y(n17655),
	.A(n22642),
	.B(n17616),
	.C(FE_OCPN27764_n22152));
   NAND3xp33_ASAP7_75t_L U17958 (.Y(n25088),
	.A(n18351),
	.B(n19072),
	.C(n19043));
   NOR3xp33_ASAP7_75t_L U17959 (.Y(n18351),
	.A(n18368),
	.B(FE_PSN8283_n22629),
	.C(n22613));
   NAND3x1_ASAP7_75t_SL U17960 (.Y(n24128),
	.A(n19072),
	.B(n18501),
	.C(n17620));
   NOR3xp33_ASAP7_75t_L U17961 (.Y(n17620),
	.A(n20446),
	.B(n21619),
	.C(n22163));
   NAND3xp33_ASAP7_75t_L U17964 (.Y(n26083),
	.A(n21371),
	.B(n21370),
	.C(n22509));
   OAI22xp33_ASAP7_75t_SRAM U17965 (.Y(n21371),
	.A1(FE_OFN28877_FE_OCPN27730_n17464),
	.A2(n21821),
	.B1(FE_OFN29061_n22505),
	.B2(n21821));
   NOR2x1_ASAP7_75t_L U17966 (.Y(n25795),
	.A(n19215),
	.B(n22511));
   NOR2xp33_ASAP7_75t_L U17967 (.Y(n19215),
	.A(n19214),
	.B(FE_OCPN28447_n23392));
   NOR3xp33_ASAP7_75t_L U17968 (.Y(n24349),
	.A(n21402),
	.B(n21401),
	.C(n24711));
   OAI21xp33_ASAP7_75t_SRAM U17970 (.Y(n25794),
	.A1(n17444),
	.A2(FE_OCPN5021_n17446),
	.B(FE_OFN29061_n22505));
   NAND2xp33_ASAP7_75t_R U17971 (.Y(n18462),
	.A(n17602),
	.B(FE_OCPN29399_sa30_3));
   NAND2xp5_ASAP7_75t_L U17972 (.Y(n18460),
	.A(n18453),
	.B(n18452));
   NOR3xp33_ASAP7_75t_SL U17973 (.Y(n24794),
	.A(n21587),
	.B(n18482),
	.C(n21628));
   INVxp33_ASAP7_75t_SRAM U17974 (.Y(n18482),
	.A(n18480));
   NOR3xp33_ASAP7_75t_L U17975 (.Y(n25084),
	.A(n21587),
	.B(n21586),
	.C(n26023));
   NAND2xp5_ASAP7_75t_SL U17976 (.Y(n21596),
	.A(n17602),
	.B(n17606));
   NOR3xp33_ASAP7_75t_L U17977 (.Y(n25120),
	.A(n21629),
	.B(n22148),
	.C(n21628));
   NAND2xp33_ASAP7_75t_L U17978 (.Y(n21624),
	.A(n21623),
	.B(n21622));
   NAND2xp33_ASAP7_75t_R U17979 (.Y(n21623),
	.A(n21618),
	.B(n21620));
   AND3x1_ASAP7_75t_SL U17980 (.Y(n23178),
	.A(n23176),
	.B(n23175),
	.C(n23174));
   NOR3xp33_ASAP7_75t_SL U17981 (.Y(n23203),
	.A(n20734),
	.B(FE_OFN29195_n22850),
	.C(FE_OCPN27933_n23328));
   NAND2xp5_ASAP7_75t_L U17982 (.Y(n20732),
	.A(n20731),
	.B(n20730));
   NAND2xp33_ASAP7_75t_SRAM U17983 (.Y(n20730),
	.A(n20729),
	.B(n20727));
   NAND3xp33_ASAP7_75t_R U17984 (.Y(n26880),
	.A(n20723),
	.B(n22271),
	.C(n18173));
   NAND2xp33_ASAP7_75t_SRAM U17985 (.Y(n18173),
	.A(n18172),
	.B(n18171));
   NAND2xp33_ASAP7_75t_SL U17986 (.Y(n18171),
	.A(n18170),
	.B(n18167));
   NAND2xp33_ASAP7_75t_R U17987 (.Y(n18172),
	.A(n18168),
	.B(n18167));
   NAND2xp5_ASAP7_75t_SL U17988 (.Y(n26874),
	.A(n18185),
	.B(n18184));
   NAND2xp33_ASAP7_75t_L U17989 (.Y(n18184),
	.A(n18183),
	.B(n22812));
   NAND2xp33_ASAP7_75t_L U17990 (.Y(n18185),
	.A(n18182),
	.B(n22812));
   NAND2xp5_ASAP7_75t_R U17992 (.Y(n24702),
	.A(n18161),
	.B(FE_OFN25952_n22312));
   NAND3x2_ASAP7_75t_L U17993 (.Y(n23329),
	.A(n23315),
	.B(n20739),
	.C(FE_OFN28680_n));
   OAI21xp33_ASAP7_75t_SRAM U17995 (.Y(n21805),
	.A1(FE_OFN25952_n22312),
	.A2(n21804),
	.B(n21803));
   NAND2xp5_ASAP7_75t_R U17996 (.Y(n21807),
	.A(n21797),
	.B(n21796));
   NOR3xp33_ASAP7_75t_SL U17997 (.Y(n21792),
	.A(n21791),
	.B(n21790),
	.C(n21789));
   NAND2xp33_ASAP7_75t_SRAM U17999 (.Y(n21791),
	.A(n21787),
	.B(n23327));
   NAND2xp33_ASAP7_75t_SRAM U18001 (.Y(n21781),
	.A(FE_RN_0_0),
	.B(FE_OCPN27721_n23336));
   NAND3xp33_ASAP7_75t_SRAM U18002 (.Y(n25191),
	.A(n23718),
	.B(n21645),
	.C(n21644));
   NOR3x1_ASAP7_75t_L U18004 (.Y(n24619),
	.A(n16439),
	.B(n16472),
	.C(FE_OCPN28141_n));
   NAND2x1_ASAP7_75t_L U18005 (.Y(n24614),
	.A(n16424),
	.B(FE_OFN28998_n16923));
   INVx1_ASAP7_75t_SL U18008 (.Y(n24624),
	.A(n16927));
   NAND2xp33_ASAP7_75t_L U18009 (.Y(n26121),
	.A(n23529),
	.B(n23528));
   NOR2xp33_ASAP7_75t_L U18010 (.Y(n18114),
	.A(n16429),
	.B(FE_OCPN27460_n16913));
   OAI222xp33_ASAP7_75t_SRAM U18011 (.Y(n25587),
	.A1(n25586),
	.A2(n25585),
	.B1(n25584),
	.B2(n25585),
	.C1(n25583),
	.C2(n25585));
   INVxp33_ASAP7_75t_SRAM U18013 (.Y(n25586),
	.A(n25578));
   NAND2xp33_ASAP7_75t_L U18014 (.Y(n25576),
	.A(n24281),
	.B(n24280));
   NOR3xp33_ASAP7_75t_L U18015 (.Y(n26155),
	.A(FE_OCPN28107_n23504),
	.B(FE_OCPN29374_FE_OFN29191_sa23_2),
	.C(n20241));
   NOR2xp33_ASAP7_75t_L U18016 (.Y(n22949),
	.A(n23514),
	.B(n22948));
   NAND3xp33_ASAP7_75t_L U18017 (.Y(n22948),
	.A(n22947),
	.B(n22946),
	.C(n23002));
   OAI21xp33_ASAP7_75t_SRAM U18018 (.Y(n22947),
	.A1(FE_OCPN28381_n26660),
	.A2(FE_OFN28787_n19000),
	.B(FE_OFN16248_n20235));
   NOR3xp33_ASAP7_75t_SL U18019 (.Y(n26553),
	.A(n18972),
	.B(n26149),
	.C(n20251));
   NOR2xp33_ASAP7_75t_L U18020 (.Y(n22018),
	.A(n25095),
	.B(n23499));
   NOR2xp33_ASAP7_75t_SRAM U18022 (.Y(n22049),
	.A(n22048),
	.B(n22047));
   NOR2xp67_ASAP7_75t_L U18023 (.Y(n22050),
	.A(n22045),
	.B(n19307));
   NAND2xp33_ASAP7_75t_L U18024 (.Y(n22047),
	.A(n22046),
	.B(n23476));
   NAND3xp33_ASAP7_75t_R U18025 (.Y(n22053),
	.A(n23475),
	.B(n22044),
	.C(n22043));
   NAND2xp33_ASAP7_75t_L U18028 (.Y(n20247),
	.A(n20246),
	.B(n20245));
   NAND2xp33_ASAP7_75t_L U18029 (.Y(n20245),
	.A(n20244),
	.B(n20243));
   NAND2xp33_ASAP7_75t_SL U18030 (.Y(n20246),
	.A(n20923),
	.B(n20243));
   NAND3xp33_ASAP7_75t_R U18031 (.Y(n17353),
	.A(n22421),
	.B(n17352),
	.C(n22422));
   INVxp67_ASAP7_75t_L U18032 (.Y(n17352),
	.A(n22601));
   NAND2xp5_ASAP7_75t_SL U18033 (.Y(n20374),
	.A(n20373),
	.B(FE_OFN26575_n20369));
   NAND2xp5_ASAP7_75t_L U18034 (.Y(n20375),
	.A(n20370),
	.B(FE_OFN26575_n20369));
   NOR3xp33_ASAP7_75t_SL U18036 (.Y(n22786),
	.A(n17922),
	.B(n25439),
	.C(FE_OFN26023_n20807));
   NAND2xp5_ASAP7_75t_L U18037 (.Y(n17913),
	.A(n17912),
	.B(FE_OFN29036_n20806));
   NAND2xp5_ASAP7_75t_L U18038 (.Y(n17914),
	.A(n17910),
	.B(FE_OFN29036_n20806));
   NOR2xp33_ASAP7_75t_L U18039 (.Y(n17912),
	.A(n24362),
	.B(n20596));
   NAND3xp33_ASAP7_75t_L U18040 (.Y(n25738),
	.A(n20817),
	.B(n23617),
	.C(n23616));
   NAND2x1_ASAP7_75t_L U18041 (.Y(n24592),
	.A(n24364),
	.B(FE_OCPN27729_n24362));
   NAND2xp5_ASAP7_75t_L U18042 (.Y(n24368),
	.A(n20815),
	.B(n20814));
   NOR3xp33_ASAP7_75t_L U18043 (.Y(n20815),
	.A(n20813),
	.B(n22718),
	.C(n23588));
   NAND3xp33_ASAP7_75t_R U18044 (.Y(n23621),
	.A(n23597),
	.B(n23596),
	.C(n23595));
   NAND3x1_ASAP7_75t_SL U18046 (.Y(n24992),
	.A(n19718),
	.B(n19697),
	.C(n18325));
   NAND2xp5_ASAP7_75t_SL U18047 (.Y(n22384),
	.A(n19743),
	.B(n17582));
   NOR2xp33_ASAP7_75t_SL U18048 (.Y(n17582),
	.A(n22369),
	.B(n19728));
   NAND2x1_ASAP7_75t_L U18050 (.Y(n19876),
	.A(n24262),
	.B(n22343));
   NOR3x1_ASAP7_75t_L U18051 (.Y(n23929),
	.A(n17832),
	.B(n17856),
	.C(n17831));
   NAND3xp33_ASAP7_75t_L U18052 (.Y(n17832),
	.A(n17830),
	.B(n17829),
	.C(n17828));
   NAND2xp33_ASAP7_75t_R U18053 (.Y(n17829),
	.A(n17827),
	.B(n17826));
   NAND2xp5_ASAP7_75t_SL U18054 (.Y(n25577),
	.A(n19868),
	.B(n19867));
   NOR2xp33_ASAP7_75t_SL U18055 (.Y(n19868),
	.A(n22708),
	.B(n23657));
   NAND3x1_ASAP7_75t_SL U18056 (.Y(n21956),
	.A(n16319),
	.B(n20832),
	.C(n25314));
   OAI22xp33_ASAP7_75t_SRAM U18057 (.Y(n16319),
	.A1(n18073),
	.A2(n18096),
	.B1(FE_OFN28669_sa31_5),
	.B2(n18096));
   OAI21xp5_ASAP7_75t_L U18058 (.Y(n21952),
	.A1(n21951),
	.A2(n21950),
	.B(n26407));
   NAND3xp33_ASAP7_75t_SL U18059 (.Y(n21950),
	.A(n21949),
	.B(n21948),
	.C(n21947));
   NAND2xp5_ASAP7_75t_L U18060 (.Y(n21991),
	.A(n16357),
	.B(n16356));
   NOR3xp33_ASAP7_75t_L U18062 (.Y(n16352),
	.A(n16347),
	.B(n26298),
	.C(n26297));
   NOR3xp33_ASAP7_75t_SL U18063 (.Y(n26307),
	.A(n16320),
	.B(FE_OCPN27316_n25849),
	.C(n21956));
   NAND2xp33_ASAP7_75t_SRAM U18064 (.Y(n16320),
	.A(n18094),
	.B(n25323));
   NOR3xp33_ASAP7_75t_L U18065 (.Y(n26306),
	.A(n16515),
	.B(n18071),
	.C(n27072));
   NOR3xp33_ASAP7_75t_SL U18067 (.Y(n26301),
	.A(n16302),
	.B(n16498),
	.C(n20858));
   NOR3xp33_ASAP7_75t_SRAM U18068 (.Y(n26300),
	.A(n18088),
	.B(n18096),
	.C(n16387));
   NOR3xp33_ASAP7_75t_SL U18070 (.Y(n24488),
	.A(n24486),
	.B(n24485),
	.C(FE_OFN16218_n18418));
   OAI222xp33_ASAP7_75t_R U18072 (.Y(n25484),
	.A1(n24594),
	.A2(n24593),
	.B1(n24592),
	.B2(n24593),
	.C1(n24591),
	.C2(n24593));
   NAND2xp33_ASAP7_75t_SRAM U18073 (.Y(n24593),
	.A(FE_OFN175_sa12_6),
	.B(FE_OFN166_sa12_7));
   NOR2xp33_ASAP7_75t_SRAM U18074 (.Y(n24594),
	.A(FE_OCPN8235_n24589),
	.B(n24588));
   OAI21xp5_ASAP7_75t_R U18076 (.Y(n26651),
	.A1(n25536),
	.A2(n25505),
	.B(n27183));
   OAI222xp33_ASAP7_75t_SRAM U18077 (.Y(n24584),
	.A1(n24218),
	.A2(n26571),
	.B1(n24217),
	.B2(n26571),
	.C1(n24216),
	.C2(n26571));
   NAND2xp33_ASAP7_75t_L U18078 (.Y(n27069),
	.A(n20051),
	.B(n21936));
   NAND3xp33_ASAP7_75t_L U18079 (.Y(n24339),
	.A(n17409),
	.B(n18406),
	.C(n17408));
   NOR3x1_ASAP7_75t_R U18080 (.Y(n25469),
	.A(n25369),
	.B(n17732),
	.C(FE_OFN25946_sa32_6));
   NAND3xp33_ASAP7_75t_L U18083 (.Y(n25216),
	.A(FE_OFN29144_n17747),
	.B(n25214),
	.C(n25213));
   NAND2xp5_ASAP7_75t_L U18084 (.Y(n26534),
	.A(n25604),
	.B(n25603));
   NAND2xp33_ASAP7_75t_SRAM U18085 (.Y(n25603),
	.A(n25602),
	.B(FE_OFN28499_sa00_6));
   NAND2xp33_ASAP7_75t_SRAM U18086 (.Y(n14193),
	.A(n15028),
	.B(FE_OCPN29500_FE_OFN28662_w3_7));
   NOR3xp33_ASAP7_75t_R U18087 (.Y(n14192),
	.A(n14191),
	.B(n14190),
	.C(n14189));
   OAI21xp33_ASAP7_75t_SRAM U18088 (.Y(n14190),
	.A1(FE_OFN26057_w3_1),
	.A2(n15808),
	.B(n14187));
   NAND2xp33_ASAP7_75t_SL U18089 (.Y(n14406),
	.A(n14346),
	.B(n14345));
   NAND2xp33_ASAP7_75t_L U18090 (.Y(n14346),
	.A(n14341),
	.B(n14343));
   NAND2xp33_ASAP7_75t_L U18091 (.Y(n14345),
	.A(n14344),
	.B(n14343));
   NOR2xp33_ASAP7_75t_SRAM U18092 (.Y(n14341),
	.A(n15534),
	.B(n14342));
   NAND3xp33_ASAP7_75t_R U18093 (.Y(n15270),
	.A(n15178),
	.B(n15177),
	.C(n15176));
   NAND2xp33_ASAP7_75t_L U18094 (.Y(n15806),
	.A(n15796),
	.B(n15795));
   NAND2xp33_ASAP7_75t_R U18095 (.Y(n15796),
	.A(n15790),
	.B(n15793));
   NAND2xp33_ASAP7_75t_R U18096 (.Y(n15795),
	.A(n15794),
	.B(n15793));
   NAND2xp33_ASAP7_75t_SRAM U18098 (.Y(n15807),
	.A(n15786),
	.B(n15785));
   NAND2xp33_ASAP7_75t_SRAM U18099 (.Y(n15786),
	.A(n15781),
	.B(n15783));
   NAND2xp33_ASAP7_75t_SRAM U18100 (.Y(n15785),
	.A(n15784),
	.B(n15783));
   NOR2xp33_ASAP7_75t_SRAM U18101 (.Y(n15781),
	.A(n15835),
	.B(n15778));
   NAND2xp33_ASAP7_75t_R U18102 (.Y(n15805),
	.A(n15804),
	.B(n15803));
   NAND2xp33_ASAP7_75t_SRAM U18103 (.Y(n15804),
	.A(n15800),
	.B(n15801));
   NAND2xp33_ASAP7_75t_R U18105 (.Y(n15889),
	.A(n15833),
	.B(n15832));
   NAND3xp33_ASAP7_75t_L U18106 (.Y(n13798),
	.A(n13740),
	.B(n15116),
	.C(n15586));
   NAND2xp33_ASAP7_75t_L U18107 (.Y(n13740),
	.A(n13738),
	.B(n13737));
   NAND2xp33_ASAP7_75t_R U18108 (.Y(n13738),
	.A(n13735),
	.B(n13734));
   OAI21xp33_ASAP7_75t_SRAM U18109 (.Y(n13939),
	.A1(FE_OFN28544_n13805),
	.A2(n15976),
	.B(n15430));
   NAND2xp33_ASAP7_75t_L U18110 (.Y(n13947),
	.A(n13945),
	.B(n13944));
   NAND2xp33_ASAP7_75t_SRAM U18111 (.Y(n13944),
	.A(n13943),
	.B(n13942));
   NAND2xp33_ASAP7_75t_SRAM U18112 (.Y(n13945),
	.A(n13940),
	.B(n13942));
   NOR2xp33_ASAP7_75t_R U18113 (.Y(n13943),
	.A(n15929),
	.B(n13941));
   OAI22xp33_ASAP7_75t_SRAM U18114 (.Y(n13946),
	.A1(n15374),
	.A2(n15449),
	.B1(FE_OFN26131_n15376),
	.B2(n15449));
   NAND2xp5_ASAP7_75t_L U18115 (.Y(n13996),
	.A(n13965),
	.B(n13964));
   NAND2xp33_ASAP7_75t_L U18116 (.Y(n13997),
	.A(n13956),
	.B(n13955));
   NAND2xp33_ASAP7_75t_L U18117 (.Y(n13627),
	.A(n13580),
	.B(n13579));
   NAND2xp33_ASAP7_75t_L U18118 (.Y(n13628),
	.A(n13573),
	.B(n13572));
   NAND3xp33_ASAP7_75t_R U18119 (.Y(n13633),
	.A(n13565),
	.B(n13564),
	.C(n13563));
   OAI222xp33_ASAP7_75t_SRAM U18120 (.Y(n13565),
	.A1(n14593),
	.A2(n13555),
	.B1(n15185),
	.B2(n13555),
	.C1(n13554),
	.C2(n13555));
   NAND2xp33_ASAP7_75t_SRAM U18121 (.Y(n13564),
	.A(n13562),
	.B(n13561));
   NAND2xp5_ASAP7_75t_L U18123 (.Y(n14878),
	.A(n14863),
	.B(n14875));
   NAND2xp33_ASAP7_75t_L U18124 (.Y(n14884),
	.A(n15802),
	.B(n14883));
   OAI21xp5_ASAP7_75t_R U18125 (.Y(n14894),
	.A1(n13741),
	.A2(n14844),
	.B(n14843));
   NAND2xp33_ASAP7_75t_R U18126 (.Y(n14841),
	.A(n14840),
	.B(n14839));
   NAND2xp33_ASAP7_75t_R U18127 (.Y(n14842),
	.A(n14836),
	.B(n14839));
   INVxp67_ASAP7_75t_SL U18128 (.Y(n14657),
	.A(n14658));
   NAND3xp33_ASAP7_75t_R U18129 (.Y(n13409),
	.A(n13347),
	.B(n13346),
	.C(n13345));
   NAND2xp33_ASAP7_75t_L U18131 (.Y(n13425),
	.A(n13419),
	.B(n13418));
   NAND2xp33_ASAP7_75t_R U18132 (.Y(n13418),
	.A(n13417),
	.B(n13416));
   NAND2xp33_ASAP7_75t_R U18133 (.Y(n13419),
	.A(n13414),
	.B(n13416));
   NOR2xp33_ASAP7_75t_SRAM U18134 (.Y(n13417),
	.A(n13677),
	.B(n13415));
   OAI22xp33_ASAP7_75t_SRAM U18135 (.Y(n13423),
	.A1(n14593),
	.A2(n13422),
	.B1(n13421),
	.B2(n13422));
   NOR2xp33_ASAP7_75t_R U18136 (.Y(n13422),
	.A(n14566),
	.B(n14504));
   INVxp33_ASAP7_75t_SRAM U18137 (.Y(n13420),
	.A(n13696));
   NAND2xp5_ASAP7_75t_R U18138 (.Y(n13474),
	.A(FE_OFN28496_n15201),
	.B(n13426));
   NOR2x1_ASAP7_75t_R U18139 (.Y(n13595),
	.A(w3_24_),
	.B(n24470));
   NAND3xp33_ASAP7_75t_SL U18140 (.Y(n15457),
	.A(FE_OFN27200_n),
	.B(n14901),
	.C(FE_PSN8271_n15924));
   NOR2xp33_ASAP7_75t_R U18141 (.Y(n14902),
	.A(n14900),
	.B(n14899));
   OAI21xp33_ASAP7_75t_SRAM U18142 (.Y(n14900),
	.A1(n15959),
	.A2(FE_OFN26007_n16010),
	.B(n14896));
   OAI21xp33_ASAP7_75t_SRAM U18143 (.Y(n14899),
	.A1(n15973),
	.A2(n16016),
	.B(n14898));
   NOR3xp33_ASAP7_75t_SRAM U18144 (.Y(n14964),
	.A(n14918),
	.B(n14917),
	.C(n14916));
   NOR3xp33_ASAP7_75t_SRAM U18145 (.Y(n14965),
	.A(n14911),
	.B(n14910),
	.C(n14909));
   NOR2x1_ASAP7_75t_L U18146 (.Y(n14971),
	.A(w3_10_),
	.B(w3_8_));
   NOR2xp33_ASAP7_75t_SRAM U18147 (.Y(n13492),
	.A(n15145),
	.B(n13708));
   OAI22xp33_ASAP7_75t_SRAM U18148 (.Y(n13496),
	.A1(FE_OFN16201_n15197),
	.A2(n13495),
	.B1(n15224),
	.B2(n13495));
   NOR3xp33_ASAP7_75t_SRAM U18149 (.Y(n13495),
	.A(FE_OFN16225_n15195),
	.B(FE_OCPN8232_FE_OFN27206_w3_30),
	.C(FE_OFN25895_n13662));
   NOR2xp33_ASAP7_75t_SRAM U18151 (.Y(n15263),
	.A(FE_OFN16412_w3_26),
	.B(FE_OFN16159_w3_24));
   NOR3xp33_ASAP7_75t_SL U18152 (.Y(n13544),
	.A(n13543),
	.B(n13542),
	.C(n13541));
   O2A1O1Ixp33_ASAP7_75t_L U18153 (.Y(n13541),
	.A1(n15200),
	.A2(n13540),
	.B(n13539),
	.C(n15259));
   OAI222xp33_ASAP7_75t_SL U18155 (.Y(n13543),
	.A1(FE_OFN16236_n13655),
	.A2(n14585),
	.B1(n13511),
	.B2(n14585),
	.C1(n13510),
	.C2(n14585));
   NOR3xp33_ASAP7_75t_L U18157 (.Y(n14421),
	.A(n14420),
	.B(n14419),
	.C(n14418));
   NAND2xp33_ASAP7_75t_R U18158 (.Y(n16041),
	.A(n15945),
	.B(n15944));
   A2O1A1Ixp33_ASAP7_75t_SL U18159 (.Y(n25765),
	.A1(n26249),
	.A2(n26248),
	.B(FE_OFN26149_n26245),
	.C(n25764));
   NAND2xp5_ASAP7_75t_L U18162 (.Y(n23935),
	.A(n23933),
	.B(n25041));
   NOR2xp33_ASAP7_75t_SRAM U18164 (.Y(n26606),
	.A(FE_OFN28503_n26596),
	.B(n26595));
   NOR3xp33_ASAP7_75t_SL U18165 (.Y(n23963),
	.A(FE_OCPN5178_n25039),
	.B(FE_OCPN27446_n24847),
	.C(n23964));
   A2O1A1Ixp33_ASAP7_75t_SL U18166 (.Y(n26037),
	.A1(n26034),
	.A2(n26033),
	.B(n26926),
	.C(n26032));
   OAI222xp33_ASAP7_75t_SRAM U18167 (.Y(n26978),
	.A1(FE_OFN28973_n25273),
	.A2(n26976),
	.B1(n26975),
	.B2(n26976),
	.C1(n26974),
	.C2(n26976));
   XNOR2xp5_ASAP7_75t_SL U18168 (.Y(n16211),
	.A(w2_9_),
	.B(n16199));
   NAND3xp33_ASAP7_75t_L U18169 (.Y(n24430),
	.A(n24431),
	.B(n24433),
	.C(n24432));
   NOR2xp33_ASAP7_75t_L U18170 (.Y(n25662),
	.A(FE_OFN16214_ld_r),
	.B(FE_OCPN27476_n26852));
   NAND2xp5_ASAP7_75t_SL U18171 (.Y(n24829),
	.A(n24826),
	.B(n24825));
   NAND3xp33_ASAP7_75t_SL U18172 (.Y(n24022),
	.A(n24023),
	.B(FE_OCPN29539_n24927),
	.C(n24024));
   A2O1A1Ixp33_ASAP7_75t_SL U18173 (.Y(n25679),
	.A1(FE_OCPN29586_n26857),
	.A2(n25044),
	.B(n25043),
	.C(n25042));
   A2O1A1Ixp33_ASAP7_75t_L U18174 (.Y(n25042),
	.A1(FE_OCPN29586_n26857),
	.A2(n25044),
	.B(FE_OFN29015_n25040),
	.C(n25144));
   NAND2xp5_ASAP7_75t_SL U18175 (.Y(n25043),
	.A(n25041),
	.B(n25145));
   O2A1O1Ixp33_ASAP7_75t_SL U18176 (.Y(n25893),
	.A1(FE_OFN16158_n26959),
	.A2(n25892),
	.B(n25891),
	.C(n25890));
   NOR2xp33_ASAP7_75t_SRAM U18177 (.Y(n25891),
	.A(w2_28_),
	.B(n25888));
   OAI22xp33_ASAP7_75t_SRAM U18178 (.Y(n25894),
	.A1(text_in_r_60_),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B1(n25895),
	.B2(FE_OFN16_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U18179 (.Y(n26094),
	.A1(text_in_r_107_),
	.A2(FE_OFN28483_ld_r),
	.B1(n26095),
	.B2(FE_OFN28483_ld_r));
   OAI222xp33_ASAP7_75t_SRAM U18180 (.Y(n24112),
	.A1(n24083),
	.A2(n17463),
	.B1(n24082),
	.B2(n17463),
	.C1(n24081),
	.C2(n17463));
   FAx1_ASAP7_75t_SL U18181 (.SN(n24295),
	.A(FE_OCPN27234_n26837),
	.B(FE_OCPN29381_n26796),
	.CI(n24290));
   NAND2xp5_ASAP7_75t_R U18182 (.Y(n24288),
	.A(FE_OFN16448_n),
	.B(n24286));
   NAND3xp33_ASAP7_75t_L U18183 (.Y(n25708),
	.A(FE_OCPN27419_n26602),
	.B(n25710),
	.C(n25709));
   A2O1A1Ixp33_ASAP7_75t_SRAM U18184 (.Y(n27198),
	.A1(FE_OFN16176_n27207),
	.A2(n27192),
	.B(n27191),
	.C(n27190));
   NAND2xp33_ASAP7_75t_SRAM U18185 (.Y(n27191),
	.A(w2_23_),
	.B(FE_OCPN29448_n27189));
   A2O1A1Ixp33_ASAP7_75t_SL U18186 (.Y(n25003),
	.A1(n26829),
	.A2(n25005),
	.B(n25002),
	.C(n25001));
   NOR2x1_ASAP7_75t_L U18189 (.Y(n26892),
	.A(FE_OFN2_ld_r),
	.B(n25982));
   NAND2xp33_ASAP7_75t_R U18190 (.Y(n25254),
	.A(n25251),
	.B(FE_OCPN27333_n25250));
   OAI22xp33_ASAP7_75t_SRAM U18192 (.Y(n25615),
	.A1(text_in_r_118_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(n25616),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U18193 (.Y(n25620),
	.A1(FE_OCPN5056_n26535),
	.A2(n26534),
	.B(n26383),
	.C(n25609));
   NOR3xp33_ASAP7_75t_L U18194 (.Y(n25609),
	.A(FE_OCPN5056_n26535),
	.B(n26383),
	.C(n26534));
   OAI22xp33_ASAP7_75t_SRAM U18195 (.Y(n26374),
	.A1(text_in_r_124_),
	.A2(FE_OFN28483_ld_r),
	.B1(n26375),
	.B2(FE_OFN28483_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SRAM U18196 (.Y(n25651),
	.A1(n26517),
	.A2(n26516),
	.B(n25646),
	.C(n25645));
   O2A1O1Ixp5_ASAP7_75t_SRAM U18197 (.Y(n25645),
	.A1(n26517),
	.A2(n26516),
	.B(FE_OCPN8261_n26513),
	.C(n25648));
   NOR2xp33_ASAP7_75t_SRAM U18198 (.Y(n25646),
	.A(w2_2_),
	.B(n26511));
   NAND2xp33_ASAP7_75t_SRAM U18199 (.Y(n26801),
	.A(n24571),
	.B(n24570));
   A2O1A1Ixp33_ASAP7_75t_L U18202 (.Y(n25241),
	.A1(n25818),
	.A2(n18101),
	.B(n27075),
	.C(n18100));
   NOR2xp33_ASAP7_75t_SRAM U18203 (.Y(n18101),
	.A(FE_OFN28984_n20851),
	.B(n18077));
   OAI22xp33_ASAP7_75t_SL U18204 (.Y(n18100),
	.A1(n26407),
	.A2(n25819),
	.B1(n25824),
	.B2(n25819));
   A2O1A1Ixp33_ASAP7_75t_SL U18206 (.Y(n25722),
	.A1(n25163),
	.A2(n25162),
	.B(n26607),
	.C(n23243));
   NAND3xp33_ASAP7_75t_R U18208 (.Y(n25725),
	.A(n25397),
	.B(n23213),
	.C(n25395));
   NOR2xp33_ASAP7_75t_SRAM U18209 (.Y(n23213),
	.A(n25160),
	.B(FE_OCPN8229_n25750));
   NOR3xp33_ASAP7_75t_SL U18210 (.Y(n19083),
	.A(n19059),
	.B(n24781),
	.C(n19057));
   NAND2xp33_ASAP7_75t_SRAM U18211 (.Y(n19057),
	.A(n19056),
	.B(n24787));
   NAND3xp33_ASAP7_75t_SRAM U18212 (.Y(n26684),
	.A(n24032),
	.B(n24031),
	.C(n24030));
   NOR3xp33_ASAP7_75t_L U18213 (.Y(n22653),
	.A(n22630),
	.B(n22629),
	.C(n22628));
   NAND3xp33_ASAP7_75t_SRAM U18214 (.Y(n22630),
	.A(n22627),
	.B(n22626),
	.C(n22625));
   NOR2xp33_ASAP7_75t_L U18216 (.Y(n22620),
	.A(n22619),
	.B(n22618));
   NOR2xp67_ASAP7_75t_SL U18217 (.Y(n16487),
	.A(n16453),
	.B(n16452));
   OAI21xp33_ASAP7_75t_SRAM U18218 (.Y(n16453),
	.A1(FE_OFN29208_n16436),
	.A2(n16673),
	.B(n16841));
   NAND3xp33_ASAP7_75t_SRAM U18219 (.Y(n26536),
	.A(n24483),
	.B(n16443),
	.C(n24484));
   OAI21xp5_ASAP7_75t_SL U18221 (.Y(n25470),
	.A1(n17736),
	.A2(n26346),
	.B(n17735));
   NOR3xp33_ASAP7_75t_L U18222 (.Y(n17736),
	.A(n17727),
	.B(n17726),
	.C(n17725));
   O2A1O1Ixp33_ASAP7_75t_SL U18223 (.Y(n17735),
	.A1(FE_OCPN28392_n22380),
	.A2(n17734),
	.B(n25367),
	.C(n17733));
   NAND3xp33_ASAP7_75t_L U18225 (.Y(n25366),
	.A(n19709),
	.B(n24853),
	.C(n24854));
   NOR3xp33_ASAP7_75t_L U18226 (.Y(n20949),
	.A(n20918),
	.B(n22999),
	.C(n20917));
   NAND2xp33_ASAP7_75t_SRAM U18227 (.Y(n20917),
	.A(n23476),
	.B(n20919));
   NAND3xp33_ASAP7_75t_R U18228 (.Y(n24037),
	.A(n24216),
	.B(n24217),
	.C(n24218));
   NOR2xp33_ASAP7_75t_L U18229 (.Y(n24038),
	.A(sa23_7_),
	.B(n26562));
   OAI21xp33_ASAP7_75t_SRAM U18230 (.Y(n19355),
	.A1(n24419),
	.A2(n26710),
	.B(n19353));
   INVxp33_ASAP7_75t_SRAM U18231 (.Y(n19353),
	.A(n24042));
   NAND2xp33_ASAP7_75t_SRAM U18232 (.Y(n19358),
	.A(n24040),
	.B(n19300));
   NOR3xp33_ASAP7_75t_SRAM U18233 (.Y(n20183),
	.A(n20135),
	.B(n25523),
	.C(n20957));
   NAND2xp5_ASAP7_75t_L U18234 (.Y(n20182),
	.A(n20148),
	.B(n20147));
   NAND3x1_ASAP7_75t_SL U18235 (.Y(n26494),
	.A(n20134),
	.B(n20133),
	.C(n20202));
   NOR3xp33_ASAP7_75t_SRAM U18236 (.Y(n20134),
	.A(n25210),
	.B(n20161),
	.C(n20996));
   NOR3xp33_ASAP7_75t_R U18237 (.Y(n20133),
	.A(n20131),
	.B(n20139),
	.C(n25201));
   NAND2xp5_ASAP7_75t_SL U18239 (.Y(n22326),
	.A(n22303),
	.B(n22302));
   NAND2xp33_ASAP7_75t_SL U18240 (.Y(n26367),
	.A(n22276),
	.B(n22275));
   NOR3xp33_ASAP7_75t_L U18241 (.Y(n22275),
	.A(n22274),
	.B(n22286),
	.C(n22273));
   NAND3xp33_ASAP7_75t_L U18242 (.Y(n24678),
	.A(n19764),
	.B(n19763),
	.C(n19762));
   NAND2xp33_ASAP7_75t_L U18243 (.Y(n19762),
	.A(n19761),
	.B(n19760));
   A2O1A1Ixp33_ASAP7_75t_SL U18244 (.Y(n24899),
	.A1(n24729),
	.A2(n24667),
	.B(n25139),
	.C(n19807));
   NAND2xp33_ASAP7_75t_L U18246 (.Y(n20699),
	.A(n20652),
	.B(n20651));
   NAND2xp5_ASAP7_75t_R U18247 (.Y(n20652),
	.A(n20648),
	.B(n20649));
   NAND3x1_ASAP7_75t_SL U18248 (.Y(n26196),
	.A(FE_OFN28649_n23802),
	.B(n20642),
	.C(n23887));
   NOR3xp33_ASAP7_75t_SL U18249 (.Y(n20642),
	.A(n20635),
	.B(n23831),
	.C(n21232));
   NAND3xp33_ASAP7_75t_L U18250 (.Y(n20635),
	.A(n20634),
	.B(n20633),
	.C(n23717));
   NAND2xp5_ASAP7_75t_R U18251 (.Y(n20634),
	.A(n20616),
	.B(n20615));
   NOR3xp33_ASAP7_75t_SRAM U18252 (.Y(n22218),
	.A(n22193),
	.B(n22192),
	.C(n22216));
   NOR3xp33_ASAP7_75t_L U18253 (.Y(n22219),
	.A(n22188),
	.B(n22187),
	.C(n22186));
   A2O1A1Ixp33_ASAP7_75t_SL U18254 (.Y(n26675),
	.A1(n25065),
	.A2(n21578),
	.B(n26464),
	.C(n21577));
   NOR3xp33_ASAP7_75t_SRAM U18255 (.Y(n21578),
	.A(n21550),
	.B(FE_OCPN28365_n21549),
	.C(n21548));
   O2A1O1Ixp5_ASAP7_75t_SL U18256 (.Y(n21577),
	.A1(n21576),
	.A2(n21575),
	.B(n26282),
	.C(n21574));
   NOR3xp33_ASAP7_75t_L U18259 (.Y(n19620),
	.A(n19597),
	.B(n27039),
	.C(n19596));
   NOR3xp33_ASAP7_75t_SRAM U18260 (.Y(n19589),
	.A(n19588),
	.B(n21147),
	.C(n17297));
   NOR3x1_ASAP7_75t_L U18261 (.Y(n19590),
	.A(n19587),
	.B(FE_OCPN28418_n19586),
	.C(n19585));
   NAND3x1_ASAP7_75t_L U18263 (.Y(n25255),
	.A(n27037),
	.B(n18626),
	.C(FE_OFN16306_n27041));
   NOR2xp33_ASAP7_75t_L U18264 (.Y(n18626),
	.A(n27040),
	.B(n27039));
   NAND2xp33_ASAP7_75t_SRAM U18265 (.Y(n23851),
	.A(n25637),
	.B(n23796));
   A2O1A1Ixp33_ASAP7_75t_SRAM U18268 (.Y(n20609),
	.A1(n20607),
	.A2(n20606),
	.B(n24377),
	.C(n20605));
   NAND2xp33_ASAP7_75t_SRAM U18269 (.Y(n20606),
	.A(n20570),
	.B(n20569));
   NOR3xp33_ASAP7_75t_R U18270 (.Y(n25337),
	.A(n27069),
	.B(n27070),
	.C(n27073));
   NAND2xp5_ASAP7_75t_R U18273 (.Y(n16627),
	.A(n16615),
	.B(n16614));
   NAND2xp33_ASAP7_75t_R U18274 (.Y(n16614),
	.A(n16613),
	.B(n16612));
   NAND3x1_ASAP7_75t_L U18279 (.Y(n26725),
	.A(FE_OFN28572_n21723),
	.B(n21722),
	.C(n21721));
   NOR3xp33_ASAP7_75t_L U18280 (.Y(n21722),
	.A(n21720),
	.B(n23448),
	.C(n23459));
   NAND2xp5_ASAP7_75t_SL U18282 (.Y(n20385),
	.A(n20384),
	.B(n20383));
   NAND2xp5_ASAP7_75t_L U18283 (.Y(n20383),
	.A(n20382),
	.B(n20381));
   NAND2xp5_ASAP7_75t_L U18284 (.Y(n20384),
	.A(n20379),
	.B(n20381));
   A2O1A1Ixp33_ASAP7_75t_SL U18285 (.Y(n25507),
	.A1(n20089),
	.A2(n20088),
	.B(n27168),
	.C(n20087));
   NAND2xp33_ASAP7_75t_L U18286 (.Y(n20088),
	.A(n20063),
	.B(n20062));
   NOR3xp33_ASAP7_75t_SRAM U18287 (.Y(n20089),
	.A(n20049),
	.B(n20048),
	.C(n20047));
   NAND2xp5_ASAP7_75t_L U18288 (.Y(n25510),
	.A(n26404),
	.B(n20046));
   NOR2xp33_ASAP7_75t_L U18289 (.Y(n20046),
	.A(n26409),
	.B(n20045));
   NAND2xp33_ASAP7_75t_SRAM U18290 (.Y(n20358),
	.A(n25354),
	.B(n24014));
   OAI21xp33_ASAP7_75t_SRAM U18294 (.Y(n19394),
	.A1(FE_OCPN5198_n25566),
	.A2(n27102),
	.B(n19392));
   NOR3xp33_ASAP7_75t_SRAM U18296 (.Y(n17180),
	.A(FE_OCPN5139_n24167),
	.B(n26235),
	.C(n17179));
   NAND2x1_ASAP7_75t_SL U18297 (.Y(n24930),
	.A(FE_OFN28533_n24995),
	.B(n24010));
   NOR2xp67_ASAP7_75t_L U18298 (.Y(n25880),
	.A(n18919),
	.B(n18918));
   NOR3xp33_ASAP7_75t_R U18299 (.Y(n17821),
	.A(n17777),
	.B(n22095),
	.C(n25212));
   INVxp33_ASAP7_75t_SRAM U18300 (.Y(n27211),
	.A(n27212));
   NAND3xp33_ASAP7_75t_SRAM U18301 (.Y(n27215),
	.A(n17767),
	.B(n17766),
	.C(n25526));
   NOR3xp33_ASAP7_75t_L U18302 (.Y(n25419),
	.A(n18865),
	.B(n23441),
	.C(n18864));
   NOR3xp33_ASAP7_75t_SRAM U18303 (.Y(n18911),
	.A(n18877),
	.B(n24244),
	.C(n21038));
   OAI21xp5_ASAP7_75t_SL U18304 (.Y(n23913),
	.A1(n23946),
	.A2(n23945),
	.B(n18058));
   NAND2xp33_ASAP7_75t_L U18306 (.Y(n23916),
	.A(n21077),
	.B(n18002));
   NAND3xp33_ASAP7_75t_L U18308 (.Y(n24178),
	.A(n25503),
	.B(n22875),
	.C(n25502));
   NOR2xp33_ASAP7_75t_SRAM U18309 (.Y(n22875),
	.A(n25536),
	.B(FE_OFN16356_n22874));
   NAND2xp5_ASAP7_75t_L U18310 (.Y(n22913),
	.A(n22886),
	.B(n22885));
   NAND2xp33_ASAP7_75t_SL U18311 (.Y(n22885),
	.A(n22884),
	.B(n22883));
   NOR3x1_ASAP7_75t_SL U18312 (.Y(n23994),
	.A(n19670),
	.B(n21893),
	.C(n21888));
   NAND3xp33_ASAP7_75t_SL U18315 (.Y(n26636),
	.A(n24345),
	.B(n21149),
	.C(n25258));
   INVxp33_ASAP7_75t_SRAM U18316 (.Y(n21459),
	.A(n24476));
   NAND2xp33_ASAP7_75t_SRAM U18317 (.Y(n21460),
	.A(n21449),
	.B(n21448));
   NOR3xp33_ASAP7_75t_SRAM U18318 (.Y(n18738),
	.A(n19089),
	.B(n26100),
	.C(FE_PSN8318_n21455));
   NAND2xp5_ASAP7_75t_L U18320 (.Y(n24100),
	.A(n17244),
	.B(n17243));
   NAND2xp5_ASAP7_75t_L U18321 (.Y(n17243),
	.A(n17242),
	.B(n17241));
   NAND2xp5_ASAP7_75t_L U18322 (.Y(n17244),
	.A(n17240),
	.B(n17241));
   INVxp33_ASAP7_75t_SRAM U18323 (.Y(n17310),
	.A(n24103));
   NOR3xp33_ASAP7_75t_SRAM U18324 (.Y(n17109),
	.A(n25557),
	.B(n17108),
	.C(n17107));
   OAI222xp33_ASAP7_75t_SRAM U18325 (.Y(n17107),
	.A1(n25541),
	.A2(n26959),
	.B1(n17106),
	.B2(n26959),
	.C1(n25562),
	.C2(n26959));
   NOR3xp33_ASAP7_75t_SL U18326 (.Y(n25551),
	.A(n17100),
	.B(n18276),
	.C(n18283));
   NAND2xp33_ASAP7_75t_SL U18328 (.Y(n25860),
	.A(n20960),
	.B(n20959));
   NOR3xp33_ASAP7_75t_SRAM U18329 (.Y(n20959),
	.A(n20958),
	.B(n20957),
	.C(n20956));
   NAND2xp33_ASAP7_75t_SRAM U18330 (.Y(n20191),
	.A(n20190),
	.B(n25301));
   NAND2xp33_ASAP7_75t_L U18332 (.Y(n22116),
	.A(n22082),
	.B(n22081));
   NOR3xp33_ASAP7_75t_SL U18333 (.Y(n22117),
	.A(n26969),
	.B(n26967),
	.C(FE_OCPN29387_n25273));
   A2O1A1Ixp33_ASAP7_75t_SL U18334 (.Y(n26911),
	.A1(n18295),
	.A2(n18294),
	.B(n27102),
	.C(n18293));
   NOR3xp33_ASAP7_75t_L U18335 (.Y(n18294),
	.A(n18274),
	.B(n25282),
	.C(n18273));
   NAND3x1_ASAP7_75t_SL U18336 (.Y(n26914),
	.A(n18255),
	.B(n18254),
	.C(n18253));
   NAND2xp33_ASAP7_75t_L U18337 (.Y(n18253),
	.A(n18252),
	.B(n18251));
   NOR3xp33_ASAP7_75t_SL U18338 (.Y(n18255),
	.A(n18246),
	.B(n20495),
	.C(n18245));
   NAND2xp33_ASAP7_75t_SRAM U18339 (.Y(n18251),
	.A(n18250),
	.B(n18249));
   NOR3xp33_ASAP7_75t_SL U18341 (.Y(n20498),
	.A(n20496),
	.B(n20495),
	.C(n20494));
   NAND2xp33_ASAP7_75t_SL U18342 (.Y(n20496),
	.A(n20493),
	.B(n20492));
   NAND2xp33_ASAP7_75t_SRAM U18343 (.Y(n20494),
	.A(n24164),
	.B(n24165));
   INVx1_ASAP7_75t_L U18347 (.Y(n24834),
	.A(n19459));
   NOR3xp33_ASAP7_75t_SL U18348 (.Y(n24835),
	.A(n19448),
	.B(n19447),
	.C(n19446));
   INVxp67_ASAP7_75t_SL U18349 (.Y(n19446),
	.A(n19445));
   A2O1A1Ixp33_ASAP7_75t_SL U18350 (.Y(n25011),
	.A1(n19694),
	.A2(n19693),
	.B(n25139),
	.C(n19692));
   NAND3xp33_ASAP7_75t_L U18354 (.Y(n17231),
	.A(n17230),
	.B(n17229),
	.C(n17228));
   NOR3xp33_ASAP7_75t_SRAM U18355 (.Y(n17230),
	.A(n17218),
	.B(n19758),
	.C(n21904));
   A2O1A1Ixp33_ASAP7_75t_SL U18356 (.Y(n26790),
	.A1(n23989),
	.A2(n21917),
	.B(n24978),
	.C(n21916));
   O2A1O1Ixp5_ASAP7_75t_SL U18357 (.Y(n21916),
	.A1(n23998),
	.A2(n21915),
	.B(n24974),
	.C(n21914));
   NAND3xp33_ASAP7_75t_L U18358 (.Y(n26793),
	.A(n21879),
	.B(n21878),
	.C(n21877));
   NOR3xp33_ASAP7_75t_SRAM U18359 (.Y(n21879),
	.A(FE_OFN28923_n21873),
	.B(n21872),
	.C(n23139));
   NAND3xp33_ASAP7_75t_R U18362 (.Y(n24939),
	.A(n23124),
	.B(n23123),
	.C(n23122));
   NOR2x1_ASAP7_75t_L U18364 (.Y(n24964),
	.A(n16651),
	.B(n16545));
   NAND2xp5_ASAP7_75t_L U18365 (.Y(n24965),
	.A(n16541),
	.B(n16540));
   NAND2xp33_ASAP7_75t_R U18366 (.Y(n16540),
	.A(n16539),
	.B(n16538));
   NAND2xp33_ASAP7_75t_L U18367 (.Y(n16541),
	.A(n16537),
	.B(n16538));
   OAI21xp5_ASAP7_75t_SRAM U18368 (.Y(n16604),
	.A1(n24979),
	.A2(n24978),
	.B(n16602));
   OAI22xp33_ASAP7_75t_R U18369 (.Y(n16602),
	.A1(n26857),
	.A2(n16601),
	.B1(n16600),
	.B2(n16601));
   NAND2xp33_ASAP7_75t_SRAM U18370 (.Y(n16600),
	.A(n24967),
	.B(n24969));
   NOR3xp33_ASAP7_75t_L U18371 (.Y(n19158),
	.A(n19130),
	.B(n19129),
	.C(n19596));
   NAND2xp33_ASAP7_75t_R U18372 (.Y(n19111),
	.A(n19110),
	.B(n19109));
   NAND2xp33_ASAP7_75t_R U18373 (.Y(n19110),
	.A(FE_OFN26172_n19609),
	.B(n19107));
   INVxp33_ASAP7_75t_SRAM U18375 (.Y(n18400),
	.A(FE_OCPN29458_n26442));
   NOR3xp33_ASAP7_75t_SL U18377 (.Y(n22171),
	.A(n26024),
	.B(n26023),
	.C(n26028));
   NAND3x1_ASAP7_75t_SL U18378 (.Y(n26583),
	.A(n22138),
	.B(n22137),
	.C(n22136));
   NOR3xp33_ASAP7_75t_L U18379 (.Y(n22137),
	.A(n22135),
	.B(n22635),
	.C(n22134));
   NAND3xp33_ASAP7_75t_L U18380 (.Y(n22135),
	.A(n22131),
	.B(n22130),
	.C(n22617));
   NAND2xp5_ASAP7_75t_L U18381 (.Y(n22131),
	.A(n22129),
	.B(n22128));
   NOR2xp33_ASAP7_75t_R U18382 (.Y(n20487),
	.A(n26028),
	.B(n20479));
   NOR3xp33_ASAP7_75t_SL U18383 (.Y(n26179),
	.A(n20484),
	.B(n20475),
	.C(n20474));
   OAI222xp33_ASAP7_75t_L U18385 (.Y(n20474),
	.A1(n22654),
	.A2(n24800),
	.B1(n20473),
	.B2(n24800),
	.C1(n20472),
	.C2(n24800));
   NAND3x1_ASAP7_75t_SL U18386 (.Y(n26183),
	.A(n20436),
	.B(n20435),
	.C(n20434));
   NAND2xp33_ASAP7_75t_SL U18387 (.Y(n20436),
	.A(n20426),
	.B(n20425));
   NOR2xp33_ASAP7_75t_SL U18388 (.Y(n20435),
	.A(n22619),
	.B(n20433));
   NAND2xp33_ASAP7_75t_SRAM U18389 (.Y(n20425),
	.A(n20424),
	.B(n20423));
   OAI222xp33_ASAP7_75t_L U18390 (.Y(n17516),
	.A1(FE_OCPN29554_n22507),
	.A2(n17506),
	.B1(n17515),
	.B2(n17506),
	.C1(n17514),
	.C2(n17506));
   NAND3xp33_ASAP7_75t_L U18392 (.Y(n24633),
	.A(n17461),
	.B(n17460),
	.C(n23371));
   NAND3xp33_ASAP7_75t_L U18395 (.Y(n24543),
	.A(n26104),
	.B(n19816),
	.C(n25258));
   NOR3xp33_ASAP7_75t_SL U18396 (.Y(n24556),
	.A(n21832),
	.B(n24079),
	.C(n24078));
   OAI22xp33_ASAP7_75t_SRAM U18397 (.Y(n21868),
	.A1(FE_OFN28877_FE_OCPN27730_n17464),
	.A2(n23267),
	.B1(FE_OFN29061_n22505),
	.B2(n23267));
   NOR3xp33_ASAP7_75t_SRAM U18398 (.Y(n21867),
	.A(n21843),
	.B(n23376),
	.C(n21842));
   NOR3xp33_ASAP7_75t_SRAM U18400 (.Y(n26739),
	.A(n22488),
	.B(n24551),
	.C(n24545));
   NOR2xp33_ASAP7_75t_R U18401 (.Y(n22522),
	.A(FE_OCPN27584_n22497),
	.B(n22496));
   NOR3xp33_ASAP7_75t_SL U18402 (.Y(n22521),
	.A(n17485),
	.B(n22498),
	.C(n24078));
   NOR3xp33_ASAP7_75t_SRAM U18403 (.Y(n21435),
	.A(n21403),
	.B(n17477),
	.C(n23274));
   NAND2xp33_ASAP7_75t_L U18404 (.Y(n21434),
	.A(n21409),
	.B(n21408));
   NAND3xp33_ASAP7_75t_L U18406 (.Y(n26372),
	.A(n25794),
	.B(n24349),
	.C(n25795));
   NAND3xp33_ASAP7_75t_SL U18407 (.Y(n23408),
	.A(n23387),
	.B(n23370),
	.C(n23369));
   NAND3xp33_ASAP7_75t_SL U18408 (.Y(n23407),
	.A(n26064),
	.B(n23372),
	.C(n23371));
   NAND2xp5_ASAP7_75t_L U18409 (.Y(n23367),
	.A(n23365),
	.B(n23364));
   NAND2xp33_ASAP7_75t_L U18410 (.Y(n23364),
	.A(n23363),
	.B(n23362));
   NOR2xp67_ASAP7_75t_L U18411 (.Y(n26082),
	.A(sa11_6_),
	.B(sa11_7_));
   NOR2xp33_ASAP7_75t_L U18412 (.Y(n25081),
	.A(FE_OFN28480_sa30_7),
	.B(n17629));
   NOR2xp33_ASAP7_75t_R U18413 (.Y(n21615),
	.A(n21602),
	.B(n21601));
   OAI222xp33_ASAP7_75t_R U18414 (.Y(n21630),
	.A1(n24579),
	.A2(n26687),
	.B1(n21588),
	.B2(n26687),
	.C1(n25084),
	.C2(n26687));
   NOR3xp33_ASAP7_75t_SRAM U18415 (.Y(n21588),
	.A(n21585),
	.B(n25082),
	.C(n25087));
   NAND2xp33_ASAP7_75t_SRAM U18416 (.Y(n21585),
	.A(n25086),
	.B(n21584));
   NAND2xp33_ASAP7_75t_SRAM U18417 (.Y(n18562),
	.A(n23716),
	.B(n20633));
   NOR3xp33_ASAP7_75t_SRAM U18419 (.Y(n18541),
	.A(n18567),
	.B(n23740),
	.C(n23691));
   NAND3xp33_ASAP7_75t_L U18420 (.Y(n25979),
	.A(n23173),
	.B(n23172),
	.C(n23171));
   NOR2xp33_ASAP7_75t_L U18421 (.Y(n23173),
	.A(n23331),
	.B(n23167));
   A2O1A1Ixp33_ASAP7_75t_L U18423 (.Y(n27113),
	.A1(n20781),
	.A2(n20780),
	.B(n23345),
	.C(n20779));
   NAND2xp33_ASAP7_75t_SRAM U18424 (.Y(n20781),
	.A(n20719),
	.B(n20718));
   NOR3xp33_ASAP7_75t_SL U18425 (.Y(n20780),
	.A(n20736),
	.B(n22304),
	.C(n20735));
   O2A1O1Ixp5_ASAP7_75t_L U18426 (.Y(n20779),
	.A1(n20778),
	.A2(n20752),
	.B(n26878),
	.C(n20777));
   NAND3xp33_ASAP7_75t_L U18427 (.Y(n27116),
	.A(n20714),
	.B(n20713),
	.C(n23334));
   NOR3xp33_ASAP7_75t_SRAM U18428 (.Y(n20714),
	.A(n20703),
	.B(n24694),
	.C(n22838));
   OAI21xp33_ASAP7_75t_SRAM U18429 (.Y(n20703),
	.A1(n20729),
	.A2(n18186),
	.B(n20702));
   NOR2xp33_ASAP7_75t_L U18430 (.Y(n21143),
	.A(n26875),
	.B(n21097));
   NAND3xp33_ASAP7_75t_SL U18431 (.Y(n21097),
	.A(n21096),
	.B(n21095),
	.C(n21094));
   NAND3xp33_ASAP7_75t_SL U18432 (.Y(n24113),
	.A(n21089),
	.B(n21088),
	.C(n24699));
   NOR2xp33_ASAP7_75t_SRAM U18433 (.Y(n21088),
	.A(n26876),
	.B(n21087));
   NOR2xp33_ASAP7_75t_SL U18434 (.Y(n22867),
	.A(n23331),
	.B(n22835));
   NAND3xp33_ASAP7_75t_L U18435 (.Y(n26482),
	.A(n22806),
	.B(n22805),
	.C(n22868));
   NOR3xp33_ASAP7_75t_L U18436 (.Y(n22805),
	.A(n22804),
	.B(n23185),
	.C(n22803));
   NOR2x1_ASAP7_75t_L U18437 (.Y(n24701),
	.A(n22838),
	.B(n18209));
   NOR2x1_ASAP7_75t_L U18438 (.Y(n24699),
	.A(FE_OFN16304_n22808),
	.B(n18179));
   NAND2xp5_ASAP7_75t_L U18439 (.Y(n18179),
	.A(n22800),
	.B(n21775));
   NOR2xp33_ASAP7_75t_L U18441 (.Y(n26878),
	.A(sa22_6_),
	.B(sa22_7_));
   NOR3xp33_ASAP7_75t_R U18442 (.Y(n21263),
	.A(n21237),
	.B(n23745),
	.C(n21236));
   NOR3xp33_ASAP7_75t_SL U18445 (.Y(n23736),
	.A(n23713),
	.B(FE_OCPN28017_n18548),
	.C(n23712));
   NAND3xp33_ASAP7_75t_SL U18447 (.Y(n27206),
	.A(n23687),
	.B(n23686),
	.C(n23685));
   NAND2xp33_ASAP7_75t_L U18448 (.Y(n23686),
	.A(n23684),
	.B(n23683));
   NAND2xp33_ASAP7_75t_L U18449 (.Y(n23683),
	.A(n23682),
	.B(n23681));
   O2A1O1Ixp5_ASAP7_75t_SL U18452 (.Y(n18448),
	.A1(n24612),
	.A2(n24611),
	.B(n24610),
	.C(n24622));
   NOR3x1_ASAP7_75t_SL U18453 (.Y(n26764),
	.A(n24622),
	.B(n18436),
	.C(n24609));
   NOR3xp33_ASAP7_75t_L U18454 (.Y(n18429),
	.A(n18428),
	.B(n24612),
	.C(n18443));
   NAND3x1_ASAP7_75t_SL U18455 (.Y(n26769),
	.A(FE_OFN25940_n24621),
	.B(n18414),
	.C(n24619));
   NOR3xp33_ASAP7_75t_L U18456 (.Y(n18414),
	.A(n24618),
	.B(n24624),
	.C(n18413));
   NAND2xp33_ASAP7_75t_R U18457 (.Y(n18413),
	.A(n18412),
	.B(n24614));
   NAND2xp33_ASAP7_75t_SRAM U18458 (.Y(n18412),
	.A(n18411),
	.B(n18410));
   NOR2xp33_ASAP7_75t_R U18459 (.Y(n17422),
	.A(n17414),
	.B(n17413));
   NAND2xp5_ASAP7_75t_L U18460 (.Y(n24309),
	.A(n17411),
	.B(n17410));
   NAND2xp33_ASAP7_75t_R U18461 (.Y(n17411),
	.A(n17403),
	.B(n17402));
   NOR3xp33_ASAP7_75t_L U18462 (.Y(n17410),
	.A(n23543),
	.B(n24339),
	.C(n23557));
   NAND2xp33_ASAP7_75t_SRAM U18463 (.Y(n17402),
	.A(n17401),
	.B(FE_OFN28935_n18104));
   A2O1A1Ixp33_ASAP7_75t_L U18466 (.Y(n16969),
	.A1(n16968),
	.A2(n16967),
	.B(n24331),
	.C(n16966));
   NAND3xp33_ASAP7_75t_R U18467 (.Y(n16970),
	.A(n16934),
	.B(n16933),
	.C(n18138));
   OA21x2_ASAP7_75t_SL U18469 (.Y(n18152),
	.A1(n18151),
	.A2(n18150),
	.B(n24610));
   NOR3xp33_ASAP7_75t_R U18471 (.Y(n26359),
	.A(n26121),
	.B(n26122),
	.C(n24612));
   NOR3xp33_ASAP7_75t_SL U18472 (.Y(n26358),
	.A(n24300),
	.B(FE_OCPN7607_n23539),
	.C(n18114));
   NOR3xp33_ASAP7_75t_R U18473 (.Y(n23566),
	.A(n23536),
	.B(n23535),
	.C(n23534));
   NOR3xp33_ASAP7_75t_SL U18474 (.Y(n24336),
	.A(n16848),
	.B(n18145),
	.C(n16867));
   NAND3xp33_ASAP7_75t_SL U18475 (.Y(n16848),
	.A(n16846),
	.B(n16845),
	.C(n16927));
   A2O1A1Ixp33_ASAP7_75t_SRAM U18476 (.Y(n16904),
	.A1(n16902),
	.A2(n16901),
	.B(n24331),
	.C(n16900));
   NOR2xp67_ASAP7_75t_R U18477 (.Y(n24610),
	.A(FE_OFN90_sa33_7),
	.B(FE_OFN174_sa33_6));
   OAI21xp5_ASAP7_75t_SL U18478 (.Y(n25593),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OFN28565_n26845),
	.B(n25594));
   NAND2xp33_ASAP7_75t_R U18479 (.Y(n18978),
	.A(n18977),
	.B(n18976));
   NOR2xp33_ASAP7_75t_L U18481 (.Y(n19026),
	.A(n26551),
	.B(n26550));
   NAND3xp33_ASAP7_75t_SL U18482 (.Y(n25736),
	.A(n22927),
	.B(n26160),
	.C(n26161));
   NOR3xp33_ASAP7_75t_L U18483 (.Y(n22927),
	.A(n22924),
	.B(n22923),
	.C(n22922));
   NAND2xp33_ASAP7_75t_L U18484 (.Y(n22921),
	.A(n22920),
	.B(n22919));
   NOR3xp33_ASAP7_75t_SL U18485 (.Y(n25701),
	.A(n20229),
	.B(FE_OCPN5109_n26551),
	.C(n24769));
   NAND3xp33_ASAP7_75t_L U18487 (.Y(n26996),
	.A(n22016),
	.B(n22015),
	.C(n22982));
   NOR3xp33_ASAP7_75t_SRAM U18488 (.Y(n22016),
	.A(n22003),
	.B(n22992),
	.C(n22002));
   NOR3xp33_ASAP7_75t_SRAM U18489 (.Y(n22015),
	.A(n22014),
	.B(n23514),
	.C(n22013));
   NOR3xp33_ASAP7_75t_SL U18491 (.Y(n22966),
	.A(n22965),
	.B(n26661),
	.C(FE_OCPN27796_n26659));
   NOR3xp33_ASAP7_75t_L U18492 (.Y(n23008),
	.A(n22977),
	.B(n22976),
	.C(n23488));
   NAND3xp33_ASAP7_75t_L U18493 (.Y(n22977),
	.A(n22969),
	.B(n22968),
	.C(n22967));
   NOR2x1_ASAP7_75t_R U18494 (.Y(n26567),
	.A(FE_OFN45_sa23_6),
	.B(FE_OFN162_sa23_7));
   NAND3xp33_ASAP7_75t_L U18495 (.Y(n25173),
	.A(n22595),
	.B(n18676),
	.C(n18675));
   NAND3xp33_ASAP7_75t_L U18496 (.Y(n18729),
	.A(n18718),
	.B(n24396),
	.C(n24395));
   NOR3xp33_ASAP7_75t_L U18497 (.Y(n18718),
	.A(n18715),
	.B(n24392),
	.C(n18722));
   NOR3xp33_ASAP7_75t_L U18501 (.Y(n23072),
	.A(n23071),
	.B(FE_OFN16341_n27008),
	.C(n23069));
   NAND3xp33_ASAP7_75t_SL U18503 (.Y(n23071),
	.A(n24222),
	.B(n23068),
	.C(n25057));
   NOR2xp33_ASAP7_75t_SL U18505 (.Y(n24122),
	.A(n24226),
	.B(n17394));
   A2O1A1Ixp33_ASAP7_75t_L U18506 (.Y(n17394),
	.A1(n24222),
	.A2(n24221),
	.B(n27004),
	.C(n17393));
   OAI21xp33_ASAP7_75t_SL U18507 (.Y(n17393),
	.A1(n24228),
	.A2(n24227),
	.B(n26679));
   NAND2xp5_ASAP7_75t_R U18508 (.Y(n24126),
	.A(n24219),
	.B(n17344));
   A2O1A1Ixp33_ASAP7_75t_SL U18510 (.Y(n25444),
	.A1(n26998),
	.A2(n22610),
	.B(n27004),
	.C(n27014));
   NOR2xp33_ASAP7_75t_SRAM U18511 (.Y(n22610),
	.A(n27001),
	.B(n22587));
   NAND3xp33_ASAP7_75t_L U18512 (.Y(n25694),
	.A(n22581),
	.B(n22580),
	.C(n27017));
   NAND2xp33_ASAP7_75t_L U18513 (.Y(n22581),
	.A(n22578),
	.B(n22577));
   NOR3xp33_ASAP7_75t_SRAM U18514 (.Y(n22580),
	.A(n22579),
	.B(n27012),
	.C(n27011));
   NAND2xp33_ASAP7_75t_SRAM U18515 (.Y(n22577),
	.A(FE_OFN25950_sa01_2),
	.B(n27008));
   OAI22xp5_ASAP7_75t_L U18516 (.Y(n22475),
	.A1(n22474),
	.A2(n27015),
	.B1(n22473),
	.B2(n27015));
   NAND3xp33_ASAP7_75t_SL U18518 (.Y(n26250),
	.A(n22430),
	.B(n22429),
	.C(n22428));
   NAND2xp33_ASAP7_75t_SRAM U18519 (.Y(n22430),
	.A(n22420),
	.B(n22419));
   NAND2xp5_ASAP7_75t_L U18520 (.Y(n22429),
	.A(n22427),
	.B(n22426));
   NAND2xp33_ASAP7_75t_R U18521 (.Y(n22420),
	.A(n22416),
	.B(n22417));
   NOR3xp33_ASAP7_75t_L U18522 (.Y(n19569),
	.A(n19537),
	.B(FE_OCPN8229_n25750),
	.C(n23572));
   NAND3xp33_ASAP7_75t_R U18523 (.Y(n19567),
	.A(n19545),
	.B(n19544),
	.C(n19543));
   NAND3xp33_ASAP7_75t_L U18524 (.Y(n25680),
	.A(n19517),
	.B(n19516),
	.C(n22786));
   NAND2xp33_ASAP7_75t_R U18525 (.Y(n19517),
	.A(n19508),
	.B(n19507));
   NOR3xp33_ASAP7_75t_R U18526 (.Y(n19516),
	.A(n19515),
	.B(n22238),
	.C(n20792));
   NAND2xp33_ASAP7_75t_R U18527 (.Y(n19507),
	.A(n19506),
	.B(n19505));
   NAND3xp33_ASAP7_75t_SL U18528 (.Y(n25178),
	.A(n17909),
	.B(n17908),
	.C(FE_OFN28560_n22749));
   NAND2xp33_ASAP7_75t_SRAM U18529 (.Y(n17908),
	.A(FE_OFN28739_n17898),
	.B(n25741));
   NOR3xp33_ASAP7_75t_SL U18530 (.Y(n17909),
	.A(n25738),
	.B(FE_OCPN8229_n25750),
	.C(n25737));
   NAND3xp33_ASAP7_75t_L U18531 (.Y(n26138),
	.A(n22733),
	.B(n22732),
	.C(n23599));
   NOR3xp33_ASAP7_75t_L U18532 (.Y(n22265),
	.A(n22243),
	.B(n22242),
	.C(n22241));
   INVx1_ASAP7_75t_L U18533 (.Y(n24210),
	.A(n25485));
   O2A1O1Ixp5_ASAP7_75t_SL U18534 (.Y(n20827),
	.A1(n24051),
	.A2(n20826),
	.B(n25682),
	.C(n20825));
   NAND3xp33_ASAP7_75t_SRAM U18535 (.Y(n20831),
	.A(n20788),
	.B(n20787),
	.C(n25442));
   NAND2xp33_ASAP7_75t_SRAM U18538 (.Y(n18346),
	.A(n25026),
	.B(n25025));
   NAND2xp33_ASAP7_75t_SL U18539 (.Y(n18319),
	.A(n18318),
	.B(n18317));
   NOR3xp33_ASAP7_75t_L U18541 (.Y(n25672),
	.A(n22376),
	.B(n22375),
	.C(FE_OFN28928_n22374));
   NAND3xp33_ASAP7_75t_SL U18542 (.Y(n24749),
	.A(n16766),
	.B(n16765),
	.C(n23639));
   NAND2xp33_ASAP7_75t_R U18543 (.Y(n16766),
	.A(n16756),
	.B(n16755));
   NOR3xp33_ASAP7_75t_SRAM U18544 (.Y(n16765),
	.A(n16759),
	.B(n20301),
	.C(n19876));
   NAND2xp33_ASAP7_75t_SRAM U18545 (.Y(n16755),
	.A(n16754),
	.B(n16753));
   NOR3xp33_ASAP7_75t_SL U18546 (.Y(n16827),
	.A(n16788),
	.B(n16787),
	.C(n16786));
   A2O1A1Ixp33_ASAP7_75t_SL U18547 (.Y(n23968),
	.A1(n17894),
	.A2(n17893),
	.B(n25585),
	.C(n17892));
   NAND2xp33_ASAP7_75t_R U18548 (.Y(n17894),
	.A(n17837),
	.B(n17836));
   NOR3xp33_ASAP7_75t_SRAM U18549 (.Y(n17893),
	.A(n17842),
	.B(n22335),
	.C(n20011));
   NOR3xp33_ASAP7_75t_SL U18551 (.Y(n19903),
	.A(n25582),
	.B(n25580),
	.C(n25578));
   NAND3xp33_ASAP7_75t_R U18552 (.Y(n25382),
	.A(n19870),
	.B(n19869),
	.C(n24281));
   NOR3xp33_ASAP7_75t_SRAM U18554 (.Y(n19869),
	.A(n24279),
	.B(n24278),
	.C(n25577));
   NAND2xp5_ASAP7_75t_L U18555 (.Y(n23673),
	.A(n23648),
	.B(n23647));
   O2A1O1Ixp5_ASAP7_75t_SL U18556 (.Y(n23672),
	.A1(n23671),
	.A2(n23670),
	.B(n25575),
	.C(n23669));
   NAND2xp33_ASAP7_75t_L U18557 (.Y(n23647),
	.A(n23646),
	.B(n23645));
   NAND3xp33_ASAP7_75t_L U18558 (.Y(n25959),
	.A(n24921),
	.B(n23637),
	.C(n24920));
   NAND2xp33_ASAP7_75t_SRAM U18559 (.Y(n23637),
	.A(n23636),
	.B(n23635));
   NAND2xp33_ASAP7_75t_R U18560 (.Y(n23635),
	.A(n23634),
	.B(n23630));
   NOR2xp33_ASAP7_75t_R U18561 (.Y(n25152),
	.A(FE_OFN16214_ld_r),
	.B(n26852));
   A2O1A1Ixp33_ASAP7_75t_L U18562 (.Y(n24846),
	.A1(n22405),
	.A2(FE_OCPN27940_n26842),
	.B(n24833),
	.C(n24832));
   NOR3xp33_ASAP7_75t_L U18563 (.Y(n21998),
	.A(n21978),
	.B(n21977),
	.C(FE_OFN26550_n16331));
   NOR3xp33_ASAP7_75t_SRAM U18564 (.Y(n21999),
	.A(n21974),
	.B(FE_OFN16367_n21973),
	.C(n21972));
   NAND3x1_ASAP7_75t_L U18565 (.Y(n26941),
	.A(n21971),
	.B(n21970),
	.C(n26296));
   NAND2xp33_ASAP7_75t_R U18566 (.Y(n21969),
	.A(n21967),
	.B(n21966));
   NAND3xp33_ASAP7_75t_SRAM U18567 (.Y(n21960),
	.A(n25314),
	.B(n21927),
	.C(n25315));
   NOR2xp33_ASAP7_75t_SRAM U18568 (.Y(n20896),
	.A(n26297),
	.B(n20848));
   NOR3xp33_ASAP7_75t_SL U18569 (.Y(n20895),
	.A(n20852),
	.B(FE_OFN28984_n20851),
	.C(FE_PSN8317_n20850));
   NAND3x1_ASAP7_75t_R U18570 (.Y(n26201),
	.A(n20846),
	.B(n20845),
	.C(n26294));
   OAI21xp33_ASAP7_75t_L U18572 (.Y(n20843),
	.A1(FE_OCPN28314_n20842),
	.A2(FE_OCPN7597_n21981),
	.B(n21992));
   NOR3xp33_ASAP7_75t_SRAM U18573 (.Y(n16411),
	.A(FE_OCPN5076_n24192),
	.B(n25856),
	.C(n16410));
   OAI222xp33_ASAP7_75t_SRAM U18574 (.Y(n16410),
	.A1(FE_OFN28521_n26007),
	.A2(n26315),
	.B1(n16409),
	.B2(n26315),
	.C1(FE_OFN25996_n26006),
	.C2(n26315));
   NOR2xp67_ASAP7_75t_L U18575 (.Y(n24191),
	.A(n21982),
	.B(n21991));
   NAND2xp33_ASAP7_75t_SRAM U18576 (.Y(n16371),
	.A(n16370),
	.B(n16369));
   NAND2xp33_ASAP7_75t_SRAM U18577 (.Y(n16369),
	.A(n16368),
	.B(n16367));
   NAND2xp33_ASAP7_75t_SRAM U18578 (.Y(n16370),
	.A(n16366),
	.B(n16367));
   NOR2xp67_ASAP7_75t_L U18579 (.Y(n26407),
	.A(sa31_6_),
	.B(sa31_7_));
   A2O1A1Ixp33_ASAP7_75t_SL U18581 (.Y(n26904),
	.A1(n26307),
	.A2(n26306),
	.B(n27168),
	.C(n16353));
   O2A1O1Ixp33_ASAP7_75t_L U18582 (.Y(n16353),
	.A1(FE_OCPN28156_n26304),
	.A2(n26303),
	.B(n26407),
	.C(n26945));
   NAND3xp33_ASAP7_75t_L U18584 (.Y(n26907),
	.A(n26300),
	.B(n26301),
	.C(n26302));
   NOR3xp33_ASAP7_75t_L U18585 (.Y(n26348),
	.A(FE_OCPN27491_n26351),
	.B(n26349),
	.C(n26350));
   OAI222xp33_ASAP7_75t_SRAM U18586 (.Y(n26350),
	.A1(n26347),
	.A2(n26346),
	.B1(n26345),
	.B2(n26346),
	.C1(n26344),
	.C2(n26346));
   NOR2x1_ASAP7_75t_SL U18587 (.Y(n26729),
	.A(FE_OFN16214_ld_r),
	.B(n25390));
   NAND3xp33_ASAP7_75t_SL U18589 (.Y(n24070),
	.A(n24071),
	.B(FE_OCPN5107_n24418),
	.C(n24147));
   NAND3xp33_ASAP7_75t_L U18590 (.Y(n24068),
	.A(FE_OCPN27815_n25769),
	.B(FE_OCPN28023_n25770),
	.C(n24069));
   OAI21xp5_ASAP7_75t_SL U18591 (.Y(n25486),
	.A1(FE_OFN16213_ld_r),
	.A2(FE_OCPN28077_n),
	.B(n25487));
   NOR3xp33_ASAP7_75t_SL U18592 (.Y(n26439),
	.A(FE_OCPN29458_n26442),
	.B(FE_OFN160_n26440),
	.C(n26441));
   NAND2xp33_ASAP7_75t_SRAM U18593 (.Y(n26827),
	.A(n26831),
	.B(n26824));
   NAND3xp33_ASAP7_75t_R U18594 (.Y(n26828),
	.A(n24888),
	.B(n22674),
	.C(n24887));
   A2O1A1Ixp33_ASAP7_75t_L U18595 (.Y(n26816),
	.A1(n26819),
	.A2(n26818),
	.B(FE_OCPN7633_n26815),
	.C(FE_OCPN27445_n26837));
   NAND2xp5_ASAP7_75t_L U18596 (.Y(n26056),
	.A(n26052),
	.B(FE_OCPN8209_n26051));
   NAND3xp33_ASAP7_75t_SL U18597 (.Y(n24660),
	.A(n24661),
	.B(FE_OCPN27991_n26336),
	.C(n26335));
   NOR3xp33_ASAP7_75t_SL U18598 (.Y(n24657),
	.A(FE_OCPN27226_n25357),
	.B(n24658),
	.C(n24659));
   A2O1A1Ixp33_ASAP7_75t_L U18599 (.Y(n26860),
	.A1(n26829),
	.A2(n26828),
	.B(n24654),
	.C(n24653));
   A2O1A1Ixp33_ASAP7_75t_SL U18600 (.Y(n24653),
	.A1(n26829),
	.A2(n26828),
	.B(n26825),
	.C(n24652));
   NAND2xp5_ASAP7_75t_SL U18601 (.Y(n24654),
	.A(n26824),
	.B(n24651));
   A2O1A1Ixp33_ASAP7_75t_SRAM U18602 (.Y(n25519),
	.A1(FE_OFN16176_n27207),
	.A2(n27192),
	.B(n25514),
	.C(n25513));
   NAND2xp33_ASAP7_75t_SRAM U18603 (.Y(n25514),
	.A(w2_6_),
	.B(FE_OCPN29448_n27189));
   NAND2xp5_ASAP7_75t_L U18604 (.Y(n24879),
	.A(FE_OFN16322_n25946),
	.B(n24876));
   NAND3xp33_ASAP7_75t_L U18606 (.Y(n24909),
	.A(n24910),
	.B(n26824),
	.C(n24911));
   OAI21xp33_ASAP7_75t_SRAM U18607 (.Y(n24911),
	.A1(FE_OCPN27458_n24891),
	.A2(n24890),
	.B(n26829));
   NAND2xp33_ASAP7_75t_L U18608 (.Y(n27055),
	.A(n27046),
	.B(n27045));
   A2O1A1Ixp33_ASAP7_75t_SRAM U18609 (.Y(n27067),
	.A1(n27062),
	.A2(n27061),
	.B(n27060),
	.C(n27059));
   NAND2xp33_ASAP7_75t_SRAM U18610 (.Y(n27060),
	.A(FE_OFN49_w0_23),
	.B(n27057));
   NOR3xp33_ASAP7_75t_SRAM U18611 (.Y(n25830),
	.A(FE_OCPN5053_n25832),
	.B(FE_OCPN27391_n27079),
	.C(n25831));
   NOR3xp33_ASAP7_75t_L U18612 (.Y(n25838),
	.A(FE_OCPN27451_n26236),
	.B(n25839),
	.C(n26235));
   A2O1A1Ixp33_ASAP7_75t_L U18613 (.Y(n25839),
	.A1(n27216),
	.A2(n25837),
	.B(n25836),
	.C(n25835));
   A2O1A1Ixp33_ASAP7_75t_R U18614 (.Y(n25835),
	.A1(n27216),
	.A2(n25837),
	.B(n25834),
	.C(w2_22_));
   A2O1A1Ixp33_ASAP7_75t_L U18616 (.Y(n25567),
	.A1(n27183),
	.A2(n27182),
	.B(n27177),
	.C(n26053));
   OAI222xp33_ASAP7_75t_R U18617 (.Y(n24333),
	.A1(FE_OFN16400_n17404),
	.A2(n24331),
	.B1(n24330),
	.B2(n24331),
	.C1(n24329),
	.C2(n24331));
   NOR2xp33_ASAP7_75t_SRAM U18618 (.Y(n24329),
	.A(n24328),
	.B(n24327));
   NOR3xp33_ASAP7_75t_SRAM U18619 (.Y(n24330),
	.A(n24326),
	.B(n24325),
	.C(n24324));
   NAND3xp33_ASAP7_75t_SL U18620 (.Y(n24500),
	.A(FE_OCPN28235_n26631),
	.B(n24502),
	.C(n24501));
   A2O1A1Ixp33_ASAP7_75t_SL U18621 (.Y(n24501),
	.A1(n27117),
	.A2(n27052),
	.B(n24499),
	.C(n24498));
   NAND2xp33_ASAP7_75t_SL U18622 (.Y(n24499),
	.A(FE_OFN29224_FE_OCPN28074_n27049),
	.B(n24506));
   NAND3xp33_ASAP7_75t_L U18623 (.Y(n24503),
	.A(n24504),
	.B(FE_OCPN28173_n27153),
	.C(FE_OCPN28150_n27152));
   OAI22xp33_ASAP7_75t_SRAM U18624 (.Y(n24505),
	.A1(text_in_r_102_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(n24506),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U18625 (.Y(n25480),
	.A1(n25575),
	.A2(n25475),
	.B(n25474),
	.C(n25473));
   O2A1O1Ixp33_ASAP7_75t_SRAM U18626 (.Y(n26695),
	.A1(FE_OFN16413_n26687),
	.A2(FE_OFN16255_n26684),
	.B(n26689),
	.C(n26688));
   NOR2xp33_ASAP7_75t_SRAM U18627 (.Y(n26689),
	.A(w1_7_),
	.B(FE_OCPN27753_n26685));
   O2A1O1Ixp33_ASAP7_75t_SRAM U18628 (.Y(n26688),
	.A1(FE_OFN16413_n26687),
	.A2(FE_OFN16255_n26684),
	.B(n26686),
	.C(n26692));
   O2A1O1Ixp33_ASAP7_75t_SRAM U18630 (.Y(n26547),
	.A1(n26542),
	.A2(n26541),
	.B(n26540),
	.C(n26539));
   NOR2xp33_ASAP7_75t_SRAM U18631 (.Y(n26540),
	.A(w0_7_),
	.B(FE_OCPN29481_n26537));
   O2A1O1Ixp33_ASAP7_75t_SRAM U18632 (.Y(n26539),
	.A1(n26542),
	.A2(n26541),
	.B(n26538),
	.C(n26544));
   XNOR2x2_ASAP7_75t_SL U18634 (.Y(n16055),
	.A(u0_rcon_31_),
	.B(n14088));
   A2O1A1Ixp33_ASAP7_75t_SL U18635 (.Y(n14088),
	.A1(n13867),
	.A2(n14087),
	.B(n14086),
	.C(n14085));
   NAND2xp33_ASAP7_75t_SL U18636 (.Y(n14086),
	.A(w0_31_),
	.B(n14083));
   NAND3xp33_ASAP7_75t_SL U18638 (.Y(n14182),
	.A(n14111),
	.B(n14110),
	.C(n14109));
   AOI22x1_ASAP7_75t_SL U18639 (.Y(n15367),
	.A1(w1_5_),
	.A2(n14004),
	.B1(FE_OFN16239_n14005),
	.B2(n24149));
   XNOR2x2_ASAP7_75t_SL U18640 (.Y(n15906),
	.A(u0_rcon_28_),
	.B(n13937));
   A2O1A1Ixp33_ASAP7_75t_SL U18641 (.Y(n13937),
	.A1(n13867),
	.A2(n13936),
	.B(n13935),
	.C(n13934));
   NAND2xp33_ASAP7_75t_SL U18642 (.Y(n13935),
	.A(w0_28_),
	.B(n13932));
   XNOR2x1_ASAP7_75t_SL U18643 (.Y(n16216),
	.A(w1_27_),
	.B(n16135));
   NAND2xp33_ASAP7_75t_SL U18644 (.Y(n15058),
	.A(n15056),
	.B(n24641));
   XNOR2x1_ASAP7_75t_SL U18646 (.Y(n16258),
	.A(w1_24_),
	.B(n16163));
   NAND2xp33_ASAP7_75t_L U18647 (.Y(n15141),
	.A(n15138),
	.B(n27160));
   NAND2xp33_ASAP7_75t_L U18648 (.Y(n15142),
	.A(n15073),
	.B(n15072));
   OAI21x1_ASAP7_75t_SL U18649 (.Y(n16172),
	.A1(n16145),
	.A2(n27135),
	.B(n16144));
   O2A1O1Ixp33_ASAP7_75t_SL U18651 (.Y(n14472),
	.A1(n13722),
	.A2(n13721),
	.B(w0_0_),
	.C(n13720));
   OAI222xp33_ASAP7_75t_L U18652 (.Y(n13721),
	.A1(n13719),
	.A2(n15259),
	.B1(n13718),
	.B2(n15259),
	.C1(n13717),
	.C2(n15259));
   OAI21x1_ASAP7_75t_SL U18653 (.Y(n16086),
	.A1(w2_0_),
	.A2(n16082),
	.B(n16081));
   NOR2xp33_ASAP7_75t_SRAM U18654 (.Y(n16168),
	.A(key_22_),
	.B(FE_OFN28458_ld));
   NOR2xp33_ASAP7_75t_SRAM U18655 (.Y(n16154),
	.A(key_7_),
	.B(FE_OFN26_n16125));
   OAI21xp5_ASAP7_75t_SL U18656 (.Y(n651),
	.A1(FE_OCPN29550_n16114),
	.A2(FE_OCPN29502_w3_23),
	.B(n16071));
   NOR2xp33_ASAP7_75t_SRAM U18657 (.Y(n16070),
	.A(key_23_),
	.B(FE_OFN26_n16125));
   OAI21xp5_ASAP7_75t_SL U18658 (.Y(n626),
	.A1(FE_OFN25892_n16264),
	.A2(FE_OFN28858_FE_OCPN27664_w3_25),
	.B(n16239));
   NOR2xp33_ASAP7_75t_SRAM U18659 (.Y(n16238),
	.A(key_25_),
	.B(FE_OFN28472_ld));
   OAI21xp33_ASAP7_75t_SL U18660 (.Y(n640),
	.A1(n16201),
	.A2(FE_OCPN29520_n24755),
	.B(n16181));
   NOR2xp33_ASAP7_75t_SRAM U18661 (.Y(n16180),
	.A(key_12_),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SL U18662 (.Y(n652),
	.A1(n16148),
	.A2(FE_OFN26129_w3_15),
	.B(n16129));
   NOR2xp33_ASAP7_75t_SRAM U18663 (.Y(n16128),
	.A(key_15_),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SL U18664 (.Y(n628),
	.A1(n16240),
	.A2(FE_OFN26163_w3_13),
	.B(n16196));
   NOR2xp33_ASAP7_75t_SRAM U18665 (.Y(n16195),
	.A(key_13_),
	.B(FE_OFN28457_ld));
   NOR2xp33_ASAP7_75t_SRAM U18666 (.Y(n16160),
	.A(key_26_),
	.B(FE_OFN28470_ld));
   NOR2xp33_ASAP7_75t_SRAM U18667 (.Y(n16245),
	.A(key_18_),
	.B(FE_OFN28461_ld));
   NOR2xp33_ASAP7_75t_SRAM U18668 (.Y(n16220),
	.A(key_10_),
	.B(FE_OFN25_n16125));
   NOR2xp33_ASAP7_75t_SRAM U18670 (.Y(n15913),
	.A(key_2_),
	.B(FE_OFN26139_n16125));
   OAI21xp33_ASAP7_75t_SL U18671 (.Y(n642),
	.A1(FE_OFN16246_n16113),
	.A2(FE_OFN27129_w3_28),
	.B(n16112));
   NOR2xp33_ASAP7_75t_SRAM U18672 (.Y(n16111),
	.A(key_28_),
	.B(FE_OFN28470_ld));
   NOR2xp33_ASAP7_75t_SRAM U18673 (.Y(n16108),
	.A(key_21_),
	.B(FE_OFN26_n16125));
   NOR2xp33_ASAP7_75t_SRAM U18675 (.Y(n16187),
	.A(key_29_),
	.B(FE_OFN28470_ld));
   NAND2xp5_ASAP7_75t_L U18676 (.Y(n14507),
	.A(n14502),
	.B(n14501));
   NAND2xp33_ASAP7_75t_L U18677 (.Y(n14501),
	.A(n14500),
	.B(FE_OFN28455_n13348));
   NAND2xp33_ASAP7_75t_SL U18678 (.Y(n14502),
	.A(n14499),
	.B(FE_OFN28455_n13348));
   NOR2xp33_ASAP7_75t_SL U18679 (.Y(n14499),
	.A(FE_OFN27206_w3_30),
	.B(n14498));
   NOR2xp33_ASAP7_75t_L U18680 (.Y(n14544),
	.A(n15182),
	.B(FE_OFN27061_n15239));
   NAND2xp5_ASAP7_75t_L U18681 (.Y(n14565),
	.A(n14561),
	.B(n14560));
   NAND2xp5_ASAP7_75t_L U18682 (.Y(n14561),
	.A(n14558),
	.B(n14559));
   INVx1_ASAP7_75t_L U18683 (.Y(n14567),
	.A(n14563));
   NOR2xp67_ASAP7_75t_L U18684 (.Y(n15229),
	.A(FE_OFN25875_n15227),
	.B(n15226));
   NOR2xp67_ASAP7_75t_L U18685 (.Y(n15225),
	.A(n15222),
	.B(n15226));
   OR2x2_ASAP7_75t_L U18686 (.Y(n15228),
	.A(FE_OFN27085_n),
	.B(n15223));
   O2A1O1Ixp33_ASAP7_75t_SL U18687 (.Y(n14118),
	.A1(FE_OFN26642_w3_14),
	.A2(FE_OFN29063_n25433),
	.B(FE_OFN27135_n15992),
	.C(FE_OFN109_n15994));
   NOR2xp33_ASAP7_75t_SL U18688 (.Y(n13603),
	.A(n14515),
	.B(n13604));
   NAND2xp33_ASAP7_75t_SL U18689 (.Y(n13607),
	.A(n13606),
	.B(n13605));
   NOR2xp33_ASAP7_75t_R U18690 (.Y(n13606),
	.A(FE_OFN25875_n15227),
	.B(n13604));
   INVx1_ASAP7_75t_L U18691 (.Y(n13599),
	.A(n13530));
   NAND2xp5_ASAP7_75t_L U18692 (.Y(n14556),
	.A(FE_OCPN29428_FE_OFN27131_w3_29),
	.B(n26355));
   INVxp67_ASAP7_75t_L U18693 (.Y(n16005),
	.A(n16001));
   NOR2xp33_ASAP7_75t_SRAM U18694 (.Y(n16014),
	.A(n16009),
	.B(n16015));
   NOR2xp33_ASAP7_75t_SRAM U18695 (.Y(n16018),
	.A(FE_OFN26131_n15376),
	.B(n16015));
   NAND2xp33_ASAP7_75t_SRAM U18696 (.Y(n14523),
	.A(n14520),
	.B(FE_OFN26112_n13288));
   NOR2xp33_ASAP7_75t_SRAM U18697 (.Y(n14520),
	.A(FE_OFN27211_w3_30),
	.B(n15200));
   NOR2xp33_ASAP7_75t_R U18698 (.Y(n14524),
	.A(n15222),
	.B(n14525));
   NOR2xp33_ASAP7_75t_R U18699 (.Y(n14506),
	.A(n15224),
	.B(n14507));
   INVxp67_ASAP7_75t_L U18700 (.Y(n14508),
	.A(n14505));
   NOR2xp33_ASAP7_75t_L U18701 (.Y(n14509),
	.A(n15223),
	.B(n14507));
   NAND2xp33_ASAP7_75t_L U18702 (.Y(n14539),
	.A(n14537),
	.B(n14536));
   NAND2xp33_ASAP7_75t_SRAM U18703 (.Y(n14537),
	.A(n14534),
	.B(FE_OFN28456_n13348));
   NOR2xp33_ASAP7_75t_SRAM U18704 (.Y(n14581),
	.A(n14579),
	.B(n14578));
   NAND2xp33_ASAP7_75t_SL U18705 (.Y(n14570),
	.A(n14564),
	.B(n14567));
   NOR2xp33_ASAP7_75t_R U18706 (.Y(n14564),
	.A(FE_OFN25875_n15227),
	.B(n14565));
   NAND2xp5_ASAP7_75t_R U18707 (.Y(n14569),
	.A(n14568),
	.B(n14567));
   NOR2xp33_ASAP7_75t_L U18708 (.Y(n14568),
	.A(n14566),
	.B(n14565));
   NAND2xp33_ASAP7_75t_R U18709 (.Y(n14583),
	.A(n14577),
	.B(n14580));
   NAND2xp33_ASAP7_75t_L U18710 (.Y(n14484),
	.A(n14478),
	.B(n14477));
   NAND2xp33_ASAP7_75t_L U18711 (.Y(n14477),
	.A(n14476),
	.B(n14475));
   NAND2xp33_ASAP7_75t_L U18712 (.Y(n14478),
	.A(n14500),
	.B(n14475));
   INVxp33_ASAP7_75t_SRAM U18713 (.Y(n14475),
	.A(n14556));
   NOR2xp33_ASAP7_75t_SRAM U18714 (.Y(n15241),
	.A(n15239),
	.B(n15238));
   NOR2xp33_ASAP7_75t_R U18715 (.Y(n14117),
	.A(n15927),
	.B(n14118));
   NAND2xp33_ASAP7_75t_L U18716 (.Y(n14121),
	.A(n14120),
	.B(n14119));
   NOR2xp33_ASAP7_75t_L U18717 (.Y(n14120),
	.A(n15934),
	.B(n14118));
   INVxp67_ASAP7_75t_L U18718 (.Y(n14145),
	.A(n14614));
   NAND2xp5_ASAP7_75t_R U18719 (.Y(n14147),
	.A(n14146),
	.B(n14145));
   NOR2xp33_ASAP7_75t_L U18720 (.Y(n14146),
	.A(n15444),
	.B(n14927));
   NAND2xp5_ASAP7_75t_L U18721 (.Y(n14797),
	.A(n14794),
	.B(n14793));
   NAND2xp33_ASAP7_75t_SL U18722 (.Y(n14793),
	.A(n14792),
	.B(FE_OFN25981_n13868));
   NAND2xp33_ASAP7_75t_SL U18723 (.Y(n14794),
	.A(n15478),
	.B(FE_OFN25981_n13868));
   NAND2xp5_ASAP7_75t_SL U18724 (.Y(n14044),
	.A(n13916),
	.B(n14042));
   NAND2xp5_ASAP7_75t_L U18725 (.Y(n13612),
	.A(n13601),
	.B(n13600));
   NAND2xp33_ASAP7_75t_L U18726 (.Y(n13600),
	.A(n13599),
	.B(FE_OFN75_n15253));
   NAND2xp33_ASAP7_75t_SL U18727 (.Y(n13601),
	.A(n13597),
	.B(FE_OFN75_n15253));
   NOR3x1_ASAP7_75t_SL U18729 (.Y(n15425),
	.A(n15375),
	.B(n15380),
	.C(FE_OFN26007_n16010));
   NAND2xp5_ASAP7_75t_SL U18730 (.Y(n13602),
	.A(n13350),
	.B(n13349));
   NAND2xp5_ASAP7_75t_L U18731 (.Y(n13349),
	.A(n13519),
	.B(FE_OFN28456_n13348));
   NOR2xp33_ASAP7_75t_SL U18732 (.Y(n15427),
	.A(FE_OCPN29509_FE_OFN16184_w3_9),
	.B(n15425));
   NOR2xp33_ASAP7_75t_SL U18733 (.Y(n15424),
	.A(FE_OCPN29583_n15422),
	.B(n15425));
   NOR3xp33_ASAP7_75t_R U18734 (.Y(n14292),
	.A(FE_OFN16210_n13876),
	.B(n15536),
	.C(n14377));
   NAND2x1_ASAP7_75t_SL U18735 (.Y(n15226),
	.A(n13430),
	.B(n13429));
   NAND2xp5_ASAP7_75t_SL U18736 (.Y(n13430),
	.A(n13599),
	.B(FE_OFN28456_n13348));
   NAND2xp5_ASAP7_75t_SL U18737 (.Y(n13429),
	.A(n14515),
	.B(FE_OFN28456_n13348));
   OA21x2_ASAP7_75t_L U18738 (.Y(n13433),
	.A1(n15217),
	.A2(n15203),
	.B(n13431));
   NAND2xp33_ASAP7_75t_R U18739 (.Y(n13431),
	.A(FE_OFN26049_w3_27),
	.B(n15188));
   INVxp67_ASAP7_75t_R U18740 (.Y(n13440),
	.A(n13438));
   OAI21xp33_ASAP7_75t_L U18741 (.Y(n15860),
	.A1(FE_OFN28695_n),
	.A2(n15862),
	.B(n15787));
   OA21x2_ASAP7_75t_L U18742 (.Y(n15521),
	.A1(n15517),
	.A2(n15480),
	.B(n15516));
   NAND3xp33_ASAP7_75t_R U18743 (.Y(n15516),
	.A(n15729),
	.B(FE_OFN26053_n25415),
	.C(FE_OFN28977_n));
   OAI21xp5_ASAP7_75t_SL U18744 (.Y(n15687),
	.A1(n15680),
	.A2(n15480),
	.B(n15679));
   O2A1O1Ixp33_ASAP7_75t_R U18745 (.Y(n15697),
	.A1(FE_OFN6_w3_22),
	.A2(n15694),
	.B(n15719),
	.C(FE_OFN27074_n13868));
   O2A1O1Ixp33_ASAP7_75t_L U18746 (.Y(n13676),
	.A1(FE_OFN27057_n13662),
	.A2(n14556),
	.B(FE_OFN25893_n15214),
	.C(n15209));
   NAND2xp5_ASAP7_75t_SL U18747 (.Y(n14426),
	.A(n15124),
	.B(n15842));
   NAND2xp33_ASAP7_75t_SL U18748 (.Y(n15962),
	.A(n15952),
	.B(n15951));
   NAND2xp33_ASAP7_75t_R U18749 (.Y(n15952),
	.A(n16009),
	.B(n15950));
   NAND2xp33_ASAP7_75t_SRAM U18750 (.Y(n15951),
	.A(n15972),
	.B(n15950));
   INVxp67_ASAP7_75t_L U18752 (.Y(n15964),
	.A(n15960));
   NAND3xp33_ASAP7_75t_SRAM U18753 (.Y(n15957),
	.A(n15956),
	.B(n15955),
	.C(n15954));
   NAND2xp33_ASAP7_75t_SRAM U18754 (.Y(n15974),
	.A(FE_OFN29017_n15921),
	.B(n15973));
   NAND2xp33_ASAP7_75t_L U18755 (.Y(n16007),
	.A(n16006),
	.B(n16005));
   NOR2xp33_ASAP7_75t_L U18756 (.Y(n16006),
	.A(n16004),
	.B(n16003));
   NAND2xp33_ASAP7_75t_L U18757 (.Y(n16008),
	.A(n16002),
	.B(n16005));
   NOR2xp33_ASAP7_75t_SRAM U18758 (.Y(n16002),
	.A(n14924),
	.B(n16003));
   NOR3xp33_ASAP7_75t_SRAM U18759 (.Y(n15996),
	.A(FE_OFN109_n15994),
	.B(n15993),
	.C(n15992));
   NAND2xp33_ASAP7_75t_L U18760 (.Y(n16021),
	.A(n16020),
	.B(n16019));
   NAND2xp5_ASAP7_75t_L U18761 (.Y(n16019),
	.A(n16018),
	.B(n16017));
   NAND2xp33_ASAP7_75t_R U18762 (.Y(n16020),
	.A(n16014),
	.B(n16017));
   INVxp33_ASAP7_75t_L U18763 (.Y(n16017),
	.A(n16013));
   NOR2xp33_ASAP7_75t_SL U18764 (.Y(n17801),
	.A(FE_OCPN27771_n19275),
	.B(n22533));
   NOR2xp33_ASAP7_75t_R U18766 (.Y(n17069),
	.A(FE_OCPN28212_n16980),
	.B(n20513));
   NAND2xp33_ASAP7_75t_SL U18774 (.Y(n14047),
	.A(n14045),
	.B(n14044));
   NAND2xp5_ASAP7_75t_R U18775 (.Y(n14045),
	.A(n14043),
	.B(n14042));
   NAND2xp33_ASAP7_75t_L U18777 (.Y(n14064),
	.A(n14062),
	.B(n14061));
   NOR2xp33_ASAP7_75t_R U18778 (.Y(n14062),
	.A(n15501),
	.B(n13875));
   INVxp33_ASAP7_75t_SRAM U18779 (.Y(n14030),
	.A(n14276));
   NAND2xp33_ASAP7_75t_SRAM U18780 (.Y(n14032),
	.A(n15347),
	.B(FE_OFN28600_n14289));
   NAND2xp5_ASAP7_75t_L U18781 (.Y(n14530),
	.A(n14529),
	.B(n14528));
   NAND2xp5_ASAP7_75t_R U18782 (.Y(n14529),
	.A(n14524),
	.B(n14526));
   NAND2xp5_ASAP7_75t_R U18783 (.Y(n14528),
	.A(n14527),
	.B(n14526));
   AND2x2_ASAP7_75t_L U18784 (.Y(n14526),
	.A(n14523),
	.B(n14522));
   NOR2xp33_ASAP7_75t_SL U18785 (.Y(n14513),
	.A(n14512),
	.B(FE_OFN16412_w3_26));
   NAND2xp5_ASAP7_75t_L U18786 (.Y(n14512),
	.A(n14511),
	.B(n14510));
   NAND2xp33_ASAP7_75t_L U18787 (.Y(n14510),
	.A(n14509),
	.B(n14508));
   NAND2xp33_ASAP7_75t_L U18788 (.Y(n14511),
	.A(n14506),
	.B(n14508));
   NOR2xp33_ASAP7_75t_R U18789 (.Y(n14483),
	.A(n15189),
	.B(n14484));
   OA21x2_ASAP7_75t_L U18790 (.Y(n14486),
	.A1(FE_OCPN27656_w3_25),
	.A2(n15200),
	.B(n14482));
   OAI22xp33_ASAP7_75t_SRAM U18791 (.Y(n14481),
	.A1(n25675),
	.A2(n14479),
	.B1(FE_OCPN29571_n26355),
	.B2(n14479));
   NOR2xp33_ASAP7_75t_R U18792 (.Y(n14487),
	.A(n14485),
	.B(n14484));
   O2A1O1Ixp5_ASAP7_75t_L U18793 (.Y(n14213),
	.A1(FE_OFN28662_w3_7),
	.A2(n13730),
	.B(FE_OFN28889_n15845),
	.C(n14210));
   O2A1O1Ixp33_ASAP7_75t_L U18794 (.Y(n14231),
	.A1(FE_OFN27156_n),
	.A2(FE_OFN28732_n),
	.B(n15842),
	.C(n13725));
   AND2x2_ASAP7_75t_SRAM U18795 (.Y(n14232),
	.A(n14229),
	.B(n14228));
   NAND2xp33_ASAP7_75t_SRAM U18796 (.Y(n14229),
	.A(n15862),
	.B(n15074));
   NAND2xp33_ASAP7_75t_R U18797 (.Y(n14228),
	.A(n15636),
	.B(n15074));
   OAI21xp5_ASAP7_75t_L U18798 (.Y(n14223),
	.A1(n15813),
	.A2(n15847),
	.B(n14220));
   NOR2xp33_ASAP7_75t_L U18799 (.Y(n14116),
	.A(n13949),
	.B(FE_OFN26007_n16010));
   NAND2xp5_ASAP7_75t_SRAM U18800 (.Y(n14373),
	.A(n15487),
	.B(FE_OFN28827_n15683));
   NAND2xp33_ASAP7_75t_R U18801 (.Y(n14372),
	.A(n14371),
	.B(FE_OFN28827_n15683));
   NOR2xp33_ASAP7_75t_SRAM U18802 (.Y(n15219),
	.A(n15217),
	.B(n15216));
   OAI21xp5_ASAP7_75t_SRAM U18803 (.Y(n15168),
	.A1(FE_OFN26049_w3_27),
	.A2(n14504),
	.B(n13582));
   NAND3xp33_ASAP7_75t_SRAM U18804 (.Y(n13582),
	.A(FE_OFN27207_w3_30),
	.B(FE_OCPN27659_w3_25),
	.C(FE_OFN16145_n15214));
   OA21x2_ASAP7_75t_SRAM U18805 (.Y(n15866),
	.A1(n15862),
	.A2(n15861),
	.B(n15860));
   NOR2xp33_ASAP7_75t_L U18807 (.Y(n15823),
	.A(n15033),
	.B(FE_OFN28792_n15787));
   NOR3xp33_ASAP7_75t_SRAM U18808 (.Y(n14126),
	.A(n14714),
	.B(FE_OFN27200_n),
	.C(FE_OCPN29570_n15423));
   NOR2xp33_ASAP7_75t_SRAM U18809 (.Y(n14161),
	.A(n15411),
	.B(n14666));
   NAND2xp33_ASAP7_75t_SL U18810 (.Y(n14163),
	.A(n14158),
	.B(n14160));
   NOR2xp33_ASAP7_75t_SRAM U18811 (.Y(n14158),
	.A(n13844),
	.B(n14666));
   NAND2xp5_ASAP7_75t_L U18812 (.Y(n14152),
	.A(n14142),
	.B(n14141));
   NAND2xp33_ASAP7_75t_L U18813 (.Y(n14142),
	.A(n14138),
	.B(FE_OFN28543_FE_OFN109_n15994));
   NAND2xp33_ASAP7_75t_L U18814 (.Y(n14141),
	.A(n14140),
	.B(FE_OFN28543_FE_OFN109_n15994));
   NOR2xp33_ASAP7_75t_R U18815 (.Y(n14151),
	.A(n14940),
	.B(n14152));
   NAND2xp5_ASAP7_75t_L U18816 (.Y(n15999),
	.A(FE_OFN27115_n),
	.B(FE_OFN26640_w3_14));
   NOR2xp33_ASAP7_75t_SL U18817 (.Y(n14796),
	.A(n15528),
	.B(n14797));
   NOR2xp33_ASAP7_75t_L U18818 (.Y(n14800),
	.A(n14798),
	.B(n14797));
   NOR2xp33_ASAP7_75t_L U18819 (.Y(n14777),
	.A(n12994),
	.B(n14779));
   NOR3xp33_ASAP7_75t_R U18820 (.Y(n14779),
	.A(n13875),
	.B(FE_OFN28551_FE_OFN26114_n),
	.C(n15714));
   OAI21xp33_ASAP7_75t_L U18821 (.Y(n13289),
	.A1(n14498),
	.A2(n15201),
	.B(FE_OFN16193_n15200));
   NOR2xp33_ASAP7_75t_R U18822 (.Y(n13747),
	.A(n15859),
	.B(n13745));
   OA21x2_ASAP7_75t_R U18823 (.Y(n13746),
	.A1(n13743),
	.A2(n15639),
	.B(n14426));
   NOR2xp33_ASAP7_75t_SRAM U18824 (.Y(n13743),
	.A(n13729),
	.B(n14996));
   NOR2xp33_ASAP7_75t_SL U18825 (.Y(n13744),
	.A(n15019),
	.B(n13745));
   NOR2xp33_ASAP7_75t_SRAM U18826 (.Y(n14194),
	.A(n15808),
	.B(n14442));
   NOR3xp33_ASAP7_75t_L U18827 (.Y(n15997),
	.A(FE_OCPN29570_n15423),
	.B(FE_OFN27200_n),
	.C(n16009));
   OA21x2_ASAP7_75t_L U18828 (.Y(n14048),
	.A1(n14795),
	.A2(n15480),
	.B(n13904));
   NAND2xp5_ASAP7_75t_L U18829 (.Y(n14068),
	.A(FE_OFN26091_n24663),
	.B(FE_OCPN28404_n13874));
   OAI21xp5_ASAP7_75t_L U18830 (.Y(n15079),
	.A1(FE_OFN28747_n),
	.A2(n15034),
	.B(n13783));
   NOR2xp33_ASAP7_75t_L U18831 (.Y(n14867),
	.A(n15829),
	.B(FE_OFN28691_n13725));
   NOR2xp33_ASAP7_75t_SL U18832 (.Y(n15107),
	.A(n15034),
	.B(n13741));
   NAND3xp33_ASAP7_75t_SRAM U18834 (.Y(n14639),
	.A(FE_OFN26642_w3_14),
	.B(n15987),
	.C(FE_OFN26624_n15376));
   O2A1O1Ixp5_ASAP7_75t_SRAM U18835 (.Y(n14638),
	.A1(FE_OFN28884_n),
	.A2(FE_OFN28856_n15450),
	.B(n13844),
	.C(n15425));
   INVxp67_ASAP7_75t_L U18836 (.Y(n15954),
	.A(n15435));
   OAI21xp5_ASAP7_75t_L U18837 (.Y(n15344),
	.A1(n13875),
	.A2(n15520),
	.B(n15342));
   NOR2xp33_ASAP7_75t_SL U18838 (.Y(n15340),
	.A(n15339),
	.B(FE_OFN28909_w3_23));
   OA21x2_ASAP7_75t_L U18839 (.Y(n15324),
	.A1(FE_OCPN8216_n13916),
	.A2(FE_OFN27074_n13868),
	.B(n15321));
   O2A1O1Ixp33_ASAP7_75t_SRAM U18841 (.Y(n15320),
	.A1(FE_OFN26091_n24663),
	.A2(n15484),
	.B(FE_PSN8334_n15539),
	.C(n13875));
   NOR2xp33_ASAP7_75t_SRAM U18842 (.Y(n15299),
	.A(n13916),
	.B(n15297));
   NOR3xp33_ASAP7_75t_SRAM U18845 (.Y(n13392),
	.A(n15223),
	.B(n15259),
	.C(n14504));
   OAI21xp33_ASAP7_75t_SRAM U18846 (.Y(n13391),
	.A1(FE_OFN26051_w3_27),
	.A2(FE_OCPN27665_w3_25),
	.B(FE_OFN27210_w3_30));
   AND2x2_ASAP7_75t_L U18847 (.Y(n13373),
	.A(n13369),
	.B(FE_OFN28456_n13348));
   NOR2xp33_ASAP7_75t_SRAM U18848 (.Y(n13369),
	.A(n14500),
	.B(n13459));
   NOR2xp33_ASAP7_75t_R U18849 (.Y(n13353),
	.A(FE_OCPN27656_w3_25),
	.B(n13602));
   NAND2xp33_ASAP7_75t_SL U18850 (.Y(n13355),
	.A(n13351),
	.B(n13352));
   NOR2xp33_ASAP7_75t_SL U18851 (.Y(n13351),
	.A(n14593),
	.B(n13602));
   NOR2xp33_ASAP7_75t_R U18852 (.Y(n15003),
	.A(FE_OFN26531_n),
	.B(n15888));
   NAND3xp33_ASAP7_75t_L U18854 (.Y(n15625),
	.A(FE_OFN28661_w3_7),
	.B(n13736),
	.C(FE_OFN28695_n));
   NAND2xp33_ASAP7_75t_SL U18856 (.Y(n15432),
	.A(n15429),
	.B(n15428));
   NAND2xp5_ASAP7_75t_SL U18857 (.Y(n15429),
	.A(n15424),
	.B(n15426));
   NAND2xp5_ASAP7_75t_L U18858 (.Y(n15428),
	.A(n15427),
	.B(n15426));
   NAND3xp33_ASAP7_75t_L U18859 (.Y(n15435),
	.A(n14924),
	.B(FE_OFN25961_w3_8),
	.C(w3_10_));
   NOR2xp33_ASAP7_75t_SRAM U18861 (.Y(n14334),
	.A(n15660),
	.B(FE_OCPN8264_n13890));
   NAND2xp5_ASAP7_75t_R U18862 (.Y(n14302),
	.A(n14288),
	.B(n14287));
   NAND2xp33_ASAP7_75t_L U18863 (.Y(n14287),
	.A(n14286),
	.B(FE_OFN27066_n13869));
   NAND2xp33_ASAP7_75t_L U18864 (.Y(n14288),
	.A(FE_OFN28769_n15478),
	.B(FE_OFN27066_n13869));
   NOR2xp33_ASAP7_75t_R U18865 (.Y(n14286),
	.A(FE_OCPN28404_n13874),
	.B(FE_PSN8280_n15660));
   INVxp67_ASAP7_75t_L U18866 (.Y(n15698),
	.A(n13891));
   NOR2xp33_ASAP7_75t_L U18867 (.Y(n14314),
	.A(FE_OCPN27987_FE_OFN4_w3_22),
	.B(n13876));
   NAND2xp5_ASAP7_75t_L U18868 (.Y(n14747),
	.A(FE_OFN4_w3_22),
	.B(n13874));
   NOR3xp33_ASAP7_75t_SRAM U18869 (.Y(n14806),
	.A(n13875),
	.B(FE_OFN28701_w3_16),
	.C(FE_OFN50_w3_18));
   NAND2xp5_ASAP7_75t_R U18870 (.Y(n13436),
	.A(n13432),
	.B(n13433));
   NOR2xp33_ASAP7_75t_SRAM U18871 (.Y(n13432),
	.A(n14593),
	.B(n15226));
   NAND2xp5_ASAP7_75t_L U18872 (.Y(n13435),
	.A(n13434),
	.B(n13433));
   NOR2xp33_ASAP7_75t_SRAM U18873 (.Y(n13434),
	.A(n15156),
	.B(n15226));
   NAND2xp33_ASAP7_75t_L U18874 (.Y(n13443),
	.A(n13439),
	.B(n13440));
   NOR2xp33_ASAP7_75t_SRAM U18875 (.Y(n13439),
	.A(n14500),
	.B(n13437));
   NAND2xp33_ASAP7_75t_R U18876 (.Y(n13442),
	.A(n13441),
	.B(n13440));
   NOR2xp33_ASAP7_75t_R U18877 (.Y(n13441),
	.A(FE_OFN16145_n15214),
	.B(n13437));
   INVxp33_ASAP7_75t_L U18878 (.Y(n13461),
	.A(n13460));
   NAND2xp5_ASAP7_75t_SL U18879 (.Y(n13464),
	.A(n13458),
	.B(n13457));
   NAND2xp33_ASAP7_75t_SL U18880 (.Y(n13458),
	.A(n13453),
	.B(n13455));
   OA21x2_ASAP7_75t_SRAM U18881 (.Y(n15611),
	.A1(n15636),
	.A2(n15607),
	.B(n15606));
   NAND2xp33_ASAP7_75t_SRAM U18882 (.Y(n15606),
	.A(FE_OFN25912_n15848),
	.B(n15636));
   O2A1O1Ixp33_ASAP7_75t_R U18884 (.Y(n15630),
	.A1(FE_OFN28695_n),
	.A2(n13771),
	.B(n15625),
	.C(FE_OFN25900_w3_4));
   INVxp67_ASAP7_75t_L U18885 (.Y(n15631),
	.A(n15628));
   OAI21xp33_ASAP7_75t_L U18886 (.Y(n15587),
	.A1(n13766),
	.A2(n15825),
	.B(n15586));
   NOR2xp33_ASAP7_75t_R U18887 (.Y(n15591),
	.A(n15829),
	.B(FE_OFN25928_n15779));
   NAND2xp5_ASAP7_75t_R U18889 (.Y(n14938),
	.A(FE_OCPN29535_FE_OFN8_w3_14),
	.B(n15972));
   NAND2xp33_ASAP7_75t_L U18890 (.Y(n15545),
	.A(n15538),
	.B(n15537));
   NAND2xp33_ASAP7_75t_SL U18891 (.Y(n15538),
	.A(n15534),
	.B(FE_OFN25981_n13868));
   INVxp67_ASAP7_75t_L U18892 (.Y(n15508),
	.A(n15504));
   INVxp67_ASAP7_75t_R U18893 (.Y(n15502),
	.A(n15715));
   OAI21xp33_ASAP7_75t_R U18894 (.Y(n15503),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(n15501),
	.B(n15729));
   NAND2xp33_ASAP7_75t_L U18895 (.Y(n15524),
	.A(n15518),
	.B(n15521));
   NOR2xp33_ASAP7_75t_SL U18896 (.Y(n15518),
	.A(n15683),
	.B(n15519));
   NAND2xp33_ASAP7_75t_L U18897 (.Y(n15523),
	.A(n15522),
	.B(n15521));
   NOR2xp33_ASAP7_75t_SL U18898 (.Y(n15522),
	.A(n15520),
	.B(n15519));
   NAND3xp33_ASAP7_75t_SL U18899 (.Y(n15513),
	.A(FE_OCPN28278_n15512),
	.B(FE_PSN8276_FE_OFN28712_n),
	.C(FE_OFN28628_n15667));
   NOR2x1_ASAP7_75t_SL U18900 (.Y(n13519),
	.A(FE_OFN26111_n13288),
	.B(n15201));
   NOR2xp33_ASAP7_75t_SRAM U18901 (.Y(n15119),
	.A(n13729),
	.B(n13741));
   OA21x2_ASAP7_75t_SL U18902 (.Y(n15120),
	.A1(n15639),
	.A2(n15626),
	.B(n15116));
   NOR3xp33_ASAP7_75t_L U18903 (.Y(n15637),
	.A(n15079),
	.B(FE_OFN28662_w3_7),
	.C(FE_OFN26073_n));
   NOR2xp33_ASAP7_75t_L U18904 (.Y(n14722),
	.A(n15936),
	.B(FE_OCPN29521_n24755));
   NAND3xp33_ASAP7_75t_SRAM U18905 (.Y(n15398),
	.A(n24755),
	.B(FE_PSN8324_n15987),
	.C(n15922));
   NOR2xp33_ASAP7_75t_SL U18906 (.Y(n14371),
	.A(FE_OFN26045_n25377),
	.B(FE_OFN26053_n25415));
   NAND2xp33_ASAP7_75t_SRAM U18907 (.Y(n15684),
	.A(FE_OFN25915_n15514),
	.B(n15683));
   INVxp33_ASAP7_75t_L U18908 (.Y(n15685),
	.A(n15682));
   NOR2xp33_ASAP7_75t_SL U18909 (.Y(n15686),
	.A(n15681),
	.B(n15687));
   NOR2xp33_ASAP7_75t_SRAM U18910 (.Y(n15681),
	.A(n15713),
	.B(FE_OCPN8264_n13890));
   NOR2xp33_ASAP7_75t_SL U18911 (.Y(n15690),
	.A(n15688),
	.B(n15687));
   NOR2xp33_ASAP7_75t_L U18912 (.Y(n15696),
	.A(n12994),
	.B(n15697));
   NOR2xp33_ASAP7_75t_L U18913 (.Y(n15700),
	.A(n15698),
	.B(n15697));
   NOR2xp33_ASAP7_75t_L U18914 (.Y(n15718),
	.A(n12994),
	.B(n15715));
   INVx1_ASAP7_75t_SL U18915 (.Y(n15721),
	.A(n15717));
   NOR3xp33_ASAP7_75t_SL U18916 (.Y(n15717),
	.A(FE_OFN29192_n13870),
	.B(FE_OFN28909_w3_23),
	.C(n15726));
   NOR2xp33_ASAP7_75t_SL U18917 (.Y(n15748),
	.A(n15729),
	.B(n15749));
   NAND2xp5_ASAP7_75t_R U18922 (.Y(n13672),
	.A(n15224),
	.B(n13670));
   NOR2xp33_ASAP7_75t_L U18923 (.Y(n13675),
	.A(FE_OFN28455_n13348),
	.B(n13676));
   NOR2xp33_ASAP7_75t_L U18924 (.Y(n13679),
	.A(n13677),
	.B(n13676));
   NOR3xp33_ASAP7_75t_SRAM U18925 (.Y(n15118),
	.A(n15639),
	.B(FE_OFN27156_n),
	.C(FE_OFN28732_n));
   NAND2xp5_ASAP7_75t_L U18926 (.Y(n15607),
	.A(n15859),
	.B(n15822));
   NOR2xp33_ASAP7_75t_SRAM U18927 (.Y(n14412),
	.A(n15838),
	.B(n15809));
   NAND2xp33_ASAP7_75t_SL U18928 (.Y(n15967),
	.A(n15961),
	.B(n15964));
   NOR2xp33_ASAP7_75t_R U18929 (.Y(n15961),
	.A(n15953),
	.B(n15962));
   NAND2xp33_ASAP7_75t_L U18930 (.Y(n15966),
	.A(n15965),
	.B(n15964));
   NOR2xp33_ASAP7_75t_R U18931 (.Y(n15965),
	.A(n15963),
	.B(n15962));
   NAND2xp33_ASAP7_75t_L U18932 (.Y(n15982),
	.A(n15977),
	.B(n15979));
   NOR2xp33_ASAP7_75t_SRAM U18933 (.Y(n15977),
	.A(FE_OFN26131_n15376),
	.B(n15978));
   NAND2xp33_ASAP7_75t_L U18934 (.Y(n15981),
	.A(n15980),
	.B(n15979));
   NOR2xp33_ASAP7_75t_SRAM U18935 (.Y(n15980),
	.A(n16009),
	.B(n15978));
   NAND2xp33_ASAP7_75t_SRAM U18936 (.Y(n15990),
	.A(n15989),
	.B(n15988));
   OAI22xp33_ASAP7_75t_SRAM U18937 (.Y(n16024),
	.A1(FE_OFN25985_n15997),
	.A2(n15996),
	.B1(FE_OFN25920_n15995),
	.B2(n15996));
   NAND2xp33_ASAP7_75t_SL U18938 (.Y(n16022),
	.A(n16008),
	.B(n16007));
   NOR2xp33_ASAP7_75t_L U18940 (.Y(n24768),
	.A(FE_OFN16248_n20235),
	.B(n24769));
   NAND2xp33_ASAP7_75t_L U18941 (.Y(n24772),
	.A(n24771),
	.B(n24770));
   NAND2xp33_ASAP7_75t_R U18942 (.Y(n25059),
	.A(n25056),
	.B(n25057));
   NAND2xp33_ASAP7_75t_R U18943 (.Y(n25058),
	.A(FE_OFN25950_sa01_2),
	.B(n25057));
   NOR2xp33_ASAP7_75t_SRAM U18944 (.Y(n24255),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(n24256));
   NAND2xp33_ASAP7_75t_L U18946 (.Y(n24188),
	.A(n24183),
	.B(n24185));
   NAND2xp5_ASAP7_75t_SL U18947 (.Y(n24971),
	.A(n24970),
	.B(FE_OFN59_sa10_7));
   NOR2x1_ASAP7_75t_SL U18948 (.Y(n24970),
	.A(n24969),
	.B(sa10_6_));
   NAND2xp5_ASAP7_75t_L U18949 (.Y(n24972),
	.A(n24968),
	.B(FE_OFN59_sa10_7));
   NOR2xp33_ASAP7_75t_L U18950 (.Y(n24968),
	.A(n24967),
	.B(sa10_6_));
   NAND2xp33_ASAP7_75t_SRAM U18951 (.Y(n24966),
	.A(n24963),
	.B(n24962));
   NAND2xp33_ASAP7_75t_R U18952 (.Y(n24962),
	.A(n24961),
	.B(n24960));
   NOR2x1_ASAP7_75t_L U18953 (.Y(n19217),
	.A(n17473),
	.B(n23255));
   NOR2xp33_ASAP7_75t_SRAM U18954 (.Y(n19996),
	.A(FE_OFN29023_n16750),
	.B(n25581));
   NAND2xp67_ASAP7_75t_SL U18955 (.Y(n16777),
	.A(n16763),
	.B(FE_OFN62_sa21_3));
   NAND2xp5_ASAP7_75t_L U18956 (.Y(n19554),
	.A(n20561),
	.B(n19552));
   NOR2xp33_ASAP7_75t_L U18957 (.Y(n19553),
	.A(FE_OFN28834_FE_OCPN28371_n17900),
	.B(n19554));
   NOR2xp33_ASAP7_75t_L U18959 (.Y(n19528),
	.A(n23603),
	.B(n24055));
   NOR2x1_ASAP7_75t_SL U18961 (.Y(n20754),
	.A(n23336),
	.B(n23161));
   OA21x2_ASAP7_75t_SL U18962 (.Y(n20755),
	.A1(n20753),
	.A2(n21785),
	.B(n21127));
   NOR2xp33_ASAP7_75t_L U18963 (.Y(n17864),
	.A(FE_OFN28779_n24257),
	.B(n22330));
   NOR2xp33_ASAP7_75t_L U18964 (.Y(n17865),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(n22330));
   NOR2xp33_ASAP7_75t_SL U18967 (.Y(n18553),
	.A(FE_OCPN27715_n23875),
	.B(FE_OCPN27532_n21643));
   INVxp33_ASAP7_75t_L U18970 (.Y(n17792),
	.A(n22560));
   NOR2xp33_ASAP7_75t_L U18973 (.Y(n17288),
	.A(n17245),
	.B(n21455));
   NOR2xp33_ASAP7_75t_L U18974 (.Y(n17290),
	.A(FE_OCPN29295_n18739),
	.B(n21455));
   NOR2x1_ASAP7_75t_SL U18975 (.Y(n17283),
	.A(n17301),
	.B(n19594));
   NOR2x1p5_ASAP7_75t_SL U18977 (.Y(n17274),
	.A(FE_OCPN29291_n17282),
	.B(n18767));
   NOR2xp33_ASAP7_75t_SL U18978 (.Y(n17260),
	.A(n18656),
	.B(n26099));
   INVxp67_ASAP7_75t_L U18979 (.Y(n17278),
	.A(n17276));
   AND3x1_ASAP7_75t_SL U18980 (.Y(n17809),
	.A(n17807),
	.B(n17806),
	.C(n20172));
   NAND2xp5_ASAP7_75t_SL U18981 (.Y(n17806),
	.A(n17805),
	.B(n17804));
   NAND2xp5_ASAP7_75t_SL U18982 (.Y(n17804),
	.A(n17803),
	.B(n17802));
   NAND2xp33_ASAP7_75t_SL U18983 (.Y(n17805),
	.A(n17801),
	.B(n17802));
   NAND2xp5_ASAP7_75t_R U18984 (.Y(n17790),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(FE_OCPN27273_sa02_3));
   NAND2x1p5_ASAP7_75t_SL U18985 (.Y(n17791),
	.A(n17799),
	.B(FE_OCPN27330_n));
   NOR2xp33_ASAP7_75t_SL U18988 (.Y(n17798),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(n26970));
   NOR2xp33_ASAP7_75t_SL U18989 (.Y(n20964),
	.A(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(n20965));
   NAND3xp33_ASAP7_75t_SL U18990 (.Y(n22088),
	.A(n20137),
	.B(n20954),
	.C(n19271));
   NOR2xp33_ASAP7_75t_SL U18991 (.Y(n19271),
	.A(n20978),
	.B(n25530));
   AND3x1_ASAP7_75t_L U18992 (.Y(n22090),
	.A(n22086),
	.B(n22085),
	.C(n22084));
   NOR2x1_ASAP7_75t_L U18993 (.Y(n17808),
	.A(FE_OCPN28158_n),
	.B(n17790));
   INVxp67_ASAP7_75t_R U18994 (.Y(n19264),
	.A(n22527));
   NAND2xp33_ASAP7_75t_L U18995 (.Y(n17145),
	.A(n16978),
	.B(n17001));
   NAND2xp5_ASAP7_75t_L U18996 (.Y(n18932),
	.A(FE_OFN27186_sa13_4),
	.B(FE_OFN16268_sa13_3));
   NAND2xp5_ASAP7_75t_SL U18997 (.Y(n17074),
	.A(n17073),
	.B(n17072));
   NAND2xp5_ASAP7_75t_L U18998 (.Y(n17072),
	.A(n17071),
	.B(n17070));
   NAND2xp5_ASAP7_75t_L U18999 (.Y(n17073),
	.A(n17069),
	.B(n17070));
   NOR2xp33_ASAP7_75t_R U19000 (.Y(n17071),
	.A(FE_OFN28801_n16978),
	.B(n20513));
   NOR2x1_ASAP7_75t_SL U19001 (.Y(n17132),
	.A(n19435),
	.B(n19409));
   NOR2x1_ASAP7_75t_L U19002 (.Y(n18900),
	.A(FE_OCPN29327_n21017),
	.B(n21729));
   NOR2xp33_ASAP7_75t_L U19005 (.Y(n16557),
	.A(n16542),
	.B(n24726));
   NOR2xp33_ASAP7_75t_L U19006 (.Y(n16559),
	.A(n24944),
	.B(n24726));
   NAND2xp33_ASAP7_75t_SL U19008 (.Y(n16587),
	.A(n16583),
	.B(n16584));
   NOR2xp33_ASAP7_75t_L U19009 (.Y(n16583),
	.A(FE_OFN28807_n24944),
	.B(n19663));
   NOR2x1_ASAP7_75t_SL U19010 (.Y(n16547),
	.A(FE_OFN28722_sa10_3),
	.B(FE_OFN25959_n23011));
   NOR3x1_ASAP7_75t_L U19011 (.Y(n17223),
	.A(FE_OFN26039_sa10_2),
	.B(FE_OFN142_sa10_0),
	.C(FE_OFN29042_n));
   NOR3xp33_ASAP7_75t_SL U19013 (.Y(n16569),
	.A(n16568),
	.B(n24734),
	.C(n16567));
   NOR2xp33_ASAP7_75t_R U19014 (.Y(n19144),
	.A(FE_OFN26651_n19573),
	.B(FE_OCPN29260_sa00_5));
   NOR2x1_ASAP7_75t_L U19015 (.Y(n18388),
	.A(n24791),
	.B(n22139));
   NAND3xp33_ASAP7_75t_SL U19016 (.Y(n18765),
	.A(FE_OCPN29542_n21151),
	.B(n21445),
	.C(FE_OCPN29463_n));
   NAND2xp5_ASAP7_75t_R U19017 (.Y(n18740),
	.A(FE_PSN8285_FE_OCPN29463_n),
	.B(FE_OCPN29295_n18739));
   NAND2x1_ASAP7_75t_SL U19018 (.Y(n21856),
	.A(FE_OFN29061_n22505),
	.B(FE_OCPN29513_n17447));
   NOR2xp33_ASAP7_75t_R U19020 (.Y(n21418),
	.A(FE_OCPN29513_n17447),
	.B(FE_OCPN28082_n21860));
   NAND2xp5_ASAP7_75t_SL U19021 (.Y(n21420),
	.A(n21416),
	.B(FE_OFN16351_n26084));
   NOR2xp33_ASAP7_75t_R U19022 (.Y(n21416),
	.A(n19162),
	.B(FE_OCPN28082_n21860));
   NAND2xp5_ASAP7_75t_L U19025 (.Y(n23390),
	.A(n19162),
	.B(n22489));
   INVx1_ASAP7_75t_R U19027 (.Y(n21394),
	.A(FE_PSN8303_n19222));
   NOR3x1_ASAP7_75t_R U19028 (.Y(n18362),
	.A(FE_OCPN27966_n18473),
	.B(FE_OFN28895_sa30_2),
	.C(n19051));
   NOR2xp33_ASAP7_75t_R U19029 (.Y(n18374),
	.A(FE_OFN25917_n21591),
	.B(n21608));
   NOR2xp33_ASAP7_75t_R U19030 (.Y(n18376),
	.A(FE_OFN28818_n17602),
	.B(n21608));
   NOR2x1_ASAP7_75t_SL U19031 (.Y(n18524),
	.A(FE_OFN29150_sa20_5),
	.B(n20636));
   NOR2xp33_ASAP7_75t_R U19032 (.Y(n21098),
	.A(n23336),
	.B(n23323));
   NOR2xp33_ASAP7_75t_SRAM U19034 (.Y(n20762),
	.A(n22828),
	.B(n21122));
   NAND2xp33_ASAP7_75t_L U19035 (.Y(n22318),
	.A(FE_OFN26141_n23307),
	.B(FE_OCPN29557_n18161));
   NOR2xp33_ASAP7_75t_SL U19037 (.Y(n20726),
	.A(n21772),
	.B(n23303));
   NAND2x1p5_ASAP7_75t_SL U19038 (.Y(n18217),
	.A(n22311),
	.B(n21105));
   NOR2x1_ASAP7_75t_SL U19040 (.Y(n18208),
	.A(n22290),
	.B(n22859));
   NAND2xp5_ASAP7_75t_SL U19041 (.Y(n21798),
	.A(n21127),
	.B(n21133));
   NOR2xp33_ASAP7_75t_SL U19042 (.Y(n18219),
	.A(FE_OFN26141_n23307),
	.B(n21122));
   NAND2xp5_ASAP7_75t_L U19044 (.Y(n18213),
	.A(FE_PSN8315_FE_OFN16135_sa22_4),
	.B(n23300));
   NAND2xp5_ASAP7_75t_SL U19045 (.Y(n21127),
	.A(n18161),
	.B(n23322));
   NOR2x1_ASAP7_75t_SL U19046 (.Y(n22811),
	.A(FE_OCPN29305_n23302),
	.B(FE_OFN25987_n23322));
   NOR2x1p5_ASAP7_75t_SL U19048 (.Y(n21224),
	.A(n18551),
	.B(n18561));
   NOR2xp33_ASAP7_75t_SL U19049 (.Y(n21219),
	.A(FE_OFN16295_n23837),
	.B(n21217));
   OAI21xp33_ASAP7_75t_L U19050 (.Y(n21215),
	.A1(n23711),
	.A2(n18530),
	.B(n23694));
   NOR2xp33_ASAP7_75t_SL U19051 (.Y(n18591),
	.A(n20685),
	.B(n23879));
   NAND2xp5_ASAP7_75t_L U19052 (.Y(n18593),
	.A(n18589),
	.B(n18590));
   NOR2xp33_ASAP7_75t_SL U19053 (.Y(n18589),
	.A(FE_OFN28988_n18597),
	.B(n23879));
   NOR2xp33_ASAP7_75t_L U19054 (.Y(n21675),
	.A(n20617),
	.B(n21676));
   NOR2xp33_ASAP7_75t_L U19055 (.Y(n21678),
	.A(n18583),
	.B(n21676));
   NAND2xp33_ASAP7_75t_L U19056 (.Y(n20689),
	.A(n20686),
	.B(n18570));
   NOR3xp33_ASAP7_75t_SL U19057 (.Y(n20666),
	.A(n18552),
	.B(n23840),
	.C(n21682));
   OAI21xp33_ASAP7_75t_L U19058 (.Y(n18552),
	.A1(FE_OFN29131_FE_OCPN27371_sa20_2),
	.A2(n21240),
	.B(n21234));
   NAND2xp5_ASAP7_75t_SL U19060 (.Y(n16457),
	.A(n16689),
	.B(FE_OFN27062_n16438));
   NAND2xp5_ASAP7_75t_L U19061 (.Y(n16684),
	.A(n16834),
	.B(n24614));
   NOR2x1p5_ASAP7_75t_L U19062 (.Y(n16689),
	.A(FE_OFN28694_sa33_4),
	.B(FE_OFN26628_n));
   OA21x2_ASAP7_75t_SL U19063 (.Y(n19309),
	.A1(FE_OCPN28266_n20920),
	.A2(n22979),
	.B(n19308));
   NOR2xp33_ASAP7_75t_L U19064 (.Y(n19310),
	.A(n19019),
	.B(n22048));
   NOR2x1_ASAP7_75t_L U19065 (.Y(n22997),
	.A(n20241),
	.B(FE_OCPN27954_n22945));
   OAI22xp33_ASAP7_75t_SL U19066 (.Y(n21564),
	.A1(n17321),
	.A2(n21563),
	.B1(FE_OCPN8219_n22197),
	.B2(n21563));
   NAND2xp33_ASAP7_75t_SRAM U19067 (.Y(n21565),
	.A(n21562),
	.B(n17321));
   INVxp33_ASAP7_75t_SRAM U19068 (.Y(n21562),
	.A(n21561));
   NOR3xp33_ASAP7_75t_SL U19070 (.Y(n21563),
	.A(n17345),
	.B(FE_OCPN27423_sa01_0),
	.C(n22598));
   NOR3xp33_ASAP7_75t_L U19072 (.Y(n22603),
	.A(n17345),
	.B(FE_OCPN27423_sa01_0),
	.C(n17318));
   NOR2x1_ASAP7_75t_SL U19073 (.Y(n20368),
	.A(FE_OCPN28380_n22433),
	.B(n18726));
   NAND3xp33_ASAP7_75t_SL U19074 (.Y(n18713),
	.A(n17359),
	.B(FE_OFN29135_n21551),
	.C(FE_OCPN27423_sa01_0));
   AND2x2_ASAP7_75t_L U19075 (.Y(n19547),
	.A(n25398),
	.B(n23235));
   NAND2xp5_ASAP7_75t_L U19076 (.Y(n19550),
	.A(n20795),
	.B(n20814));
   NAND2xp33_ASAP7_75t_L U19077 (.Y(n19549),
	.A(n20545),
	.B(n19547));
   NOR2xp33_ASAP7_75t_R U19079 (.Y(n19523),
	.A(n24362),
	.B(n22718));
   NAND2x1_ASAP7_75t_SL U19080 (.Y(n17970),
	.A(n20593),
	.B(n23220));
   NAND2xp5_ASAP7_75t_SL U19081 (.Y(n22236),
	.A(FE_OFN25908_sa12_2),
	.B(n23206));
   NAND2xp5_ASAP7_75t_SL U19082 (.Y(n22222),
	.A(FE_OCPN29559_n17900),
	.B(n23587));
   NAND3xp33_ASAP7_75t_SL U19083 (.Y(n19503),
	.A(n22745),
	.B(n17906),
	.C(FE_OCPN29485_sa12_3));
   NOR2xp33_ASAP7_75t_L U19084 (.Y(n20545),
	.A(FE_OFN29075_n22745),
	.B(n23582));
   NOR2xp33_ASAP7_75t_L U19086 (.Y(n20546),
	.A(n19546),
	.B(n23582));
   NOR2x1_ASAP7_75t_L U19087 (.Y(n20571),
	.A(FE_OCPN28232_n17949),
	.B(n19502));
   NAND3xp33_ASAP7_75t_L U19088 (.Y(n17163),
	.A(n17162),
	.B(n17161),
	.C(n17160));
   NOR2xp33_ASAP7_75t_SRAM U19089 (.Y(n17167),
	.A(n16980),
	.B(n17165));
   NAND2xp5_ASAP7_75t_SL U19090 (.Y(n17535),
	.A(n17533),
	.B(n17532));
   NAND2xp5_ASAP7_75t_L U19091 (.Y(n17532),
	.A(n17531),
	.B(n17530));
   NAND3xp33_ASAP7_75t_SL U19093 (.Y(n19943),
	.A(FE_OCPN29449_n17521),
	.B(n17560),
	.C(FE_OCPN29420_FE_OFN16128_sa32_2));
   NOR2x1_ASAP7_75t_SL U19094 (.Y(n17581),
	.A(n19740),
	.B(n24869));
   NOR2xp33_ASAP7_75t_SRAM U19096 (.Y(n19731),
	.A(n17560),
	.B(n19732));
   NAND2x1p5_ASAP7_75t_L U19098 (.Y(n18836),
	.A(FE_OCPN29420_FE_OFN16128_sa32_2),
	.B(n17521));
   NOR3x1_ASAP7_75t_L U19100 (.Y(n20345),
	.A(n23633),
	.B(FE_OCPN29414_n),
	.C(n16801));
   NOR3xp33_ASAP7_75t_SL U19101 (.Y(n16789),
	.A(n16777),
	.B(FE_OCPN27328_sa21_2),
	.C(FE_OCPN27556_n17843));
   NAND2x1p5_ASAP7_75t_SL U19102 (.Y(n20344),
	.A(n25351),
	.B(n22661));
   NAND2x1_ASAP7_75t_L U19103 (.Y(n19872),
	.A(FE_OFN28779_n24257),
	.B(FE_OCPN27642_n16758));
   NOR2xp33_ASAP7_75t_SL U19104 (.Y(n22351),
	.A(n17882),
	.B(n19871));
   NAND2xp33_ASAP7_75t_SL U19106 (.Y(n20032),
	.A(n20026),
	.B(FE_OFN25972_n20056));
   NOR2xp33_ASAP7_75t_SL U19107 (.Y(n20026),
	.A(n20841),
	.B(n20027));
   NOR2xp33_ASAP7_75t_SRAM U19108 (.Y(n20879),
	.A(n21989),
	.B(n21922));
   NAND2xp33_ASAP7_75t_SL U19109 (.Y(n20881),
	.A(n20877),
	.B(n20878));
   NOR2xp33_ASAP7_75t_R U19110 (.Y(n20877),
	.A(FE_OCPN27516_n26292),
	.B(n21922));
   NOR3xp33_ASAP7_75t_SL U19111 (.Y(n16490),
	.A(n21981),
	.B(FE_OCPN29482_FE_OFN26014_sa31_3),
	.C(n16340));
   NOR3xp33_ASAP7_75t_L U19112 (.Y(n16345),
	.A(n16321),
	.B(FE_OFN28669_sa31_5),
	.C(n16329));
   NOR2x1_ASAP7_75t_SL U19113 (.Y(n20033),
	.A(n20074),
	.B(FE_OCPN7597_n21981));
   NOR2xp33_ASAP7_75t_SL U19117 (.Y(n16516),
	.A(FE_OFN29047_n21980),
	.B(FE_OCPN28334_n16497));
   NAND2xp5_ASAP7_75t_SL U19118 (.Y(n16374),
	.A(n18068),
	.B(n16326));
   NAND3xp33_ASAP7_75t_L U19119 (.Y(n16502),
	.A(n20868),
	.B(n16300),
	.C(FE_OCPN29526_sa31_4));
   NOR2xp33_ASAP7_75t_SL U19120 (.Y(n18308),
	.A(n17679),
	.B(n18827));
   NOR2xp33_ASAP7_75t_SL U19122 (.Y(n17045),
	.A(FE_OCPN5143_n19361),
	.B(FE_OFN28738_n16989));
   NOR2x1_ASAP7_75t_L U19123 (.Y(n19871),
	.A(FE_OCPN5082_n22663),
	.B(n23633));
   NOR2x1_ASAP7_75t_L U19125 (.Y(n20028),
	.A(FE_OFN29147_sa31_1),
	.B(FE_OFN28492_sa31_0));
   NOR2xp33_ASAP7_75t_L U19126 (.Y(n20053),
	.A(n21922),
	.B(n20027));
   NAND3xp33_ASAP7_75t_R U19127 (.Y(n16922),
	.A(FE_OFN29164_sa33_2),
	.B(FE_OCPN27555_n16422),
	.C(n16427));
   NOR2xp33_ASAP7_75t_R U19128 (.Y(n16838),
	.A(FE_OCPN29487_FE_OFN28694_sa33_4),
	.B(n16851));
   NAND2x1p5_ASAP7_75t_SL U19129 (.Y(n16894),
	.A(n16464),
	.B(n16463));
   NAND2x1_ASAP7_75t_L U19130 (.Y(n16463),
	.A(n16462),
	.B(n16461));
   NOR2xp67_ASAP7_75t_L U19131 (.Y(n16462),
	.A(FE_OFN29101_n16418),
	.B(n24613));
   NAND2xp33_ASAP7_75t_L U19132 (.Y(n14057),
	.A(n14052),
	.B(n14054));
   NOR2xp33_ASAP7_75t_SRAM U19133 (.Y(n14052),
	.A(n12994),
	.B(n14053));
   NAND2xp33_ASAP7_75t_L U19134 (.Y(n14056),
	.A(n14055),
	.B(n14054));
   NOR2xp33_ASAP7_75t_L U19135 (.Y(n14055),
	.A(n15349),
	.B(n14053));
   NAND2xp33_ASAP7_75t_SL U19136 (.Y(n14051),
	.A(n14046),
	.B(n14048));
   NOR2xp33_ASAP7_75t_L U19137 (.Y(n14046),
	.A(n15729),
	.B(n14047));
   NAND2xp33_ASAP7_75t_SL U19138 (.Y(n14050),
	.A(n14049),
	.B(n14048));
   NOR2xp33_ASAP7_75t_L U19139 (.Y(n14049),
	.A(FE_OFN28769_n15478),
	.B(n14047));
   NOR3xp33_ASAP7_75t_L U19140 (.Y(n14041),
	.A(n13870),
	.B(n14377),
	.C(n15541));
   NAND2xp33_ASAP7_75t_R U19141 (.Y(n14067),
	.A(n14063),
	.B(n14064));
   NOR2xp33_ASAP7_75t_R U19142 (.Y(n14063),
	.A(n15487),
	.B(n14250));
   NAND2xp33_ASAP7_75t_R U19143 (.Y(n14066),
	.A(n14065),
	.B(n14064));
   NOR2xp33_ASAP7_75t_R U19144 (.Y(n14065),
	.A(FE_OFN27066_n13869),
	.B(n14250));
   NAND2xp33_ASAP7_75t_SL U19145 (.Y(n14072),
	.A(n14070),
	.B(n14069));
   NOR2xp33_ASAP7_75t_L U19146 (.Y(n14070),
	.A(FE_OCPN29329_n15517),
	.B(n15749));
   NAND2xp5_ASAP7_75t_L U19147 (.Y(n14071),
	.A(n15748),
	.B(n14069));
   NOR2xp33_ASAP7_75t_SRAM U19148 (.Y(n14074),
	.A(n15536),
	.B(FE_OFN16210_n13876));
   NOR2xp33_ASAP7_75t_SRAM U19149 (.Y(n14073),
	.A(FE_OFN27074_n13868),
	.B(n15719));
   NOR2xp33_ASAP7_75t_SRAM U19150 (.Y(n14016),
	.A(n15484),
	.B(n15347));
   NOR2xp33_ASAP7_75t_L U19151 (.Y(n14774),
	.A(FE_OFN28_w3_23),
	.B(FE_OFN25909_w3_20));
   NAND2xp5_ASAP7_75t_L U19152 (.Y(n14532),
	.A(n14531),
	.B(FE_OFN25880_w3_24));
   NAND2xp5_ASAP7_75t_L U19153 (.Y(n14533),
	.A(n14513),
	.B(FE_OFN25880_w3_24));
   NOR2xp33_ASAP7_75t_L U19154 (.Y(n14531),
	.A(n14530),
	.B(FE_OFN16412_w3_26));
   NOR2xp33_ASAP7_75t_L U19155 (.Y(n14591),
	.A(n15158),
	.B(n14595));
   INVx1_ASAP7_75t_SL U19156 (.Y(n14597),
	.A(n14590));
   NAND2xp33_ASAP7_75t_L U19157 (.Y(n14589),
	.A(n14543),
	.B(n14542));
   NAND2xp33_ASAP7_75t_L U19158 (.Y(n14588),
	.A(n14555),
	.B(n14554));
   NOR2xp33_ASAP7_75t_SRAM U19159 (.Y(n14492),
	.A(n14498),
	.B(n14474));
   NOR3xp33_ASAP7_75t_SRAM U19160 (.Y(n14474),
	.A(FE_OFN16451_n),
	.B(FE_OFN27208_w3_30),
	.C(FE_OFN28890_n));
   OA21x2_ASAP7_75t_R U19161 (.Y(n14494),
	.A1(n14491),
	.A2(FE_OFN25893_n15214),
	.B(n14490));
   NAND2xp33_ASAP7_75t_L U19162 (.Y(n14490),
	.A(n14489),
	.B(n14488));
   NAND2xp33_ASAP7_75t_R U19163 (.Y(n14488),
	.A(n14487),
	.B(n14486));
   NAND2xp33_ASAP7_75t_L U19164 (.Y(n14489),
	.A(n14483),
	.B(n14486));
   NOR2xp33_ASAP7_75t_L U19165 (.Y(n14216),
	.A(n14214),
	.B(n14213));
   NOR2xp67_ASAP7_75t_SL U19167 (.Y(n14211),
	.A(n15782),
	.B(FE_OFN26084_n15106));
   NOR2xp33_ASAP7_75t_L U19168 (.Y(n14212),
	.A(n15792),
	.B(n14213));
   NOR2xp33_ASAP7_75t_SL U19169 (.Y(n14225),
	.A(n15856),
	.B(n14223));
   OA21x2_ASAP7_75t_R U19170 (.Y(n14224),
	.A1(n15814),
	.A2(n15808),
	.B(n14221));
   NAND2xp5_ASAP7_75t_R U19171 (.Y(n14235),
	.A(n14230),
	.B(n14232));
   NOR2xp33_ASAP7_75t_SRAM U19172 (.Y(n14230),
	.A(n14410),
	.B(n14231));
   NAND2xp5_ASAP7_75t_R U19173 (.Y(n14234),
	.A(n14233),
	.B(n14232));
   NOR2xp33_ASAP7_75t_SRAM U19174 (.Y(n14233),
	.A(n15779),
	.B(n14231));
   NAND2xp33_ASAP7_75t_SL U19175 (.Y(n14227),
	.A(n14222),
	.B(n14224));
   NOR2xp33_ASAP7_75t_L U19176 (.Y(n14222),
	.A(n15838),
	.B(n14223));
   INVx1_ASAP7_75t_L U19177 (.Y(n14210),
	.A(n15020));
   NOR3xp33_ASAP7_75t_SRAM U19178 (.Y(n14197),
	.A(FE_OFN25928_n15779),
	.B(FE_OFN28747_n),
	.C(FE_OFN16195_n13771));
   NOR2xp33_ASAP7_75t_SRAM U19180 (.Y(n13819),
	.A(n14116),
	.B(n13820));
   NAND2xp33_ASAP7_75t_SL U19181 (.Y(n13818),
	.A(n13817),
	.B(FE_OFN25920_n15995));
   NOR3xp33_ASAP7_75t_SRAM U19182 (.Y(n13817),
	.A(FE_OCPN29570_n15423),
	.B(n14941),
	.C(FE_OFN27200_n));
   OAI21xp33_ASAP7_75t_R U19183 (.Y(n13842),
	.A1(n15973),
	.A2(FE_OFN28898_n13805),
	.B(n13841));
   OAI21xp33_ASAP7_75t_SRAM U19184 (.Y(n13841),
	.A1(FE_OFN26641_w3_14),
	.A2(FE_OFN28813_n15414),
	.B(n15934));
   NAND2xp33_ASAP7_75t_L U19185 (.Y(n13850),
	.A(n13846),
	.B(n13847));
   NOR2xp33_ASAP7_75t_R U19186 (.Y(n13846),
	.A(n13843),
	.B(n14610));
   NAND2xp33_ASAP7_75t_R U19187 (.Y(n13849),
	.A(n13848),
	.B(n13847));
   INVxp33_ASAP7_75t_SRAM U19188 (.Y(n13848),
	.A(n15446));
   NOR2xp33_ASAP7_75t_SRAM U19189 (.Y(n13829),
	.A(n15451),
	.B(n14712));
   NOR2xp33_ASAP7_75t_SRAM U19190 (.Y(n13831),
	.A(n13830),
	.B(n14712));
   NAND2xp33_ASAP7_75t_SRAM U19191 (.Y(n13830),
	.A(n15999),
	.B(n14159));
   OAI21xp33_ASAP7_75t_L U19192 (.Y(n14362),
	.A1(FE_OFN26614_n),
	.A2(n14760),
	.B(n14357));
   NOR2xp33_ASAP7_75t_SRAM U19193 (.Y(n14360),
	.A(n12994),
	.B(n14362));
   OA21x2_ASAP7_75t_SRAM U19194 (.Y(n14363),
	.A1(FE_OCPN29329_n15517),
	.A2(n13875),
	.B(n14359));
   O2A1O1Ixp33_ASAP7_75t_SL U19195 (.Y(n14359),
	.A1(FE_OFN6_w3_22),
	.A2(n15694),
	.B(n15729),
	.C(n14358));
   NOR2xp33_ASAP7_75t_SL U19196 (.Y(n14358),
	.A(FE_OFN28683_w3_21),
	.B(n14749));
   NAND2xp33_ASAP7_75t_L U19197 (.Y(n14368),
	.A(FE_OFN27082_n25377),
	.B(n15339));
   NAND2xp5_ASAP7_75t_L U19198 (.Y(n14367),
	.A(FE_OFN6_w3_22),
	.B(n15479));
   OAI222xp33_ASAP7_75t_L U19199 (.Y(n14381),
	.A1(n15528),
	.A2(n14380),
	.B1(n15694),
	.B2(n14380),
	.C1(FE_OFN28551_FE_OFN26114_n),
	.C2(n14380));
   NAND2xp5_ASAP7_75t_L U19200 (.Y(n14379),
	.A(n15680),
	.B(FE_OFN25981_n13868));
   NAND2xp33_ASAP7_75t_L U19201 (.Y(n14378),
	.A(n14377),
	.B(FE_OFN25981_n13868));
   NOR3xp33_ASAP7_75t_L U19202 (.Y(n14382),
	.A(n14376),
	.B(n14375),
	.C(n14374));
   NAND2xp33_ASAP7_75t_L U19203 (.Y(n14374),
	.A(n14373),
	.B(n14372));
   OAI21xp33_ASAP7_75t_SL U19204 (.Y(n14376),
	.A1(n14748),
	.A2(FE_OCPN8264_n13890),
	.B(n14370));
   NOR2xp33_ASAP7_75t_R U19205 (.Y(n14384),
	.A(FE_OFN28977_n),
	.B(FE_OCPN28278_n15512));
   OA21x2_ASAP7_75t_L U19206 (.Y(n14337),
	.A1(FE_OFN27151_n),
	.A2(FE_OFN16210_n13876),
	.B(n14335));
   O2A1O1Ixp33_ASAP7_75t_SRAM U19207 (.Y(n14335),
	.A1(FE_OFN27151_n),
	.A2(n13874),
	.B(n12994),
	.C(n15333));
   NOR2xp33_ASAP7_75t_R U19208 (.Y(n14336),
	.A(n14334),
	.B(n14333));
   O2A1O1Ixp33_ASAP7_75t_SRAM U19209 (.Y(n14333),
	.A1(FE_OFN27151_n),
	.A2(n15694),
	.B(n15484),
	.C(FE_OFN16352_n14289));
   OAI21xp5_ASAP7_75t_L U19210 (.Y(n15283),
	.A1(FE_OFN26539_w3_19),
	.A2(FE_OFN26091_n24663),
	.B(n14068));
   NAND2xp5_ASAP7_75t_SL U19211 (.Y(n15250),
	.A(n15244),
	.B(n15247));
   NAND2xp33_ASAP7_75t_SL U19212 (.Y(n15261),
	.A(n15213),
	.B(n15212));
   NAND2xp33_ASAP7_75t_R U19213 (.Y(n15213),
	.A(n15207),
	.B(n15210));
   NAND2xp33_ASAP7_75t_R U19214 (.Y(n15212),
	.A(n15211),
	.B(n15210));
   NAND2xp33_ASAP7_75t_R U19215 (.Y(n15260),
	.A(n15221),
	.B(n15220));
   NAND2xp33_ASAP7_75t_SRAM U19216 (.Y(n15221),
	.A(n15215),
	.B(n15218));
   NAND2xp33_ASAP7_75t_SRAM U19217 (.Y(n15220),
	.A(n15219),
	.B(n15218));
   NOR2xp33_ASAP7_75t_SRAM U19218 (.Y(n15215),
	.A(FE_OFN16437_n),
	.B(n15216));
   NAND2xp33_ASAP7_75t_SRAM U19219 (.Y(n15194),
	.A(n15193),
	.B(n15192));
   NAND2xp33_ASAP7_75t_R U19220 (.Y(n15193),
	.A(FE_OFN28929_n15182),
	.B(n15190));
   NAND2xp33_ASAP7_75t_R U19221 (.Y(n15192),
	.A(n15191),
	.B(n15190));
   NAND2xp5_ASAP7_75t_R U19222 (.Y(n15179),
	.A(FE_OFN25966_n13646),
	.B(FE_OFN28817_n));
   INVxp33_ASAP7_75t_SRAM U19223 (.Y(n15172),
	.A(n15168));
   NOR3xp33_ASAP7_75t_SRAM U19224 (.Y(n15791),
	.A(FE_OFN28889_n15845),
	.B(n15862),
	.C(n13741));
   NAND2xp33_ASAP7_75t_SL U19225 (.Y(n15869),
	.A(n15863),
	.B(n15866));
   NOR2xp33_ASAP7_75t_L U19226 (.Y(n15863),
	.A(n15859),
	.B(n15864));
   NAND2xp33_ASAP7_75t_L U19227 (.Y(n15868),
	.A(n15867),
	.B(n15866));
   NOR2xp33_ASAP7_75t_SL U19228 (.Y(n15867),
	.A(n15865),
	.B(n15864));
   NAND2xp33_ASAP7_75t_R U19229 (.Y(n15878),
	.A(n15874),
	.B(n15873));
   NOR2xp33_ASAP7_75t_R U19230 (.Y(n15874),
	.A(n15871),
	.B(n15875));
   NOR3xp33_ASAP7_75t_SRAM U19232 (.Y(n15816),
	.A(n15808),
	.B(FE_OFN16195_n13771),
	.C(n14996));
   OA21x2_ASAP7_75t_R U19233 (.Y(n15818),
	.A1(n15814),
	.A2(n15813),
	.B(n15812));
   OAI222xp33_ASAP7_75t_L U19234 (.Y(n15812),
	.A1(FE_OFN25897_w3_4),
	.A2(n15811),
	.B1(n15810),
	.B2(n15811),
	.C1(n15857),
	.C2(n15811));
   NOR2xp33_ASAP7_75t_L U19235 (.Y(n15828),
	.A(n15822),
	.B(n13730));
   NOR2xp33_ASAP7_75t_L U19237 (.Y(n14099),
	.A(n14913),
	.B(n14938));
   OAI21xp33_ASAP7_75t_R U19238 (.Y(n14805),
	.A1(FE_OCPN28404_n13874),
	.A2(FE_OCPN4685_n15658),
	.B(n14803));
   NAND2xp33_ASAP7_75t_SRAM U19239 (.Y(n14803),
	.A(FE_OCPN29578_FE_OFN27214_w3_17),
	.B(n15729));
   NAND2xp5_ASAP7_75t_SL U19240 (.Y(n14809),
	.A(n14802),
	.B(n14801));
   NAND2xp33_ASAP7_75t_SL U19241 (.Y(n14801),
	.A(n14800),
	.B(n14799));
   NAND2xp5_ASAP7_75t_SL U19242 (.Y(n14802),
	.A(n14796),
	.B(n14799));
   OA21x2_ASAP7_75t_SL U19243 (.Y(n14799),
	.A1(FE_OFN16210_n13876),
	.A2(n15709),
	.B(n15711));
   NAND3xp33_ASAP7_75t_SRAM U19244 (.Y(n14807),
	.A(n15694),
	.B(n15719),
	.C(n14806));
   NOR2xp33_ASAP7_75t_SL U19245 (.Y(n14792),
	.A(FE_OFN26538_w3_19),
	.B(n15660));
   NAND2xp5_ASAP7_75t_SL U19246 (.Y(n14749),
	.A(n14377),
	.B(FE_PSN8276_FE_OFN28712_n));
   NOR2xp33_ASAP7_75t_R U19247 (.Y(n14754),
	.A(n12994),
	.B(n14775));
   NAND2xp5_ASAP7_75t_SRAM U19249 (.Y(n15252),
	.A(n15205),
	.B(n15158));
   NOR2xp33_ASAP7_75t_R U19251 (.Y(n13303),
	.A(FE_OFN26059_n),
	.B(n15216));
   INVxp67_ASAP7_75t_L U19252 (.Y(n13309),
	.A(n13691));
   NAND3xp33_ASAP7_75t_SRAM U19253 (.Y(n13308),
	.A(FE_OFN28604_n14534),
	.B(n15257),
	.C(n13447));
   NOR2xp33_ASAP7_75t_R U19254 (.Y(n13317),
	.A(n25675),
	.B(n13318));
   INVx1_ASAP7_75t_L U19255 (.Y(n13320),
	.A(n13316));
   NAND2xp33_ASAP7_75t_SL U19256 (.Y(n13315),
	.A(n13314),
	.B(n13313));
   OR2x2_ASAP7_75t_SRAM U19257 (.Y(n13313),
	.A(n14572),
	.B(n13312));
   NOR2xp33_ASAP7_75t_SRAM U19258 (.Y(n14480),
	.A(FE_OFN27130_w3_28),
	.B(FE_OCPN29428_FE_OFN27131_w3_29));
   NOR2xp33_ASAP7_75t_R U19260 (.Y(n13296),
	.A(FE_OFN25875_n15227),
	.B(n13294));
   NOR2xp33_ASAP7_75t_SRAM U19261 (.Y(n13293),
	.A(n14498),
	.B(n13294));
   NAND2xp33_ASAP7_75t_SRAM U19263 (.Y(n13758),
	.A(n14423),
	.B(n13757));
   O2A1O1Ixp33_ASAP7_75t_SL U19264 (.Y(n13760),
	.A1(n15813),
	.A2(n15856),
	.B(n13750),
	.C(n15888));
   NAND2xp33_ASAP7_75t_SL U19265 (.Y(n13750),
	.A(n13749),
	.B(n13748));
   NAND2xp33_ASAP7_75t_L U19266 (.Y(n13749),
	.A(n13744),
	.B(n13746));
   NAND2xp33_ASAP7_75t_L U19267 (.Y(n13748),
	.A(n13747),
	.B(n13746));
   NOR2xp33_ASAP7_75t_R U19268 (.Y(n13780),
	.A(n25140),
	.B(n13778));
   NAND2xp33_ASAP7_75t_L U19269 (.Y(n13782),
	.A(n13777),
	.B(n13779));
   NOR2xp33_ASAP7_75t_L U19270 (.Y(n13777),
	.A(n14194),
	.B(n13778));
   NOR3xp33_ASAP7_75t_SRAM U19271 (.Y(n13784),
	.A(n15079),
	.B(FE_OFN28662_w3_7),
	.C(n13730));
   NOR2xp33_ASAP7_75t_L U19272 (.Y(n15858),
	.A(n15842),
	.B(n15808));
   NAND2xp33_ASAP7_75t_L U19274 (.Y(n13972),
	.A(n13968),
	.B(n13967));
   OA21x2_ASAP7_75t_R U19275 (.Y(n13953),
	.A1(FE_OFN109_n15994),
	.A2(n14615),
	.B(n13950));
   NAND2xp33_ASAP7_75t_SRAM U19276 (.Y(n13959),
	.A(n14140),
	.B(FE_OFN26624_n15376));
   NAND2xp33_ASAP7_75t_SRAM U19277 (.Y(n13958),
	.A(n15438),
	.B(FE_OFN26624_n15376));
   NOR2xp33_ASAP7_75t_SRAM U19278 (.Y(n13903),
	.A(n15713),
	.B(n13902));
   NAND2xp5_ASAP7_75t_L U19279 (.Y(n14798),
	.A(FE_PSN8334_n15539),
	.B(n15714));
   NAND2xp5_ASAP7_75t_R U19280 (.Y(n13911),
	.A(n13910),
	.B(n13909));
   NOR2xp33_ASAP7_75t_R U19281 (.Y(n13910),
	.A(FE_OFN27066_n13869),
	.B(n14315));
   OR2x2_ASAP7_75t_L U19282 (.Y(n13909),
	.A(FE_OCPN29329_n15517),
	.B(FE_OFN16352_n14289));
   NAND2xp33_ASAP7_75t_L U19283 (.Y(n13907),
	.A(n13905),
	.B(n14048));
   NOR2xp33_ASAP7_75t_L U19284 (.Y(n13905),
	.A(n14025),
	.B(n14271));
   NAND2xp33_ASAP7_75t_L U19285 (.Y(n13906),
	.A(FE_OFN25915_n15514),
	.B(n14048));
   NAND3xp33_ASAP7_75t_L U19286 (.Y(n15296),
	.A(FE_OFN16426_w3_20),
	.B(n14766),
	.C(FE_OFN28628_n15667));
   NOR2xp33_ASAP7_75t_SRAM U19287 (.Y(n13897),
	.A(n15660),
	.B(n13875));
   OAI21xp33_ASAP7_75t_L U19288 (.Y(n15747),
	.A1(n14068),
	.A2(n13875),
	.B(n13877));
   NAND2xp5_ASAP7_75t_L U19289 (.Y(n13877),
	.A(FE_OFN28976_n),
	.B(n14314));
   O2A1O1Ixp5_ASAP7_75t_SRAM U19291 (.Y(n13591),
	.A1(FE_OFN28456_n13348),
	.A2(FE_OFN28530_n14593),
	.B(n15171),
	.C(n13590));
   NAND2xp33_ASAP7_75t_L U19292 (.Y(n13592),
	.A(n13587),
	.B(n13586));
   OAI222xp33_ASAP7_75t_R U19293 (.Y(n13619),
	.A1(n13595),
	.A2(n13594),
	.B1(n15181),
	.B2(n13594),
	.C1(FE_OFN16206_n15240),
	.C2(n13594));
   NAND2xp5_ASAP7_75t_SL U19294 (.Y(n13618),
	.A(n13617),
	.B(n13616));
   NOR3xp33_ASAP7_75t_L U19295 (.Y(n13594),
	.A(FE_OFN28453_n13348),
	.B(n15235),
	.C(n15259));
   NAND2xp33_ASAP7_75t_SRAM U19297 (.Y(n13567),
	.A(FE_OFN26567_n),
	.B(FE_OCPN27665_w3_25));
   NOR3xp33_ASAP7_75t_SL U19298 (.Y(n13566),
	.A(n14504),
	.B(FE_OFN26112_n13288),
	.C(FE_OFN27207_w3_30));
   OA21x2_ASAP7_75t_SRAM U19299 (.Y(n13559),
	.A1(FE_OFN27057_n13662),
	.A2(n15199),
	.B(n13557));
   NAND2xp33_ASAP7_75t_L U19300 (.Y(n14854),
	.A(n14882),
	.B(n14890));
   NAND2xp5_ASAP7_75t_L U19301 (.Y(n14880),
	.A(n14860),
	.B(n14859));
   OR2x2_ASAP7_75t_L U19302 (.Y(n14860),
	.A(n14856),
	.B(n15045));
   NAND2xp5_ASAP7_75t_L U19303 (.Y(n14859),
	.A(n14858),
	.B(n14857));
   NOR2xp33_ASAP7_75t_L U19304 (.Y(n14882),
	.A(FE_OFN28831_n15838),
	.B(n14851));
   NOR2xp33_ASAP7_75t_L U19305 (.Y(n14851),
	.A(n15865),
	.B(FE_OFN28792_n15787));
   NAND2xp33_ASAP7_75t_SRAM U19306 (.Y(n14830),
	.A(n15033),
	.B(FE_OFN16269_n15808));
   NAND2xp33_ASAP7_75t_L U19307 (.Y(n14829),
	.A(n15107),
	.B(FE_OFN16269_n15808));
   NOR2xp67_ASAP7_75t_L U19308 (.Y(n15811),
	.A(n14986),
	.B(FE_OFN25928_n15779));
   NAND2xp5_ASAP7_75t_R U19309 (.Y(n14629),
	.A(n14939),
	.B(n15983));
   OAI21xp33_ASAP7_75t_L U19310 (.Y(n15998),
	.A1(FE_OFN29125_n),
	.A2(FE_OFN26638_w3_14),
	.B(n15422));
   NOR3xp33_ASAP7_75t_L U19311 (.Y(n14635),
	.A(n14634),
	.B(n24755),
	.C(n14913));
   OAI21xp33_ASAP7_75t_L U19312 (.Y(n14634),
	.A1(FE_OCPN29534_FE_OFN8_w3_14),
	.A2(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(n15948));
   NOR2xp33_ASAP7_75t_SL U19313 (.Y(n14632),
	.A(n14929),
	.B(FE_OFN109_n15994));
   NOR2xp33_ASAP7_75t_SL U19314 (.Y(n14647),
	.A(n15379),
	.B(n14646));
   NAND2xp33_ASAP7_75t_SRAM U19315 (.Y(n14642),
	.A(n15936),
	.B(n15959));
   A2O1A1Ixp33_ASAP7_75t_L U19316 (.Y(n14641),
	.A1(FE_OFN26642_w3_14),
	.A2(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(n15927),
	.C(n16032));
   NAND2xp33_ASAP7_75t_SL U19317 (.Y(n14649),
	.A(n14644),
	.B(n14643));
   NOR2xp33_ASAP7_75t_SL U19318 (.Y(n14644),
	.A(n15954),
	.B(n14646));
   OAI222xp33_ASAP7_75t_SRAM U19319 (.Y(n15351),
	.A1(FE_OFN5_w3_22),
	.A2(n15338),
	.B1(FE_OFN28706_n),
	.B2(n15338),
	.C1(FE_OFN26539_w3_19),
	.C2(n15338));
   NAND2xp33_ASAP7_75t_L U19320 (.Y(n15327),
	.A(n15322),
	.B(n15324));
   NOR2xp33_ASAP7_75t_R U19321 (.Y(n15322),
	.A(n15319),
	.B(n15323));
   NAND2xp33_ASAP7_75t_L U19322 (.Y(n15326),
	.A(n15325),
	.B(n15324));
   NOR2xp33_ASAP7_75t_R U19323 (.Y(n15325),
	.A(FE_OFN27066_n13869),
	.B(n15323));
   NAND2xp33_ASAP7_75t_L U19324 (.Y(n15337),
	.A(n15335),
	.B(n15334));
   NOR2xp33_ASAP7_75t_L U19325 (.Y(n15335),
	.A(n15333),
	.B(n15332));
   NAND2xp33_ASAP7_75t_L U19326 (.Y(n15332),
	.A(n15331),
	.B(n15330));
   NAND2xp33_ASAP7_75t_SRAM U19327 (.Y(n15336),
	.A(FE_OFN37_w3_23),
	.B(n15334));
   NAND2xp33_ASAP7_75t_R U19328 (.Y(n15306),
	.A(n15295),
	.B(n15294));
   NAND2xp33_ASAP7_75t_SRAM U19329 (.Y(n15295),
	.A(FE_OFN28769_n15478),
	.B(n15683));
   NAND2xp33_ASAP7_75t_SRAM U19330 (.Y(n15294),
	.A(n15536),
	.B(n15683));
   OAI22xp33_ASAP7_75t_SRAM U19331 (.Y(n13390),
	.A1(FE_OFN26049_w3_27),
	.A2(n15155),
	.B1(FE_OCPN27665_w3_25),
	.B2(n15155));
   NAND2xp33_ASAP7_75t_SL U19332 (.Y(n13389),
	.A(n13388),
	.B(n13387));
   NAND2xp33_ASAP7_75t_SL U19333 (.Y(n13387),
	.A(n13484),
	.B(n13386));
   INVxp67_ASAP7_75t_L U19334 (.Y(n15181),
	.A(n13499));
   NAND3xp33_ASAP7_75t_R U19335 (.Y(n13613),
	.A(FE_OFN26051_w3_27),
	.B(FE_OCPN27665_w3_25),
	.C(FE_OFN27210_w3_30));
   OA21x2_ASAP7_75t_SL U19336 (.Y(n13374),
	.A1(FE_OFN16225_n15195),
	.A2(n13421),
	.B(n13371));
   O2A1O1Ixp33_ASAP7_75t_SL U19337 (.Y(n13371),
	.A1(FE_OFN27057_n13662),
	.A2(n15171),
	.B(FE_OFN16206_n15240),
	.C(n13370));
   NOR3xp33_ASAP7_75t_SL U19338 (.Y(n13370),
	.A(n15203),
	.B(n14498),
	.C(FE_OFN26552_n14545));
   NOR2xp33_ASAP7_75t_R U19339 (.Y(n13375),
	.A(n13540),
	.B(n13373));
   NAND2xp33_ASAP7_75t_SL U19340 (.Y(n13377),
	.A(n13372),
	.B(n13374));
   NOR2xp33_ASAP7_75t_SRAM U19341 (.Y(n13372),
	.A(FE_OFN16437_n),
	.B(n13373));
   NAND2xp33_ASAP7_75t_SL U19343 (.Y(n13356),
	.A(n13355),
	.B(n13354));
   NAND2xp33_ASAP7_75t_SRAM U19344 (.Y(n13357),
	.A(FE_OFN25966_n13646),
	.B(n15217));
   NAND2xp33_ASAP7_75t_L U19345 (.Y(n13354),
	.A(n13353),
	.B(n13352));
   O2A1O1Ixp33_ASAP7_75t_L U19346 (.Y(n15009),
	.A1(n15589),
	.A2(n15888),
	.B(n15001),
	.C(FE_OFN25928_n15779));
   NAND2xp33_ASAP7_75t_SRAM U19347 (.Y(n15001),
	.A(FE_OCPN27985_n24831),
	.B(n15884));
   NOR2xp33_ASAP7_75t_SL U19348 (.Y(n15008),
	.A(n15619),
	.B(n15009));
   AND2x2_ASAP7_75t_L U19349 (.Y(n15011),
	.A(n15007),
	.B(n15006));
   NAND2xp33_ASAP7_75t_L U19350 (.Y(n15006),
	.A(n15005),
	.B(n15004));
   NAND2xp33_ASAP7_75t_L U19351 (.Y(n15007),
	.A(n15003),
	.B(n15004));
   NOR2xp33_ASAP7_75t_R U19352 (.Y(n15005),
	.A(FE_OFN25887_w3_3),
	.B(n15888));
   O2A1O1Ixp5_ASAP7_75t_SRAM U19353 (.Y(n15023),
	.A1(FE_OFN28661_w3_7),
	.A2(n15019),
	.B(n15625),
	.C(n13730));
   NOR2xp33_ASAP7_75t_R U19354 (.Y(n15022),
	.A(n15779),
	.B(n15023));
   NOR2xp33_ASAP7_75t_SL U19355 (.Y(n15440),
	.A(n15438),
	.B(n15437));
   NOR2xp33_ASAP7_75t_SL U19356 (.Y(n15436),
	.A(n16032),
	.B(n15437));
   NAND2xp5_ASAP7_75t_L U19357 (.Y(n15445),
	.A(FE_OFN26131_n15376),
	.B(n15983));
   O2A1O1Ixp33_ASAP7_75t_R U19358 (.Y(n15454),
	.A1(FE_OFN109_n15994),
	.A2(n15453),
	.B(n15452),
	.C(n16026));
   OAI21xp5_ASAP7_75t_L U19359 (.Y(n15402),
	.A1(FE_OFN28883_n),
	.A2(n15972),
	.B(n14159));
   NOR2xp33_ASAP7_75t_L U19361 (.Y(n15417),
	.A(n15411),
	.B(FE_OFN29018_n15921));
   NOR2xp33_ASAP7_75t_L U19362 (.Y(n14250),
	.A(n14289),
	.B(FE_OFN28624_n13874));
   NOR3xp33_ASAP7_75t_SRAM U19363 (.Y(n15273),
	.A(n14276),
	.B(FE_OFN28_w3_23),
	.C(n15658));
   NOR2xp33_ASAP7_75t_R U19364 (.Y(n14255),
	.A(n14334),
	.B(n15496));
   NOR2xp33_ASAP7_75t_SRAM U19365 (.Y(n14257),
	.A(FE_PSN8334_n15539),
	.B(n15496));
   NOR2xp33_ASAP7_75t_SRAM U19366 (.Y(n14301),
	.A(n15528),
	.B(n14302));
   AND3x1_ASAP7_75t_SL U19367 (.Y(n14304),
	.A(n14300),
	.B(n14299),
	.C(n14298));
   NAND3xp33_ASAP7_75t_SRAM U19368 (.Y(n14299),
	.A(n15347),
	.B(FE_OFN28712_n),
	.C(FE_OFN28_w3_23));
   NAND2xp5_ASAP7_75t_SL U19369 (.Y(n14300),
	.A(n14296),
	.B(n14295));
   NOR2xp33_ASAP7_75t_SRAM U19370 (.Y(n14305),
	.A(n14303),
	.B(n14302));
   OAI222xp33_ASAP7_75t_SRAM U19371 (.Y(n14789),
	.A1(n14315),
	.A2(n14314),
	.B1(FE_OFN37_w3_23),
	.B2(n14314),
	.C1(FE_OCPN27987_FE_OFN4_w3_22),
	.C2(n14314));
   OAI21xp5_ASAP7_75t_L U19372 (.Y(n15520),
	.A1(FE_OFN27214_w3_17),
	.A2(FE_OFN4_w3_22),
	.B(n14747));
   NOR2xp33_ASAP7_75t_R U19373 (.Y(n14279),
	.A(n15683),
	.B(n14790));
   INVxp67_ASAP7_75t_L U19374 (.Y(n14280),
	.A(n14278));
   NAND2xp33_ASAP7_75t_SL U19375 (.Y(n14277),
	.A(n14398),
	.B(n15339));
   INVxp33_ASAP7_75t_SRAM U19376 (.Y(n14281),
	.A(n14795));
   NOR2xp33_ASAP7_75t_R U19377 (.Y(n13447),
	.A(n15259),
	.B(n15195));
   NAND2xp5_ASAP7_75t_R U19378 (.Y(n15605),
	.A(n15599),
	.B(n15602));
   NOR2xp33_ASAP7_75t_R U19379 (.Y(n15599),
	.A(n15595),
	.B(n15600));
   NAND2xp5_ASAP7_75t_R U19380 (.Y(n15604),
	.A(n15603),
	.B(n15602));
   NOR2xp33_ASAP7_75t_R U19381 (.Y(n15603),
	.A(n15601),
	.B(n15600));
   NAND2xp33_ASAP7_75t_L U19382 (.Y(n15614),
	.A(n15608),
	.B(n15611));
   NOR2xp33_ASAP7_75t_SRAM U19383 (.Y(n15608),
	.A(n15838),
	.B(n15609));
   NAND2xp33_ASAP7_75t_L U19384 (.Y(n15613),
	.A(n15612),
	.B(n15611));
   NOR2xp33_ASAP7_75t_R U19385 (.Y(n15612),
	.A(n15610),
	.B(n15609));
   NAND2xp33_ASAP7_75t_L U19387 (.Y(n15643),
	.A(n15638),
	.B(n15640));
   NOR2xp33_ASAP7_75t_SL U19388 (.Y(n15638),
	.A(n15636),
	.B(n15789));
   NAND2xp33_ASAP7_75t_L U19389 (.Y(n15642),
	.A(n15641),
	.B(n15640));
   NOR2xp33_ASAP7_75t_R U19390 (.Y(n15641),
	.A(FE_OFN25912_n15848),
	.B(n15789));
   NAND2xp33_ASAP7_75t_SRAM U19391 (.Y(n15634),
	.A(n15629),
	.B(n15631));
   NOR2xp33_ASAP7_75t_L U19392 (.Y(n15629),
	.A(n15838),
	.B(n15630));
   NAND2xp33_ASAP7_75t_R U19393 (.Y(n15633),
	.A(n15632),
	.B(n15631));
   NOR2xp33_ASAP7_75t_L U19394 (.Y(n15632),
	.A(n15847),
	.B(n15630));
   NAND2x1p5_ASAP7_75t_L U19395 (.Y(n15948),
	.A(FE_OFN16417_n),
	.B(n15386));
   NOR2xp33_ASAP7_75t_SL U19396 (.Y(n14952),
	.A(n14951),
	.B(n14950));
   NAND3xp33_ASAP7_75t_SL U19397 (.Y(n14950),
	.A(n14949),
	.B(n14948),
	.C(n14947));
   NAND2xp5_ASAP7_75t_L U19398 (.Y(n14948),
	.A(FE_OFN27200_n),
	.B(n14943));
   NAND2xp33_ASAP7_75t_SRAM U19399 (.Y(n14954),
	.A(n13844),
	.B(n15444));
   NOR2xp33_ASAP7_75t_SL U19400 (.Y(n14906),
	.A(n15386),
	.B(n16009));
   NAND2xp33_ASAP7_75t_L U19401 (.Y(n15413),
	.A(FE_OFN26624_n15376),
	.B(n14938));
   NOR3xp33_ASAP7_75t_SL U19402 (.Y(n15715),
	.A(FE_OFN16210_n13876),
	.B(FE_OFN26535_w3_19),
	.C(FE_OFN28551_FE_OFN26114_n));
   NOR2xp33_ASAP7_75t_L U19403 (.Y(n15540),
	.A(n13875),
	.B(FE_PSN8334_n15539));
   NAND2xp5_ASAP7_75t_L U19404 (.Y(n15549),
	.A(n15544),
	.B(n15546));
   NOR2xp33_ASAP7_75t_R U19405 (.Y(n15544),
	.A(n12994),
	.B(n15545));
   OAI21xp5_ASAP7_75t_R U19406 (.Y(n15688),
	.A1(FE_OFN28977_n),
	.A2(FE_OFN26053_n25415),
	.B(FE_OFN6_w3_22));
   NAND2xp33_ASAP7_75t_L U19407 (.Y(n15500),
	.A(n15495),
	.B(n15497));
   NOR2xp33_ASAP7_75t_SRAM U19408 (.Y(n15495),
	.A(n15492),
	.B(n15496));
   NOR2xp33_ASAP7_75t_R U19409 (.Y(n15498),
	.A(n15714),
	.B(n15496));
   NAND2xp33_ASAP7_75t_L U19410 (.Y(n15511),
	.A(n15505),
	.B(n15508));
   NOR2xp33_ASAP7_75t_SRAM U19411 (.Y(n15505),
	.A(n12994),
	.B(n15507));
   NAND2xp5_ASAP7_75t_L U19412 (.Y(n15510),
	.A(n15509),
	.B(n15508));
   NOR2xp33_ASAP7_75t_SL U19413 (.Y(n15509),
	.A(FE_OFN72_n15506),
	.B(n15507));
   NAND2xp5_ASAP7_75t_L U19414 (.Y(n15526),
	.A(n15515),
	.B(n15525));
   NAND2xp33_ASAP7_75t_SL U19415 (.Y(n15525),
	.A(n15524),
	.B(n15523));
   NAND2xp5_ASAP7_75t_L U19417 (.Y(n13486),
	.A(n13485),
	.B(n13482));
   AND3x1_ASAP7_75t_L U19418 (.Y(n13506),
	.A(n13503),
	.B(n13502),
	.C(n13501));
   NOR3xp33_ASAP7_75t_SL U19420 (.Y(n13655),
	.A(n15200),
	.B(FE_OFN27212_w3_30),
	.C(FE_OFN28890_n));
   INVxp67_ASAP7_75t_R U19421 (.Y(n15234),
	.A(n13519));
   OAI21xp33_ASAP7_75t_L U19422 (.Y(n13520),
	.A1(n14559),
	.A2(FE_OFN16225_n15195),
	.B(n13515));
   NAND2xp33_ASAP7_75t_SRAM U19423 (.Y(n13515),
	.A(FE_OFN28530_n14593),
	.B(n15185));
   NOR2xp33_ASAP7_75t_SRAM U19424 (.Y(n13518),
	.A(FE_OFN16193_n15200),
	.B(n13520));
   OA21x2_ASAP7_75t_SRAM U19425 (.Y(n13521),
	.A1(FE_OFN28453_n13348),
	.A2(n15196),
	.B(n13517));
   OAI222xp33_ASAP7_75t_L U19426 (.Y(n13517),
	.A1(FE_OCPN27656_w3_25),
	.A2(n13516),
	.B1(FE_OFN25966_n13646),
	.B2(n13516),
	.C1(FE_OFN27044_n15236),
	.C2(n13516));
   NAND2xp33_ASAP7_75t_SRAM U19427 (.Y(n13531),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN25966_n13646));
   OAI22xp33_ASAP7_75t_R U19428 (.Y(n13529),
	.A1(FE_OFN27044_n15236),
	.A2(n13528),
	.B1(n14493),
	.B2(n13528));
   NOR2xp33_ASAP7_75t_SRAM U19429 (.Y(n13536),
	.A(FE_OFN16437_n),
	.B(n13534));
   NOR2xp33_ASAP7_75t_SRAM U19430 (.Y(n13533),
	.A(n14566),
	.B(n13534));
   NOR2xp33_ASAP7_75t_SRAM U19431 (.Y(n15103),
	.A(n15859),
	.B(n15101));
   OA21x2_ASAP7_75t_L U19432 (.Y(n15102),
	.A1(n24831),
	.A2(n15099),
	.B(n15098));
   NAND2xp33_ASAP7_75t_L U19433 (.Y(n15098),
	.A(n15097),
	.B(n15096));
   NAND2xp33_ASAP7_75t_L U19434 (.Y(n15097),
	.A(n15095),
	.B(n15094));
   O2A1O1Ixp33_ASAP7_75t_R U19435 (.Y(n15592),
	.A1(FE_OFN28732_n),
	.A2(n25140),
	.B(n13736),
	.C(FE_OFN28695_n));
   NOR2xp33_ASAP7_75t_L U19436 (.Y(n15082),
	.A(n15637),
	.B(n15081));
   NOR2xp33_ASAP7_75t_SRAM U19437 (.Y(n15081),
	.A(n15598),
	.B(FE_OCPN28398_n15808));
   NAND2xp33_ASAP7_75t_L U19438 (.Y(n14726),
	.A(n14725),
	.B(n14724));
   NAND2xp33_ASAP7_75t_SRAM U19439 (.Y(n14724),
	.A(n15380),
	.B(n14723));
   NAND2xp33_ASAP7_75t_SL U19440 (.Y(n14725),
	.A(n14722),
	.B(n14723));
   NAND2xp5_ASAP7_75t_SL U19442 (.Y(n14728),
	.A(n14721),
	.B(n14720));
   NAND2xp33_ASAP7_75t_SL U19443 (.Y(n14721),
	.A(n14718),
	.B(n14717));
   OAI21xp33_ASAP7_75t_SRAM U19445 (.Y(n14729),
	.A1(FE_OCPN29583_n15422),
	.A2(n14712),
	.B(n15955));
   NOR2xp33_ASAP7_75t_R U19446 (.Y(n14702),
	.A(n15972),
	.B(n14694));
   OA21x2_ASAP7_75t_L U19447 (.Y(n14703),
	.A1(n13805),
	.A2(FE_OFN25920_n15995),
	.B(n14700));
   NAND2xp5_ASAP7_75t_L U19448 (.Y(n14699),
	.A(n14698),
	.B(n14697));
   NAND2xp5_ASAP7_75t_R U19449 (.Y(n14698),
	.A(n14696),
	.B(n14919));
   NOR3xp33_ASAP7_75t_SRAM U19450 (.Y(n14707),
	.A(FE_OFN112_n15994),
	.B(FE_OFN26639_w3_14),
	.C(FE_OFN16459_n));
   OR3x1_ASAP7_75t_SRAM U19451 (.Y(n14709),
	.A(n14901),
	.B(n16009),
	.C(n16016));
   NOR2xp33_ASAP7_75t_SL U19452 (.Y(n14686),
	.A(n15380),
	.B(n13805));
   NAND2xp5_ASAP7_75t_L U19453 (.Y(n14685),
	.A(n14683),
	.B(n14682));
   NAND2xp33_ASAP7_75t_SRAM U19454 (.Y(n14682),
	.A(n14681),
	.B(FE_OFN29017_n15921));
   NAND2xp33_ASAP7_75t_SRAM U19455 (.Y(n14683),
	.A(n14680),
	.B(FE_OFN29017_n15921));
   NAND2xp5_ASAP7_75t_SL U19456 (.Y(n15705),
	.A(n15692),
	.B(n15691));
   NAND2xp5_ASAP7_75t_L U19457 (.Y(n15691),
	.A(n15690),
	.B(n15689));
   NAND2xp5_ASAP7_75t_L U19458 (.Y(n15692),
	.A(n15686),
	.B(n15689));
   AND2x2_ASAP7_75t_L U19459 (.Y(n15689),
	.A(n15685),
	.B(n15684));
   NAND2xp5_ASAP7_75t_L U19460 (.Y(n15703),
	.A(n15702),
	.B(n15701));
   NAND2xp33_ASAP7_75t_L U19461 (.Y(n15701),
	.A(n15700),
	.B(n15699));
   NAND2xp33_ASAP7_75t_L U19462 (.Y(n15702),
	.A(n15696),
	.B(n15699));
   INVxp67_ASAP7_75t_L U19463 (.Y(n15699),
	.A(n15695));
   NOR2xp33_ASAP7_75t_SRAM U19464 (.Y(n15731),
	.A(n15729),
	.B(n15728));
   OA21x2_ASAP7_75t_L U19465 (.Y(n15730),
	.A1(n15726),
	.A2(FE_OFN16352_n14289),
	.B(n15724));
   NAND2xp5_ASAP7_75t_L U19466 (.Y(n15724),
	.A(n15723),
	.B(n15722));
   NAND2xp33_ASAP7_75t_SL U19467 (.Y(n15722),
	.A(n15720),
	.B(n15721));
   NAND2xp33_ASAP7_75t_SL U19468 (.Y(n15723),
	.A(n15718),
	.B(n15721));
   NOR2xp33_ASAP7_75t_SRAM U19469 (.Y(n15727),
	.A(n15712),
	.B(n15728));
   NAND2xp33_ASAP7_75t_R U19470 (.Y(n15742),
	.A(n15741),
	.B(FE_OFN28600_n14289));
   NOR2xp33_ASAP7_75t_SRAM U19471 (.Y(n15741),
	.A(FE_OFN28624_n13874),
	.B(n15739));
   NAND2xp5_ASAP7_75t_L U19472 (.Y(n15754),
	.A(n15748),
	.B(n15751));
   NAND2xp33_ASAP7_75t_R U19473 (.Y(n15753),
	.A(n15752),
	.B(n15751));
   NOR2xp33_ASAP7_75t_L U19474 (.Y(n15752),
	.A(n15750),
	.B(n15749));
   NOR2xp33_ASAP7_75t_SL U19475 (.Y(n15746),
	.A(FE_OFN28769_n15478),
	.B(FE_OFN27074_n13868));
   NOR2xp33_ASAP7_75t_SL U19477 (.Y(n13663),
	.A(n13657),
	.B(n13656));
   NOR2xp33_ASAP7_75t_R U19478 (.Y(n13657),
	.A(FE_OFN26552_n14545),
	.B(FE_OFN25893_n15214));
   OA21x2_ASAP7_75t_L U19480 (.Y(n13664),
	.A1(FE_OFN25895_n13662),
	.A2(n14504),
	.B(n13661));
   NAND2xp5_ASAP7_75t_L U19481 (.Y(n13661),
	.A(n15197),
	.B(n13660));
   NAND2xp5_ASAP7_75t_SL U19482 (.Y(n13688),
	.A(n13687),
	.B(n13686));
   NAND2xp33_ASAP7_75t_L U19483 (.Y(n13686),
	.A(n13685),
	.B(n13684));
   NOR2xp33_ASAP7_75t_SRAM U19484 (.Y(n13685),
	.A(n25675),
	.B(n15162));
   NAND2xp33_ASAP7_75t_SL U19485 (.Y(n13690),
	.A(n13681),
	.B(n13680));
   NAND2xp33_ASAP7_75t_L U19486 (.Y(n13680),
	.A(n13679),
	.B(n13678));
   NAND2xp33_ASAP7_75t_L U19487 (.Y(n13681),
	.A(n13675),
	.B(n13678));
   INVxp67_ASAP7_75t_L U19488 (.Y(n13678),
	.A(n13674));
   NOR2xp33_ASAP7_75t_SL U19489 (.Y(n13691),
	.A(n15200),
	.B(n15259));
   NAND3xp33_ASAP7_75t_L U19490 (.Y(n13695),
	.A(FE_OFN25966_n13646),
	.B(FE_OFN16159_w3_24),
	.C(FE_OFN16412_w3_26));
   NOR2xp33_ASAP7_75t_L U19491 (.Y(n14455),
	.A(n14453),
	.B(n14452));
   NAND2xp33_ASAP7_75t_SRAM U19492 (.Y(n14453),
	.A(FE_OFN25928_n15779),
	.B(n15825));
   NAND2xp33_ASAP7_75t_L U19493 (.Y(n14457),
	.A(n14451),
	.B(n14454));
   NOR2xp33_ASAP7_75t_L U19494 (.Y(n14833),
	.A(n14458),
	.B(n15118));
   NOR2xp33_ASAP7_75t_R U19495 (.Y(n14458),
	.A(n14989),
	.B(n15813));
   NOR2xp33_ASAP7_75t_SRAM U19496 (.Y(n14423),
	.A(FE_OFN25886_w3_3),
	.B(n14996));
   NOR2xp33_ASAP7_75t_L U19497 (.Y(n14411),
	.A(FE_OCPN29537_FE_OFN28699_w3_6),
	.B(n14412));
   NOR2xp33_ASAP7_75t_L U19498 (.Y(n14414),
	.A(FE_OFN28732_n),
	.B(n14412));
   A2O1A1Ixp33_ASAP7_75t_SL U19499 (.Y(n16031),
	.A1(n15971),
	.A2(n15970),
	.B(n15969),
	.C(n15968));
   NAND2xp33_ASAP7_75t_SL U19501 (.Y(n15968),
	.A(n15967),
	.B(n15966));
   OAI21xp33_ASAP7_75t_L U19502 (.Y(n15947),
	.A1(FE_OCPN29564_n16012),
	.A2(n16010),
	.B(n15946));
   NOR2xp33_ASAP7_75t_SL U19503 (.Y(n16030),
	.A(n15972),
	.B(n16031));
   INVxp67_ASAP7_75t_L U19504 (.Y(n16033),
	.A(n16029));
   A2O1A1Ixp33_ASAP7_75t_L U19505 (.Y(n16029),
	.A1(n16028),
	.A2(n16027),
	.B(n16026),
	.C(n16025));
   NAND2xp5_ASAP7_75t_R U19506 (.Y(n16027),
	.A(n15991),
	.B(n15990));
   NAND2xp33_ASAP7_75t_L U19507 (.Y(n16028),
	.A(n15982),
	.B(n15981));
   NOR2x1_ASAP7_75t_L U19508 (.Y(n16032),
	.A(FE_OFN109_n15994),
	.B(n15969));
   NOR2xp33_ASAP7_75t_R U19509 (.Y(n15928),
	.A(n15993),
	.B(FE_OFN29017_n15921));
   OAI22xp33_ASAP7_75t_SRAM U19510 (.Y(n15926),
	.A1(n15922),
	.A2(FE_OFN26131_n15376),
	.B1(n15987),
	.B2(FE_OFN26131_n15376));
   NAND2xp33_ASAP7_75t_SRAM U19511 (.Y(n15925),
	.A(FE_PSN8271_n15924),
	.B(n15923));
   NOR2xp33_ASAP7_75t_R U19512 (.Y(n15938),
	.A(n15934),
	.B(n15939));
   INVxp33_ASAP7_75t_R U19513 (.Y(n15940),
	.A(n15937));
   NAND3xp33_ASAP7_75t_SL U19514 (.Y(n24518),
	.A(n24100),
	.B(FE_OCPN29376_n24099),
	.C(n24098));
   NAND2xp33_ASAP7_75t_R U19516 (.Y(n25744),
	.A(n25743),
	.B(n25742));
   NOR2xp33_ASAP7_75t_SRAM U19517 (.Y(n25743),
	.A(n25741),
	.B(n25740));
   NAND2xp33_ASAP7_75t_R U19518 (.Y(n25745),
	.A(n25739),
	.B(n25742));
   NAND3xp33_ASAP7_75t_L U19519 (.Y(n24777),
	.A(n24776),
	.B(n24775),
	.C(n24774));
   NAND2xp5_ASAP7_75t_R U19520 (.Y(n24776),
	.A(n24773),
	.B(n24772));
   NAND2xp33_ASAP7_75t_L U19521 (.Y(n24773),
	.A(n24768),
	.B(n24770));
   A2O1A1Ixp33_ASAP7_75t_SL U19522 (.Y(n24628),
	.A1(n24626),
	.A2(n24625),
	.B(n26777),
	.C(n26773));
   NAND2xp5_ASAP7_75t_SL U19525 (.Y(n25096),
	.A(FE_OCPN28098_n20907),
	.B(n19329));
   NOR2x1_ASAP7_75t_L U19526 (.Y(n24739),
	.A(n23119),
	.B(n24956));
   NAND2xp5_ASAP7_75t_SL U19527 (.Y(n26598),
	.A(n25442),
	.B(n25441));
   NAND3xp33_ASAP7_75t_L U19528 (.Y(n25068),
	.A(n25062),
	.B(n25061),
	.C(n25060));
   NAND3xp33_ASAP7_75t_L U19529 (.Y(n25067),
	.A(n25065),
	.B(FE_OCPN28427_n25064),
	.C(n25063));
   NAND2xp33_ASAP7_75t_L U19530 (.Y(n25061),
	.A(n25059),
	.B(n25058));
   NAND3xp33_ASAP7_75t_R U19532 (.Y(n25260),
	.A(n25259),
	.B(n26104),
	.C(n25258));
   NAND2xp33_ASAP7_75t_SRAM U19533 (.Y(n25257),
	.A(FE_OFN30_n25256),
	.B(FE_OFN28767_n26103));
   NAND2xp5_ASAP7_75t_L U19535 (.Y(n26072),
	.A(n26070),
	.B(n26069));
   NAND2xp33_ASAP7_75t_L U19536 (.Y(n26069),
	.A(n26068),
	.B(n26067));
   NAND2xp5_ASAP7_75t_R U19537 (.Y(n26070),
	.A(n26066),
	.B(n26067));
   NAND2xp5_ASAP7_75t_SL U19538 (.Y(n25550),
	.A(n25548),
	.B(n25547));
   NAND2xp33_ASAP7_75t_L U19539 (.Y(n25548),
	.A(n25543),
	.B(n17058));
   NAND2xp33_ASAP7_75t_SL U19540 (.Y(n25547),
	.A(n25546),
	.B(n17058));
   NOR2xp33_ASAP7_75t_L U19541 (.Y(n25543),
	.A(FE_OFN28584_n17001),
	.B(n25544));
   O2A1O1Ixp5_ASAP7_75t_SL U19544 (.Y(n25851),
	.A1(n24194),
	.A2(n24193),
	.B(n26407),
	.C(n24192));
   NAND3xp33_ASAP7_75t_SL U19545 (.Y(n24193),
	.A(n24191),
	.B(n24190),
	.C(n24189));
   NAND2xp5_ASAP7_75t_R U19546 (.Y(n24190),
	.A(n24188),
	.B(n24187));
   NAND2xp33_ASAP7_75t_L U19547 (.Y(n24187),
	.A(n24186),
	.B(n24185));
   NAND2xp33_ASAP7_75t_L U19549 (.Y(n26564),
	.A(n26563),
	.B(n26562));
   NOR2xp33_ASAP7_75t_L U19550 (.Y(n26563),
	.A(n26561),
	.B(sa23_7_));
   INVx1_ASAP7_75t_L U19551 (.Y(n26706),
	.A(n26703));
   NAND2xp33_ASAP7_75t_L U19552 (.Y(n25713),
	.A(n26663),
	.B(n20912));
   INVxp33_ASAP7_75t_SRAM U19553 (.Y(n20912),
	.A(n22971));
   NOR3xp33_ASAP7_75t_SL U19555 (.Y(n25138),
	.A(n24954),
	.B(n24953),
	.C(n24952));
   NAND2xp33_ASAP7_75t_L U19556 (.Y(n24950),
	.A(n24948),
	.B(n24947));
   NAND2xp33_ASAP7_75t_L U19557 (.Y(n24947),
	.A(n24946),
	.B(n24945));
   NAND2xp33_ASAP7_75t_SRAM U19558 (.Y(n19208),
	.A(n23391),
	.B(n19207));
   OAI22xp33_ASAP7_75t_SRAM U19559 (.Y(n19207),
	.A1(n17444),
	.A2(n21817),
	.B1(n19206),
	.B2(n21817));
   NAND2xp5_ASAP7_75t_SL U19560 (.Y(n23283),
	.A(n19234),
	.B(n19233));
   NAND2xp5_ASAP7_75t_L U19561 (.Y(n19234),
	.A(n19230),
	.B(n19231));
   NOR2xp33_ASAP7_75t_SRAM U19564 (.Y(n19212),
	.A(n21821),
	.B(FE_OCPN27496_n21820));
   NOR2xp33_ASAP7_75t_SL U19565 (.Y(n20010),
	.A(FE_OFN28914_n20007),
	.B(n20011));
   AND3x1_ASAP7_75t_SRAM U19566 (.Y(n20012),
	.A(n20009),
	.B(n23656),
	.C(n20008));
   NAND2xp5_ASAP7_75t_SL U19567 (.Y(n20014),
	.A(n20013),
	.B(n20012));
   NOR2xp33_ASAP7_75t_SL U19568 (.Y(n20013),
	.A(FE_OFN29023_n16750),
	.B(n20011));
   NAND2xp5_ASAP7_75t_R U19569 (.Y(n19992),
	.A(n16771),
	.B(FE_OCPN28298_n));
   NOR2x1_ASAP7_75t_L U19570 (.Y(n19967),
	.A(FE_OCPN27556_n17843),
	.B(n16777));
   NAND2xp5_ASAP7_75t_L U19572 (.Y(n18084),
	.A(FE_PSN8293_n25317),
	.B(n26399));
   NOR2xp33_ASAP7_75t_L U19573 (.Y(n18086),
	.A(n18085),
	.B(n18084));
   NAND2xp5_ASAP7_75t_SL U19574 (.Y(n18087),
	.A(n24181),
	.B(n16348));
   NAND2xp5_ASAP7_75t_SL U19575 (.Y(n23233),
	.A(n19558),
	.B(n19557));
   NAND2xp5_ASAP7_75t_L U19576 (.Y(n19557),
	.A(n19556),
	.B(n19555));
   NAND2xp5_ASAP7_75t_L U19577 (.Y(n19558),
	.A(n19553),
	.B(n19555));
   NOR2xp33_ASAP7_75t_R U19578 (.Y(n19556),
	.A(n23587),
	.B(n19554));
   NOR2xp33_ASAP7_75t_R U19579 (.Y(n23228),
	.A(FE_OCPN5137_n23600),
	.B(n23588));
   NAND2xp33_ASAP7_75t_SL U19580 (.Y(n23230),
	.A(n23226),
	.B(n23227));
   NOR2xp33_ASAP7_75t_SRAM U19581 (.Y(n23226),
	.A(n24364),
	.B(n23588));
   INVx1_ASAP7_75t_L U19582 (.Y(n23221),
	.A(n23218));
   NAND2xp33_ASAP7_75t_R U19584 (.Y(n22770),
	.A(n22766),
	.B(n22767));
   NAND2xp5_ASAP7_75t_SL U19585 (.Y(n23268),
	.A(n19170),
	.B(n19225));
   NOR2xp33_ASAP7_75t_L U19586 (.Y(n17495),
	.A(n21365),
	.B(n19192));
   OAI21xp5_ASAP7_75t_L U19587 (.Y(n21395),
	.A1(FE_OCPN27313_n21845),
	.A2(FE_OCPN28006_n17454),
	.B(n19210));
   NOR2xp33_ASAP7_75t_R U19588 (.Y(n21827),
	.A(n21819),
	.B(FE_OCPN28175_n21818));
   AND3x1_ASAP7_75t_SL U19589 (.Y(n21828),
	.A(n21825),
	.B(n21846),
	.C(n21824));
   NOR2xp33_ASAP7_75t_R U19591 (.Y(n22157),
	.A(FE_OCPN29398_sa30_3),
	.B(n18503));
   NOR2x1_ASAP7_75t_SL U19592 (.Y(n23323),
	.A(FE_OCPN29305_n23302),
	.B(n23160));
   NAND2xp5_ASAP7_75t_SL U19593 (.Y(n23343),
	.A(n20758),
	.B(n20757));
   NAND2xp33_ASAP7_75t_SL U19594 (.Y(n20757),
	.A(n20756),
	.B(n20755));
   NAND2xp33_ASAP7_75t_SL U19595 (.Y(n20758),
	.A(n20754),
	.B(n20755));
   NOR2x1_ASAP7_75t_L U19596 (.Y(n20756),
	.A(FE_OFN25952_n22312),
	.B(n23161));
   AND3x1_ASAP7_75t_R U19597 (.Y(n23316),
	.A(n23312),
	.B(n23311),
	.C(n23310));
   NAND3xp33_ASAP7_75t_SL U19599 (.Y(n22709),
	.A(n20299),
	.B(n22657),
	.C(n22689));
   NOR2x1_ASAP7_75t_L U19600 (.Y(n16710),
	.A(n26122),
	.B(n16852));
   NAND2xp5_ASAP7_75t_SL U19601 (.Y(n16726),
	.A(n16424),
	.B(n16425));
   NOR2xp33_ASAP7_75t_R U19602 (.Y(n16425),
	.A(n23556),
	.B(FE_OFN27062_n16438));
   NAND2xp33_ASAP7_75t_L U19604 (.Y(n16480),
	.A(n16840),
	.B(n16686));
   NOR2xp33_ASAP7_75t_L U19606 (.Y(n16471),
	.A(n24328),
	.B(n18431));
   OAI22xp33_ASAP7_75t_SRAM U19607 (.Y(n16440),
	.A1(FE_OFN29101_n16418),
	.A2(n17405),
	.B1(n16430),
	.B2(n17405));
   NOR2x1_ASAP7_75t_SL U19608 (.Y(n23750),
	.A(n23719),
	.B(n21648));
   NAND2xp5_ASAP7_75t_L U19609 (.Y(n19704),
	.A(n18299),
	.B(n18335));
   NOR2xp33_ASAP7_75t_SL U19610 (.Y(n17680),
	.A(FE_OFN69_sa32_4),
	.B(n19701));
   NOR2xp33_ASAP7_75t_SL U19611 (.Y(n17682),
	.A(n19712),
	.B(n19701));
   NAND2xp33_ASAP7_75t_SL U19612 (.Y(n17013),
	.A(n17010),
	.B(n18955));
   NOR2xp33_ASAP7_75t_SL U19613 (.Y(n17010),
	.A(FE_OCPN28212_n16980),
	.B(n20490));
   NAND2xp33_ASAP7_75t_SL U19614 (.Y(n17012),
	.A(n17011),
	.B(n18955));
   NOR2xp33_ASAP7_75t_L U19615 (.Y(n17011),
	.A(FE_OCPN27859_n25868),
	.B(n20490));
   NAND3xp33_ASAP7_75t_SL U19617 (.Y(n17019),
	.A(n25223),
	.B(n17018),
	.C(n17017));
   NAND2xp33_ASAP7_75t_SRAM U19618 (.Y(n17024),
	.A(n18946),
	.B(FE_OFN25977_n18922));
   NAND3xp33_ASAP7_75t_SRAM U19619 (.Y(n19263),
	.A(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(FE_OCPN27384_n22888),
	.C(FE_OFN28703_FE_OCPN27740_sa02_4));
   NOR2x1_ASAP7_75t_SL U19620 (.Y(n17565),
	.A(FE_OFN26035_n),
	.B(FE_OCPN27812_FE_OFN16463_sa32_0));
   NOR2x1p5_ASAP7_75t_SL U19621 (.Y(n19740),
	.A(FE_OCPN27882_n18829),
	.B(FE_OCPN27420_n18794));
   NAND2x1_ASAP7_75t_L U19622 (.Y(n19741),
	.A(FE_OCPN27230_sa32_3),
	.B(FE_OCPN27792_n18333));
   INVxp33_ASAP7_75t_SRAM U19623 (.Y(n19714),
	.A(n19710));
   NAND2xp33_ASAP7_75t_SRAM U19624 (.Y(n17567),
	.A(n18309),
	.B(n22372));
   NOR3x1_ASAP7_75t_SL U19625 (.Y(n24861),
	.A(n19732),
	.B(FE_OCPN7586_n17693),
	.C(n17675));
   NOR2x1p5_ASAP7_75t_R U19627 (.Y(n19703),
	.A(FE_OCPN27267_n18794),
	.B(FE_OCPN29323_n19721));
   AND3x2_ASAP7_75t_SL U19628 (.Y(n22022),
	.A(n20925),
	.B(n22006),
	.C(n20924));
   O2A1O1Ixp33_ASAP7_75t_SL U19629 (.Y(n20925),
	.A1(n19019),
	.A2(FE_OFN16248_n20235),
	.B(FE_OFN28752_n),
	.C(n22997));
   NAND2xp5_ASAP7_75t_R U19630 (.Y(n20915),
	.A(FE_OCPN29489_sa23_3),
	.B(n19337));
   NAND2xp33_ASAP7_75t_L U19633 (.Y(n19335),
	.A(n20258),
	.B(n22046));
   NAND2xp5_ASAP7_75t_L U19634 (.Y(n19319),
	.A(n19318),
	.B(n19317));
   NOR2xp33_ASAP7_75t_L U19635 (.Y(n19318),
	.A(FE_OFN27056_n22995),
	.B(n22035));
   NAND2xp5_ASAP7_75t_L U19636 (.Y(n19320),
	.A(n19316),
	.B(n19317));
   NOR2xp33_ASAP7_75t_R U19638 (.Y(n19288),
	.A(FE_OFN28752_n),
	.B(n20931));
   NOR2x1_ASAP7_75t_L U19639 (.Y(n20943),
	.A(FE_OCPN28086_n22034),
	.B(n19002));
   NOR2x1_ASAP7_75t_L U19640 (.Y(n19302),
	.A(n22952),
	.B(FE_OCPN28289_n20235));
   NAND2xp33_ASAP7_75t_SL U19641 (.Y(n20160),
	.A(n20156),
	.B(n20157));
   NOR2xp33_ASAP7_75t_SL U19642 (.Y(n20156),
	.A(FE_OFN108_n26971),
	.B(n20175));
   NAND2xp33_ASAP7_75t_SL U19643 (.Y(n20159),
	.A(n20158),
	.B(n20157));
   NOR2xp33_ASAP7_75t_SL U19644 (.Y(n20158),
	.A(FE_OFN28626_n22094),
	.B(n20175));
   NAND2xp33_ASAP7_75t_R U19645 (.Y(n20151),
	.A(n20149),
	.B(n21004));
   NOR2xp33_ASAP7_75t_L U19646 (.Y(n20143),
	.A(n17757),
	.B(n20144));
   NOR2xp67_ASAP7_75t_L U19647 (.Y(n20129),
	.A(FE_OCPN27624_n26971),
	.B(FE_OCPN29341_FE_OFN29148_n));
   NAND2xp5_ASAP7_75t_L U19648 (.Y(n22553),
	.A(n22552),
	.B(n22551));
   NAND2xp33_ASAP7_75t_L U19649 (.Y(n22552),
	.A(n22548),
	.B(n22549));
   NAND2xp33_ASAP7_75t_SL U19650 (.Y(n22551),
	.A(n22550),
	.B(n22549));
   NOR3xp33_ASAP7_75t_SRAM U19651 (.Y(n22559),
	.A(n25531),
	.B(FE_OCPN27972_n20988),
	.C(n25523));
   NAND3x1_ASAP7_75t_SL U19652 (.Y(n22565),
	.A(n20174),
	.B(n20173),
	.C(FE_OCPN27689_n20172));
   NOR3x1_ASAP7_75t_L U19653 (.Y(n20173),
	.A(n20212),
	.B(n20978),
	.C(FE_OFN28924_n25912));
   NAND2xp5_ASAP7_75t_SL U19654 (.Y(n22562),
	.A(n22110),
	.B(n20153));
   NOR2xp33_ASAP7_75t_SL U19655 (.Y(n22564),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(n19263));
   NAND2xp5_ASAP7_75t_SL U19656 (.Y(n20142),
	.A(FE_OCPN27261_sa02_0),
	.B(n17749));
   NOR2xp33_ASAP7_75t_SL U19657 (.Y(n20136),
	.A(n20962),
	.B(FE_OFN29184_n17744));
   NOR3x1_ASAP7_75t_SL U19658 (.Y(n20203),
	.A(n20140),
	.B(n20139),
	.C(n20138));
   NAND3xp33_ASAP7_75t_SL U19659 (.Y(n20140),
	.A(n20137),
	.B(n22892),
	.C(n25204));
   NOR3xp33_ASAP7_75t_L U19660 (.Y(n23346),
	.A(n22288),
	.B(n22287),
	.C(n22286));
   NAND2xp5_ASAP7_75t_L U19661 (.Y(n22288),
	.A(n22285),
	.B(n22284));
   NOR3xp33_ASAP7_75t_SL U19662 (.Y(n22284),
	.A(n22283),
	.B(n22282),
	.C(n22281));
   NAND2xp5_ASAP7_75t_L U19663 (.Y(n22283),
	.A(n22280),
	.B(n22279));
   NOR2x1_ASAP7_75t_L U19664 (.Y(n22296),
	.A(n26871),
	.B(n22850));
   OAI21xp33_ASAP7_75t_L U19666 (.Y(n22836),
	.A1(n23160),
	.A2(FE_OCPN29305_n23302),
	.B(n22311));
   NAND3xp33_ASAP7_75t_SL U19667 (.Y(n22313),
	.A(n20766),
	.B(n23337),
	.C(n18181));
   NOR2xp33_ASAP7_75t_L U19668 (.Y(n18181),
	.A(n22321),
	.B(n21114));
   NAND2xp5_ASAP7_75t_R U19669 (.Y(n23342),
	.A(n22318),
	.B(n22317));
   NAND2xp33_ASAP7_75t_L U19670 (.Y(n21785),
	.A(FE_OFN16135_sa22_4),
	.B(n23308));
   NAND2xp33_ASAP7_75t_R U19671 (.Y(n19795),
	.A(n19790),
	.B(n19792));
   NAND3xp33_ASAP7_75t_SL U19672 (.Y(n24893),
	.A(n19801),
	.B(n23126),
	.C(n21884));
   NAND2xp5_ASAP7_75t_L U19673 (.Y(n19801),
	.A(n19800),
	.B(n19799));
   NAND2xp5_ASAP7_75t_L U19674 (.Y(n19800),
	.A(n19796),
	.B(n19797));
   NAND2xp5_ASAP7_75t_L U19675 (.Y(n19799),
	.A(n19798),
	.B(n19797));
   NOR2xp33_ASAP7_75t_L U19676 (.Y(n19802),
	.A(n19774),
	.B(n16617));
   NAND2xp33_ASAP7_75t_L U19677 (.Y(n16617),
	.A(n16616),
	.B(n19669));
   NAND2xp5_ASAP7_75t_L U19678 (.Y(n19777),
	.A(FE_OFN29204_sa10_2),
	.B(n17221));
   NAND2xp33_ASAP7_75t_R U19679 (.Y(n20665),
	.A(n20661),
	.B(n20662));
   NOR2xp33_ASAP7_75t_SRAM U19680 (.Y(n20661),
	.A(n20617),
	.B(n23775));
   NAND2xp33_ASAP7_75t_R U19681 (.Y(n20664),
	.A(n20663),
	.B(n20662));
   NAND2xp5_ASAP7_75t_L U19682 (.Y(n20673),
	.A(n20668),
	.B(n20667));
   NOR2xp33_ASAP7_75t_L U19683 (.Y(n20668),
	.A(FE_OFN29112_FE_OCPN27870_n18527),
	.B(n20669));
   NAND2x1_ASAP7_75t_L U19685 (.Y(n21684),
	.A(FE_OCPN27606_n23869),
	.B(FE_OFN16295_n23837));
   NAND2xp5_ASAP7_75t_L U19686 (.Y(n22210),
	.A(n22209),
	.B(n22208));
   OAI21xp5_ASAP7_75t_SL U19687 (.Y(n22205),
	.A1(FE_OFN26648_n22197),
	.A2(FE_OFN25878_n17329),
	.B(n18706));
   NAND2xp5_ASAP7_75t_SL U19688 (.Y(n21569),
	.A(n20368),
	.B(n22183));
   NAND2xp33_ASAP7_75t_L U19689 (.Y(n17373),
	.A(FE_OCPN8219_n22197),
	.B(n17321));
   OAI21xp5_ASAP7_75t_L U19690 (.Y(n21537),
	.A1(FE_OCPN27423_sa01_0),
	.A2(FE_OFN27150_n22175),
	.B(n22605));
   NOR2x1_ASAP7_75t_L U19691 (.Y(n19592),
	.A(n19150),
	.B(n21148));
   NOR2xp33_ASAP7_75t_SRAM U19692 (.Y(n19577),
	.A(FE_OCPN28389_n21479),
	.B(n19578));
   NAND2x1p5_ASAP7_75t_L U19693 (.Y(n18640),
	.A(FE_OFN28744_FE_OCPN27908),
	.B(FE_OFN28514_sa00_1));
   NAND2xp33_ASAP7_75t_L U19694 (.Y(n18628),
	.A(FE_OCPN29553_n19602),
	.B(n18742));
   NOR2x1p5_ASAP7_75t_SL U19695 (.Y(n18744),
	.A(n19578),
	.B(n19845));
   NAND2xp33_ASAP7_75t_SL U19697 (.Y(n23797),
	.A(n23765),
	.B(n18537));
   NOR2xp33_ASAP7_75t_SRAM U19699 (.Y(n23813),
	.A(FE_OCPN27715_n23875),
	.B(n23814));
   NAND2xp33_ASAP7_75t_SL U19700 (.Y(n23826),
	.A(n23822),
	.B(FE_OFN16328_n23821));
   NAND2xp33_ASAP7_75t_SL U19701 (.Y(n23825),
	.A(n23824),
	.B(FE_OFN16328_n23821));
   NAND3xp33_ASAP7_75t_SL U19702 (.Y(n25627),
	.A(n23834),
	.B(n23833),
	.C(n23832));
   NAND2xp5_ASAP7_75t_L U19703 (.Y(n25630),
	.A(n23844),
	.B(n23843));
   NAND2xp33_ASAP7_75t_L U19704 (.Y(n23843),
	.A(n23842),
	.B(FE_OFN16328_n23821));
   NAND2xp33_ASAP7_75t_L U19705 (.Y(n23844),
	.A(n23839),
	.B(FE_OFN16328_n23821));
   OAI21xp5_ASAP7_75t_SL U19706 (.Y(n21217),
	.A1(n23688),
	.A2(FE_OCPN28257_n23689),
	.B(n18570));
   NOR2xp33_ASAP7_75t_R U19707 (.Y(n20681),
	.A(FE_OFN29081_n18526),
	.B(FE_OCPN29567_n23806));
   NOR2xp33_ASAP7_75t_R U19709 (.Y(n20679),
	.A(FE_OFN16295_n23837),
	.B(FE_OCPN29567_n23806));
   NAND2xp33_ASAP7_75t_SRAM U19710 (.Y(n20594),
	.A(FE_OCPN28386_n17899),
	.B(FE_OCPN29555_n20593));
   NAND2x1_ASAP7_75t_SL U19711 (.Y(n20555),
	.A(FE_OCPN27429_sa12_3),
	.B(n17906));
   NAND2xp5_ASAP7_75t_SL U19712 (.Y(n18093),
	.A(n20050),
	.B(n20060));
   NAND3xp33_ASAP7_75t_L U19713 (.Y(n16398),
	.A(n16300),
	.B(n16348),
	.C(FE_OFN26060_sa31_4));
   NAND2xp33_ASAP7_75t_SRAM U19714 (.Y(n16504),
	.A(n26291),
	.B(FE_OFN29016_n16512));
   NAND2xp5_ASAP7_75t_SL U19715 (.Y(n16521),
	.A(n16376),
	.B(n16375));
   NOR3xp33_ASAP7_75t_L U19716 (.Y(n16376),
	.A(n26298),
	.B(n20876),
	.C(n16372));
   NOR2xp33_ASAP7_75t_SL U19717 (.Y(n16375),
	.A(n21965),
	.B(n16374));
   NAND2xp5_ASAP7_75t_SL U19718 (.Y(n18095),
	.A(n25816),
	.B(n16520));
   NOR2xp33_ASAP7_75t_SL U19719 (.Y(n16520),
	.A(n27070),
	.B(n20067));
   NAND2x1p5_ASAP7_75t_SL U19720 (.Y(n16594),
	.A(FE_OFN26587_n23011),
	.B(FE_OCPN28323_FE_OFN16427_sa10_3));
   NAND2xp5_ASAP7_75t_SL U19721 (.Y(n16652),
	.A(n16609),
	.B(n16608));
   NAND2xp33_ASAP7_75t_R U19722 (.Y(n16609),
	.A(FE_OFN28916_sa10_4),
	.B(n16631));
   NAND2xp33_ASAP7_75t_L U19723 (.Y(n16608),
	.A(n23024),
	.B(n16631));
   NAND3xp33_ASAP7_75t_SL U19724 (.Y(n23030),
	.A(n16652),
	.B(n21886),
	.C(n19683));
   NOR2xp33_ASAP7_75t_R U19725 (.Y(n21051),
	.A(FE_OFN28588_n21048),
	.B(FE_OCPN27405_sa03_4));
   NOR2xp33_ASAP7_75t_SRAM U19726 (.Y(n21053),
	.A(FE_OFN28614_n21715),
	.B(n21051));
   OR2x2_ASAP7_75t_SL U19727 (.Y(n21046),
	.A(n21706),
	.B(FE_OFN28588_n21048));
   NAND2xp5_ASAP7_75t_L U19729 (.Y(n19469),
	.A(n19465),
	.B(n19466));
   OR3x1_ASAP7_75t_SRAM U19730 (.Y(n21756),
	.A(n21730),
	.B(n21729),
	.C(n21728));
   NAND2xp5_ASAP7_75t_L U19731 (.Y(n21730),
	.A(n21727),
	.B(n21726));
   NOR3xp33_ASAP7_75t_L U19732 (.Y(n23497),
	.A(n20920),
	.B(FE_OCPN29374_FE_OFN29191_sa23_2),
	.C(n23504));
   AND3x1_ASAP7_75t_SL U19733 (.Y(n20937),
	.A(n20935),
	.B(n22019),
	.C(n20934));
   NOR2xp33_ASAP7_75t_SL U19735 (.Y(n20926),
	.A(n22998),
	.B(n23490));
   NAND3xp33_ASAP7_75t_L U19736 (.Y(n26146),
	.A(n18971),
	.B(FE_OFN27056_n22995),
	.C(FE_OCPN27627_sa23_1));
   NAND2xp33_ASAP7_75t_SRAM U19737 (.Y(n20412),
	.A(n20411),
	.B(n20410));
   NOR3xp33_ASAP7_75t_SL U19738 (.Y(n26465),
	.A(n20407),
	.B(FE_OFN26649_n22206),
	.C(n24392));
   NOR2xp33_ASAP7_75t_SL U19739 (.Y(n20360),
	.A(n22598),
	.B(n17345));
   NOR2xp33_ASAP7_75t_L U19740 (.Y(n25060),
	.A(n21560),
	.B(n23087));
   NAND2xp5_ASAP7_75t_R U19741 (.Y(n20380),
	.A(n25057),
	.B(n20367));
   NOR2xp33_ASAP7_75t_L U19742 (.Y(n20073),
	.A(FE_OCPN27786_n16490),
	.B(n20023));
   NOR2xp67_ASAP7_75t_R U19744 (.Y(n16499),
	.A(FE_OFN16415_sa31_2),
	.B(FE_PSN8293_n25317));
   NOR2xp33_ASAP7_75t_L U19745 (.Y(n18083),
	.A(n16496),
	.B(n16495));
   NAND2xp5_ASAP7_75t_L U19747 (.Y(n20343),
	.A(n20338),
	.B(n20340));
   NAND2xp5_ASAP7_75t_SL U19748 (.Y(n20342),
	.A(n20341),
	.B(n20340));
   NAND2xp33_ASAP7_75t_R U19749 (.Y(n20348),
	.A(n22682),
	.B(n20346));
   NAND2xp5_ASAP7_75t_SL U19750 (.Y(n16723),
	.A(n23533),
	.B(n18405));
   NAND2x1_ASAP7_75t_L U19751 (.Y(n16707),
	.A(n16427),
	.B(n16424));
   NOR2xp33_ASAP7_75t_SL U19753 (.Y(n17624),
	.A(n17622),
	.B(n18458));
   NAND2xp33_ASAP7_75t_SRAM U19755 (.Y(n17668),
	.A(n17664),
	.B(n17665));
   NAND3xp33_ASAP7_75t_R U19756 (.Y(n19387),
	.A(n19386),
	.B(n19385),
	.C(n25864));
   NAND3xp33_ASAP7_75t_SL U19757 (.Y(n19388),
	.A(n19384),
	.B(n19383),
	.C(n25228));
   NOR2xp33_ASAP7_75t_SRAM U19758 (.Y(n19383),
	.A(n19382),
	.B(n19381));
   NOR2xp33_ASAP7_75t_SRAM U19759 (.Y(n19384),
	.A(n19380),
	.B(FE_OCPN8231_n20522));
   NAND2xp33_ASAP7_75t_SL U19760 (.Y(n19369),
	.A(n19365),
	.B(n19366));
   NOR2xp33_ASAP7_75t_L U19761 (.Y(n19365),
	.A(FE_OFN28584_n17001),
	.B(FE_OCPN29437_n25864));
   NAND2xp5_ASAP7_75t_L U19762 (.Y(n19368),
	.A(n19367),
	.B(n19366));
   NOR2xp33_ASAP7_75t_SL U19763 (.Y(n19367),
	.A(FE_OCPN8213_FE_OFN29234_n16996),
	.B(FE_OCPN29437_n25864));
   OAI21xp5_ASAP7_75t_SL U19764 (.Y(n17139),
	.A1(n16989),
	.A2(n17002),
	.B(n17161));
   NAND2xp33_ASAP7_75t_SRAM U19765 (.Y(n17174),
	.A(n25995),
	.B(n18254));
   AND3x1_ASAP7_75t_SL U19766 (.Y(n17175),
	.A(n27088),
	.B(n18260),
	.C(n17172));
   NAND3xp33_ASAP7_75t_SL U19768 (.Y(n17162),
	.A(n19376),
	.B(FE_OCPN28121_n16975),
	.C(FE_OFN28491_sa13_3));
   NOR2x1_ASAP7_75t_SL U19769 (.Y(n20111),
	.A(n19932),
	.B(n19710));
   NAND3x1_ASAP7_75t_SL U19770 (.Y(n25988),
	.A(n25868),
	.B(FE_OCPN27761_n16977),
	.C(FE_OFN28809_n));
   NAND2xp33_ASAP7_75t_L U19771 (.Y(n18951),
	.A(n18950),
	.B(n18949));
   NAND2xp33_ASAP7_75t_SRAM U19772 (.Y(n18949),
	.A(n18948),
	.B(FE_OCPN29569_n18947));
   NAND2xp33_ASAP7_75t_SL U19773 (.Y(n18950),
	.A(n18946),
	.B(FE_OCPN29569_n18947));
   NOR2x1_ASAP7_75t_L U19774 (.Y(n18926),
	.A(n19430),
	.B(n17171));
   NOR2xp33_ASAP7_75t_SL U19775 (.Y(n18923),
	.A(n18921),
	.B(n20513));
   NOR2xp33_ASAP7_75t_SL U19776 (.Y(n18934),
	.A(FE_OCPN27859_n25868),
	.B(FE_OFN28622_n25870));
   NAND2xp33_ASAP7_75t_SL U19778 (.Y(n18937),
	.A(n18936),
	.B(FE_OFN25999_n25875));
   NOR2xp33_ASAP7_75t_R U19779 (.Y(n18936),
	.A(FE_OFN28584_n17001),
	.B(FE_OFN28622_n25870));
   NAND3xp33_ASAP7_75t_SL U19780 (.Y(n17077),
	.A(FE_OCPN29369_n16982),
	.B(n17170),
	.C(FE_OFN16444_sa13_1));
   NOR2x1_ASAP7_75t_L U19781 (.Y(n20168),
	.A(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(n17759));
   NAND2xp5_ASAP7_75t_L U19782 (.Y(n17759),
	.A(n22543),
	.B(n17758));
   INVxp67_ASAP7_75t_L U19783 (.Y(n17758),
	.A(n22529));
   NAND2xp5_ASAP7_75t_SL U19785 (.Y(n17740),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(FE_OCPN27740_sa02_4));
   NOR2x2_ASAP7_75t_SL U19786 (.Y(n25530),
	.A(FE_OFN28800_n22526),
	.B(n17780));
   NOR2x1_ASAP7_75t_L U19787 (.Y(n20172),
	.A(n20161),
	.B(n22894));
   NOR2xp33_ASAP7_75t_SRAM U19788 (.Y(n19925),
	.A(FE_OCPN29524_n25029),
	.B(n19926));
   AND3x1_ASAP7_75t_SL U19789 (.Y(n19927),
	.A(n19924),
	.B(n19923),
	.C(n19922));
   NOR2x1_ASAP7_75t_SL U19790 (.Y(n19932),
	.A(FE_OCPN27882_n18829),
	.B(n18828));
   NOR2xp33_ASAP7_75t_SRAM U19791 (.Y(n19944),
	.A(n18298),
	.B(n20107));
   NOR2xp33_ASAP7_75t_SRAM U19793 (.Y(n19946),
	.A(n22392),
	.B(n20107));
   NOR3x1_ASAP7_75t_L U19794 (.Y(n19700),
	.A(n19907),
	.B(n19740),
	.C(n19739));
   NOR2xp33_ASAP7_75t_R U19795 (.Y(n21283),
	.A(sa03_3_),
	.B(n21284));
   NAND3xp33_ASAP7_75t_SL U19796 (.Y(n21034),
	.A(n21304),
	.B(n18016),
	.C(FE_OCPN27726_n));
   NAND2xp5_ASAP7_75t_L U19797 (.Y(n21032),
	.A(n21030),
	.B(n21029));
   INVx1_ASAP7_75t_L U19798 (.Y(n21328),
	.A(n21325));
   NAND2xp33_ASAP7_75t_SL U19799 (.Y(n21324),
	.A(n21323),
	.B(n21322));
   NAND2xp5_ASAP7_75t_L U19800 (.Y(n21322),
	.A(n21321),
	.B(n21320));
   OAI21xp33_ASAP7_75t_L U19801 (.Y(n21284),
	.A1(FE_OFN28677_n17998),
	.A2(FE_OCPN27733_n17996),
	.B(n21044));
   NOR2xp33_ASAP7_75t_SRAM U19802 (.Y(n21044),
	.A(n21043),
	.B(FE_OCPN27918_n21042));
   NAND3xp33_ASAP7_75t_R U19803 (.Y(n21074),
	.A(n21047),
	.B(n21046),
	.C(n21045));
   OAI21x1_ASAP7_75t_SL U19804 (.Y(n23451),
	.A1(FE_OCPN27990_FE_OFN16132_sa03_5),
	.A2(n21726),
	.B(n23417));
   NAND2xp5_ASAP7_75t_L U19806 (.Y(n19457),
	.A(n19455),
	.B(n19454));
   NAND2xp33_ASAP7_75t_SL U19807 (.Y(n19455),
	.A(n19451),
	.B(n19452));
   NOR2xp33_ASAP7_75t_L U19808 (.Y(n21746),
	.A(FE_OCPN27393_sa03_0),
	.B(n18035));
   NAND2xp33_ASAP7_75t_SRAM U19809 (.Y(n18035),
	.A(n21295),
	.B(n18034));
   NAND3xp33_ASAP7_75t_R U19810 (.Y(n19449),
	.A(FE_OCPN28001_n21310),
	.B(n21708),
	.C(FE_OCPN29349_FE_OCPN27405_sa03_4));
   NOR2x1_ASAP7_75t_SL U19811 (.Y(n21714),
	.A(n21279),
	.B(n18888));
   NAND3xp33_ASAP7_75t_SL U19812 (.Y(n18888),
	.A(n21064),
	.B(n18892),
	.C(n18887));
   NAND3xp33_ASAP7_75t_L U19814 (.Y(n23943),
	.A(n17991),
	.B(n17990),
	.C(n18887));
   NOR2xp33_ASAP7_75t_SRAM U19815 (.Y(n17991),
	.A(n18904),
	.B(n21023));
   NOR2xp33_ASAP7_75t_SRAM U19816 (.Y(n17990),
	.A(FE_OCPN27628_n23455),
	.B(n21502));
   NOR2x1_ASAP7_75t_SL U19817 (.Y(n22873),
	.A(FE_OFN27058_n22094),
	.B(FE_OCPN27503_n20195));
   NOR2xp33_ASAP7_75t_SL U19818 (.Y(n22876),
	.A(FE_OCPN29318_n25524),
	.B(n20952));
   NOR2x1_ASAP7_75t_SL U19819 (.Y(n22906),
	.A(n19253),
	.B(n19252));
   NAND3xp33_ASAP7_75t_L U19820 (.Y(n19253),
	.A(n19249),
	.B(n19248),
	.C(n19256));
   OAI21xp5_ASAP7_75t_SL U19821 (.Y(n23015),
	.A1(FE_OFN28832_n19789),
	.A2(n23982),
	.B(n19662));
   NAND3xp33_ASAP7_75t_SRAM U19822 (.Y(n21175),
	.A(FE_OCPN29542_n21151),
	.B(n21166),
	.C(FE_OCPN29396_n19149));
   NAND2xp5_ASAP7_75t_L U19823 (.Y(n21165),
	.A(FE_OFN28522_n17261),
	.B(n18770));
   NAND2xp5_ASAP7_75t_R U19824 (.Y(n21173),
	.A(n21169),
	.B(n21170));
   OAI21xp5_ASAP7_75t_L U19827 (.Y(n21477),
	.A1(FE_OCPN28270_n17237),
	.A2(FE_OFN26172_n19609),
	.B(n21155));
   NAND2xp33_ASAP7_75t_SRAM U19828 (.Y(n21478),
	.A(n21474),
	.B(n21473));
   NAND2xp33_ASAP7_75t_SRAM U19829 (.Y(n21484),
	.A(n21483),
	.B(n21482));
   NAND2xp33_ASAP7_75t_R U19830 (.Y(n18779),
	.A(n18775),
	.B(n19123));
   NOR2xp33_ASAP7_75t_SRAM U19831 (.Y(n18775),
	.A(FE_OCPN28021_n21445),
	.B(n18776));
   NAND3xp33_ASAP7_75t_SL U19832 (.Y(n19848),
	.A(n24085),
	.B(n18759),
	.C(n18765));
   NOR3xp33_ASAP7_75t_SRAM U19833 (.Y(n18758),
	.A(n18757),
	.B(n21439),
	.C(FE_OFN28958_n17261));
   NAND2xp5_ASAP7_75t_R U19835 (.Y(n19094),
	.A(n21154),
	.B(FE_OCPN27819_n17245));
   OAI21xp33_ASAP7_75t_L U19836 (.Y(n18627),
	.A1(FE_OCPN27908_FE_OFN16156_sa00_2),
	.A2(n21473),
	.B(n19603));
   NOR2x1_ASAP7_75t_L U19837 (.Y(n17082),
	.A(n16992),
	.B(n20527));
   OAI21xp33_ASAP7_75t_R U19838 (.Y(n19381),
	.A1(FE_OCPN28202_n16991),
	.A2(FE_OCPN5143_n19361),
	.B(n18940));
   NOR2xp33_ASAP7_75t_L U19840 (.Y(n17144),
	.A(FE_OCPN5143_n19361),
	.B(FE_OCPN28202_n16991));
   OAI222xp33_ASAP7_75t_SL U19841 (.Y(n17152),
	.A1(FE_OFN28809_n),
	.A2(n20513),
	.B1(FE_OCPN27761_n16977),
	.B2(n20513),
	.C1(FE_OFN16319_n20527),
	.C2(n20513));
   NOR2x1_ASAP7_75t_L U19842 (.Y(n19256),
	.A(FE_OFN26033_n20197),
	.B(n20973));
   NOR2x1_ASAP7_75t_L U19843 (.Y(n20973),
	.A(n20962),
	.B(FE_OCPN27919_n20155));
   NOR2x1_ASAP7_75t_SL U19846 (.Y(n20952),
	.A(FE_OCPN27919_n20155),
	.B(FE_OFN28800_n22526));
   OAI21xp5_ASAP7_75t_L U19847 (.Y(n25525),
	.A1(FE_OCPN27919_n20155),
	.A2(FE_OCPN27574_n20196),
	.B(n22892));
   NOR2x1_ASAP7_75t_L U19848 (.Y(n25296),
	.A(FE_OCPN27624_n26971),
	.B(n17780));
   OAI21xp33_ASAP7_75t_L U19849 (.Y(n20162),
	.A1(FE_OCPN27566_FE_OFN16138_sa02_5),
	.A2(FE_OCPN29423_n26970),
	.B(n22112));
   NOR2x1_ASAP7_75t_L U19850 (.Y(n22084),
	.A(n20136),
	.B(n22539));
   NOR3xp33_ASAP7_75t_SL U19852 (.Y(n20969),
	.A(n20199),
	.B(n25523),
	.C(FE_OCPN27424_n22560));
   NOR3xp33_ASAP7_75t_SL U19853 (.Y(n22878),
	.A(n20211),
	.B(n20995),
	.C(n26972));
   NAND2xp5_ASAP7_75t_L U19858 (.Y(n20205),
	.A(n20127),
	.B(n22075));
   NOR2xp33_ASAP7_75t_SL U19859 (.Y(n20987),
	.A(FE_OCPN27624_n26971),
	.B(n22083));
   NOR2xp33_ASAP7_75t_L U19860 (.Y(n25274),
	.A(n20973),
	.B(n20987));
   OAI22xp33_ASAP7_75t_R U19861 (.Y(n25275),
	.A1(FE_PSN8330_n17761),
	.A2(n20985),
	.B1(FE_OFN28844_FE_OCPN27570_n17791),
	.B2(n20985));
   NAND3xp33_ASAP7_75t_SRAM U19862 (.Y(n25276),
	.A(n20214),
	.B(n22110),
	.C(n20213));
   NOR2x1p5_ASAP7_75t_SL U19864 (.Y(n25297),
	.A(FE_OFN28800_n22526),
	.B(n22083));
   NOR2x1_ASAP7_75t_SL U19865 (.Y(n20194),
	.A(FE_OCPN27573_n20196),
	.B(n22083));
   NOR2x1_ASAP7_75t_L U19866 (.Y(n22872),
	.A(n20962),
	.B(FE_OFN27058_n22094));
   NOR2xp33_ASAP7_75t_SL U19867 (.Y(n22557),
	.A(FE_OFN28897_n20132),
	.B(n26972));
   NOR2x1p5_ASAP7_75t_L U19868 (.Y(n22871),
	.A(n22083),
	.B(n20195));
   NAND3xp33_ASAP7_75t_SL U19869 (.Y(n22067),
	.A(n17761),
	.B(FE_OFN28844_FE_OCPN27570_n17791),
	.C(FE_OFN27202_n));
   NAND3xp33_ASAP7_75t_SL U19870 (.Y(n22115),
	.A(FE_OFN41_n20971),
	.B(n20970),
	.C(n20969));
   NAND2xp5_ASAP7_75t_SL U19871 (.Y(n20970),
	.A(n20968),
	.B(n20967));
   NAND2xp5_ASAP7_75t_L U19872 (.Y(n20967),
	.A(n20966),
	.B(n20963));
   NAND2xp5_ASAP7_75t_L U19873 (.Y(n20968),
	.A(n20964),
	.B(n20963));
   NAND2xp33_ASAP7_75t_R U19874 (.Y(n22101),
	.A(n22096),
	.B(n22098));
   NAND2xp33_ASAP7_75t_SRAM U19875 (.Y(n22100),
	.A(n22099),
	.B(n22098));
   NOR2x1_ASAP7_75t_L U19876 (.Y(n20152),
	.A(FE_OFN28961_n17744),
	.B(n20195));
   NOR2xp33_ASAP7_75t_SL U19877 (.Y(n22111),
	.A(n22109),
	.B(n22108));
   NAND3xp33_ASAP7_75t_SL U19878 (.Y(n22108),
	.A(n22107),
	.B(n22106),
	.C(n22105));
   NAND2xp5_ASAP7_75t_SL U19879 (.Y(n22104),
	.A(n22093),
	.B(n22092));
   NAND2xp5_ASAP7_75t_L U19880 (.Y(n22092),
	.A(n22091),
	.B(n22090));
   NAND2xp5_ASAP7_75t_L U19881 (.Y(n22093),
	.A(n22087),
	.B(n22090));
   NOR2xp33_ASAP7_75t_L U19882 (.Y(n22091),
	.A(n22089),
	.B(n22088));
   NAND2xp5_ASAP7_75t_L U19883 (.Y(n22103),
	.A(n19264),
	.B(n17808));
   OA21x2_ASAP7_75t_SRAM U19884 (.Y(n19265),
	.A1(FE_OFN28730_FE_OCPN28416_sa02_3),
	.A2(n20961),
	.B(n22065));
   NOR3xp33_ASAP7_75t_L U19885 (.Y(n22560),
	.A(FE_OFN29148_n),
	.B(FE_OFN29102_FE_OCPN27261_sa02_0),
	.C(FE_OCPN27624_n26971));
   NAND2xp33_ASAP7_75t_L U19886 (.Y(n19268),
	.A(FE_OFN152_n20170),
	.B(n19265));
   NOR2xp67_ASAP7_75t_L U19888 (.Y(n22074),
	.A(n22900),
	.B(n20952));
   NAND2xp5_ASAP7_75t_SL U19889 (.Y(n18278),
	.A(n17068),
	.B(n18254));
   NOR2x1_ASAP7_75t_SL U19890 (.Y(n17068),
	.A(n18919),
	.B(n25991));
   NAND2xp5_ASAP7_75t_SL U19891 (.Y(n18275),
	.A(n17064),
	.B(n17162));
   NOR2xp33_ASAP7_75t_SL U19892 (.Y(n17064),
	.A(FE_OFN16220_n25219),
	.B(n19429));
   NAND2xp5_ASAP7_75t_L U19893 (.Y(n18279),
	.A(n17120),
	.B(FE_OFN28913_n18247));
   NOR2xp33_ASAP7_75t_L U19894 (.Y(n17120),
	.A(n18283),
	.B(n25990));
   NAND2xp5_ASAP7_75t_SL U19895 (.Y(n19433),
	.A(n19428),
	.B(n20492));
   NOR2xp33_ASAP7_75t_SL U19896 (.Y(n19428),
	.A(n20522),
	.B(n25996));
   NOR3xp33_ASAP7_75t_L U19897 (.Y(n19434),
	.A(FE_OCPN5143_n19361),
	.B(FE_OCPN29369_n16982),
	.C(FE_OFN29243_n17065));
   NAND2xp5_ASAP7_75t_L U19898 (.Y(n19422),
	.A(n19418),
	.B(n19419));
   NOR3x1_ASAP7_75t_SL U19899 (.Y(n19435),
	.A(FE_OCPN29340_n17079),
	.B(FE_OFN28809_n),
	.C(FE_OCPN29544_n20527));
   NOR2x1_ASAP7_75t_SL U19900 (.Y(n25227),
	.A(n19430),
	.B(n18267));
   NOR3x1_ASAP7_75t_SL U19901 (.Y(n18269),
	.A(n18932),
	.B(FE_OFN16181_sa13_5),
	.C(n16992));
   NOR2xp33_ASAP7_75t_SL U19902 (.Y(n18268),
	.A(n17045),
	.B(n18922));
   NOR2x1p5_ASAP7_75t_R U19903 (.Y(n19410),
	.A(n20527),
	.B(FE_OCPN28202_n16991));
   OAI222xp33_ASAP7_75t_SL U19905 (.Y(n19431),
	.A1(FE_OFN29173_n),
	.A2(n18921),
	.B1(FE_OCPN28137_n17170),
	.B2(n18921),
	.C1(FE_OCPN27761_n16977),
	.C2(n18921));
   NOR2xp33_ASAP7_75t_SRAM U19906 (.Y(n18956),
	.A(FE_OFN16162_n25869),
	.B(n18954));
   INVx1_ASAP7_75t_L U19907 (.Y(n18955),
	.A(n18286));
   NOR2x1p5_ASAP7_75t_SL U19908 (.Y(n17171),
	.A(FE_OFN28738_n16989),
	.B(FE_OCPN27836_n16976));
   NOR2xp33_ASAP7_75t_L U19909 (.Y(n17123),
	.A(n25869),
	.B(n18279));
   NOR2xp33_ASAP7_75t_L U19910 (.Y(n17124),
	.A(FE_OFN29234_n16996),
	.B(n18279));
   OAI21xp5_ASAP7_75t_SL U19911 (.Y(n17129),
	.A1(n18932),
	.A2(FE_OCPN29490_n17001),
	.B(n17034));
   NAND3xp33_ASAP7_75t_SL U19912 (.Y(n17128),
	.A(n17088),
	.B(n18263),
	.C(n18939));
   NAND3xp33_ASAP7_75t_SL U19913 (.Y(n20507),
	.A(n17132),
	.B(n27090),
	.C(n17131));
   NAND3x1_ASAP7_75t_SL U19914 (.Y(n20506),
	.A(n25285),
	.B(n25221),
	.C(n17009));
   NOR3x1_ASAP7_75t_SL U19915 (.Y(n17009),
	.A(n17008),
	.B(n18919),
	.C(n25990));
   OAI222xp33_ASAP7_75t_R U19917 (.Y(n18260),
	.A1(FE_OFN16445_sa13_1),
	.A2(n17171),
	.B1(FE_OFN29074_n17170),
	.B2(n17171),
	.C1(FE_OCPN27902_n20514),
	.C2(n17171));
   NOR2xp33_ASAP7_75t_L U19918 (.Y(n18261),
	.A(FE_OCPN28189_n20491),
	.B(FE_OCPN27589_n25987));
   NOR2x1_ASAP7_75t_SL U19919 (.Y(n21023),
	.A(FE_OCPN27675_n17986),
	.B(n21706));
   NOR2xp33_ASAP7_75t_SL U19921 (.Y(n21513),
	.A(FE_OFN29109_n),
	.B(n19489));
   NAND2xp5_ASAP7_75t_SL U19922 (.Y(n21509),
	.A(n21022),
	.B(n21709));
   NAND2xp33_ASAP7_75t_L U19923 (.Y(n21020),
	.A(n21019),
	.B(n21018));
   NAND2xp33_ASAP7_75t_L U19924 (.Y(n21021),
	.A(n21016),
	.B(n21018));
   NAND3x1_ASAP7_75t_SL U19925 (.Y(n18024),
	.A(n18018),
	.B(n18017),
	.C(n18871));
   NOR2xp67_ASAP7_75t_L U19926 (.Y(n21505),
	.A(FE_OFN28997_sa03_4),
	.B(n17997));
   NAND2xp5_ASAP7_75t_L U19927 (.Y(n17997),
	.A(FE_OCPN28001_n21310),
	.B(n21708));
   NOR2x1_ASAP7_75t_L U19928 (.Y(n21502),
	.A(FE_OFN27133_n21725),
	.B(FE_OFN28588_n21048));
   NAND2xp5_ASAP7_75t_L U19929 (.Y(n21503),
	.A(n18026),
	.B(n21035));
   NAND2xp33_ASAP7_75t_SRAM U19930 (.Y(n18025),
	.A(n21719),
	.B(n21718));
   NOR2x1_ASAP7_75t_L U19932 (.Y(n21296),
	.A(n23457),
	.B(FE_OFN26581_n21317));
   NOR2x1_ASAP7_75t_L U19933 (.Y(n19478),
	.A(FE_OCPN28184_n18020),
	.B(n21012));
   NOR3xp33_ASAP7_75t_SL U19934 (.Y(n19689),
	.A(n19765),
	.B(n21894),
	.C(n17190));
   NAND2x1_ASAP7_75t_SL U19935 (.Y(n19686),
	.A(n23121),
	.B(FE_OCPN5153_n23127));
   NAND2xp5_ASAP7_75t_SL U19936 (.Y(n23028),
	.A(FE_OFN130_sa10_5),
	.B(n16577));
   NAND3x1_ASAP7_75t_L U19937 (.Y(n19789),
	.A(FE_OCPN28053_sa10_1),
	.B(FE_OCPN28145_n16535),
	.C(FE_OFN28749_n));
   NAND2xp33_ASAP7_75t_SRAM U19939 (.Y(n19668),
	.A(FE_OFN28807_n24944),
	.B(n16542));
   NAND2xp5_ASAP7_75t_R U19940 (.Y(n17209),
	.A(n17208),
	.B(n17207));
   NAND2xp33_ASAP7_75t_R U19941 (.Y(n17207),
	.A(n17206),
	.B(n17205));
   NAND2xp33_ASAP7_75t_R U19942 (.Y(n17208),
	.A(n17204),
	.B(n17205));
   INVxp33_ASAP7_75t_SRAM U19943 (.Y(n17206),
	.A(n23148));
   INVx1_ASAP7_75t_L U19945 (.Y(n17217),
	.A(n16653));
   NAND2xp33_ASAP7_75t_L U19946 (.Y(n16623),
	.A(n16622),
	.B(n16621));
   NOR2x1_ASAP7_75t_SL U19948 (.Y(n19663),
	.A(n23982),
	.B(n23036));
   NOR3xp33_ASAP7_75t_SL U19949 (.Y(n19765),
	.A(FE_OFN25956_n16575),
	.B(FE_OFN27196_n),
	.C(n16647));
   NAND2xp33_ASAP7_75t_R U19950 (.Y(n21910),
	.A(n21905),
	.B(n21907));
   NOR2xp33_ASAP7_75t_SRAM U19951 (.Y(n21905),
	.A(n21903),
	.B(n21906));
   INVxp33_ASAP7_75t_SRAM U19952 (.Y(n21903),
	.A(n21902));
   NAND2xp33_ASAP7_75t_SL U19953 (.Y(n21909),
	.A(n21908),
	.B(n21907));
   NOR2xp33_ASAP7_75t_SRAM U19954 (.Y(n21908),
	.A(n23035),
	.B(n21906));
   NAND2xp33_ASAP7_75t_SRAM U19955 (.Y(n19768),
	.A(n17223),
	.B(n24955));
   NOR3xp33_ASAP7_75t_SRAM U19956 (.Y(n24951),
	.A(n24726),
	.B(n19774),
	.C(n16640));
   NOR2xp33_ASAP7_75t_L U19957 (.Y(n24949),
	.A(n23131),
	.B(FE_OFN29154_n19753));
   NOR2x1_ASAP7_75t_SL U19958 (.Y(n19672),
	.A(n23982),
	.B(n16648));
   NAND2xp5_ASAP7_75t_SRAM U19960 (.Y(n23151),
	.A(n23150),
	.B(n23149));
   NAND2xp5_ASAP7_75t_SRAM U19961 (.Y(n23152),
	.A(n23147),
	.B(n23149));
   NAND2xp5_ASAP7_75t_SL U19964 (.Y(n23128),
	.A(n23148),
	.B(n23980));
   NOR3xp33_ASAP7_75t_SL U19965 (.Y(n21899),
	.A(n16556),
	.B(FE_OFN28749_n),
	.C(n23981));
   INVx1_ASAP7_75t_L U19966 (.Y(n19641),
	.A(n19789));
   NAND3xp33_ASAP7_75t_SL U19967 (.Y(n19788),
	.A(n17216),
	.B(n19630),
	.C(FE_OFN29255_n));
   NOR2x1_ASAP7_75t_SL U19968 (.Y(n17226),
	.A(FE_OCPN28358_n21899),
	.B(n16549));
   NAND2xp5_ASAP7_75t_SL U19969 (.Y(n16549),
	.A(n16632),
	.B(n17200));
   NOR3xp33_ASAP7_75t_SRAM U19970 (.Y(n17210),
	.A(n19672),
	.B(n16640),
	.C(n19670));
   NOR3x1_ASAP7_75t_SL U19971 (.Y(n19687),
	.A(n16592),
	.B(n19672),
	.C(n16633));
   NAND3xp33_ASAP7_75t_L U19972 (.Y(n16592),
	.A(n17217),
	.B(n16582),
	.C(n24739));
   NOR2xp33_ASAP7_75t_L U19973 (.Y(n16572),
	.A(FE_OCPN27900_n23949),
	.B(n23119));
   NAND3xp33_ASAP7_75t_SRAM U19974 (.Y(n24952),
	.A(n17194),
	.B(n19769),
	.C(n16663));
   NAND3xp33_ASAP7_75t_L U19975 (.Y(n24941),
	.A(n19647),
	.B(n19646),
	.C(n17197));
   NOR2xp33_ASAP7_75t_L U19976 (.Y(n19118),
	.A(n17275),
	.B(FE_OCPN27968_n21154));
   OAI21xp33_ASAP7_75t_SRAM U19977 (.Y(n19138),
	.A1(FE_OFN26172_n19609),
	.A2(n17275),
	.B(n18756));
   NAND2xp5_ASAP7_75t_SL U19978 (.Y(n22623),
	.A(n22166),
	.B(n25104));
   NAND2xp5_ASAP7_75t_SL U19979 (.Y(n18369),
	.A(n20456),
	.B(n18360));
   NAND2xp33_ASAP7_75t_SRAM U19980 (.Y(n19035),
	.A(n22125),
	.B(n18483));
   NAND2xp33_ASAP7_75t_L U19981 (.Y(n18372),
	.A(n18392),
	.B(FE_PSN8333_n18478));
   NAND2xp33_ASAP7_75t_SRAM U19982 (.Y(n22146),
	.A(FE_OCPN28057_n17603),
	.B(FE_OFN25917_n21591));
   NAND2xp5_ASAP7_75t_R U19983 (.Y(n24792),
	.A(n22151),
	.B(n24127));
   NOR2x1_ASAP7_75t_L U19984 (.Y(n22152),
	.A(FE_OCPN27829_n25102),
	.B(FE_OCPN27428_n26027));
   NOR2x1_ASAP7_75t_L U19985 (.Y(n22159),
	.A(FE_OCPN27829_n25102),
	.B(n18473));
   NAND3xp33_ASAP7_75t_SL U19986 (.Y(n22163),
	.A(n21584),
	.B(n18471),
	.C(n17619));
   NOR2x1_ASAP7_75t_L U19987 (.Y(n22161),
	.A(FE_OCPN28027_n22125),
	.B(n18473));
   NAND2xp33_ASAP7_75t_L U19988 (.Y(n18475),
	.A(n17606),
	.B(n22125));
   NAND2xp5_ASAP7_75t_L U19989 (.Y(n22166),
	.A(n21607),
	.B(n24780));
   NAND3xp33_ASAP7_75t_SL U19990 (.Y(n22144),
	.A(n19047),
	.B(n19046),
	.C(n19045));
   NOR2xp33_ASAP7_75t_SL U19991 (.Y(n17645),
	.A(FE_PSN8270_n26027),
	.B(FE_OFN25901_n22133));
   NAND3xp33_ASAP7_75t_SL U19993 (.Y(n20446),
	.A(n19046),
	.B(n22643),
	.C(n17617));
   NOR2xp33_ASAP7_75t_L U19994 (.Y(n17617),
	.A(n17616),
	.B(n20450));
   NOR2x1_ASAP7_75t_L U19996 (.Y(n20456),
	.A(n26029),
	.B(n22159));
   INVxp33_ASAP7_75t_SRAM U19997 (.Y(n20455),
	.A(n21586));
   NAND2xp5_ASAP7_75t_L U19998 (.Y(n18478),
	.A(n22125),
	.B(FE_OFN25917_n21591));
   NAND2x1_ASAP7_75t_SL U19999 (.Y(n19198),
	.A(n21847),
	.B(n21362));
   NAND2xp5_ASAP7_75t_L U20000 (.Y(n19210),
	.A(n21366),
	.B(n17453));
   NAND3xp33_ASAP7_75t_SL U20002 (.Y(n17500),
	.A(n24567),
	.B(n23356),
	.C(n23256));
   NOR3xp33_ASAP7_75t_L U20003 (.Y(n17502),
	.A(n23262),
	.B(n21422),
	.C(FE_OFN28627_n21377));
   NAND2xp33_ASAP7_75t_L U20004 (.Y(n23269),
	.A(n19162),
	.B(FE_OCPN5021_n17446));
   NAND3xp33_ASAP7_75t_L U20005 (.Y(n18759),
	.A(n17254),
	.B(FE_OFN28835_n),
	.C(FE_OFN28744_FE_OCPN27908));
   NOR2xp33_ASAP7_75t_R U20007 (.Y(n19850),
	.A(FE_OCPN27703_n19847),
	.B(n24087));
   NAND2x1p5_ASAP7_75t_SL U20008 (.Y(n19844),
	.A(n19591),
	.B(n19132));
   NOR2xp33_ASAP7_75t_SL U20009 (.Y(n21450),
	.A(n19839),
	.B(n19838));
   NOR2x1_ASAP7_75t_SL U20010 (.Y(n21438),
	.A(FE_OFN29062_n18651),
	.B(n17275));
   NOR3x1_ASAP7_75t_SL U20011 (.Y(n21439),
	.A(n17298),
	.B(FE_OCPN29396_n19149),
	.C(FE_OFN26651_n19573));
   OAI22xp5_ASAP7_75t_L U20012 (.Y(n19833),
	.A1(FE_OCPN28389_n21479),
	.A2(n26099),
	.B1(FE_OFN16216_n19573),
	.B2(n26099));
   NOR2xp33_ASAP7_75t_L U20013 (.Y(n19831),
	.A(FE_OFN28958_n17261),
	.B(n19593));
   NAND2xp5_ASAP7_75t_SL U20014 (.Y(n17262),
	.A(FE_OCPN29260_sa00_5),
	.B(n17248));
   NOR3xp33_ASAP7_75t_SL U20016 (.Y(n19813),
	.A(FE_OCPN29292_n18640),
	.B(FE_OCPN27818_n17267),
	.C(FE_OCPN27951_n19098));
   NAND3xp33_ASAP7_75t_L U20017 (.Y(n18635),
	.A(FE_OCPN27500_n19834),
	.B(FE_PSN8282_n21154),
	.C(FE_OFN29172_sa00_4));
   NOR2xp33_ASAP7_75t_SL U20018 (.Y(n21162),
	.A(n18634),
	.B(n18633));
   NAND2xp33_ASAP7_75t_L U20019 (.Y(n18633),
	.A(n18632),
	.B(n19595));
   NAND3x1_ASAP7_75t_L U20020 (.Y(n21858),
	.A(n17447),
	.B(FE_OCPN27903_n19223),
	.C(n17473));
   NOR2xp33_ASAP7_75t_L U20021 (.Y(n21846),
	.A(n21823),
	.B(n21822));
   AND2x2_ASAP7_75t_SL U20022 (.Y(n21378),
	.A(n21412),
	.B(n21411));
   NAND2xp5_ASAP7_75t_SL U20023 (.Y(n21837),
	.A(n23259),
	.B(n21851));
   NAND2xp33_ASAP7_75t_SL U20024 (.Y(n21836),
	.A(n17445),
	.B(n17446));
   NOR2xp33_ASAP7_75t_SL U20025 (.Y(n21833),
	.A(FE_PSN8303_n19222),
	.B(n22500));
   NAND2x1_ASAP7_75t_SL U20026 (.Y(n21838),
	.A(n19164),
	.B(n17468));
   NAND3x1_ASAP7_75t_SL U20027 (.Y(n21363),
	.A(n21858),
	.B(n23357),
	.C(n23259));
   NOR2x1_ASAP7_75t_SL U20028 (.Y(n21821),
	.A(FE_OFN28570_n19172),
	.B(FE_OFN29033_FE_OCPN27414_n23359));
   NOR2xp33_ASAP7_75t_L U20029 (.Y(n24546),
	.A(FE_OCPN27313_n21845),
	.B(FE_OFN28508_sa11_0));
   NOR2xp33_ASAP7_75t_L U20030 (.Y(n22510),
	.A(n21406),
	.B(n21356));
   OAI21xp5_ASAP7_75t_L U20031 (.Y(n21356),
	.A1(FE_OCPN28006_n17454),
	.A2(n21355),
	.B(n21428));
   NOR2xp67_ASAP7_75t_L U20032 (.Y(n22514),
	.A(n21422),
	.B(n21395));
   NOR2xp67_ASAP7_75t_L U20033 (.Y(n22509),
	.A(FE_OCPN27807_n23375),
	.B(n21369));
   NAND2xp33_ASAP7_75t_L U20034 (.Y(n21369),
	.A(n21856),
	.B(n21851));
   NAND2xp5_ASAP7_75t_L U20035 (.Y(n21848),
	.A(n21856),
	.B(n21858));
   NAND2x1_ASAP7_75t_SL U20036 (.Y(n21411),
	.A(FE_PSN8310_n17473),
	.B(n21349));
   O2A1O1Ixp33_ASAP7_75t_SL U20037 (.Y(n21410),
	.A1(FE_OFN29061_n22505),
	.A2(n19162),
	.B(FE_OCPN5021_n17446),
	.C(n21352));
   NAND2xp33_ASAP7_75t_SL U20038 (.Y(n19214),
	.A(FE_OFN28811_n19170),
	.B(FE_OFN28874_FE_OCPN27551_sa11_4));
   NAND2x1_ASAP7_75t_SL U20039 (.Y(n22511),
	.A(n23250),
	.B(n21383));
   NAND3xp33_ASAP7_75t_L U20040 (.Y(n25792),
	.A(n17446),
	.B(FE_OCPN27241_sa11_1),
	.C(n17473));
   NAND2xp33_ASAP7_75t_SRAM U20041 (.Y(n24711),
	.A(n21824),
	.B(n21411));
   NAND2x1_ASAP7_75t_SL U20042 (.Y(n23402),
	.A(n21833),
	.B(n19228));
   NOR2x1_ASAP7_75t_SL U20043 (.Y(n19228),
	.A(n21363),
	.B(n19227));
   NAND3xp33_ASAP7_75t_SL U20044 (.Y(n19227),
	.A(n23268),
	.B(n23249),
	.C(n19226));
   NOR2xp33_ASAP7_75t_L U20045 (.Y(n19226),
	.A(n23374),
	.B(n21377));
   NAND2xp5_ASAP7_75t_SL U20046 (.Y(n24544),
	.A(n26064),
	.B(n23254));
   NAND2xp33_ASAP7_75t_SL U20047 (.Y(n23394),
	.A(n21847),
	.B(n21367));
   NAND2xp33_ASAP7_75t_SRAM U20048 (.Y(n21367),
	.A(n21366),
	.B(n21365));
   NAND2xp5_ASAP7_75t_SL U20049 (.Y(n23373),
	.A(n21398),
	.B(n21397));
   NAND3xp33_ASAP7_75t_L U20050 (.Y(n23272),
	.A(n24567),
	.B(n17458),
	.C(n21859));
   NAND2xp5_ASAP7_75t_L U20051 (.Y(n17462),
	.A(n21394),
	.B(n23378));
   NAND2xp5_ASAP7_75t_SL U20052 (.Y(n23391),
	.A(n19171),
	.B(n17447));
   NAND2xp5_ASAP7_75t_L U20053 (.Y(n21398),
	.A(n19191),
	.B(n19190));
   NAND2xp5_ASAP7_75t_L U20054 (.Y(n19190),
	.A(n19189),
	.B(n19188));
   NAND2xp5_ASAP7_75t_R U20055 (.Y(n19191),
	.A(n19187),
	.B(n19188));
   NOR2x1_ASAP7_75t_SL U20057 (.Y(n19200),
	.A(FE_OCPN27757_n21819),
	.B(FE_OCPN28447_n23392));
   NOR2x1_ASAP7_75t_L U20058 (.Y(n18452),
	.A(n18362),
	.B(n20421));
   NAND3xp33_ASAP7_75t_SL U20059 (.Y(n18459),
	.A(n20476),
	.B(FE_OCPN28172_n20449),
	.C(n20453));
   NAND2x1p5_ASAP7_75t_SL U20060 (.Y(n18352),
	.A(n17601),
	.B(n18379));
   NOR3xp33_ASAP7_75t_SL U20061 (.Y(n25083),
	.A(n18352),
	.B(n17618),
	.C(n18381));
   NOR2x1_ASAP7_75t_L U20062 (.Y(n21590),
	.A(n20428),
	.B(n20429));
   NOR2x1_ASAP7_75t_L U20064 (.Y(n21676),
	.A(n23838),
	.B(n23677));
   NOR2x1_ASAP7_75t_L U20065 (.Y(n23811),
	.A(n21224),
	.B(n23740));
   NOR2x1_ASAP7_75t_L U20066 (.Y(n23809),
	.A(n20653),
	.B(n23792));
   AND3x1_ASAP7_75t_SL U20067 (.Y(n18575),
	.A(n25188),
	.B(n18573),
	.C(n18572));
   NOR2xp67_ASAP7_75t_SL U20068 (.Y(n18572),
	.A(n23831),
	.B(n21232));
   NAND2x1p5_ASAP7_75t_L U20069 (.Y(n20766),
	.A(n18159),
	.B(FE_OCPN27947_n18177));
   NOR2xp33_ASAP7_75t_SRAM U20072 (.Y(n20769),
	.A(n18162),
	.B(FE_OFN29241_n22811));
   NOR3xp33_ASAP7_75t_SL U20073 (.Y(n23189),
	.A(n20775),
	.B(n22821),
	.C(n26870));
   NAND2x1_ASAP7_75t_L U20074 (.Y(n21779),
	.A(n22270),
	.B(n20751));
   NOR3xp33_ASAP7_75t_L U20075 (.Y(n20751),
	.A(n20750),
	.B(n21804),
	.C(n20749));
   NAND2xp33_ASAP7_75t_L U20076 (.Y(n20750),
	.A(FE_OCPN28016_n21124),
	.B(FE_OFN28939_n21129));
   INVxp67_ASAP7_75t_L U20077 (.Y(n20740),
	.A(n20737));
   OAI21xp33_ASAP7_75t_L U20078 (.Y(n20749),
	.A1(FE_OCPN29305_n23302),
	.A2(n23303),
	.B(n20723));
   NAND3xp33_ASAP7_75t_R U20079 (.Y(n21103),
	.A(FE_PSN8320_n18176),
	.B(n18162),
	.C(FE_OCPN27979_FE_OFN16147_sa22_1));
   NAND2x1p5_ASAP7_75t_SL U20080 (.Y(n21105),
	.A(FE_OFN27173_n),
	.B(FE_OCPN27721_n23336));
   OAI22xp33_ASAP7_75t_SRAM U20081 (.Y(n20759),
	.A1(n18159),
	.A2(n20720),
	.B1(FE_OCPN29557_n18161),
	.B2(n20720));
   AND3x1_ASAP7_75t_SL U20082 (.Y(n20709),
	.A(n23174),
	.B(n20707),
	.C(n22285));
   NOR3xp33_ASAP7_75t_L U20083 (.Y(n20707),
	.A(n21115),
	.B(n20706),
	.C(n23300));
   NAND2x1p5_ASAP7_75t_SL U20085 (.Y(n22311),
	.A(n18159),
	.B(n18162));
   NOR2xp33_ASAP7_75t_SL U20087 (.Y(n20746),
	.A(FE_OFN26548_n18206),
	.B(n18178));
   NAND2x1_ASAP7_75t_SL U20088 (.Y(n22281),
	.A(n20766),
	.B(n23182));
   NAND2xp33_ASAP7_75t_R U20089 (.Y(n21110),
	.A(n21106),
	.B(n21108));
   NOR2x1_ASAP7_75t_L U20090 (.Y(n21085),
	.A(FE_OFN29238_n22811),
	.B(n18217));
   NOR2xp33_ASAP7_75t_L U20091 (.Y(n21771),
	.A(FE_OFN25987_n23322),
	.B(FE_OCPN27719_n23306));
   NOR2xp33_ASAP7_75t_R U20093 (.Y(n20706),
	.A(FE_OCPN29305_n23302),
	.B(n23303));
   NAND2xp5_ASAP7_75t_SL U20094 (.Y(n24692),
	.A(n23329),
	.B(n20773));
   NOR2xp33_ASAP7_75t_SRAM U20095 (.Y(n18168),
	.A(FE_RN_0_0),
	.B(n18217));
   NOR2x1p5_ASAP7_75t_SL U20096 (.Y(n23322),
	.A(n18160),
	.B(n18174));
   INVxp67_ASAP7_75t_L U20097 (.Y(n18160),
	.A(FE_OCPN29269_sa22_1));
   NOR3xp33_ASAP7_75t_SL U20098 (.Y(n18232),
	.A(n18230),
	.B(n22309),
	.C(n18229));
   NAND2xp33_ASAP7_75t_SRAM U20099 (.Y(n18211),
	.A(n18200),
	.B(n18203));
   NAND2xp33_ASAP7_75t_R U20100 (.Y(n18203),
	.A(n18202),
	.B(n18201));
   NOR3x1_ASAP7_75t_SL U20101 (.Y(n22827),
	.A(n18178),
	.B(FE_OCPN27521_n18163),
	.C(FE_OFN29080_n22310));
   NOR2x1p5_ASAP7_75t_L U20103 (.Y(n21801),
	.A(n22277),
	.B(n18187));
   NAND2x1_ASAP7_75t_SL U20104 (.Y(n18187),
	.A(n18216),
	.B(n23329));
   NAND3xp33_ASAP7_75t_L U20105 (.Y(n21119),
	.A(n23336),
	.B(n18176),
	.C(FE_OCPN29269_sa22_1));
   NOR3xp33_ASAP7_75t_L U20106 (.Y(n24705),
	.A(n18195),
	.B(n21130),
	.C(n23168));
   OAI21xp33_ASAP7_75t_SRAM U20107 (.Y(n18195),
	.A1(FE_OCPN29478_n23306),
	.A2(FE_OFN25987_n23322),
	.B(n22272));
   NAND2x1p5_ASAP7_75t_SL U20108 (.Y(n22320),
	.A(n21801),
	.B(n21800));
   NOR3x1_ASAP7_75t_SL U20109 (.Y(n21800),
	.A(n21799),
	.B(n23297),
	.C(n21798));
   NAND2xp33_ASAP7_75t_R U20110 (.Y(n21796),
	.A(n21795),
	.B(n23328));
   NOR2xp33_ASAP7_75t_SRAM U20111 (.Y(n21795),
	.A(n22828),
	.B(FE_OFN29195_n22850));
   NAND2xp33_ASAP7_75t_R U20112 (.Y(n21797),
	.A(n21794),
	.B(n23328));
   NOR2xp33_ASAP7_75t_SRAM U20113 (.Y(n21794),
	.A(n21793),
	.B(FE_OFN29195_n22850));
   NOR2x1_ASAP7_75t_SL U20114 (.Y(n21804),
	.A(FE_OCPN27673_n18163),
	.B(n23312));
   NOR3x1_ASAP7_75t_SL U20116 (.Y(n21130),
	.A(n21785),
	.B(FE_OFN55_sa22_5),
	.C(n18186));
   NAND2xp5_ASAP7_75t_SL U20119 (.Y(n25632),
	.A(n21655),
	.B(n25189));
   NOR2x1_ASAP7_75t_L U20120 (.Y(n20685),
	.A(FE_OFN29021_sa20_3),
	.B(FE_OCPN28257_n23689));
   NAND2xp33_ASAP7_75t_SRAM U20121 (.Y(n21249),
	.A(n18599),
	.B(n21247));
   NAND2xp33_ASAP7_75t_R U20122 (.Y(n21248),
	.A(n21242),
	.B(n21247));
   NAND2xp33_ASAP7_75t_SL U20123 (.Y(n21244),
	.A(n21243),
	.B(n23715));
   NAND2xp33_ASAP7_75t_R U20124 (.Y(n21245),
	.A(n21242),
	.B(n23715));
   NAND2xp33_ASAP7_75t_L U20125 (.Y(n21227),
	.A(n21226),
	.B(FE_OCPN27531_n21643));
   NOR2xp33_ASAP7_75t_SRAM U20126 (.Y(n21226),
	.A(FE_OCPN27606_n23869),
	.B(n21224));
   NAND2xp33_ASAP7_75t_L U20127 (.Y(n21228),
	.A(n21223),
	.B(FE_OCPN27531_n21643));
   NOR2xp33_ASAP7_75t_R U20128 (.Y(n21223),
	.A(n18583),
	.B(n21224));
   NOR2xp33_ASAP7_75t_L U20129 (.Y(n21230),
	.A(n23831),
	.B(n23884));
   NOR2xp33_ASAP7_75t_R U20130 (.Y(n23778),
	.A(FE_OFN28868_FE_OCPN27715_n23875),
	.B(n23840));
   NOR2x1_ASAP7_75t_L U20131 (.Y(n21204),
	.A(FE_OFN26150_n21253),
	.B(n21674));
   NOR2xp33_ASAP7_75t_R U20132 (.Y(n23839),
	.A(FE_OCPN27606_n23869),
	.B(n23840));
   NOR3xp33_ASAP7_75t_SL U20133 (.Y(n21643),
	.A(n23837),
	.B(n18522),
	.C(n18582));
   NAND3xp33_ASAP7_75t_SL U20134 (.Y(n21638),
	.A(FE_OFN28988_n18597),
	.B(n21195),
	.C(FE_OCPN27633_sa20_5));
   NOR3xp33_ASAP7_75t_SL U20135 (.Y(n21238),
	.A(n18596),
	.B(FE_OFN28510_n21215),
	.C(n21256));
   NAND2xp5_ASAP7_75t_SL U20137 (.Y(n18594),
	.A(n18593),
	.B(n18592));
   NAND2xp5_ASAP7_75t_SL U20138 (.Y(n18592),
	.A(n18591),
	.B(n18590));
   NOR2xp33_ASAP7_75t_L U20139 (.Y(n21673),
	.A(FE_OCPN27633_sa20_5),
	.B(n23688));
   NOR2xp33_ASAP7_75t_L U20140 (.Y(n21685),
	.A(FE_OFN29251_n18536),
	.B(n23865));
   NOR2xp67_ASAP7_75t_L U20141 (.Y(n23835),
	.A(FE_OFN28815_n18523),
	.B(n23677));
   NAND2xp33_ASAP7_75t_L U20142 (.Y(n21688),
	.A(n21687),
	.B(n21686));
   NOR2xp33_ASAP7_75t_SL U20143 (.Y(n21687),
	.A(n23855),
	.B(n23865));
   NOR3x2_ASAP7_75t_SL U20144 (.Y(n23830),
	.A(n18534),
	.B(FE_OFN29246_n),
	.C(n18582));
   NOR2x1_ASAP7_75t_L U20145 (.Y(n18585),
	.A(FE_OCPN27606_n23869),
	.B(n23830));
   NOR3x1_ASAP7_75t_SL U20147 (.Y(n23718),
	.A(n21641),
	.B(n21682),
	.C(n21640));
   OAI21xp33_ASAP7_75t_SRAM U20148 (.Y(n21640),
	.A1(FE_OFN28815_n18523),
	.A2(n21639),
	.B(n23721));
   NAND3xp33_ASAP7_75t_SL U20149 (.Y(n21641),
	.A(n21638),
	.B(n21637),
	.C(n21636));
   NOR2x1_ASAP7_75t_L U20150 (.Y(n23779),
	.A(n21648),
	.B(n20675));
   NAND2xp33_ASAP7_75t_L U20151 (.Y(n23715),
	.A(n18522),
	.B(n18540));
   NOR2xp33_ASAP7_75t_R U20152 (.Y(n23706),
	.A(n18583),
	.B(n23792));
   AND3x1_ASAP7_75t_SL U20153 (.Y(n23705),
	.A(n23703),
	.B(n23702),
	.C(n23781));
   NOR3xp33_ASAP7_75t_SL U20154 (.Y(n23703),
	.A(n23691),
	.B(n23740),
	.C(n23690));
   NAND2xp5_ASAP7_75t_L U20155 (.Y(n23702),
	.A(n23697),
	.B(n23696));
   NAND2xp5_ASAP7_75t_L U20156 (.Y(n23678),
	.A(n20617),
	.B(FE_OFN28869_FE_OCPN27715_n23875));
   NAND2xp5_ASAP7_75t_SL U20157 (.Y(n21654),
	.A(n23852),
	.B(n18564));
   NOR2xp33_ASAP7_75t_L U20159 (.Y(n21649),
	.A(FE_OCPN28353_n18534),
	.B(n18530));
   NOR3x1_ASAP7_75t_SL U20160 (.Y(n23776),
	.A(n21693),
	.B(n23863),
	.C(n23680));
   NOR2xp33_ASAP7_75t_R U20161 (.Y(n23874),
	.A(FE_OCPN27606_n23869),
	.B(n23885));
   NOR2xp33_ASAP7_75t_L U20162 (.Y(n23876),
	.A(FE_OFN28868_FE_OCPN27715_n23875),
	.B(n23885));
   NOR2x1_ASAP7_75t_L U20164 (.Y(n23856),
	.A(FE_OFN16385_n18525),
	.B(FE_OFN31_sa20_0));
   NAND2x1_ASAP7_75t_L U20166 (.Y(n20644),
	.A(n20636),
	.B(n18580));
   NAND3xp33_ASAP7_75t_L U20167 (.Y(n16919),
	.A(FE_OFN28999_n16923),
	.B(FE_OCPN27555_n16422),
	.C(FE_OCPN29391_FE_OFN29162_sa33_2));
   NOR2xp33_ASAP7_75t_L U20168 (.Y(n18421),
	.A(FE_OFN25960_n),
	.B(FE_OCPN27460_n16913));
   NOR2x1_ASAP7_75t_SL U20169 (.Y(n18416),
	.A(n24613),
	.B(n16709));
   NAND2xp5_ASAP7_75t_SL U20170 (.Y(n16709),
	.A(n16924),
	.B(n23528));
   OAI21xp33_ASAP7_75t_L U20171 (.Y(n16469),
	.A1(FE_OCPN27460_n16913),
	.A2(FE_OCPN27604_n16421),
	.B(n16855));
   NOR2x1_ASAP7_75t_L U20173 (.Y(n16959),
	.A(n18109),
	.B(n16871));
   NAND3xp33_ASAP7_75t_SL U20174 (.Y(n17426),
	.A(n16881),
	.B(n16880),
	.C(n18424));
   NAND2xp5_ASAP7_75t_SL U20175 (.Y(n16879),
	.A(n16877),
	.B(FE_OFN27089_n23558));
   NOR2x1p5_ASAP7_75t_L U20176 (.Y(n18430),
	.A(n16457),
	.B(n16436));
   OAI21xp33_ASAP7_75t_L U20177 (.Y(n16912),
	.A1(FE_OCPN28127_n16872),
	.A2(FE_OCPN27604_n16421),
	.B(n16726));
   NOR2xp33_ASAP7_75t_R U20178 (.Y(n16956),
	.A(FE_OFN29101_n16418),
	.B(n18145));
   NOR2xp33_ASAP7_75t_R U20179 (.Y(n16954),
	.A(n16430),
	.B(n18145));
   NAND2xp33_ASAP7_75t_SRAM U20181 (.Y(n17432),
	.A(n16418),
	.B(n16430));
   NAND2xp33_ASAP7_75t_SL U20182 (.Y(n16961),
	.A(n16959),
	.B(n18406));
   NAND2xp33_ASAP7_75t_L U20183 (.Y(n16957),
	.A(n16956),
	.B(n16955));
   NAND3xp33_ASAP7_75t_SL U20184 (.Y(n16965),
	.A(n24614),
	.B(n16884),
	.C(n16883));
   NAND2xp33_ASAP7_75t_SRAM U20185 (.Y(n16884),
	.A(n16427),
	.B(FE_OCPN27782_n16873));
   NOR3xp33_ASAP7_75t_SL U20186 (.Y(n16883),
	.A(n18146),
	.B(n16882),
	.C(n17426));
   NOR3x1_ASAP7_75t_L U20188 (.Y(n16472),
	.A(n16676),
	.B(FE_OFN26055_n),
	.C(FE_OCPN27666_n17418));
   NOR3xp33_ASAP7_75t_SL U20189 (.Y(n18109),
	.A(FE_OCPN27604_n16421),
	.B(FE_OCPN29391_FE_OFN29162_sa33_2),
	.C(FE_OCPN27539_n16875));
   NOR3xp33_ASAP7_75t_L U20190 (.Y(n18124),
	.A(n16911),
	.B(n23530),
	.C(n24617));
   NOR2xp67_ASAP7_75t_L U20191 (.Y(n17412),
	.A(FE_OCPN28322_n18141),
	.B(n16718));
   NOR2x1_ASAP7_75t_L U20192 (.Y(n16720),
	.A(n16457),
	.B(FE_OCPN27460_n16913));
   OAI21xp33_ASAP7_75t_L U20193 (.Y(n16837),
	.A1(n16429),
	.A2(FE_OCPN27460_n16913),
	.B(n16690));
   NAND2xp33_ASAP7_75t_R U20194 (.Y(n16690),
	.A(n16689),
	.B(n16424));
   NAND2x1_ASAP7_75t_SL U20195 (.Y(n18129),
	.A(FE_OCPN27546_sa33_4),
	.B(n18108));
   NAND3xp33_ASAP7_75t_L U20196 (.Y(n23532),
	.A(FE_PSN8337_n16909),
	.B(n16946),
	.C(FE_OCPN29487_FE_OFN28694_sa33_4));
   NAND3xp33_ASAP7_75t_SL U20197 (.Y(n23533),
	.A(n16424),
	.B(n16417),
	.C(FE_OFN28771_n));
   OAI21xp33_ASAP7_75t_SRAM U20198 (.Y(n23531),
	.A1(FE_OCPN27555_n16422),
	.A2(n16852),
	.B(FE_OFN28999_n16923));
   NAND2x1p5_ASAP7_75t_SL U20199 (.Y(n16676),
	.A(FE_OFN28694_sa33_4),
	.B(FE_OCPN27568_sa33_3));
   NOR3xp33_ASAP7_75t_R U20200 (.Y(n16908),
	.A(n16913),
	.B(FE_OFN25938_sa33_3),
	.C(n16677));
   NOR2xp33_ASAP7_75t_L U20201 (.Y(n18149),
	.A(n16838),
	.B(n16837));
   NOR2x1_ASAP7_75t_L U20202 (.Y(n16840),
	.A(n18415),
	.B(n18433));
   NOR2x1_ASAP7_75t_SL U20203 (.Y(n23529),
	.A(n24328),
	.B(n16859));
   NAND3xp33_ASAP7_75t_L U20204 (.Y(n16880),
	.A(n16831),
	.B(n16417),
	.C(FE_OFN25938_sa33_3));
   NOR2x1_ASAP7_75t_L U20205 (.Y(n20934),
	.A(n25095),
	.B(n25096));
   NOR2x1_ASAP7_75t_SL U20206 (.Y(n18988),
	.A(FE_OCPN27288_n25091),
	.B(n25092));
   NOR3xp33_ASAP7_75t_SL U20207 (.Y(n22943),
	.A(n18985),
	.B(n20224),
	.C(n25711));
   NOR2x1_ASAP7_75t_L U20208 (.Y(n20257),
	.A(n22925),
	.B(n23490));
   NAND2xp33_ASAP7_75t_SL U20210 (.Y(n18994),
	.A(n18991),
	.B(FE_OFN16250_n26165));
   NOR2xp33_ASAP7_75t_L U20211 (.Y(n18991),
	.A(FE_OFN27056_n22995),
	.B(n22033));
   NAND2xp33_ASAP7_75t_L U20212 (.Y(n18993),
	.A(n18992),
	.B(FE_OFN16250_n26165));
   NOR3xp33_ASAP7_75t_SL U20215 (.Y(n22945),
	.A(FE_OCPN27956_n),
	.B(FE_OFN29189_sa23_0),
	.C(n22951));
   NOR2xp33_ASAP7_75t_L U20216 (.Y(n20232),
	.A(FE_OCPN28381_n26660),
	.B(n20928));
   NAND3xp33_ASAP7_75t_SL U20217 (.Y(n19331),
	.A(n18986),
	.B(n26146),
	.C(n26147));
   NOR2xp33_ASAP7_75t_SL U20218 (.Y(n18986),
	.A(n26149),
	.B(n26148));
   NOR2xp33_ASAP7_75t_L U20219 (.Y(n19015),
	.A(FE_OFN28580_n23491),
	.B(n22935));
   NAND2xp33_ASAP7_75t_SL U20220 (.Y(n19305),
	.A(n19304),
	.B(n19303));
   NAND2xp33_ASAP7_75t_SL U20221 (.Y(n22045),
	.A(n19338),
	.B(n20930));
   OAI21xp5_ASAP7_75t_SL U20222 (.Y(n22041),
	.A1(FE_OCPN27288_n25091),
	.A2(FE_OFN28841_n22980),
	.B(n19001));
   NAND3xp33_ASAP7_75t_SL U20223 (.Y(n22035),
	.A(n22985),
	.B(n19315),
	.C(n20234));
   NAND2xp5_ASAP7_75t_L U20224 (.Y(n19315),
	.A(n19312),
	.B(n19311));
   NAND2xp5_ASAP7_75t_L U20225 (.Y(n19311),
	.A(n19310),
	.B(n19309));
   NAND2xp5_ASAP7_75t_L U20226 (.Y(n19312),
	.A(n22952),
	.B(n19309));
   NOR2xp33_ASAP7_75t_SL U20227 (.Y(n22034),
	.A(n22010),
	.B(n20235));
   NOR2xp33_ASAP7_75t_SL U20228 (.Y(n20923),
	.A(FE_OFN28752_n),
	.B(n23472));
   OA21x2_ASAP7_75t_L U20229 (.Y(n20243),
	.A1(n22010),
	.A2(FE_OFN25889_n20913),
	.B(n20242));
   NOR2xp33_ASAP7_75t_SRAM U20230 (.Y(n20244),
	.A(FE_OFN29026_n20911),
	.B(n23472));
   NOR3xp33_ASAP7_75t_SL U20231 (.Y(n22004),
	.A(n22010),
	.B(FE_OCPN29374_FE_OFN29191_sa23_2),
	.C(FE_OCPN28107_n23504));
   AND3x1_ASAP7_75t_SL U20232 (.Y(n22025),
	.A(n22022),
	.B(n22021),
	.C(n22020));
   NOR2x1_ASAP7_75t_L U20233 (.Y(n19343),
	.A(n22033),
	.B(n23472));
   NOR3xp33_ASAP7_75t_L U20234 (.Y(n23000),
	.A(n22999),
	.B(n22998),
	.C(n22997));
   NOR2x1_ASAP7_75t_SL U20235 (.Y(n19344),
	.A(n23473),
	.B(n20909));
   NAND2xp33_ASAP7_75t_L U20236 (.Y(n22592),
	.A(n21534),
	.B(n23104));
   NAND2xp5_ASAP7_75t_L U20237 (.Y(n21540),
	.A(FE_OFN16208_n23101),
	.B(n17382));
   NOR3x1_ASAP7_75t_SL U20238 (.Y(n24389),
	.A(n22459),
	.B(n23087),
	.C(FE_OFN78_n22457));
   NOR2xp33_ASAP7_75t_SRAM U20240 (.Y(n26997),
	.A(n22597),
	.B(n22584));
   NAND2xp5_ASAP7_75t_L U20241 (.Y(n18687),
	.A(n18683),
	.B(FE_OFN26054_sa01_3));
   NAND2xp5_ASAP7_75t_L U20242 (.Y(n18683),
	.A(n18682),
	.B(n23078));
   NOR3x1_ASAP7_75t_L U20243 (.Y(n21552),
	.A(n18686),
	.B(n18714),
	.C(n20378));
   NAND2xp5_ASAP7_75t_SL U20244 (.Y(n18686),
	.A(n22431),
	.B(n20389));
   NOR2xp33_ASAP7_75t_SRAM U20245 (.Y(n18688),
	.A(FE_OFN29254_n),
	.B(n22584));
   OAI21xp5_ASAP7_75t_L U20246 (.Y(n22459),
	.A1(FE_OFN27072_n18671),
	.A2(n17318),
	.B(n18713));
   NOR2x1_ASAP7_75t_L U20247 (.Y(n25062),
	.A(n20391),
	.B(n20378));
   NAND2xp5_ASAP7_75t_SL U20248 (.Y(n17351),
	.A(n17350),
	.B(n17349));
   NAND2xp5_ASAP7_75t_L U20249 (.Y(n17349),
	.A(n17348),
	.B(n22198));
   NAND2xp5_ASAP7_75t_L U20250 (.Y(n17350),
	.A(n17347),
	.B(n22198));
   NAND2xp5_ASAP7_75t_L U20251 (.Y(n22421),
	.A(FE_OFN28594_n26454),
	.B(FE_OFN29135_n21551));
   NAND2xp5_ASAP7_75t_L U20252 (.Y(n20366),
	.A(n22469),
	.B(n22458));
   NAND2xp33_ASAP7_75t_SRAM U20253 (.Y(n17366),
	.A(n17363),
	.B(n20361));
   NAND2xp33_ASAP7_75t_R U20254 (.Y(n17365),
	.A(n17364),
	.B(n20361));
   NAND2xp5_ASAP7_75t_R U20255 (.Y(n17362),
	.A(n17358),
	.B(n23088));
   NOR2x1_ASAP7_75t_SL U20256 (.Y(n21554),
	.A(n17391),
	.B(n17390));
   NAND2xp33_ASAP7_75t_L U20257 (.Y(n17325),
	.A(n17320),
	.B(n17322));
   NAND2x1p5_ASAP7_75t_L U20258 (.Y(n18685),
	.A(n17386),
	.B(FE_OFN29135_n21551));
   NAND2xp5_ASAP7_75t_L U20259 (.Y(n17339),
	.A(n17338),
	.B(n17337));
   NAND3xp33_ASAP7_75t_SL U20260 (.Y(n17355),
	.A(n22183),
	.B(n17334),
	.C(n22588));
   NOR3xp33_ASAP7_75t_SL U20261 (.Y(n22606),
	.A(n22600),
	.B(FE_OCPN28397_n23082),
	.C(n22599));
   NOR3xp33_ASAP7_75t_SRAM U20262 (.Y(n22604),
	.A(n22603),
	.B(n22602),
	.C(n22601));
   NOR2xp33_ASAP7_75t_L U20263 (.Y(n22590),
	.A(n23093),
	.B(n23092));
   NAND2xp5_ASAP7_75t_R U20264 (.Y(n22589),
	.A(n17385),
	.B(n17384));
   NAND2xp33_ASAP7_75t_R U20265 (.Y(n17384),
	.A(n22418),
	.B(n17369));
   NAND2xp33_ASAP7_75t_SRAM U20266 (.Y(n17385),
	.A(n22416),
	.B(n17369));
   NOR3xp33_ASAP7_75t_SL U20267 (.Y(n27010),
	.A(n22599),
	.B(n23076),
	.C(n23075));
   NAND2xp5_ASAP7_75t_SL U20268 (.Y(n21535),
	.A(FE_OFN26054_sa01_3),
	.B(n20404));
   NAND3x1_ASAP7_75t_SL U20269 (.Y(n22458),
	.A(FE_OCPN27887_n17331),
	.B(FE_OFN29135_n21551),
	.C(FE_OFN29254_n));
   NAND3xp33_ASAP7_75t_SL U20270 (.Y(n22414),
	.A(n17331),
	.B(n23059),
	.C(FE_OCPN8251_FE_OFN28672_sa01_2));
   NOR3xp33_ASAP7_75t_SL U20271 (.Y(n22433),
	.A(n23101),
	.B(FE_OCPN29429_FE_OFN16141_sa01_3),
	.C(n17389));
   NOR2x1_ASAP7_75t_L U20272 (.Y(n22431),
	.A(FE_OCPN28301_n22448),
	.B(n20387));
   NAND3xp33_ASAP7_75t_SL U20273 (.Y(n22453),
	.A(FE_OCPN29309_n26452),
	.B(n17375),
	.C(n17374));
   OAI21xp33_ASAP7_75t_L U20274 (.Y(n20369),
	.A1(n18667),
	.A2(n17318),
	.B(n18713));
   NOR2xp33_ASAP7_75t_SL U20275 (.Y(n20373),
	.A(n20371),
	.B(n21569));
   NOR2xp33_ASAP7_75t_SL U20277 (.Y(n17958),
	.A(FE_OFN28834_FE_OCPN28371_n17900),
	.B(n20784));
   NAND2xp33_ASAP7_75t_SL U20278 (.Y(n17960),
	.A(n17957),
	.B(n22735));
   NOR2xp33_ASAP7_75t_L U20279 (.Y(n17957),
	.A(n23587),
	.B(n20784));
   NOR2x1p5_ASAP7_75t_L U20280 (.Y(n19539),
	.A(FE_OFN27070_n),
	.B(FE_OCPN27253_n17923));
   NAND3xp33_ASAP7_75t_SL U20281 (.Y(n20562),
	.A(n25399),
	.B(n25398),
	.C(n23236));
   NAND3xp33_ASAP7_75t_L U20282 (.Y(n20543),
	.A(FE_OCPN28198_n22776),
	.B(FE_OCPN5137_n23600),
	.C(FE_OFN25907_sa12_2));
   NAND3xp33_ASAP7_75t_SL U20283 (.Y(n20584),
	.A(n19560),
	.B(n19559),
	.C(n23233));
   NAND2xp5_ASAP7_75t_L U20284 (.Y(n19560),
	.A(n19549),
	.B(n19548));
   NOR3xp33_ASAP7_75t_L U20285 (.Y(n19559),
	.A(n19551),
	.B(n20793),
	.C(n19550));
   NAND2xp33_ASAP7_75t_L U20286 (.Y(n19548),
	.A(n20546),
	.B(n19547));
   NOR2xp33_ASAP7_75t_L U20288 (.Y(n20598),
	.A(n23582),
	.B(n19511));
   NAND2xp5_ASAP7_75t_L U20289 (.Y(n19511),
	.A(n20543),
	.B(n22222));
   INVxp67_ASAP7_75t_R U20290 (.Y(n19510),
	.A(n25741));
   NAND3xp33_ASAP7_75t_SRAM U20291 (.Y(n17975),
	.A(n19540),
	.B(n20797),
	.C(n23617));
   NOR3xp33_ASAP7_75t_L U20292 (.Y(n17977),
	.A(n17939),
	.B(n23582),
	.C(n22233));
   NAND2xp5_ASAP7_75t_SL U20293 (.Y(n19534),
	.A(n17933),
	.B(n17932));
   NAND2xp5_ASAP7_75t_SL U20294 (.Y(n17933),
	.A(n17930),
	.B(n17931));
   NOR2xp33_ASAP7_75t_SL U20295 (.Y(n17930),
	.A(n17954),
	.B(n20556));
   NOR2xp33_ASAP7_75t_L U20296 (.Y(n17910),
	.A(n19539),
	.B(n20596));
   NOR2x1_ASAP7_75t_SL U20298 (.Y(n23206),
	.A(FE_OCPN27253_n17923),
	.B(FE_OCPN29324_n23216));
   NAND2xp5_ASAP7_75t_L U20300 (.Y(n22739),
	.A(n19561),
	.B(n23617));
   OAI21xp33_ASAP7_75t_SRAM U20301 (.Y(n22777),
	.A1(FE_OCPN28198_n22776),
	.A2(n24364),
	.B(FE_OCPN27729_n24362));
   NAND2x1_ASAP7_75t_SL U20302 (.Y(n22256),
	.A(n19539),
	.B(n23600));
   NOR2xp33_ASAP7_75t_R U20303 (.Y(n22746),
	.A(FE_OFN29075_n22745),
	.B(n25439));
   NAND2xp33_ASAP7_75t_L U20305 (.Y(n22748),
	.A(n22744),
	.B(n20814));
   NOR2xp33_ASAP7_75t_SRAM U20307 (.Y(n22245),
	.A(n25741),
	.B(n25439));
   AND2x2_ASAP7_75t_L U20308 (.Y(n23227),
	.A(n22244),
	.B(n23617));
   NAND2xp5_ASAP7_75t_SL U20309 (.Y(n22248),
	.A(n20597),
	.B(n20790));
   NAND3xp33_ASAP7_75t_SRAM U20310 (.Y(n20597),
	.A(FE_OCPN29477_sa12_5),
	.B(FE_OFN29075_n22745),
	.C(FE_OCPN27429_sa12_3));
   NAND2xp33_ASAP7_75t_SL U20311 (.Y(n22252),
	.A(n24367),
	.B(FE_OCPN27729_n24362));
   NOR2xp33_ASAP7_75t_L U20312 (.Y(n20602),
	.A(n20784),
	.B(n20583));
   NOR2x1_ASAP7_75t_L U20313 (.Y(n22730),
	.A(FE_OCPN27804_sa12_1),
	.B(n20805));
   NOR2xp33_ASAP7_75t_SRAM U20315 (.Y(n17942),
	.A(n22745),
	.B(n20583));
   NAND2xp33_ASAP7_75t_L U20316 (.Y(n22774),
	.A(n23612),
	.B(n19562));
   NOR2xp33_ASAP7_75t_SL U20317 (.Y(n19514),
	.A(n19502),
	.B(FE_OCPN29324_n23216));
   NOR2x1_ASAP7_75t_L U20318 (.Y(n22250),
	.A(n23602),
	.B(n17946));
   NAND3xp33_ASAP7_75t_SL U20319 (.Y(n17946),
	.A(n20558),
	.B(n20595),
	.C(n24585));
   NAND2xp5_ASAP7_75t_SL U20320 (.Y(n23583),
	.A(n22758),
	.B(n22759));
   NOR2x1_ASAP7_75t_SL U20321 (.Y(n23582),
	.A(n19502),
	.B(n20555));
   NAND2xp5_ASAP7_75t_L U20322 (.Y(n20813),
	.A(n22256),
	.B(n19503));
   NOR3xp33_ASAP7_75t_SL U20323 (.Y(n23618),
	.A(n23615),
	.B(n24589),
	.C(n23614));
   NAND3xp33_ASAP7_75t_SL U20324 (.Y(n23615),
	.A(n23610),
	.B(n23609),
	.C(n23608));
   NAND2xp5_ASAP7_75t_SL U20325 (.Y(n23610),
	.A(n23607),
	.B(n23606));
   NAND2xp33_ASAP7_75t_L U20326 (.Y(n23597),
	.A(n23594),
	.B(n23593));
   NAND2xp33_ASAP7_75t_R U20327 (.Y(n23593),
	.A(n23592),
	.B(FE_OFN85_n23588));
   NOR2xp33_ASAP7_75t_L U20328 (.Y(n23595),
	.A(FE_OFN26023_n20807),
	.B(n20806));
   NAND2xp33_ASAP7_75t_L U20329 (.Y(n22255),
	.A(n22254),
	.B(n22253));
   NAND2xp5_ASAP7_75t_L U20330 (.Y(n24363),
	.A(n22759),
	.B(n22779));
   NAND2xp5_ASAP7_75t_L U20332 (.Y(n23574),
	.A(n20785),
	.B(n22778));
   NAND2xp5_ASAP7_75t_L U20333 (.Y(n20805),
	.A(FE_OCPN28386_n17899),
	.B(n19546));
   NAND2xp33_ASAP7_75t_SL U20334 (.Y(n20802),
	.A(n20801),
	.B(n20800));
   NOR2xp33_ASAP7_75t_R U20335 (.Y(n17963),
	.A(n20796),
	.B(n22734));
   NAND2xp5_ASAP7_75t_SL U20336 (.Y(n20790),
	.A(FE_OCPN29492_sa12_4),
	.B(n20571));
   NAND3xp33_ASAP7_75t_SL U20337 (.Y(n20793),
	.A(n23612),
	.B(n20565),
	.C(n22722));
   NAND2xp5_ASAP7_75t_SL U20339 (.Y(n17921),
	.A(FE_OCPN29555_n20593),
	.B(n24367));
   INVx1_ASAP7_75t_L U20340 (.Y(n20785),
	.A(n23590));
   NAND2xp5_ASAP7_75t_L U20341 (.Y(n20558),
	.A(FE_OCPN5137_n23600),
	.B(n24364));
   OAI22x1_ASAP7_75t_L U20342 (.Y(n20789),
	.A1(FE_OFN25907_sa12_2),
	.A2(n23238),
	.B1(n23206),
	.B2(n23238));
   NOR2xp33_ASAP7_75t_R U20343 (.Y(n20585),
	.A(n23587),
	.B(n22734));
   OAI21xp33_ASAP7_75t_SL U20345 (.Y(n17585),
	.A1(n18832),
	.A2(FE_OCPN27420_n18794),
	.B(n18839));
   NOR2xp33_ASAP7_75t_L U20346 (.Y(n17587),
	.A(FE_OFN69_sa32_4),
	.B(n18320));
   NAND2x1p5_ASAP7_75t_SL U20347 (.Y(n17566),
	.A(FE_OFN16463_sa32_0),
	.B(FE_OFN26035_n));
   NOR2x1_ASAP7_75t_L U20348 (.Y(n18340),
	.A(n19926),
	.B(n17574));
   NAND2xp5_ASAP7_75t_L U20349 (.Y(n17574),
	.A(n18321),
	.B(n25025));
   NOR3xp33_ASAP7_75t_SL U20350 (.Y(n18341),
	.A(n18339),
	.B(n19936),
	.C(n18795));
   NAND2xp33_ASAP7_75t_SRAM U20351 (.Y(n18339),
	.A(n18336),
	.B(n18335));
   NAND3xp33_ASAP7_75t_SL U20352 (.Y(n18328),
	.A(n18851),
	.B(n18326),
	.C(n18325));
   NAND2xp33_ASAP7_75t_SRAM U20353 (.Y(n18326),
	.A(n18324),
	.B(n19940));
   NAND2xp5_ASAP7_75t_R U20354 (.Y(n18327),
	.A(n24646),
	.B(FE_OFN28965_n24869));
   NOR2x1_ASAP7_75t_SL U20355 (.Y(n18338),
	.A(n20096),
	.B(n19740));
   NOR3x1_ASAP7_75t_L U20356 (.Y(n19956),
	.A(n17558),
	.B(n17557),
	.C(n17556));
   NAND3xp33_ASAP7_75t_SL U20357 (.Y(n17558),
	.A(n17555),
	.B(n17713),
	.C(n24647));
   NOR2xp33_ASAP7_75t_L U20358 (.Y(n17555),
	.A(n18846),
	.B(n17571));
   NOR2x1_ASAP7_75t_SL U20359 (.Y(n19732),
	.A(FE_OCPN28423_n18836),
	.B(n18828));
   NAND2xp5_ASAP7_75t_R U20360 (.Y(n18805),
	.A(n24867),
	.B(n18306));
   NOR3xp33_ASAP7_75t_SL U20361 (.Y(n18814),
	.A(n18322),
	.B(n18830),
	.C(n20103));
   NAND2xp5_ASAP7_75t_L U20362 (.Y(n18322),
	.A(n22396),
	.B(n18320));
   NAND2xp5_ASAP7_75t_SL U20363 (.Y(n18793),
	.A(FE_OFN26035_n),
	.B(FE_OCPN27812_FE_OFN16463_sa32_0));
   NAND2xp33_ASAP7_75t_L U20364 (.Y(n17571),
	.A(n24867),
	.B(n20094));
   NAND2xp5_ASAP7_75t_L U20365 (.Y(n17700),
	.A(FE_OCPN29459_n),
	.B(n17529));
   NAND2xp5_ASAP7_75t_SL U20366 (.Y(n18330),
	.A(FE_OFN69_sa32_4),
	.B(n19712));
   NAND3xp33_ASAP7_75t_R U20367 (.Y(n22390),
	.A(n19938),
	.B(n19725),
	.C(FE_OFN69_sa32_4));
   NOR2x1_ASAP7_75t_SL U20368 (.Y(n22377),
	.A(n18841),
	.B(n19703));
   NOR2xp33_ASAP7_75t_L U20369 (.Y(n19743),
	.A(n20095),
	.B(FE_OCPN27490_n18798));
   NAND2xp5_ASAP7_75t_R U20370 (.Y(n18320),
	.A(n19725),
	.B(n19940));
   NOR2x1_ASAP7_75t_SL U20371 (.Y(n16763),
	.A(n16783),
	.B(FE_OCPN29307_FE_OFN25989_sa21_4));
   NOR3xp33_ASAP7_75t_L U20372 (.Y(n17876),
	.A(FE_OFN28820_n),
	.B(FE_OFN25989_sa21_4),
	.C(n16801));
   NOR2x1_ASAP7_75t_SL U20373 (.Y(n20304),
	.A(n23633),
	.B(n16785));
   NAND2xp33_ASAP7_75t_L U20374 (.Y(n16785),
	.A(n16784),
	.B(FE_OFN28985_sa21_5));
   NAND2xp33_ASAP7_75t_L U20375 (.Y(n16816),
	.A(n17838),
	.B(n16814));
   NAND2xp33_ASAP7_75t_R U20376 (.Y(n16821),
	.A(n16818),
	.B(n23662));
   NOR2xp33_ASAP7_75t_SRAM U20377 (.Y(n16818),
	.A(n16758),
	.B(n19890));
   NOR2x1_ASAP7_75t_L U20378 (.Y(n16808),
	.A(FE_OFN62_sa21_3),
	.B(n22329));
   NAND2xp5_ASAP7_75t_R U20380 (.Y(n16796),
	.A(FE_OFN27155_sa21_4),
	.B(n16795));
   NOR3xp33_ASAP7_75t_L U20382 (.Y(n17838),
	.A(n19896),
	.B(n22330),
	.C(n20345));
   NAND2xp33_ASAP7_75t_R U20384 (.Y(n17827),
	.A(n17825),
	.B(n17824));
   NOR2x1_ASAP7_75t_L U20385 (.Y(n17828),
	.A(FE_OCPN27508_n20339),
	.B(n19877));
   NOR2x1_ASAP7_75t_L U20386 (.Y(n20298),
	.A(FE_OCPN29294_n23925),
	.B(n24881));
   NAND3xp33_ASAP7_75t_L U20387 (.Y(n20333),
	.A(n19979),
	.B(n16757),
	.C(FE_OCPN27289_sa21_5));
   INVx1_ASAP7_75t_L U20388 (.Y(n19878),
	.A(n19875));
   NOR2x1_ASAP7_75t_L U20389 (.Y(n17872),
	.A(FE_OCPN27289_sa21_5),
	.B(n19981));
   NOR3x1_ASAP7_75t_SL U20390 (.Y(n22694),
	.A(FE_OCPN27246_n22663),
	.B(FE_OCPN27328_sa21_2),
	.C(FE_OCPN29418_n));
   NAND2x1_ASAP7_75t_SL U20391 (.Y(n20335),
	.A(n19897),
	.B(n22343));
   NOR2x1_ASAP7_75t_L U20392 (.Y(n19897),
	.A(n22658),
	.B(n19896));
   NAND2xp5_ASAP7_75t_SL U20393 (.Y(n17857),
	.A(n16815),
	.B(n17873));
   NOR3xp33_ASAP7_75t_SL U20394 (.Y(n16815),
	.A(n20004),
	.B(n23925),
	.C(n19871));
   NOR3x1_ASAP7_75t_SL U20395 (.Y(n20326),
	.A(n19866),
	.B(n24881),
	.C(FE_OCPN5079_n20287));
   O2A1O1Ixp33_ASAP7_75t_L U20396 (.Y(n19865),
	.A1(FE_OFN28778_FE_OCPN28352_n16748),
	.A2(FE_OFN27157_n23928),
	.B(FE_OCPN28299_n),
	.C(n25353));
   OAI22xp5_ASAP7_75t_L U20397 (.Y(n19863),
	.A1(n16757),
	.A2(FE_OFN28970_n19890),
	.B1(FE_OFN28529_n16774),
	.B2(FE_OFN28970_n19890));
   NAND2xp5_ASAP7_75t_SL U20398 (.Y(n22708),
	.A(FE_OCPN27774_n25351),
	.B(n19992));
   NAND2x1_ASAP7_75t_SL U20399 (.Y(n22355),
	.A(n20337),
	.B(n25350));
   NOR3x1_ASAP7_75t_SL U20400 (.Y(n20337),
	.A(n20336),
	.B(n20335),
	.C(n20334));
   NAND2xp5_ASAP7_75t_L U20401 (.Y(n20336),
	.A(n20333),
	.B(n20332));
   NOR2xp33_ASAP7_75t_SL U20403 (.Y(n20308),
	.A(n22675),
	.B(n22679));
   NAND2xp33_ASAP7_75t_SL U20404 (.Y(n20310),
	.A(n20306),
	.B(n20307));
   NOR2xp33_ASAP7_75t_SL U20405 (.Y(n20306),
	.A(FE_OCPN5126_sa21_2),
	.B(n22679));
   NOR2xp33_ASAP7_75t_L U20407 (.Y(n19892),
	.A(n17860),
	.B(FE_OFN27140_n20007));
   NAND2x1_ASAP7_75t_L U20408 (.Y(n22333),
	.A(FE_OCPN29414_n),
	.B(n19975));
   NAND2xp5_ASAP7_75t_R U20409 (.Y(n22340),
	.A(FE_OCPN27642_n16758),
	.B(FE_OFN16447_n16749));
   NOR2x1_ASAP7_75t_SL U20410 (.Y(n20003),
	.A(n16800),
	.B(n16799));
   NAND2xp5_ASAP7_75t_SL U20411 (.Y(n16799),
	.A(n23649),
	.B(n20324));
   NAND3xp33_ASAP7_75t_L U20412 (.Y(n16800),
	.A(n19988),
	.B(n20333),
	.C(n17828));
   NAND3x1_ASAP7_75t_SL U20413 (.Y(n20004),
	.A(FE_OFN29215_n24262),
	.B(n23625),
	.C(n22665));
   NAND3xp33_ASAP7_75t_SL U20415 (.Y(n16773),
	.A(n23650),
	.B(n19889),
	.C(n16772));
   NAND3xp33_ASAP7_75t_SL U20416 (.Y(n23659),
	.A(n23656),
	.B(n24918),
	.C(n24269));
   NAND2xp33_ASAP7_75t_SRAM U20417 (.Y(n23665),
	.A(n23660),
	.B(n23662));
   NAND3x1_ASAP7_75t_SL U20418 (.Y(n23658),
	.A(n22351),
	.B(n25355),
	.C(n22350));
   NOR2x1_ASAP7_75t_L U20420 (.Y(n19988),
	.A(n22330),
	.B(FE_OFN27163_n20304));
   NOR2xp33_ASAP7_75t_L U20421 (.Y(n19984),
	.A(FE_OFN16447_n16749),
	.B(n23925));
   NAND2xp5_ASAP7_75t_L U20422 (.Y(n19986),
	.A(n19985),
	.B(n19983));
   NOR2xp33_ASAP7_75t_L U20423 (.Y(n19985),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(n23925));
   NAND2xp5_ASAP7_75t_L U20424 (.Y(n20054),
	.A(n20841),
	.B(n16348));
   NAND2xp5_ASAP7_75t_L U20425 (.Y(n16349),
	.A(FE_OCPN27877_n21980),
	.B(n20028));
   NAND3xp33_ASAP7_75t_L U20426 (.Y(n21965),
	.A(n20882),
	.B(n24182),
	.C(n16373));
   NOR2xp33_ASAP7_75t_L U20427 (.Y(n16373),
	.A(n18072),
	.B(n18096));
   NAND3xp33_ASAP7_75t_SL U20428 (.Y(n16309),
	.A(FE_OFN29136_n),
	.B(FE_OFN28492_sa31_0),
	.C(FE_OFN29147_sa31_1));
   NAND2x1_ASAP7_75t_SL U20429 (.Y(n20076),
	.A(FE_OFN28753_sa31_2),
	.B(FE_OFN28492_sa31_0));
   NOR2xp33_ASAP7_75t_L U20430 (.Y(n20873),
	.A(n18072),
	.B(n16496));
   NOR2xp33_ASAP7_75t_SL U20431 (.Y(n20867),
	.A(n21989),
	.B(n25849));
   NOR2xp33_ASAP7_75t_SRAM U20432 (.Y(n20870),
	.A(n20868),
	.B(n25849));
   NAND2xp5_ASAP7_75t_SL U20433 (.Y(n18069),
	.A(n26291),
	.B(n16348));
   NAND3xp33_ASAP7_75t_SL U20434 (.Y(n21951),
	.A(n16502),
	.B(FE_OCPN27780_n20083),
	.C(n16501));
   NOR3xp33_ASAP7_75t_L U20435 (.Y(n16501),
	.A(n26409),
	.B(n20840),
	.C(n21988));
   NOR2xp33_ASAP7_75t_SL U20436 (.Y(n20885),
	.A(FE_OFN28808_n26291),
	.B(n21930));
   NAND2xp33_ASAP7_75t_L U20437 (.Y(n20883),
	.A(n20881),
	.B(n20880));
   NAND2xp33_ASAP7_75t_R U20438 (.Y(n20880),
	.A(n20879),
	.B(n20878));
   NOR2xp33_ASAP7_75t_SL U20439 (.Y(n20887),
	.A(FE_OFN29032_FE_OCPN27728_n21981),
	.B(n21930));
   NOR2xp33_ASAP7_75t_SL U20440 (.Y(n20857),
	.A(n16295),
	.B(n20858));
   NOR2xp33_ASAP7_75t_R U20441 (.Y(n20860),
	.A(n16299),
	.B(n20858));
   OAI21x1_ASAP7_75t_SL U20442 (.Y(n16391),
	.A1(n21981),
	.A2(FE_OCPN28314_n20842),
	.B(n18087));
   NAND2x1_ASAP7_75t_SL U20443 (.Y(n20856),
	.A(n16303),
	.B(n20050));
   NOR2xp33_ASAP7_75t_L U20445 (.Y(n16372),
	.A(n20854),
	.B(n20853));
   NOR2x1_ASAP7_75t_SL U20447 (.Y(n16513),
	.A(n21968),
	.B(n16358));
   OAI21xp33_ASAP7_75t_L U20448 (.Y(n16358),
	.A1(n20853),
	.A2(FE_OCPN28334_n16497),
	.B(n20054));
   NAND2x1_ASAP7_75t_L U20449 (.Y(n18068),
	.A(FE_OFN28710_n20841),
	.B(FE_OFN29032_FE_OCPN27728_n21981));
   NOR2xp33_ASAP7_75t_SL U20450 (.Y(n16359),
	.A(n20059),
	.B(FE_OCPN27786_n16490));
   NAND2xp33_ASAP7_75t_L U20451 (.Y(n20838),
	.A(FE_OFN16415_sa31_2),
	.B(n16345));
   NOR2xp33_ASAP7_75t_L U20452 (.Y(n18082),
	.A(n26402),
	.B(n20033));
   NOR3xp33_ASAP7_75t_L U20453 (.Y(n20849),
	.A(FE_OCPN27316_n25849),
	.B(n21982),
	.C(n16395));
   NOR3xp33_ASAP7_75t_L U20454 (.Y(n25846),
	.A(n20858),
	.B(n26290),
	.C(n18061));
   OAI21xp5_ASAP7_75t_SL U20455 (.Y(n20043),
	.A1(FE_OFN26060_sa31_4),
	.A2(n16350),
	.B(n20874));
   NAND2xp5_ASAP7_75t_L U20456 (.Y(n26298),
	.A(n16406),
	.B(n20838));
   NAND2xp33_ASAP7_75t_SL U20457 (.Y(n16515),
	.A(n21936),
	.B(n16331));
   NOR2x1_ASAP7_75t_L U20458 (.Y(n18071),
	.A(FE_OFN29047_n21980),
	.B(n16290));
   NAND2x1_ASAP7_75t_SL U20459 (.Y(n20858),
	.A(n16301),
	.B(n16502));
   NOR3xp33_ASAP7_75t_SL U20460 (.Y(n16301),
	.A(n16374),
	.B(n16516),
	.C(n16361));
   NAND2xp5_ASAP7_75t_SL U20461 (.Y(n16498),
	.A(n25316),
	.B(n20066));
   NAND2xp5_ASAP7_75t_L U20462 (.Y(n18088),
	.A(n21948),
	.B(n20856));
   NOR3x1_ASAP7_75t_SL U20463 (.Y(n19916),
	.A(n17575),
	.B(n19728),
	.C(n19704));
   NAND3x1_ASAP7_75t_SL U20464 (.Y(n17575),
	.A(n20100),
	.B(n18340),
	.C(n22377));
   NOR2xp33_ASAP7_75t_L U20465 (.Y(n19917),
	.A(FE_OFN28564_n18308),
	.B(n22370));
   NAND3xp33_ASAP7_75t_SRAM U20467 (.Y(n25230),
	.A(n25228),
	.B(n25290),
	.C(n25227));
   NAND2xp33_ASAP7_75t_SRAM U20468 (.Y(n25226),
	.A(n25222),
	.B(n25221));
   NAND2xp33_ASAP7_75t_SRAM U20470 (.Y(n24058),
	.A(n24057),
	.B(n24056));
   NOR2xp33_ASAP7_75t_SRAM U20471 (.Y(n24057),
	.A(FE_OCPN27729_n24362),
	.B(n24055));
   NOR3xp33_ASAP7_75t_SL U20472 (.Y(n24062),
	.A(n20560),
	.B(n20559),
	.C(n26599));
   NAND3xp33_ASAP7_75t_SL U20473 (.Y(n20560),
	.A(n20557),
	.B(n20595),
	.C(n23234));
   AND2x2_ASAP7_75t_L U20474 (.Y(n20557),
	.A(n20790),
	.B(n20795));
   NOR3xp33_ASAP7_75t_SL U20475 (.Y(n22670),
	.A(n19871),
	.B(n22330),
	.C(FE_OFN27163_n20304));
   NAND2xp5_ASAP7_75t_SL U20476 (.Y(n22665),
	.A(FE_OCPN27631_n16774),
	.B(FE_OCPN27642_n16758));
   NAND3xp33_ASAP7_75t_R U20477 (.Y(n22657),
	.A(n19979),
	.B(FE_OFN28981_n16767),
	.C(FE_OCPN27289_sa21_5));
   NAND2xp33_ASAP7_75t_SRAM U20478 (.Y(n17845),
	.A(FE_OFN28529_n16774),
	.B(n16771));
   NAND2xp5_ASAP7_75t_SL U20479 (.Y(n22658),
	.A(n22333),
	.B(n23650));
   NOR2xp33_ASAP7_75t_SRAM U20480 (.Y(n24676),
	.A(n26857),
	.B(FE_OCPN5099_n24677));
   NOR2xp33_ASAP7_75t_SRAM U20481 (.Y(n24680),
	.A(n24678),
	.B(FE_OCPN5099_n24677));
   NAND2xp33_ASAP7_75t_R U20482 (.Y(n23991),
	.A(n23988),
	.B(n23987));
   NAND2xp33_ASAP7_75t_R U20483 (.Y(n23987),
	.A(n23986),
	.B(n23985));
   NAND2xp33_ASAP7_75t_R U20484 (.Y(n23988),
	.A(n23984),
	.B(n23985));
   INVxp33_ASAP7_75t_L U20485 (.Y(n23985),
	.A(n23983));
   NOR3xp33_ASAP7_75t_SL U20486 (.Y(n24001),
	.A(n23999),
	.B(n23998),
	.C(n23997));
   OAI21xp33_ASAP7_75t_SRAM U20487 (.Y(n24002),
	.A1(n23996),
	.A2(n23995),
	.B(FE_OCPN27636_sa10_4));
   NOR2x1_ASAP7_75t_SL U20488 (.Y(n23044),
	.A(n16533),
	.B(n16610));
   NAND2x1_ASAP7_75t_SL U20489 (.Y(n23048),
	.A(n19659),
	.B(n19658));
   NAND2xp5_ASAP7_75t_L U20490 (.Y(n19658),
	.A(n19657),
	.B(n19656));
   NAND2xp33_ASAP7_75t_L U20492 (.Y(n23042),
	.A(n23037),
	.B(n23039));
   NAND2xp33_ASAP7_75t_L U20493 (.Y(n23041),
	.A(n23040),
	.B(n23039));
   NAND2xp33_ASAP7_75t_L U20495 (.Y(n18061),
	.A(n21932),
	.B(n16519));
   NAND2xp5_ASAP7_75t_SL U20496 (.Y(n25236),
	.A(n26620),
	.B(n26621));
   NAND2xp33_ASAP7_75t_R U20497 (.Y(n24162),
	.A(n24161),
	.B(n24160));
   NAND2xp33_ASAP7_75t_R U20498 (.Y(n24161),
	.A(n24158),
	.B(n24159));
   NAND2xp33_ASAP7_75t_R U20499 (.Y(n24160),
	.A(FE_OFN28479_sa13_2),
	.B(n24159));
   NAND2xp33_ASAP7_75t_L U20500 (.Y(n19378),
	.A(n17148),
	.B(n17147));
   NOR2xp33_ASAP7_75t_SRAM U20501 (.Y(n17148),
	.A(n18919),
	.B(n17144));
   NOR2xp33_ASAP7_75t_L U20502 (.Y(n17147),
	.A(n19364),
	.B(n19429));
   NOR2x1_ASAP7_75t_L U20503 (.Y(n18954),
	.A(n20527),
	.B(FE_OFN28583_n17001));
   NAND3xp33_ASAP7_75t_L U20504 (.Y(n17142),
	.A(n20514),
	.B(FE_OCPN29358_n17159),
	.C(FE_OFN16444_sa13_1));
   OAI21xp33_ASAP7_75t_L U20505 (.Y(n16508),
	.A1(FE_OFN28516_FE_OFN27192_sa31_2),
	.A2(n25317),
	.B(n20053));
   INVx1_ASAP7_75t_L U20506 (.Y(n16952),
	.A(n24296));
   NAND2xp5_ASAP7_75t_L U20507 (.Y(n16851),
	.A(n17416),
	.B(FE_PSN8337_n16909));
   NAND3xp33_ASAP7_75t_SL U20508 (.Y(n16850),
	.A(n16417),
	.B(n16479),
	.C(FE_OFN16430_sa33_3));
   NAND2xp5_ASAP7_75t_L U20509 (.Y(n17415),
	.A(n16924),
	.B(n16707));
   NAND2xp5_ASAP7_75t_SL U20510 (.Y(n16882),
	.A(n18445),
	.B(n16922));
   NOR2xp33_ASAP7_75t_L U20511 (.Y(n16868),
	.A(n24297),
	.B(n16937));
   NAND2x1_ASAP7_75t_SL U20512 (.Y(n16875),
	.A(FE_OFN29134_sa33_0),
	.B(FE_OFN28727_sa33_1));
   AND2x2_ASAP7_75t_SL U20513 (.Y(n18123),
	.A(n16886),
	.B(n16885));
   NAND2xp33_ASAP7_75t_SRAM U20514 (.Y(n16885),
	.A(n16418),
	.B(FE_OFN28999_n16923));
   NOR2xp67_ASAP7_75t_SL U20515 (.Y(n16886),
	.A(n17414),
	.B(n16965));
   NOR2x1_ASAP7_75t_SL U20516 (.Y(n16870),
	.A(n16853),
	.B(n16711));
   NAND3x1_ASAP7_75t_SL U20517 (.Y(n16711),
	.A(n18416),
	.B(n16725),
	.C(n16710));
   NOR2xp33_ASAP7_75t_L U20518 (.Y(n17407),
	.A(FE_OCPN28127_n16872),
	.B(n16874));
   NOR2xp33_ASAP7_75t_L U20519 (.Y(n17424),
	.A(FE_OCPN27460_n16913),
	.B(n16432));
   NAND2xp33_ASAP7_75t_SRAM U20520 (.Y(n16432),
	.A(FE_OFN25938_sa33_3),
	.B(FE_OCPN27544_sa33_4));
   NOR2x1p5_ASAP7_75t_L U20521 (.Y(n17405),
	.A(FE_OCPN27604_n16421),
	.B(FE_OFN26545_n16447));
   NOR2x1_ASAP7_75t_L U20522 (.Y(n16893),
	.A(n18433),
	.B(n16445));
   NAND2xp5_ASAP7_75t_L U20523 (.Y(n16445),
	.A(n16444),
	.B(n16855));
   NAND2xp33_ASAP7_75t_SRAM U20524 (.Y(n16444),
	.A(n17416),
	.B(n16854));
   NAND2x1_ASAP7_75t_L U20525 (.Y(n23528),
	.A(n17416),
	.B(n16430));
   NAND2xp33_ASAP7_75t_SRAM U20526 (.Y(n16896),
	.A(n16895),
	.B(n16894));
   OAI222xp33_ASAP7_75t_R U20528 (.Y(n14060),
	.A1(FE_OFN28769_n15478),
	.A2(n14041),
	.B1(n15514),
	.B2(n14041),
	.C1(FE_OFN27066_n13869),
	.C2(n14041));
   NAND2xp5_ASAP7_75t_R U20529 (.Y(n14059),
	.A(n14051),
	.B(n14050));
   NAND2xp33_ASAP7_75t_L U20530 (.Y(n14058),
	.A(n14057),
	.B(n14056));
   NAND3xp33_ASAP7_75t_L U20531 (.Y(n14078),
	.A(n14077),
	.B(n14076),
	.C(n14075));
   O2A1O1Ixp33_ASAP7_75t_SRAM U20532 (.Y(n14075),
	.A1(FE_OFN26091_n24663),
	.A2(n15694),
	.B(n14074),
	.C(n14073));
   NAND2xp33_ASAP7_75t_SL U20533 (.Y(n14076),
	.A(n14072),
	.B(n14071));
   NAND2xp33_ASAP7_75t_L U20534 (.Y(n14077),
	.A(n14067),
	.B(n14066));
   OAI22xp33_ASAP7_75t_SRAM U20535 (.Y(n14029),
	.A1(FE_OCPN27987_FE_OFN4_w3_22),
	.A2(n13889),
	.B1(FE_OFN25915_n15514),
	.B2(n13889));
   NAND2xp33_ASAP7_75t_R U20536 (.Y(n14039),
	.A(n14038),
	.B(n14037));
   NOR2xp33_ASAP7_75t_SRAM U20537 (.Y(n14038),
	.A(n15507),
	.B(n14036));
   NAND2xp33_ASAP7_75t_R U20538 (.Y(n14040),
	.A(n14035),
	.B(n14037));
   NAND3xp33_ASAP7_75t_SRAM U20539 (.Y(n14187),
	.A(FE_OFN28695_n),
	.B(n15859),
	.C(FE_OCPN27978_w3_3));
   OAI21xp33_ASAP7_75t_SRAM U20540 (.Y(n14189),
	.A1(n15870),
	.A2(n14831),
	.B(n14188));
   OAI21xp33_ASAP7_75t_L U20541 (.Y(n14191),
	.A1(n14410),
	.A2(n15861),
	.B(n14186));
   NAND2xp33_ASAP7_75t_SL U20542 (.Y(n13825),
	.A(n13824),
	.B(n13823));
   NAND2xp33_ASAP7_75t_L U20543 (.Y(n13823),
	.A(n13822),
	.B(n13821));
   NAND2xp33_ASAP7_75t_L U20544 (.Y(n13824),
	.A(n13819),
	.B(n13821));
   NOR2xp33_ASAP7_75t_SRAM U20545 (.Y(n13822),
	.A(n14159),
	.B(n13820));
   A2O1A1Ixp33_ASAP7_75t_L U20546 (.Y(n13855),
	.A1(FE_OFN29017_n15921),
	.A2(n14959),
	.B(n13854),
	.C(n14183));
   NAND3xp33_ASAP7_75t_SL U20547 (.Y(n13854),
	.A(n13853),
	.B(n13852),
	.C(n14612));
   NAND2xp33_ASAP7_75t_SL U20548 (.Y(n13852),
	.A(n13850),
	.B(n13849));
   OAI22xp33_ASAP7_75t_L U20549 (.Y(n13853),
	.A1(FE_OCPN28296_n15386),
	.A2(n13842),
	.B1(n14626),
	.B2(n13842));
   NAND2xp33_ASAP7_75t_L U20550 (.Y(n13857),
	.A(n13833),
	.B(n13832));
   NAND2xp33_ASAP7_75t_R U20551 (.Y(n13832),
	.A(n13831),
	.B(n13828));
   NAND2xp33_ASAP7_75t_L U20552 (.Y(n13833),
	.A(n13829),
	.B(n13828));
   NAND2xp33_ASAP7_75t_R U20553 (.Y(n13856),
	.A(n13840),
	.B(n13839));
   NAND2xp33_ASAP7_75t_SRAM U20554 (.Y(n13840),
	.A(n13836),
	.B(n13835));
   NAND2xp33_ASAP7_75t_SRAM U20555 (.Y(n13839),
	.A(n13838),
	.B(n13835));
   NAND2xp33_ASAP7_75t_SRAM U20556 (.Y(n14640),
	.A(n14941),
	.B(FE_PSN8271_n15924));
   INVxp33_ASAP7_75t_SRAM U20557 (.Y(n13815),
	.A(n16015));
   NOR2xp33_ASAP7_75t_L U20558 (.Y(n14959),
	.A(n15380),
	.B(n15375));
   NAND3xp33_ASAP7_75t_R U20559 (.Y(n14396),
	.A(n14395),
	.B(n15679),
	.C(n14394));
   OAI22xp33_ASAP7_75t_L U20560 (.Y(n14394),
	.A1(n15514),
	.A2(n14392),
	.B1(n14393),
	.B2(n14392));
   OAI22xp33_ASAP7_75t_SRAM U20561 (.Y(n14393),
	.A1(FE_OFN27082_n25377),
	.A2(n15480),
	.B1(FE_PSN8298_FE_OFN27151_n),
	.B2(n15480));
   NOR2xp33_ASAP7_75t_SRAM U20562 (.Y(n14397),
	.A(n13916),
	.B(FE_OCPN8264_n13890));
   NAND2xp33_ASAP7_75t_SL U20563 (.Y(n14390),
	.A(n14366),
	.B(n14365));
   NAND2xp33_ASAP7_75t_L U20564 (.Y(n14365),
	.A(n14364),
	.B(n14363));
   NAND2xp33_ASAP7_75t_L U20565 (.Y(n14366),
	.A(n14360),
	.B(n14363));
   NOR2xp33_ASAP7_75t_SRAM U20566 (.Y(n14364),
	.A(n14773),
	.B(n14362));
   NAND2xp33_ASAP7_75t_L U20567 (.Y(n14387),
	.A(n14386),
	.B(n14385));
   NAND3xp33_ASAP7_75t_SRAM U20568 (.Y(n14388),
	.A(n14382),
	.B(n15711),
	.C(n14381));
   NAND2xp33_ASAP7_75t_SRAM U20569 (.Y(n14386),
	.A(n15713),
	.B(n14383));
   NAND2xp33_ASAP7_75t_L U20570 (.Y(n14391),
	.A(n14356),
	.B(n14355));
   NAND2xp33_ASAP7_75t_SRAM U20571 (.Y(n14355),
	.A(n14354),
	.B(n14353));
   NAND2xp33_ASAP7_75t_R U20572 (.Y(n14356),
	.A(n14352),
	.B(n14353));
   NAND2xp33_ASAP7_75t_L U20573 (.Y(n14342),
	.A(n14332),
	.B(n14331));
   NAND2xp33_ASAP7_75t_SRAM U20574 (.Y(n14331),
	.A(n14330),
	.B(FE_OFN25981_n13868));
   NAND2xp33_ASAP7_75t_SRAM U20575 (.Y(n14332),
	.A(n15739),
	.B(FE_OFN25981_n13868));
   NOR2xp33_ASAP7_75t_R U20576 (.Y(n14344),
	.A(FE_OFN27066_n13869),
	.B(n14342));
   OA21x2_ASAP7_75t_L U20577 (.Y(n14343),
	.A1(n13875),
	.A2(n15283),
	.B(n14340));
   NAND2xp5_ASAP7_75t_L U20578 (.Y(n14340),
	.A(n14339),
	.B(n14338));
   NAND2xp5_ASAP7_75t_R U20579 (.Y(n14339),
	.A(n14336),
	.B(n14337));
   NAND2xp5_ASAP7_75t_R U20580 (.Y(n14338),
	.A(FE_OFN25915_n15514),
	.B(n14337));
   OAI21xp33_ASAP7_75t_SRAM U20581 (.Y(n15265),
	.A1(n15181),
	.A2(n15200),
	.B(n15179));
   OAI21xp33_ASAP7_75t_SRAM U20582 (.Y(n15264),
	.A1(n15196),
	.A2(FE_OFN16225_n15195),
	.B(n15194));
   NAND2xp33_ASAP7_75t_SRAM U20583 (.Y(n15178),
	.A(n15153),
	.B(n15152));
   NAND2xp33_ASAP7_75t_SRAM U20584 (.Y(n15152),
	.A(n15151),
	.B(n15150));
   NAND2xp33_ASAP7_75t_SRAM U20585 (.Y(n15177),
	.A(n15166),
	.B(n15165));
   NAND2xp33_ASAP7_75t_R U20586 (.Y(n15166),
	.A(n15161),
	.B(n15163));
   NAND2xp33_ASAP7_75t_R U20587 (.Y(n15165),
	.A(n15164),
	.B(n15163));
   NAND2xp33_ASAP7_75t_SRAM U20588 (.Y(n15176),
	.A(n15175),
	.B(n15174));
   NAND2xp33_ASAP7_75t_SRAM U20589 (.Y(n15175),
	.A(n15169),
	.B(n15172));
   NAND2xp33_ASAP7_75t_SRAM U20590 (.Y(n15174),
	.A(n15173),
	.B(n15172));
   INVxp33_ASAP7_75t_SRAM U20591 (.Y(n15169),
	.A(n15167));
   NOR2xp33_ASAP7_75t_SL U20592 (.Y(n15789),
	.A(FE_OFN26084_n15106),
	.B(n15635));
   NOR3xp33_ASAP7_75t_L U20593 (.Y(n15778),
	.A(n15813),
	.B(FE_OFN28671_FE_OCPN28076),
	.C(n13771));
   INVxp33_ASAP7_75t_SRAM U20594 (.Y(n15784),
	.A(n15782));
   INVxp33_ASAP7_75t_L U20595 (.Y(n15799),
	.A(n15797));
   OAI21xp33_ASAP7_75t_SRAM U20597 (.Y(n15882),
	.A1(n14996),
	.A2(n15858),
	.B(n15857));
   NAND2xp33_ASAP7_75t_L U20598 (.Y(n15879),
	.A(n15878),
	.B(n15877));
   NAND2xp5_ASAP7_75t_R U20599 (.Y(n15880),
	.A(n15869),
	.B(n15868));
   NAND2xp5_ASAP7_75t_R U20600 (.Y(n15855),
	.A(n15854),
	.B(n15853));
   NAND2xp33_ASAP7_75t_L U20601 (.Y(n15853),
	.A(n15852),
	.B(n15849));
   NAND2xp5_ASAP7_75t_L U20602 (.Y(n15854),
	.A(n15850),
	.B(n15849));
   INVxp33_ASAP7_75t_L U20603 (.Y(n15886),
	.A(n15839));
   NOR2xp33_ASAP7_75t_SRAM U20604 (.Y(n15837),
	.A(FE_OFN25928_n15779),
	.B(n15834));
   NAND2xp33_ASAP7_75t_R U20605 (.Y(n15821),
	.A(n15815),
	.B(n15818));
   NOR2xp33_ASAP7_75t_SRAM U20606 (.Y(n15815),
	.A(n15809),
	.B(n15816));
   NAND2xp5_ASAP7_75t_SRAM U20607 (.Y(n15820),
	.A(n15819),
	.B(n15818));
   NOR2xp33_ASAP7_75t_R U20608 (.Y(n15819),
	.A(n15817),
	.B(n15816));
   NAND2xp33_ASAP7_75t_R U20609 (.Y(n15833),
	.A(n15827),
	.B(n15830));
   NOR2xp33_ASAP7_75t_SRAM U20610 (.Y(n15827),
	.A(n15859),
	.B(n15828));
   NAND2xp33_ASAP7_75t_R U20611 (.Y(n15832),
	.A(n15831),
	.B(n15830));
   NOR2xp33_ASAP7_75t_SRAM U20612 (.Y(n15831),
	.A(n15829),
	.B(n15828));
   OAI22xp33_ASAP7_75t_L U20613 (.Y(n14135),
	.A1(n15953),
	.A2(n14134),
	.B1(n14133),
	.B2(n14134));
   NAND2xp33_ASAP7_75t_L U20614 (.Y(n14136),
	.A(n14130),
	.B(n14129));
   NOR2xp33_ASAP7_75t_SL U20616 (.Y(n14175),
	.A(n16032),
	.B(n14173));
   A2O1A1Ixp33_ASAP7_75t_SL U20618 (.Y(n14171),
	.A1(n14170),
	.A2(n14169),
	.B(n14168),
	.C(n14167));
   NAND2xp33_ASAP7_75t_SRAM U20619 (.Y(n14168),
	.A(w3_8_),
	.B(n25051));
   NOR2xp33_ASAP7_75t_SRAM U20620 (.Y(n14102),
	.A(n14932),
	.B(n14098));
   NOR2xp33_ASAP7_75t_SRAM U20621 (.Y(n14101),
	.A(n14099),
	.B(n14102));
   OAI21xp5_ASAP7_75t_SL U20622 (.Y(n14812),
	.A1(n15347),
	.A2(n15710),
	.B(n14811));
   A2O1A1Ixp33_ASAP7_75t_SL U20623 (.Y(n14810),
	.A1(n14809),
	.A2(n14808),
	.B(n15704),
	.C(n14807));
   NOR3xp33_ASAP7_75t_SL U20624 (.Y(n14808),
	.A(n14805),
	.B(n14804),
	.C(n12994));
   OAI21xp33_ASAP7_75t_L U20625 (.Y(n14813),
	.A1(FE_OFN16352_n14289),
	.A2(n15527),
	.B(n14791));
   NAND2xp33_ASAP7_75t_SL U20626 (.Y(n14788),
	.A(n14783),
	.B(n14785));
   NOR2xp33_ASAP7_75t_R U20627 (.Y(n14783),
	.A(n14772),
	.B(n14784));
   NAND2xp33_ASAP7_75t_SL U20628 (.Y(n14787),
	.A(n14786),
	.B(n14785));
   NOR2xp33_ASAP7_75t_R U20629 (.Y(n14786),
	.A(n15528),
	.B(n14784));
   NAND2xp5_ASAP7_75t_SRAM U20630 (.Y(n14768),
	.A(n14765),
	.B(n14764));
   NAND2xp33_ASAP7_75t_SRAM U20631 (.Y(n14764),
	.A(n14792),
	.B(n15683));
   NAND2xp33_ASAP7_75t_SRAM U20632 (.Y(n14765),
	.A(n15713),
	.B(n15683));
   OAI21xp33_ASAP7_75t_SRAM U20633 (.Y(n14767),
	.A1(FE_OFN6_w3_22),
	.A2(n15714),
	.B(n14766));
   NAND2xp5_ASAP7_75t_R U20634 (.Y(n13325),
	.A(n13307),
	.B(n13306));
   NAND2xp33_ASAP7_75t_L U20635 (.Y(n13306),
	.A(n13305),
	.B(n13304));
   NAND2xp33_ASAP7_75t_L U20636 (.Y(n13307),
	.A(n13303),
	.B(n13304));
   NOR2xp33_ASAP7_75t_R U20637 (.Y(n13305),
	.A(n15252),
	.B(n15216));
   NAND2xp5_ASAP7_75t_SL U20638 (.Y(n13324),
	.A(n13323),
	.B(n13322));
   NAND2xp33_ASAP7_75t_L U20639 (.Y(n13322),
	.A(n13321),
	.B(n13320));
   NAND2xp33_ASAP7_75t_L U20640 (.Y(n13323),
	.A(n13317),
	.B(n13320));
   NOR2xp33_ASAP7_75t_R U20641 (.Y(n13321),
	.A(n13319),
	.B(n13318));
   OAI22xp33_ASAP7_75t_SRAM U20642 (.Y(n13326),
	.A1(n14480),
	.A2(n13300),
	.B1(FE_OFN26111_n13288),
	.B2(n13300));
   NOR2xp33_ASAP7_75t_SRAM U20643 (.Y(n13300),
	.A(FE_OFN27061_n15239),
	.B(n14535));
   NAND2xp33_ASAP7_75t_L U20644 (.Y(n13299),
	.A(n13298),
	.B(n13297));
   NAND2xp33_ASAP7_75t_L U20645 (.Y(n13298),
	.A(n13293),
	.B(n13295));
   NAND2xp33_ASAP7_75t_L U20646 (.Y(n13297),
	.A(n13296),
	.B(n13295));
   INVxp67_ASAP7_75t_R U20647 (.Y(n13295),
	.A(n13292));
   INVx2_ASAP7_75t_L U20648 (.Y(n14515),
	.A(n13673));
   NOR2xp33_ASAP7_75t_SRAM U20649 (.Y(n13282),
	.A(n15167),
	.B(n13280));
   OAI22xp33_ASAP7_75t_SRAM U20650 (.Y(n13277),
	.A1(n15188),
	.A2(n13290),
	.B1(FE_OFN26049_w3_27),
	.B2(n13290));
   A2O1A1Ixp33_ASAP7_75t_L U20652 (.Y(n13276),
	.A1(FE_OCPN8232_FE_OFN27206_w3_30),
	.A2(FE_OFN25895_n13662),
	.B(n15203),
	.C(n13275));
   OAI21x1_ASAP7_75t_L U20653 (.Y(n15116),
	.A1(FE_OFN28695_n),
	.A2(n15817),
	.B(n15595));
   NOR2xp33_ASAP7_75t_R U20654 (.Y(n13739),
	.A(n24831),
	.B(n15813));
   NOR2xp33_ASAP7_75t_SRAM U20655 (.Y(n13735),
	.A(n15792),
	.B(n13728));
   OAI21xp33_ASAP7_75t_SRAM U20656 (.Y(n13728),
	.A1(n15092),
	.A2(FE_OFN28889_n15845),
	.B(n13727));
   INVxp33_ASAP7_75t_L U20657 (.Y(n13734),
	.A(n13733));
   NOR3xp33_ASAP7_75t_L U20658 (.Y(n13775),
	.A(n14838),
	.B(FE_OFN28662_w3_7),
	.C(n13726));
   NAND2xp33_ASAP7_75t_SRAM U20659 (.Y(n15976),
	.A(n15447),
	.B(n15446));
   OAI21xp33_ASAP7_75t_R U20661 (.Y(n15929),
	.A1(n13804),
	.A2(n15921),
	.B(n15975));
   NOR3xp33_ASAP7_75t_SRAM U20662 (.Y(n13941),
	.A(n14913),
	.B(FE_OCPN29521_n24755),
	.C(n14957));
   OR3x1_ASAP7_75t_SRAM U20663 (.Y(n13942),
	.A(FE_OFN26007_n16010),
	.B(n15438),
	.C(n15374));
   NAND2xp5_ASAP7_75t_L U20665 (.Y(n13991),
	.A(n13983),
	.B(n13982));
   NAND3xp33_ASAP7_75t_R U20666 (.Y(n13993),
	.A(n14693),
	.B(n13974),
	.C(n13973));
   NAND2xp33_ASAP7_75t_SRAM U20667 (.Y(n13974),
	.A(n13844),
	.B(n14607));
   NAND2xp5_ASAP7_75t_R U20668 (.Y(n13973),
	.A(n13972),
	.B(n13971));
   NAND2xp33_ASAP7_75t_L U20669 (.Y(n13971),
	.A(n13970),
	.B(n13967));
   NAND2xp33_ASAP7_75t_L U20670 (.Y(n13956),
	.A(n13951),
	.B(n13953));
   NOR2xp33_ASAP7_75t_SRAM U20671 (.Y(n13951),
	.A(n15934),
	.B(n13952));
   NAND2xp33_ASAP7_75t_R U20672 (.Y(n13955),
	.A(n13954),
	.B(n13953));
   NOR2xp33_ASAP7_75t_SRAM U20673 (.Y(n13954),
	.A(n15375),
	.B(n13952));
   NAND2xp33_ASAP7_75t_R U20674 (.Y(n13964),
	.A(n13963),
	.B(n13962));
   NOR2xp33_ASAP7_75t_SRAM U20675 (.Y(n13963),
	.A(FE_OCPN29583_n15422),
	.B(n13961));
   NAND2xp33_ASAP7_75t_L U20676 (.Y(n13965),
	.A(n13960),
	.B(n13962));
   NOR2xp33_ASAP7_75t_SRAM U20677 (.Y(n13960),
	.A(n13957),
	.B(n13961));
   NAND2xp33_ASAP7_75t_L U20679 (.Y(n13913),
	.A(n13907),
	.B(n13906));
   NAND2xp33_ASAP7_75t_SL U20680 (.Y(n13912),
	.A(n13908),
	.B(n13911));
   NAND3xp33_ASAP7_75t_SL U20681 (.Y(n13927),
	.A(n13926),
	.B(n14316),
	.C(n13925));
   O2A1O1Ixp5_ASAP7_75t_SRAM U20682 (.Y(n13925),
	.A1(FE_OFN6_w3_22),
	.A2(FE_OFN28623_n13874),
	.B(n15528),
	.C(n13924));
   O2A1O1Ixp5_ASAP7_75t_SRAM U20683 (.Y(n13924),
	.A1(FE_OFN6_w3_22),
	.A2(n15536),
	.B(n15719),
	.C(FE_OCPN8264_n13890));
   NAND2xp33_ASAP7_75t_R U20684 (.Y(n13900),
	.A(n13896),
	.B(n13895));
   NOR2xp33_ASAP7_75t_SRAM U20685 (.Y(n13896),
	.A(n14377),
	.B(n13897));
   NAND2xp33_ASAP7_75t_SRAM U20686 (.Y(n13899),
	.A(n13898),
	.B(n13895));
   NOR2xp33_ASAP7_75t_SRAM U20687 (.Y(n13898),
	.A(FE_OFN27066_n13869),
	.B(n13897));
   NOR2xp33_ASAP7_75t_SRAM U20688 (.Y(n13884),
	.A(n13882),
	.B(n13881));
   NOR2xp33_ASAP7_75t_SRAM U20690 (.Y(n13880),
	.A(n15275),
	.B(n13881));
   NAND2xp5_ASAP7_75t_L U20691 (.Y(n13625),
	.A(n13620),
	.B(n13622));
   NOR2xp33_ASAP7_75t_L U20692 (.Y(n13620),
	.A(n15246),
	.B(n13621));
   NAND2xp5_ASAP7_75t_L U20693 (.Y(n13624),
	.A(n13623),
	.B(n13622));
   NOR2xp33_ASAP7_75t_SL U20694 (.Y(n13623),
	.A(n13650),
	.B(n13621));
   NAND2xp33_ASAP7_75t_R U20695 (.Y(n13572),
	.A(n13571),
	.B(n13570));
   NOR2xp33_ASAP7_75t_SRAM U20696 (.Y(n13571),
	.A(FE_OFN28603_n14534),
	.B(n13569));
   NAND2xp33_ASAP7_75t_R U20697 (.Y(n13573),
	.A(n13568),
	.B(n13570));
   NOR2xp33_ASAP7_75t_SRAM U20698 (.Y(n13568),
	.A(n14572),
	.B(n13569));
   NAND2xp33_ASAP7_75t_SRAM U20699 (.Y(n13580),
	.A(n13576),
	.B(n13577));
   NOR2xp33_ASAP7_75t_SRAM U20700 (.Y(n13576),
	.A(FE_OFN26567_n),
	.B(FE_OCPN29573_n15184));
   NAND2xp33_ASAP7_75t_SRAM U20701 (.Y(n13579),
	.A(n13578),
	.B(n13577));
   OAI21xp33_ASAP7_75t_SRAM U20702 (.Y(n14485),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OFN27212_w3_30),
	.B(n15205));
   NAND2xp33_ASAP7_75t_SRAM U20703 (.Y(n13562),
	.A(n13558),
	.B(n13559));
   NOR2xp33_ASAP7_75t_SRAM U20704 (.Y(n13558),
	.A(FE_OFN26567_n),
	.B(n13566));
   NAND2xp33_ASAP7_75t_R U20705 (.Y(n13561),
	.A(n13560),
	.B(n13559));
   NOR2xp33_ASAP7_75t_SRAM U20706 (.Y(n13560),
	.A(n14479),
	.B(n13566));
   INVx1_ASAP7_75t_SL U20707 (.Y(n15185),
	.A(n13459));
   NAND2xp33_ASAP7_75t_SRAM U20708 (.Y(n13552),
	.A(n13551),
	.B(FE_OFN25966_n13646));
   NAND2xp33_ASAP7_75t_R U20709 (.Y(n13553),
	.A(n13550),
	.B(FE_OFN25966_n13646));
   OA21x2_ASAP7_75t_L U20710 (.Y(n14883),
	.A1(n14881),
	.A2(n15808),
	.B(n14880));
   INVxp33_ASAP7_75t_L U20712 (.Y(n15802),
	.A(n15626));
   NAND2xp33_ASAP7_75t_R U20713 (.Y(n14885),
	.A(n14882),
	.B(n14883));
   NOR2xp33_ASAP7_75t_L U20715 (.Y(n14850),
	.A(n14849),
	.B(n14848));
   A2O1A1Ixp33_ASAP7_75t_R U20716 (.Y(n14848),
	.A1(n15825),
	.A2(n15870),
	.B(n25140),
	.C(n14847));
   NAND3xp33_ASAP7_75t_SL U20717 (.Y(n14886),
	.A(n14874),
	.B(n14873),
	.C(n14872));
   OAI222xp33_ASAP7_75t_L U20718 (.Y(n14874),
	.A1(FE_OFN29052_w3_5),
	.A2(n14865),
	.B1(n15627),
	.B2(n14865),
	.C1(FE_OFN25897_w3_4),
	.C2(n14865));
   NAND2xp33_ASAP7_75t_R U20719 (.Y(n14873),
	.A(n14871),
	.B(n14870));
   NOR2xp33_ASAP7_75t_SRAM U20720 (.Y(n14836),
	.A(n15838),
	.B(n14837));
   AND3x1_ASAP7_75t_L U20721 (.Y(n14839),
	.A(n14835),
	.B(n14834),
	.C(n14833));
   OAI222xp33_ASAP7_75t_SRAM U20722 (.Y(n14834),
	.A1(n15859),
	.A2(n15778),
	.B1(n13771),
	.B2(n15778),
	.C1(FE_OFN28671_FE_OCPN28076),
	.C2(n15778));
   OAI22xp33_ASAP7_75t_L U20723 (.Y(n14835),
	.A1(n15811),
	.A2(n14832),
	.B1(n14831),
	.B2(n14832));
   NAND2xp33_ASAP7_75t_L U20724 (.Y(n14832),
	.A(n14830),
	.B(n14829));
   NOR2xp33_ASAP7_75t_SRAM U20725 (.Y(n14840),
	.A(n14838),
	.B(n14837));
   NAND2xp33_ASAP7_75t_R U20726 (.Y(n15289),
	.A(n15285),
	.B(n15284));
   NAND2xp33_ASAP7_75t_R U20727 (.Y(n15288),
	.A(n15287),
	.B(n15284));
   NOR2xp33_ASAP7_75t_R U20728 (.Y(n15287),
	.A(n15528),
	.B(n15286));
   NAND2xp33_ASAP7_75t_SRAM U20729 (.Y(n15279),
	.A(n15276),
	.B(n15277));
   NOR2xp33_ASAP7_75t_R U20730 (.Y(n15276),
	.A(n15274),
	.B(n15273));
   NOR2xp33_ASAP7_75t_SRAM U20731 (.Y(n15274),
	.A(n13916),
	.B(FE_OFN27074_n13868));
   NAND2xp33_ASAP7_75t_SRAM U20732 (.Y(n15278),
	.A(n15536),
	.B(n15277));
   NOR2xp33_ASAP7_75t_L U20733 (.Y(n15661),
	.A(FE_OFN28769_n15478),
	.B(n13875));
   NAND2xp33_ASAP7_75t_SRAM U20734 (.Y(n13342),
	.A(n13337),
	.B(n13339));
   NAND2xp33_ASAP7_75t_L U20735 (.Y(n13341),
	.A(n13340),
	.B(n13339));
   NAND2xp33_ASAP7_75t_SRAM U20737 (.Y(n13343),
	.A(FE_OFN28452_w3_29),
	.B(FE_OFN27129_w3_28));
   NOR3x1_ASAP7_75t_SL U20738 (.Y(n15240),
	.A(FE_OFN28571_w3_28),
	.B(FE_OFN28452_w3_29),
	.C(FE_OCPN28096_w3_31));
   NAND2xp5_ASAP7_75t_SL U20739 (.Y(n15017),
	.A(n15014),
	.B(n15013));
   NAND2xp33_ASAP7_75t_L U20740 (.Y(n15013),
	.A(n15012),
	.B(n15011));
   NAND2xp33_ASAP7_75t_L U20741 (.Y(n15014),
	.A(n15008),
	.B(n15011));
   NOR2xp33_ASAP7_75t_L U20742 (.Y(n15012),
	.A(n15010),
	.B(n15009));
   NOR2xp33_ASAP7_75t_SRAM U20743 (.Y(n15015),
	.A(n13736),
	.B(FE_OFN28682_n15888));
   NAND2xp33_ASAP7_75t_SRAM U20744 (.Y(n14999),
	.A(n14996),
	.B(n15787));
   NAND2xp33_ASAP7_75t_SRAM U20745 (.Y(n14998),
	.A(n14997),
	.B(n15787));
   NAND2xp5_ASAP7_75t_R U20746 (.Y(n15049),
	.A(n15884),
	.B(n15048));
   NAND3xp33_ASAP7_75t_SL U20747 (.Y(n15048),
	.A(n15047),
	.B(n15046),
	.C(n15073));
   NAND2xp5_ASAP7_75t_SRAM U20748 (.Y(n15051),
	.A(n15039),
	.B(n15626));
   NAND2xp33_ASAP7_75t_R U20749 (.Y(n15039),
	.A(n15038),
	.B(n15037));
   NAND2xp33_ASAP7_75t_SRAM U20750 (.Y(n15050),
	.A(n15044),
	.B(n15842));
   NAND2xp33_ASAP7_75t_SRAM U20751 (.Y(n15044),
	.A(n15043),
	.B(n15042));
   NAND2xp33_ASAP7_75t_L U20752 (.Y(n15031),
	.A(n15027),
	.B(n15026));
   NAND2xp33_ASAP7_75t_L U20753 (.Y(n15026),
	.A(n15025),
	.B(n15024));
   NAND2xp33_ASAP7_75t_L U20754 (.Y(n15027),
	.A(n15022),
	.B(n15024));
   NOR2xp33_ASAP7_75t_R U20755 (.Y(n15025),
	.A(n15788),
	.B(n15023));
   OAI222xp33_ASAP7_75t_R U20756 (.Y(n15030),
	.A1(n15843),
	.A2(n15029),
	.B1(FE_OFN25900_w3_4),
	.B2(n15029),
	.C1(FE_OCPN8252_FE_OFN28661_w3_7),
	.C2(n15029));
   NAND3xp33_ASAP7_75t_L U20757 (.Y(n15040),
	.A(FE_OFN25900_w3_4),
	.B(n15601),
	.C(n15857));
   NOR2xp33_ASAP7_75t_SRAM U20758 (.Y(n15381),
	.A(n15380),
	.B(FE_OFN112_n15994));
   NAND2xp33_ASAP7_75t_L U20759 (.Y(n15384),
	.A(n15383),
	.B(n15382));
   INVxp33_ASAP7_75t_SRAM U20760 (.Y(n15379),
	.A(n14645));
   NAND2xp5_ASAP7_75t_SL U20761 (.Y(n14308),
	.A(n14307),
	.B(n14306));
   NAND2xp5_ASAP7_75t_L U20762 (.Y(n14306),
	.A(n14305),
	.B(n14304));
   NAND2xp33_ASAP7_75t_SL U20763 (.Y(n14307),
	.A(n14301),
	.B(n14304));
   NAND3xp33_ASAP7_75t_SRAM U20764 (.Y(n14318),
	.A(n14317),
	.B(n14316),
	.C(n14789));
   NAND2xp33_ASAP7_75t_L U20765 (.Y(n14317),
	.A(n14313),
	.B(n14312));
   NAND2xp33_ASAP7_75t_SRAM U20766 (.Y(n14312),
	.A(n14311),
	.B(n13892));
   NAND2xp33_ASAP7_75t_SL U20767 (.Y(n14313),
	.A(n14309),
	.B(n13892));
   NAND2xp5_ASAP7_75t_L U20768 (.Y(n14284),
	.A(n14283),
	.B(n14282));
   NAND2xp33_ASAP7_75t_SL U20769 (.Y(n14282),
	.A(n14281),
	.B(n14280));
   NAND2xp33_ASAP7_75t_SL U20770 (.Y(n14283),
	.A(n14279),
	.B(n14280));
   OAI21xp33_ASAP7_75t_SRAM U20771 (.Y(n15527),
	.A1(FE_OFN26114_n),
	.A2(FE_OFN28623_n13874),
	.B(n14276));
   NAND2xp33_ASAP7_75t_L U20772 (.Y(n14275),
	.A(n14269),
	.B(n14272));
   NOR2xp33_ASAP7_75t_R U20773 (.Y(n14269),
	.A(n15757),
	.B(n14270));
   NOR2xp33_ASAP7_75t_R U20774 (.Y(n14273),
	.A(n14271),
	.B(n14270));
   NAND2xp33_ASAP7_75t_R U20775 (.Y(n13415),
	.A(n13450),
	.B(n13412));
   NAND2xp33_ASAP7_75t_R U20776 (.Y(n13412),
	.A(n13411),
	.B(FE_OFN28455_n13348));
   NOR2xp33_ASAP7_75t_SRAM U20777 (.Y(n13411),
	.A(FE_OFN26111_n13288),
	.B(n14479));
   NAND2xp5_ASAP7_75t_L U20778 (.Y(n13677),
	.A(n15185),
	.B(n13596));
   NOR2xp33_ASAP7_75t_R U20779 (.Y(n13414),
	.A(FE_OFN16193_n15200),
	.B(n13415));
   OA21x2_ASAP7_75t_R U20780 (.Y(n13416),
	.A1(FE_OFN16451_n),
	.A2(n15196),
	.B(n13563));
   OAI21xp33_ASAP7_75t_SRAM U20781 (.Y(n13696),
	.A1(FE_OCPN29350_w3_25),
	.A2(FE_OFN28891_n),
	.B(FE_OFN27206_w3_30));
   NOR2xp33_ASAP7_75t_L U20782 (.Y(n13469),
	.A(n14491),
	.B(n13467));
   NAND2xp5_ASAP7_75t_SL U20783 (.Y(n13471),
	.A(n13466),
	.B(n13468));
   NOR2xp33_ASAP7_75t_L U20784 (.Y(n13466),
	.A(n13447),
	.B(n13467));
   OAI21xp5_ASAP7_75t_L U20787 (.Y(n15973),
	.A1(FE_OCPN29536_FE_OFN8_w3_14),
	.A2(n14912),
	.B(n15955));
   OAI21xp33_ASAP7_75t_SL U20788 (.Y(n14960),
	.A1(n14959),
	.A2(FE_OFN16348_n15949),
	.B(n14958));
   NOR3xp33_ASAP7_75t_SRAM U20789 (.Y(n14955),
	.A(FE_OFN109_n15994),
	.B(w3_10_),
	.C(w3_8_));
   NOR3xp33_ASAP7_75t_SL U20791 (.Y(n14926),
	.A(n14925),
	.B(n14924),
	.C(n14923));
   NOR2xp33_ASAP7_75t_SRAM U20792 (.Y(n14925),
	.A(n16016),
	.B(n15983));
   OAI21xp33_ASAP7_75t_L U20793 (.Y(n14961),
	.A1(n14941),
	.A2(n14937),
	.B(n14936));
   NOR3xp33_ASAP7_75t_L U20794 (.Y(n14936),
	.A(n14935),
	.B(n14934),
	.C(n15978));
   NAND2xp33_ASAP7_75t_R U20795 (.Y(n14909),
	.A(n14908),
	.B(n14907));
   NAND2xp33_ASAP7_75t_SRAM U20796 (.Y(n14908),
	.A(n14906),
	.B(n14919));
   NAND2xp33_ASAP7_75t_SRAM U20797 (.Y(n14903),
	.A(FE_OCPN29583_n15422),
	.B(n15956));
   NAND2xp33_ASAP7_75t_SRAM U20798 (.Y(n14904),
	.A(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(n14924));
   OAI22xp33_ASAP7_75t_SRAM U20799 (.Y(n14905),
	.A1(FE_OFN27115_n),
	.A2(n15455),
	.B1(FE_OCPN29535_FE_OFN8_w3_14),
	.B2(n15455));
   NOR2xp33_ASAP7_75t_SRAM U20800 (.Y(n14918),
	.A(n14912),
	.B(n15413));
   NOR3xp33_ASAP7_75t_SRAM U20801 (.Y(n14917),
	.A(n14914),
	.B(FE_OCPN29521_n24755),
	.C(n14913));
   NOR3xp33_ASAP7_75t_SRAM U20802 (.Y(n14916),
	.A(n14915),
	.B(FE_OCPN29427_w3_15),
	.C(n15423));
   NAND3xp33_ASAP7_75t_L U20803 (.Y(n15554),
	.A(n15552),
	.B(n15551),
	.C(n15550));
   OAI21xp33_ASAP7_75t_SRAM U20804 (.Y(n15550),
	.A1(n15739),
	.A2(n15715),
	.B(FE_OFN26614_n));
   NAND2xp33_ASAP7_75t_SL U20805 (.Y(n15552),
	.A(n15549),
	.B(n15548));
   NAND2xp5_ASAP7_75t_L U20806 (.Y(n15548),
	.A(n15547),
	.B(n15546));
   O2A1O1Ixp5_ASAP7_75t_SRAM U20807 (.Y(n15553),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(n15501),
	.B(n15688),
	.C(n15491));
   NOR2xp33_ASAP7_75t_SRAM U20808 (.Y(n15533),
	.A(n13867),
	.B(n15553));
   INVx1_ASAP7_75t_SL U20809 (.Y(n15555),
	.A(n15532));
   NAND2xp33_ASAP7_75t_SL U20810 (.Y(n15530),
	.A(n15511),
	.B(n15510));
   NAND2xp33_ASAP7_75t_SL U20811 (.Y(n15531),
	.A(n15500),
	.B(n15499));
   NOR2xp33_ASAP7_75t_SRAM U20812 (.Y(n13490),
	.A(n15162),
	.B(n13708));
   INVx1_ASAP7_75t_SL U20813 (.Y(n13491),
	.A(n13489));
   O2A1O1Ixp33_ASAP7_75t_L U20814 (.Y(n13489),
	.A1(FE_OFN28929_n15182),
	.A2(FE_OFN28453_n13348),
	.B(n14559),
	.C(n13488));
   NAND2xp5_ASAP7_75t_L U20815 (.Y(n13488),
	.A(n13487),
	.B(n13486));
   NAND2xp5_ASAP7_75t_L U20816 (.Y(n13487),
	.A(n13483),
	.B(n13482));
   NAND2xp33_ASAP7_75t_L U20817 (.Y(n13510),
	.A(n13509),
	.B(n13508));
   NAND2xp33_ASAP7_75t_R U20818 (.Y(n13508),
	.A(n13507),
	.B(n13506));
   NAND2xp33_ASAP7_75t_L U20819 (.Y(n13509),
	.A(n13504),
	.B(n13506));
   NOR2xp33_ASAP7_75t_R U20820 (.Y(n13507),
	.A(FE_OFN26059_n),
	.B(n13505));
   NAND3xp33_ASAP7_75t_R U20821 (.Y(n13511),
	.A(n13556),
	.B(n15156),
	.C(FE_OFN25875_n15227));
   NAND2xp5_ASAP7_75t_L U20823 (.Y(n13525),
	.A(n13524),
	.B(n13523));
   NAND2xp5_ASAP7_75t_R U20824 (.Y(n13523),
	.A(n13522),
	.B(n13521));
   NAND2xp5_ASAP7_75t_L U20825 (.Y(n13524),
	.A(n13518),
	.B(n13521));
   NOR2xp33_ASAP7_75t_SRAM U20826 (.Y(n13522),
	.A(n15234),
	.B(n13520));
   NOR3xp33_ASAP7_75t_L U20827 (.Y(n13514),
	.A(FE_OFN25893_n15214),
	.B(FE_OFN28603_n14534),
	.C(FE_OFN16201_n15197));
   NAND2xp33_ASAP7_75t_L U20828 (.Y(n13539),
	.A(n13538),
	.B(n13537));
   NAND2xp33_ASAP7_75t_L U20829 (.Y(n13538),
	.A(n13533),
	.B(n13535));
   NAND2xp33_ASAP7_75t_R U20830 (.Y(n13537),
	.A(n13536),
	.B(n13535));
   NAND2xp67_ASAP7_75t_SL U20832 (.Y(n15834),
	.A(FE_OCPN29537_FE_OFN28699_w3_6),
	.B(n25140));
   NAND2xp33_ASAP7_75t_SRAM U20834 (.Y(n15077),
	.A(n15075),
	.B(n15074));
   NOR2xp33_ASAP7_75t_SRAM U20835 (.Y(n15075),
	.A(n15578),
	.B(FE_OFN28662_w3_7));
   NOR3xp33_ASAP7_75t_SRAM U20836 (.Y(n15780),
	.A(n13730),
	.B(FE_OCPN8252_FE_OFN28661_w3_7),
	.C(n15814));
   OAI21xp33_ASAP7_75t_SRAM U20837 (.Y(n15132),
	.A1(n13766),
	.A2(n13730),
	.B(n15115));
   NOR2xp33_ASAP7_75t_L U20838 (.Y(n15130),
	.A(n15843),
	.B(n15129));
   NAND3xp33_ASAP7_75t_L U20839 (.Y(n15131),
	.A(n15127),
	.B(n15126),
	.C(n15125));
   NAND2xp33_ASAP7_75t_L U20840 (.Y(n15135),
	.A(n15105),
	.B(n15104));
   NAND2xp33_ASAP7_75t_L U20841 (.Y(n15105),
	.A(n15100),
	.B(n15102));
   NAND2xp33_ASAP7_75t_L U20842 (.Y(n15104),
	.A(n15103),
	.B(n15102));
   INVxp33_ASAP7_75t_R U20843 (.Y(n15100),
	.A(n15092));
   NAND2xp33_ASAP7_75t_L U20844 (.Y(n15134),
	.A(n15114),
	.B(n15113));
   NAND2xp33_ASAP7_75t_R U20845 (.Y(n15113),
	.A(n15112),
	.B(n15111));
   NAND2xp33_ASAP7_75t_R U20846 (.Y(n15114),
	.A(n15110),
	.B(n15111));
   NAND2xp33_ASAP7_75t_L U20847 (.Y(n15090),
	.A(n15085),
	.B(n15084));
   NAND2xp33_ASAP7_75t_SRAM U20848 (.Y(n15084),
	.A(FE_OFN29052_w3_5),
	.B(n15083));
   NAND2xp33_ASAP7_75t_L U20849 (.Y(n15085),
	.A(n15082),
	.B(n15083));
   OR2x2_ASAP7_75t_R U20850 (.Y(n15083),
	.A(n15592),
	.B(n15861));
   NAND2xp33_ASAP7_75t_SRAM U20851 (.Y(n15089),
	.A(n15589),
	.B(n15088));
   NAND2xp33_ASAP7_75t_SRAM U20852 (.Y(n15088),
	.A(n15087),
	.B(n15086));
   NOR2xp33_ASAP7_75t_SRAM U20853 (.Y(n15087),
	.A(n15835),
	.B(n15093));
   NOR2x1_ASAP7_75t_R U20854 (.Y(n15809),
	.A(FE_OFN28721_n),
	.B(n15639));
   NOR2x1_ASAP7_75t_L U20855 (.Y(n15627),
	.A(n24831),
	.B(n25140));
   NAND2xp5_ASAP7_75t_SL U20856 (.Y(n15635),
	.A(FE_OFN28671_FE_OCPN28076),
	.B(n13771));
   NAND2xp33_ASAP7_75t_R U20857 (.Y(n15068),
	.A(n15063),
	.B(n15065));
   NAND2xp33_ASAP7_75t_R U20858 (.Y(n15067),
	.A(n15066),
	.B(n15065));
   NOR2xp33_ASAP7_75t_L U20859 (.Y(n14666),
	.A(n14157),
	.B(FE_OFN26007_n16010));
   NOR3xp33_ASAP7_75t_L U20860 (.Y(n15383),
	.A(FE_OCPN29570_n15423),
	.B(FE_OFN27200_n),
	.C(n15374));
   NAND2xp33_ASAP7_75t_R U20861 (.Y(n15664),
	.A(n15663),
	.B(n15662));
   NAND2xp33_ASAP7_75t_SRAM U20862 (.Y(n15663),
	.A(FE_PSN8280_n15660),
	.B(n15659));
   NOR2xp33_ASAP7_75t_SRAM U20865 (.Y(n15676),
	.A(n15674),
	.B(n15673));
   AND3x1_ASAP7_75t_L U20866 (.Y(n15675),
	.A(n15671),
	.B(n15670),
	.C(n15669));
   OAI222xp33_ASAP7_75t_L U20867 (.Y(n15671),
	.A1(FE_OFN26045_n25377),
	.A2(n15666),
	.B1(n15729),
	.B2(n15666),
	.C1(FE_OFN26091_n24663),
	.C2(n15666));
   NOR2xp33_ASAP7_75t_L U20869 (.Y(n13708),
	.A(FE_OFN16225_n15195),
	.B(FE_OFN28717_n15158));
   NAND2xp33_ASAP7_75t_SRAM U20871 (.Y(n14459),
	.A(n15859),
	.B(n15810));
   NAND2xp33_ASAP7_75t_SL U20872 (.Y(n14460),
	.A(n14457),
	.B(n14456));
   NAND2xp33_ASAP7_75t_SL U20873 (.Y(n14456),
	.A(n14455),
	.B(n14454));
   O2A1O1Ixp33_ASAP7_75t_R U20874 (.Y(n14462),
	.A1(n15782),
	.A2(n15639),
	.B(n14447),
	.C(n15881));
   NAND3xp33_ASAP7_75t_L U20876 (.Y(n14446),
	.A(n14844),
	.B(n14445),
	.C(n14444));
   NAND2xp5_ASAP7_75t_L U20877 (.Y(n14435),
	.A(n14434),
	.B(n14433));
   NAND2xp33_ASAP7_75t_SL U20878 (.Y(n14434),
	.A(n14428),
	.B(n14431));
   NAND2xp33_ASAP7_75t_R U20879 (.Y(n14438),
	.A(n14425),
	.B(n14424));
   NAND2xp33_ASAP7_75t_SRAM U20880 (.Y(n14425),
	.A(n14422),
	.B(n15787));
   NAND2xp33_ASAP7_75t_SRAM U20881 (.Y(n14424),
	.A(n14423),
	.B(n15787));
   NOR2xp33_ASAP7_75t_SRAM U20882 (.Y(n14422),
	.A(FE_OCPN27985_n24831),
	.B(n14996));
   OAI21xp33_ASAP7_75t_SRAM U20883 (.Y(n14437),
	.A1(FE_OCPN27985_n24831),
	.A2(FE_OFN25887_w3_3),
	.B(FE_OFN26531_n));
   NOR2x1_ASAP7_75t_L U20884 (.Y(n15033),
	.A(FE_OFN26645_n),
	.B(FE_OFN28732_n));
   NOR2x2_ASAP7_75t_SL U20885 (.Y(n15862),
	.A(FE_OCPN27978_w3_3),
	.B(FE_OFN27124_w3_1));
   NOR3xp33_ASAP7_75t_L U20886 (.Y(n15619),
	.A(n15808),
	.B(w3_0_),
	.C(w3_2_));
   NAND2xp33_ASAP7_75t_L U20887 (.Y(n14419),
	.A(n14416),
	.B(n14415));
   NAND2xp33_ASAP7_75t_R U20888 (.Y(n14415),
	.A(n14414),
	.B(n14413));
   NAND2xp33_ASAP7_75t_SRAM U20889 (.Y(n14416),
	.A(n14411),
	.B(n14413));
   INVxp33_ASAP7_75t_SRAM U20890 (.Y(n14413),
	.A(n14846));
   OAI21xp5_ASAP7_75t_L U20892 (.Y(n15610),
	.A1(FE_OFN28747_n),
	.A2(n15034),
	.B(n15834));
   NAND2xp5_ASAP7_75t_SL U20893 (.Y(n16037),
	.A(n16036),
	.B(n16035));
   NAND2xp5_ASAP7_75t_L U20894 (.Y(n16035),
	.A(n16034),
	.B(n16033));
   NAND2xp33_ASAP7_75t_SL U20895 (.Y(n16036),
	.A(n16030),
	.B(n16033));
   NOR2xp33_ASAP7_75t_L U20896 (.Y(n16034),
	.A(n16032),
	.B(n16031));
   NAND2xp33_ASAP7_75t_R U20897 (.Y(n15945),
	.A(n15933),
	.B(n15932));
   NAND2xp33_ASAP7_75t_R U20898 (.Y(n15932),
	.A(n15931),
	.B(n15930));
   NAND2xp33_ASAP7_75t_R U20899 (.Y(n15933),
	.A(n15928),
	.B(n15930));
   NAND2xp33_ASAP7_75t_SRAM U20901 (.Y(n15944),
	.A(n15943),
	.B(n15942));
   NAND2xp33_ASAP7_75t_SRAM U20902 (.Y(n15942),
	.A(n15941),
	.B(n15940));
   NAND2xp33_ASAP7_75t_SRAM U20903 (.Y(n15943),
	.A(n15938),
	.B(n15940));
   NOR2xp33_ASAP7_75t_R U20904 (.Y(n15941),
	.A(FE_OFN27115_n),
	.B(n15939));
   NAND2xp5_ASAP7_75t_SRAM U20907 (.Y(n26582),
	.A(n26580),
	.B(n26578));
   O2A1O1Ixp5_ASAP7_75t_SL U20908 (.Y(n24283),
	.A1(n25577),
	.A2(n25576),
	.B(n25575),
	.C(n25379));
   NOR2x1_ASAP7_75t_L U20909 (.Y(n25764),
	.A(FE_OCPN5119_n25762),
	.B(n25761));
   NAND2xp5_ASAP7_75t_L U20911 (.Y(n23915),
	.A(FE_OFN140_w3_2),
	.B(FE_OCPN28089_n23913));
   NAND2xp5_ASAP7_75t_R U20912 (.Y(n23920),
	.A(n23910),
	.B(n23909));
   NAND2xp33_ASAP7_75t_R U20913 (.Y(n23909),
	.A(n23908),
	.B(n23907));
   NAND2xp33_ASAP7_75t_SRAM U20914 (.Y(n23910),
	.A(n23905),
	.B(n23907));
   INVxp33_ASAP7_75t_SRAM U20915 (.Y(n23919),
	.A(n23911));
   OAI21xp5_ASAP7_75t_SL U20916 (.Y(n26011),
	.A1(n25852),
	.A2(n27168),
	.B(n25851));
   NOR3xp33_ASAP7_75t_SL U20917 (.Y(n25852),
	.A(n25850),
	.B(FE_OCPN27316_n25849),
	.C(n25848));
   NAND2xp33_ASAP7_75t_L U20918 (.Y(n25850),
	.A(n25847),
	.B(n25846));
   NOR3xp33_ASAP7_75t_R U20919 (.Y(n26000),
	.A(n25998),
	.B(FE_OCPN29437_n25864),
	.C(n25996));
   O2A1O1Ixp5_ASAP7_75t_SL U20920 (.Y(n26903),
	.A1(n26900),
	.A2(n26899),
	.B(n27207),
	.C(n26898));
   NAND3xp33_ASAP7_75t_L U20922 (.Y(n25330),
	.A(n25899),
	.B(n25902),
	.C(FE_OCPN28366_n25329));
   NAND2xp33_ASAP7_75t_SL U20924 (.Y(n26883),
	.A(n26882),
	.B(n26881));
   NAND2xp33_ASAP7_75t_L U20925 (.Y(n26869),
	.A(FE_OFN29024_n),
	.B(n26866));
   O2A1O1Ixp33_ASAP7_75t_L U20926 (.Y(n26886),
	.A1(n26889),
	.A2(n26888),
	.B(n26885),
	.C(n26884));
   NAND2xp5_ASAP7_75t_L U20930 (.Y(n27115),
	.A(FE_OFN29011_n27113),
	.B(FE_OFN16331_n27151));
   NAND2xp33_ASAP7_75t_L U20933 (.Y(n18054),
	.A(n18053),
	.B(n18892));
   NAND3xp33_ASAP7_75t_SL U20936 (.Y(n26979),
	.A(n25915),
	.B(n25914),
	.C(n25913));
   A2O1A1Ixp33_ASAP7_75t_SL U20937 (.Y(n25752),
	.A1(n26250),
	.A2(n26282),
	.B(n26251),
	.C(n26277));
   NAND2xp33_ASAP7_75t_SL U20938 (.Y(n25753),
	.A(FE_OFN28990_n26276),
	.B(FE_OFN28525_n25751));
   NOR2xp33_ASAP7_75t_R U20939 (.Y(n25659),
	.A(FE_OFN28582_n25657),
	.B(n25667));
   NAND2xp5_ASAP7_75t_L U20940 (.Y(n25655),
	.A(FE_OFN25899_w3_4),
	.B(FE_OFN28504_n25956));
   NAND2x1_ASAP7_75t_SL U20941 (.Y(n24006),
	.A(n26335),
	.B(FE_OCPN27991_n26336));
   A2O1A1Ixp33_ASAP7_75t_SL U20942 (.Y(n24021),
	.A1(n26819),
	.A2(n26725),
	.B(n24019),
	.C(n24018));
   NAND2xp33_ASAP7_75t_SRAM U20943 (.Y(n24019),
	.A(n26721),
	.B(FE_OFN16276_w3_5));
   NAND2xp33_ASAP7_75t_SRAM U20945 (.Y(n25036),
	.A(n25035),
	.B(n25034));
   NAND2xp33_ASAP7_75t_SRAM U20946 (.Y(n25037),
	.A(n25023),
	.B(n25034));
   NAND2xp33_ASAP7_75t_SRAM U20947 (.Y(n25886),
	.A(n25879),
	.B(n25878));
   NAND2xp5_ASAP7_75t_SL U20949 (.Y(n24743),
	.A(n25953),
	.B(n25954));
   NAND2xp33_ASAP7_75t_SRAM U20950 (.Y(n26170),
	.A(n26158),
	.B(n26562));
   NAND2xp33_ASAP7_75t_SRAM U20951 (.Y(n26169),
	.A(n26168),
	.B(n26562));
   NAND2xp33_ASAP7_75t_SL U20952 (.Y(n26174),
	.A(FE_OFN25939_n26275),
	.B(FE_OFN135_n26172));
   A2O1A1Ixp33_ASAP7_75t_SL U20954 (.Y(n24353),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(n24351),
	.C(n24350));
   NAND2xp33_ASAP7_75t_R U20955 (.Y(n24351),
	.A(n26362),
	.B(n24358));
   NAND2xp5_ASAP7_75t_SL U20956 (.Y(n24340),
	.A(n27152),
	.B(n27153));
   OAI222xp33_ASAP7_75t_SRAM U20957 (.Y(n24379),
	.A1(FE_OFN28651_FE_OFN26140_n23585),
	.A2(n24377),
	.B1(n24376),
	.B2(n24377),
	.C1(n24375),
	.C2(n24377));
   NAND2xp33_ASAP7_75t_SRAM U20958 (.Y(n24376),
	.A(n24374),
	.B(n24373));
   NAND2xp33_ASAP7_75t_SRAM U20959 (.Y(n24373),
	.A(n24372),
	.B(n24371));
   NAND2xp33_ASAP7_75t_SRAM U20960 (.Y(n24374),
	.A(n24369),
	.B(n24371));
   A2O1A1Ixp33_ASAP7_75t_SL U20961 (.Y(n25761),
	.A1(n24137),
	.A2(n24136),
	.B(n24800),
	.C(n24135));
   O2A1O1Ixp5_ASAP7_75t_SL U20962 (.Y(n24135),
	.A1(n24134),
	.A2(n24133),
	.B(FE_OFN16163_n26584),
	.C(n24132));
   NOR3xp33_ASAP7_75t_L U20964 (.Y(n24130),
	.A(n24129),
	.B(n25082),
	.C(n24128));
   A2O1A1Ixp33_ASAP7_75t_SL U20965 (.Y(n24144),
	.A1(n26282),
	.A2(n24142),
	.B(n24141),
	.C(n24140));
   NAND2xp33_ASAP7_75t_SL U20966 (.Y(n24141),
	.A(FE_OCPN29528_n24138),
	.B(n24149));
   A2O1A1Ixp33_ASAP7_75t_L U20967 (.Y(n24140),
	.A1(n26282),
	.A2(n24142),
	.B(n24139),
	.C(w1_5_));
   NAND2xp5_ASAP7_75t_L U20968 (.Y(n24997),
	.A(FE_OFN28533_n24995),
	.B(n24994));
   A2O1A1Ixp33_ASAP7_75t_R U20970 (.Y(n24311),
	.A1(FE_PSN8300_n26482),
	.A2(n27117),
	.B(FE_PSN8287_FE_OCPN27494_n26479),
	.C(FE_OFN26546_n24537));
   NAND2xp33_ASAP7_75t_L U20971 (.Y(n24312),
	.A(FE_OCPN29263_n24537),
	.B(n26477));
   O2A1O1Ixp33_ASAP7_75t_L U20972 (.Y(n24307),
	.A1(FE_OFN16180_n26542),
	.A2(n26431),
	.B(FE_OCPN27637_n26428),
	.C(n24320));
   NOR2xp33_ASAP7_75t_SL U20975 (.Y(n25857),
	.A(n25856),
	.B(n25855));
   OAI21xp5_ASAP7_75t_SL U20978 (.Y(n26697),
	.A1(n26465),
	.A2(n26464),
	.B(n26463));
   NAND2xp33_ASAP7_75t_R U20980 (.Y(n24445),
	.A(n24444),
	.B(FE_OFN118_sa03_7));
   O2A1O1Ixp33_ASAP7_75t_SRAM U20983 (.Y(n24554),
	.A1(n17463),
	.A2(n24556),
	.B(n24553),
	.C(n25970));
   NOR2xp33_ASAP7_75t_SRAM U20984 (.Y(n24555),
	.A(n25971),
	.B(FE_OFN28934_n24552));
   NAND2xp33_ASAP7_75t_R U20985 (.Y(n24542),
	.A(w0_25_),
	.B(n24540));
   NAND2xp33_ASAP7_75t_R U20987 (.Y(n26110),
	.A(n24515),
	.B(FE_OFN163_sa00_7));
   NOR2xp33_ASAP7_75t_SRAM U20988 (.Y(n24515),
	.A(n25258),
	.B(FE_OFN28499_sa00_6));
   O2A1O1Ixp5_ASAP7_75t_SRAM U20990 (.Y(n24302),
	.A1(n16946),
	.A2(n24300),
	.B(FE_OCPN27544_sa33_4),
	.C(n24299));
   NOR3xp33_ASAP7_75t_SRAM U20991 (.Y(n24303),
	.A(FE_OCPN29577_n24298),
	.B(n24297),
	.C(FE_OCPN28078_n24296));
   NAND2x1_ASAP7_75t_L U20992 (.Y(n25386),
	.A(FE_OCPN27538_n25383),
	.B(FE_OCPN27435_n26790));
   NAND2xp33_ASAP7_75t_SRAM U20993 (.Y(n25381),
	.A(n25378),
	.B(FE_OFN28674_n));
   A2O1A1Ixp33_ASAP7_75t_SL U20995 (.Y(n25936),
	.A1(n27206),
	.A2(FE_OFN16177_n27207),
	.B(FE_OCPN29445_n27203),
	.C(n25935));
   NAND2xp5_ASAP7_75t_SL U20996 (.Y(n25937),
	.A(FE_OCPN29267_n25935),
	.B(n27201));
   NOR2x1_ASAP7_75t_SRAM U20997 (.Y(n25933),
	.A(w2_1_),
	.B(FE_OFN26650_n27164));
   INVxp33_ASAP7_75t_SRAM U20998 (.Y(n25907),
	.A(sa20_7_));
   NAND2xp33_ASAP7_75t_SRAM U20999 (.Y(n25909),
	.A(n25908),
	.B(n25907));
   NOR2xp33_ASAP7_75t_SRAM U21000 (.Y(n25908),
	.A(n25906),
	.B(sa20_6_));
   NOR3x1_ASAP7_75t_SL U21002 (.Y(n27167),
	.A(n25326),
	.B(n25325),
	.C(n25324));
   NAND2xp33_ASAP7_75t_L U21003 (.Y(n25326),
	.A(n25315),
	.B(n25314));
   NOR3xp33_ASAP7_75t_SL U21004 (.Y(n27139),
	.A(n25278),
	.B(n25277),
	.C(n25276));
   NAND3xp33_ASAP7_75t_R U21005 (.Y(n25278),
	.A(FE_OFN28973_n25273),
	.B(n25275),
	.C(n25274));
   NAND2xp5_ASAP7_75t_R U21007 (.Y(n26510),
	.A(FE_OFN26558_n26911),
	.B(n26507));
   NOR2xp33_ASAP7_75t_SL U21008 (.Y(n26515),
	.A(w2_19_),
	.B(n26511));
   NOR2xp33_ASAP7_75t_R U21009 (.Y(n25142),
	.A(FE_OCPN8254_w3_3),
	.B(FE_OFN28902_n25414));
   NOR2xp33_ASAP7_75t_R U21010 (.Y(n25148),
	.A(n25144),
	.B(n25143));
   NAND2xp5_ASAP7_75t_L U21011 (.Y(n25623),
	.A(n26936),
	.B(FE_OCPN27778_n25621));
   INVxp67_ASAP7_75t_SL U21012 (.Y(n26511),
	.A(n26513));
   NAND2x1_ASAP7_75t_SL U21013 (.Y(n25922),
	.A(n25342),
	.B(n25341));
   NAND2xp5_ASAP7_75t_SL U21014 (.Y(n25342),
	.A(n26407),
	.B(n26046));
   INVx1_ASAP7_75t_SL U21015 (.Y(n25341),
	.A(n25340));
   A2O1A1Ixp33_ASAP7_75t_SL U21016 (.Y(n26990),
	.A1(n24802),
	.A2(n24801),
	.B(n24800),
	.C(n24799));
   NOR2xp33_ASAP7_75t_SL U21017 (.Y(n24801),
	.A(FE_OCPN29496_n24789),
	.B(n24788));
   O2A1O1Ixp5_ASAP7_75t_SL U21018 (.Y(n24799),
	.A1(n24798),
	.A2(n24797),
	.B(n26584),
	.C(n24796));
   O2A1O1Ixp33_ASAP7_75t_R U21019 (.Y(n27024),
	.A1(n27027),
	.A2(FE_RN_213_0),
	.B(n27023),
	.C(n27022));
   O2A1O1Ixp33_ASAP7_75t_L U21022 (.Y(n26993),
	.A1(n26926),
	.A2(n26995),
	.B(n26992),
	.C(n26991));
   NAND2xp33_ASAP7_75t_SRAM U21023 (.Y(n26321),
	.A(n26318),
	.B(FE_OFN26019_n26319));
   NOR2xp33_ASAP7_75t_SL U21024 (.Y(n26313),
	.A(w2_3_),
	.B(n26946));
   NOR3x1_ASAP7_75t_L U21025 (.Y(n26776),
	.A(n24095),
	.B(n24094),
	.C(n24093));
   NAND2xp5_ASAP7_75t_L U21027 (.Y(n26768),
	.A(n26764),
	.B(FE_OFN29039_n26763));
   O2A1O1Ixp33_ASAP7_75t_SRAM U21028 (.Y(n26774),
	.A1(n26777),
	.A2(n26776),
	.B(FE_OCPN27935_n26773),
	.C(n26772));
   NAND2xp5_ASAP7_75t_L U21030 (.Y(n26493),
	.A(FE_OFN25911_n26491),
	.B(FE_OFN70_w2_20));
   A2O1A1Ixp33_ASAP7_75t_SL U21031 (.Y(n26492),
	.A1(n27216),
	.A2(n26494),
	.B(FE_OCPN28307_n26491),
	.C(w2_20_));
   O2A1O1Ixp5_ASAP7_75t_L U21032 (.Y(n26497),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(FE_OCPN28119_n26955),
	.C(n26496));
   O2A1O1Ixp33_ASAP7_75t_SL U21033 (.Y(n25807),
	.A1(FE_OFN16180_n26542),
	.A2(n18158),
	.B(n26088),
	.C(n25806));
   NOR2xp33_ASAP7_75t_SL U21034 (.Y(n25808),
	.A(n25805),
	.B(FE_OFN25973_n26087));
   A2O1A1Ixp33_ASAP7_75t_SL U21035 (.Y(n25803),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(FE_OCPN27744_n26362),
	.C(w0_4_));
   NOR3x1_ASAP7_75t_R U21036 (.Y(n26702),
	.A(n26462),
	.B(n26461),
	.C(n26460));
   NAND3xp33_ASAP7_75t_R U21037 (.Y(n26462),
	.A(FE_OCPN29330_n26459),
	.B(n26458),
	.C(n26457));
   NOR2xp33_ASAP7_75t_L U21038 (.Y(n26701),
	.A(w1_20_),
	.B(n26697));
   O2A1O1Ixp5_ASAP7_75t_L U21039 (.Y(n26707),
	.A1(n26710),
	.A2(n26709),
	.B(n26706),
	.C(n26705));
   O2A1O1Ixp5_ASAP7_75t_SL U21040 (.Y(n25721),
	.A1(n26661),
	.A2(n25718),
	.B(n26567),
	.C(n26683));
   NAND3xp33_ASAP7_75t_SL U21041 (.Y(n25718),
	.A(FE_OCPN29548_n25717),
	.B(n25716),
	.C(n25715));
   NOR3xp33_ASAP7_75t_L U21042 (.Y(n25715),
	.A(n25714),
	.B(n26154),
	.C(FE_OCPN27796_n26659));
   NAND2xp33_ASAP7_75t_SRAM U21043 (.Y(n25714),
	.A(n25713),
	.B(n25712));
   NAND2xp33_ASAP7_75t_SRAM U21044 (.Y(n25352),
	.A(FE_OCPN27774_n25351),
	.B(n25350));
   NAND2xp5_ASAP7_75t_SL U21045 (.Y(n24562),
	.A(n22507),
	.B(FE_OCPN7649_n23259));
   NAND2xp33_ASAP7_75t_R U21046 (.Y(n19186),
	.A(n19182),
	.B(n19183));
   NAND2xp33_ASAP7_75t_R U21047 (.Y(n19185),
	.A(n19184),
	.B(n19183));
   NOR3x1_ASAP7_75t_L U21048 (.Y(n25787),
	.A(n17474),
	.B(n23267),
	.C(FE_OCPN27807_n23375));
   NAND3xp33_ASAP7_75t_L U21049 (.Y(n24561),
	.A(n23269),
	.B(n23391),
	.C(n21351));
   NAND2xp33_ASAP7_75t_SRAM U21051 (.Y(n20016),
	.A(FE_OFN28981_n16767),
	.B(FE_OFN16267_sa21_4));
   NAND2xp5_ASAP7_75t_SL U21052 (.Y(n20017),
	.A(n20015),
	.B(n20014));
   NAND2xp5_ASAP7_75t_SL U21053 (.Y(n20015),
	.A(n20010),
	.B(n20012));
   NAND3xp33_ASAP7_75t_R U21054 (.Y(n24266),
	.A(n20312),
	.B(n24918),
	.C(n22348));
   NAND3xp33_ASAP7_75t_L U21055 (.Y(n24267),
	.A(n20002),
	.B(n20001),
	.C(n20296));
   NAND2xp33_ASAP7_75t_SRAM U21056 (.Y(n20001),
	.A(n16771),
	.B(FE_OFN16267_sa21_4));
   NAND3xp33_ASAP7_75t_SL U21057 (.Y(n24252),
	.A(n23668),
	.B(n20326),
	.C(n24921));
   NAND3xp33_ASAP7_75t_R U21058 (.Y(n24253),
	.A(n19993),
	.B(n19992),
	.C(n23654));
   NAND3xp33_ASAP7_75t_SRAM U21059 (.Y(n24272),
	.A(n22703),
	.B(n20327),
	.C(n20300));
   NOR3xp33_ASAP7_75t_SL U21060 (.Y(n23232),
	.A(n23237),
	.B(n23225),
	.C(n23224));
   NAND2xp5_ASAP7_75t_SL U21061 (.Y(n23231),
	.A(n23230),
	.B(n23229));
   NAND2xp33_ASAP7_75t_L U21062 (.Y(n23229),
	.A(n23228),
	.B(n23227));
   NAND3xp33_ASAP7_75t_L U21063 (.Y(n25164),
	.A(n23242),
	.B(n23241),
	.C(n23240));
   NOR3xp33_ASAP7_75t_SRAM U21064 (.Y(n23241),
	.A(n23239),
	.B(n23238),
	.C(n23237));
   NAND2xp33_ASAP7_75t_SRAM U21065 (.Y(n25160),
	.A(n25399),
	.B(n25398));
   NOR3xp33_ASAP7_75t_R U21067 (.Y(n19071),
	.A(n19069),
	.B(n19068),
	.C(n19067));
   NAND2xp33_ASAP7_75t_L U21068 (.Y(n19069),
	.A(n22141),
	.B(n19063));
   NAND3xp33_ASAP7_75t_L U21069 (.Y(n19079),
	.A(n19078),
	.B(n19077),
	.C(n20434));
   NOR3xp33_ASAP7_75t_L U21070 (.Y(n19077),
	.A(n19076),
	.B(n22628),
	.C(n19075));
   NAND2xp33_ASAP7_75t_L U21071 (.Y(n19076),
	.A(n22167),
	.B(n19074));
   OAI222xp33_ASAP7_75t_SL U21072 (.Y(n23290),
	.A1(FE_OCPN29422_n23397),
	.A2(n26078),
	.B1(n23276),
	.B2(n26078),
	.C1(n23275),
	.C2(n26078));
   NOR3xp33_ASAP7_75t_SRAM U21073 (.Y(n23276),
	.A(n23274),
	.B(n23273),
	.C(n23272));
   NAND3xp33_ASAP7_75t_L U21074 (.Y(n23289),
	.A(n23280),
	.B(n23287),
	.C(n23288));
   NAND3xp33_ASAP7_75t_SL U21075 (.Y(n23270),
	.A(FE_OCPN27848_n23255),
	.B(n23254),
	.C(n23253));
   OAI22xp33_ASAP7_75t_L U21076 (.Y(n23253),
	.A1(FE_OCPN28038_n23252),
	.A2(n23251),
	.B1(n17447),
	.B2(n23251));
   NAND3xp33_ASAP7_75t_SL U21077 (.Y(n23251),
	.A(n23250),
	.B(n23249),
	.C(n23248));
   NAND2xp33_ASAP7_75t_L U21078 (.Y(n24564),
	.A(n21375),
	.B(n23380));
   NOR2xp33_ASAP7_75t_SRAM U21079 (.Y(n23277),
	.A(FE_OCPN28006_n17454),
	.B(FE_OCPN29378_n23266));
   NAND2xp5_ASAP7_75t_SL U21080 (.Y(n23256),
	.A(n17499),
	.B(n17498));
   NAND2xp33_ASAP7_75t_SL U21081 (.Y(n17499),
	.A(n17495),
	.B(n17496));
   NAND2xp33_ASAP7_75t_L U21082 (.Y(n17498),
	.A(n17497),
	.B(n17496));
   NOR2x1p5_ASAP7_75t_L U21086 (.Y(n23262),
	.A(n21819),
	.B(n21814));
   NAND2xp33_ASAP7_75t_SRAM U21087 (.Y(n22637),
	.A(n22634),
	.B(n22633));
   NAND2xp33_ASAP7_75t_SRAM U21088 (.Y(n22634),
	.A(n17602),
	.B(FE_OCPN28378_n22632));
   OAI222xp33_ASAP7_75t_R U21089 (.Y(n22649),
	.A1(n22648),
	.A2(n26687),
	.B1(n22647),
	.B2(n26687),
	.C1(n22646),
	.C2(n26687));
   NOR3xp33_ASAP7_75t_SRAM U21090 (.Y(n22648),
	.A(n22642),
	.B(n22641),
	.C(n22640));
   NOR2xp33_ASAP7_75t_L U21091 (.Y(n22647),
	.A(n22645),
	.B(n22644));
   NOR2x1_ASAP7_75t_L U21093 (.Y(n22614),
	.A(n18473),
	.B(FE_OFN29121_n26026));
   NOR2x1_ASAP7_75t_R U21094 (.Y(n22615),
	.A(n18368),
	.B(FE_OCPN27764_n22152));
   NOR2x1_ASAP7_75t_L U21095 (.Y(n23324),
	.A(n22287),
	.B(n21125));
   NOR2xp33_ASAP7_75t_R U21097 (.Y(n23344),
	.A(n23342),
	.B(n20748));
   NAND2xp5_ASAP7_75t_L U21098 (.Y(n23349),
	.A(n23334),
	.B(n23333));
   NAND3xp33_ASAP7_75t_L U21099 (.Y(n23348),
	.A(n23341),
	.B(n23339),
	.C(FE_PSN8336_n23340));
   NOR2xp33_ASAP7_75t_SL U21100 (.Y(n23338),
	.A(FE_OCPN27721_n23336),
	.B(n23335));
   NAND3xp33_ASAP7_75t_L U21101 (.Y(n23298),
	.A(n23172),
	.B(n18198),
	.C(n21118));
   NAND2xp33_ASAP7_75t_SRAM U21102 (.Y(n18198),
	.A(n22828),
	.B(FE_OFN27173_n));
   NOR2xp33_ASAP7_75t_R U21103 (.Y(n23299),
	.A(FE_RN_0_0),
	.B(n21107));
   INVxp33_ASAP7_75t_SRAM U21104 (.Y(n23301),
	.A(n23300));
   NOR2x1_ASAP7_75t_L U21105 (.Y(n22715),
	.A(FE_OFN27179_n20327),
	.B(n17855));
   NAND3xp33_ASAP7_75t_SL U21106 (.Y(n17855),
	.A(n25355),
	.B(n24919),
	.C(n22346));
   NOR3x1_ASAP7_75t_L U21107 (.Y(n24268),
	.A(n19978),
	.B(n19977),
	.C(n20288));
   NOR3xp33_ASAP7_75t_SRAM U21110 (.Y(n22702),
	.A(n22693),
	.B(n22692),
	.C(FE_OFN26038_n24887));
   NAND2xp33_ASAP7_75t_SRAM U21111 (.Y(n22699),
	.A(n22698),
	.B(n22697));
   NAND2xp5_ASAP7_75t_L U21112 (.Y(n16673),
	.A(FE_OCPN29487_FE_OFN28694_sa33_4),
	.B(FE_OFN27062_n16438));
   NAND3xp33_ASAP7_75t_L U21113 (.Y(n16485),
	.A(n16730),
	.B(n16467),
	.C(n16679));
   NOR3xp33_ASAP7_75t_L U21115 (.Y(n16482),
	.A(n16481),
	.B(n17415),
	.C(n16480));
   NOR3xp33_ASAP7_75t_SL U21116 (.Y(n16483),
	.A(n16478),
	.B(n16938),
	.C(n16477));
   NAND2xp33_ASAP7_75t_SRAM U21117 (.Y(n16481),
	.A(n16726),
	.B(n23550));
   NAND3xp33_ASAP7_75t_SL U21118 (.Y(n16452),
	.A(n23533),
	.B(FE_OCPN29561_n23532),
	.C(n23562));
   NOR2xp33_ASAP7_75t_SL U21119 (.Y(n16841),
	.A(n18421),
	.B(n17405));
   NAND3xp33_ASAP7_75t_SL U21121 (.Y(n23761),
	.A(n21196),
	.B(n23871),
	.C(n23720));
   NOR2xp33_ASAP7_75t_SL U21122 (.Y(n23782),
	.A(n23892),
	.B(n23780));
   NAND2xp5_ASAP7_75t_L U21123 (.Y(n23780),
	.A(n23779),
	.B(n23778));
   NOR2xp33_ASAP7_75t_L U21124 (.Y(n23783),
	.A(n23841),
	.B(n23775));
   NAND2xp5_ASAP7_75t_SL U21125 (.Y(n23770),
	.A(n23769),
	.B(n23768));
   NAND2xp5_ASAP7_75t_SL U21126 (.Y(n23741),
	.A(n23700),
	.B(n23699));
   NOR2xp33_ASAP7_75t_L U21127 (.Y(n23744),
	.A(FE_OFN28729_n20617),
	.B(n23745));
   INVxp33_ASAP7_75t_L U21128 (.Y(n23746),
	.A(n23743));
   NAND2xp33_ASAP7_75t_L U21129 (.Y(n23748),
	.A(n23747),
	.B(n23746));
   NOR2xp33_ASAP7_75t_L U21130 (.Y(n23747),
	.A(FE_OFN28869_FE_OCPN27715_n23875),
	.B(n23745));
   OAI22xp33_ASAP7_75t_L U21131 (.Y(n17728),
	.A1(n17527),
	.A2(n24868),
	.B1(n18847),
	.B2(n24868));
   AND3x1_ASAP7_75t_SRAM U21132 (.Y(n17731),
	.A(n18335),
	.B(n18329),
	.C(n18825));
   NAND2xp5_ASAP7_75t_SL U21134 (.Y(n17043),
	.A(FE_OFN26572_n19405),
	.B(n20492));
   NAND2xp5_ASAP7_75t_SL U21135 (.Y(n17149),
	.A(n16987),
	.B(n16986));
   NOR2xp33_ASAP7_75t_SRAM U21136 (.Y(n16987),
	.A(n19409),
	.B(n17027));
   NOR3xp33_ASAP7_75t_SL U21137 (.Y(n16986),
	.A(n16985),
	.B(n20502),
	.C(n25225));
   NOR2x1_ASAP7_75t_SL U21138 (.Y(n25204),
	.A(n22900),
	.B(n22899));
   NOR2xp33_ASAP7_75t_SRAM U21139 (.Y(n25206),
	.A(FE_OCPN27652_n20176),
	.B(n22871));
   NAND2xp5_ASAP7_75t_SL U21140 (.Y(n25202),
	.A(n20200),
	.B(n19263));
   NAND3xp33_ASAP7_75t_SL U21141 (.Y(n25211),
	.A(n22086),
	.B(n17772),
	.C(n19274));
   NAND3xp33_ASAP7_75t_SL U21142 (.Y(n19747),
	.A(FE_OFN28535_n19738),
	.B(n19737),
	.C(n22401));
   NOR2xp33_ASAP7_75t_SRAM U21144 (.Y(n19745),
	.A(n19740),
	.B(n19739));
   NOR2xp33_ASAP7_75t_SL U21145 (.Y(n19744),
	.A(n24998),
	.B(n19742));
   NAND3xp33_ASAP7_75t_SL U21146 (.Y(n19742),
	.A(n22378),
	.B(n19741),
	.C(n25024));
   NAND3xp33_ASAP7_75t_R U21147 (.Y(n19748),
	.A(n19727),
	.B(n19951),
	.C(n19726));
   NAND2xp33_ASAP7_75t_SRAM U21148 (.Y(n19727),
	.A(n19725),
	.B(n17529));
   NAND3xp33_ASAP7_75t_L U21149 (.Y(n19724),
	.A(n19719),
	.B(FE_OFN28965_n24869),
	.C(n19718));
   NAND2xp33_ASAP7_75t_SRAM U21150 (.Y(n19719),
	.A(n19717),
	.B(n19716));
   NAND2xp33_ASAP7_75t_R U21151 (.Y(n19716),
	.A(n19715),
	.B(n19714));
   NAND2xp33_ASAP7_75t_R U21152 (.Y(n19717),
	.A(n19711),
	.B(n19714));
   NAND2x1_ASAP7_75t_SL U21153 (.Y(n19701),
	.A(n24861),
	.B(n17678));
   NAND3xp33_ASAP7_75t_SL U21156 (.Y(n20919),
	.A(n20933),
	.B(FE_OCPN29480_n20913),
	.C(FE_OCPN27482_sa23_5));
   NOR3xp33_ASAP7_75t_SL U21157 (.Y(n20944),
	.A(n23484),
	.B(n20942),
	.C(n23479));
   NAND3xp33_ASAP7_75t_R U21158 (.Y(n20946),
	.A(n22022),
	.B(n20929),
	.C(n23475));
   NOR2xp33_ASAP7_75t_R U21159 (.Y(n20929),
	.A(n19341),
	.B(FE_OFN29151_n22988));
   NAND2xp33_ASAP7_75t_R U21160 (.Y(n20947),
	.A(n20923),
	.B(n26159));
   NAND2xp5_ASAP7_75t_L U21161 (.Y(n22999),
	.A(n20916),
	.B(n22007));
   A2O1A1Ixp33_ASAP7_75t_L U21162 (.Y(n24042),
	.A1(n19352),
	.A2(n19351),
	.B(n26571),
	.C(n19350));
   NOR3xp33_ASAP7_75t_SRAM U21163 (.Y(n19352),
	.A(n25711),
	.B(FE_PSN8328_n20260),
	.C(n25093));
   NOR3xp33_ASAP7_75t_SL U21164 (.Y(n19351),
	.A(n19336),
	.B(n22923),
	.C(n19335));
   OAI21xp5_ASAP7_75t_L U21165 (.Y(n19350),
	.A1(n19341),
	.A2(n19349),
	.B(n26567));
   NAND3xp33_ASAP7_75t_SRAM U21166 (.Y(n24044),
	.A(n20926),
	.B(n26146),
	.C(n20943));
   NOR2x1_ASAP7_75t_SL U21167 (.Y(n25097),
	.A(n22048),
	.B(n19302));
   NAND3xp33_ASAP7_75t_R U21168 (.Y(n20250),
	.A(FE_OCPN29331_n20933),
	.B(FE_OFN29026_n20911),
	.C(FE_OFN27078_sa23_5));
   NAND3xp33_ASAP7_75t_L U21169 (.Y(n20180),
	.A(n20167),
	.B(n20166),
	.C(n25299));
   NAND2xp5_ASAP7_75t_R U21170 (.Y(n20167),
	.A(n20151),
	.B(n20150));
   NAND2xp5_ASAP7_75t_SL U21171 (.Y(n20166),
	.A(n20160),
	.B(n20159));
   NAND2xp33_ASAP7_75t_R U21172 (.Y(n20150),
	.A(FE_OCPN27579_FE_OFN16138_sa02_5),
	.B(n21004));
   NOR3xp33_ASAP7_75t_SRAM U21174 (.Y(n20177),
	.A(n22881),
	.B(FE_OCPN27972_n20988),
	.C(FE_OCPN27652_n20176));
   NOR3xp33_ASAP7_75t_SL U21175 (.Y(n20178),
	.A(n25277),
	.B(n22565),
	.C(n20175));
   NAND2xp33_ASAP7_75t_SL U21176 (.Y(n20148),
	.A(n20143),
	.B(n20145));
   NAND2xp33_ASAP7_75t_SL U21177 (.Y(n20147),
	.A(n20146),
	.B(n20145));
   OAI21xp33_ASAP7_75t_L U21178 (.Y(n20135),
	.A1(FE_OCPN27574_n20196),
	.A2(FE_OFN28961_n17744),
	.B(n20954));
   NAND3xp33_ASAP7_75t_L U21179 (.Y(n20127),
	.A(n20170),
	.B(FE_OCPN27634_n20169),
	.C(FE_OFN26159_n22080));
   NAND3xp33_ASAP7_75t_SL U21180 (.Y(n25201),
	.A(n19259),
	.B(FE_OCPN28303_n20961),
	.C(n20960));
   NAND2xp5_ASAP7_75t_L U21181 (.Y(n20139),
	.A(n22876),
	.B(n20130));
   NOR2xp33_ASAP7_75t_SL U21182 (.Y(n20130),
	.A(n20129),
	.B(n22060));
   NAND2xp33_ASAP7_75t_SL U21183 (.Y(n22904),
	.A(n25502),
	.B(n22542));
   NOR2xp33_ASAP7_75t_L U21184 (.Y(n22542),
	.A(n25530),
	.B(n22541));
   NOR2xp33_ASAP7_75t_SRAM U21185 (.Y(n22545),
	.A(FE_OCPN29318_n25524),
	.B(n25523));
   NAND2xp33_ASAP7_75t_SRAM U21186 (.Y(n22544),
	.A(FE_PSN8323_n22543),
	.B(FE_OCPN27384_n22888));
   NAND3xp33_ASAP7_75t_SL U21187 (.Y(n22569),
	.A(n22568),
	.B(n22567),
	.C(n22566));
   NOR3xp33_ASAP7_75t_SRAM U21188 (.Y(n22568),
	.A(n22562),
	.B(n22561),
	.C(FE_OCPN27424_n22560));
   NOR3xp33_ASAP7_75t_L U21190 (.Y(n22567),
	.A(n25217),
	.B(n22564),
	.C(n22563));
   NAND2xp5_ASAP7_75t_L U21191 (.Y(n22541),
	.A(n22535),
	.B(n22534));
   NOR2xp33_ASAP7_75t_L U21192 (.Y(n22535),
	.A(n22533),
	.B(n22561));
   NAND3xp33_ASAP7_75t_SL U21193 (.Y(n22536),
	.A(n20142),
	.B(n20141),
	.C(n20203));
   NOR3xp33_ASAP7_75t_SRAM U21194 (.Y(n20141),
	.A(n20186),
	.B(n20136),
	.C(n20176));
   NOR2xp33_ASAP7_75t_SRAM U21195 (.Y(n22531),
	.A(n22527),
	.B(FE_OFN28800_n22526));
   NAND2xp33_ASAP7_75t_R U21196 (.Y(n22303),
	.A(n22289),
	.B(n22300));
   NOR2xp33_ASAP7_75t_SL U21197 (.Y(n22289),
	.A(n23346),
	.B(sa22_6_));
   NAND2xp5_ASAP7_75t_L U21198 (.Y(n22302),
	.A(n22301),
	.B(n22300));
   NOR2xp33_ASAP7_75t_SL U21199 (.Y(n22301),
	.A(n22299),
	.B(sa22_6_));
   NOR3xp33_ASAP7_75t_SL U21200 (.Y(n22299),
	.A(n22298),
	.B(n23297),
	.C(n22297));
   NAND2xp33_ASAP7_75t_L U21201 (.Y(n22297),
	.A(n23187),
	.B(n22296));
   NOR3xp33_ASAP7_75t_SL U21202 (.Y(n22316),
	.A(n22309),
	.B(n23200),
	.C(n22308));
   NOR3xp33_ASAP7_75t_R U21203 (.Y(n22314),
	.A(FE_OFN28930_n22836),
	.B(n23161),
	.C(FE_OFN16203_n22313));
   NAND3xp33_ASAP7_75t_SRAM U21204 (.Y(n22315),
	.A(FE_OFN28798_FE_OCPN27947_n18177),
	.B(FE_PSN8294_n22310),
	.C(FE_OCPN27673_n18163));
   NOR3xp33_ASAP7_75t_L U21205 (.Y(n22323),
	.A(n23342),
	.B(n22320),
	.C(n22319));
   NAND2xp33_ASAP7_75t_L U21206 (.Y(n22286),
	.A(n22272),
	.B(n22271));
   NAND2xp33_ASAP7_75t_SRAM U21208 (.Y(n19761),
	.A(n19796),
	.B(n19759));
   NAND2xp33_ASAP7_75t_SRAM U21209 (.Y(n19760),
	.A(n19798),
	.B(n19759));
   NOR2xp33_ASAP7_75t_L U21210 (.Y(n19753),
	.A(n23982),
	.B(FE_OFN28832_n19789));
   NAND2xp33_ASAP7_75t_SRAM U21211 (.Y(n24895),
	.A(n21885),
	.B(n23128));
   NOR2x1_ASAP7_75t_L U21212 (.Y(n24671),
	.A(n19786),
	.B(n19785));
   NAND3xp33_ASAP7_75t_L U21213 (.Y(n19786),
	.A(n19783),
	.B(n19782),
	.C(n19781));
   OAI22xp33_ASAP7_75t_SRAM U21214 (.Y(n19783),
	.A1(n24959),
	.A2(FE_OCPN28157_n16534),
	.B1(n24955),
	.B2(FE_OCPN28157_n16534));
   NOR2xp33_ASAP7_75t_SRAM U21216 (.Y(n20695),
	.A(n20678),
	.B(n23724));
   NAND3xp33_ASAP7_75t_SL U21218 (.Y(n20697),
	.A(n20677),
	.B(n20676),
	.C(n23779));
   NAND2xp5_ASAP7_75t_R U21219 (.Y(n20676),
	.A(n20673),
	.B(n20672));
   NAND2xp33_ASAP7_75t_L U21220 (.Y(n20677),
	.A(n20665),
	.B(n20664));
   NAND2xp33_ASAP7_75t_L U21221 (.Y(n20672),
	.A(n20671),
	.B(n20667));
   NOR2xp33_ASAP7_75t_SRAM U21222 (.Y(n20650),
	.A(FE_OFN28868_FE_OCPN27715_n23875),
	.B(n23763));
   NOR3xp33_ASAP7_75t_SL U21224 (.Y(n20658),
	.A(n20657),
	.B(FE_OFN27088_n23754),
	.C(FE_OCPN5147_n18548));
   NAND2xp33_ASAP7_75t_L U21225 (.Y(n20616),
	.A(n20613),
	.B(n20693));
   NAND2xp5_ASAP7_75t_SL U21228 (.Y(n22212),
	.A(n22211),
	.B(n22210));
   NAND2xp5_ASAP7_75t_L U21229 (.Y(n22211),
	.A(n22207),
	.B(n22208));
   NAND3xp33_ASAP7_75t_L U21230 (.Y(n22215),
	.A(n22204),
	.B(n22203),
	.C(n22202));
   NAND2xp33_ASAP7_75t_L U21232 (.Y(n22203),
	.A(n22201),
	.B(n22200));
   NAND2xp33_ASAP7_75t_SRAM U21233 (.Y(n22201),
	.A(n22195),
	.B(n22198));
   NAND2xp33_ASAP7_75t_SRAM U21235 (.Y(n22188),
	.A(n22184),
	.B(n22183));
   NAND3xp33_ASAP7_75t_SL U21236 (.Y(n22216),
	.A(n23074),
	.B(n20398),
	.C(n20397));
   NOR3xp33_ASAP7_75t_L U21237 (.Y(n20398),
	.A(n20396),
	.B(n22436),
	.C(n23075));
   OAI22xp33_ASAP7_75t_SRAM U21239 (.Y(n22190),
	.A1(n23059),
	.A2(n22189),
	.B1(n17331),
	.B2(n22189));
   INVxp33_ASAP7_75t_L U21241 (.Y(n22179),
	.A(n22178));
   NOR2xp33_ASAP7_75t_SRAM U21242 (.Y(n22184),
	.A(n21546),
	.B(n21545));
   NAND3xp33_ASAP7_75t_L U21243 (.Y(n22422),
	.A(n21553),
	.B(FE_OCPN8219_n22197),
	.C(n17326));
   NAND3xp33_ASAP7_75t_SL U21244 (.Y(n21575),
	.A(n21557),
	.B(n25057),
	.C(n22202));
   NAND2xp33_ASAP7_75t_R U21245 (.Y(n21576),
	.A(n21552),
	.B(n12999));
   NOR2xp33_ASAP7_75t_SRAM U21246 (.Y(n12999),
	.A(FE_OFN29135_n21551),
	.B(n23099));
   NOR3xp33_ASAP7_75t_SL U21248 (.Y(n19613),
	.A(n19612),
	.B(n19611),
	.C(n19610));
   NAND3xp33_ASAP7_75t_R U21249 (.Y(n19617),
	.A(n19608),
	.B(n19607),
	.C(n21177));
   NOR3xp33_ASAP7_75t_SRAM U21250 (.Y(n19608),
	.A(n19600),
	.B(FE_OFN26644_n19599),
	.C(n21444));
   NAND3xp33_ASAP7_75t_R U21252 (.Y(n19618),
	.A(n19592),
	.B(n21152),
	.C(n19591));
   NAND2x1_ASAP7_75t_SL U21253 (.Y(n19588),
	.A(n18766),
	.B(n17264));
   NAND2xp5_ASAP7_75t_L U21254 (.Y(n17264),
	.A(FE_OCPN27908_FE_OFN16156_sa00_2),
	.B(FE_OCPN27703_n19847));
   NOR3xp33_ASAP7_75t_SRAM U21255 (.Y(n18630),
	.A(n21477),
	.B(n18746),
	.C(n18628));
   NOR3xp33_ASAP7_75t_SL U21258 (.Y(n18658),
	.A(n18657),
	.B(n18656),
	.C(n19145));
   OAI21xp33_ASAP7_75t_R U21259 (.Y(n18657),
	.A1(n19097),
	.A2(FE_OCPN28270_n17237),
	.B(n19131));
   NAND3xp33_ASAP7_75t_L U21260 (.Y(n18661),
	.A(n18649),
	.B(n18652),
	.C(n18653));
   NAND2xp33_ASAP7_75t_R U21261 (.Y(n18647),
	.A(n18646),
	.B(n18645));
   NAND3x1_ASAP7_75t_L U21262 (.Y(n19611),
	.A(n18763),
	.B(n18643),
	.C(n18642));
   NOR3xp33_ASAP7_75t_L U21263 (.Y(n18643),
	.A(FE_PSN8284_n21438),
	.B(n19593),
	.C(n19139));
   NOR3xp33_ASAP7_75t_L U21264 (.Y(n25642),
	.A(n23799),
	.B(n23798),
	.C(n23797));
   NOR3xp33_ASAP7_75t_SL U21265 (.Y(n25643),
	.A(n23807),
	.B(FE_OCPN29567_n23806),
	.C(n23805));
   NAND2xp33_ASAP7_75t_SL U21266 (.Y(n23805),
	.A(n23804),
	.B(n23803));
   NAND3xp33_ASAP7_75t_SL U21267 (.Y(n25638),
	.A(n23828),
	.B(n23827),
	.C(n25329));
   NAND2xp33_ASAP7_75t_R U21268 (.Y(n23828),
	.A(n23818),
	.B(n23817));
   NAND2xp33_ASAP7_75t_SL U21269 (.Y(n23827),
	.A(n23826),
	.B(n23825));
   NAND2xp33_ASAP7_75t_R U21270 (.Y(n23818),
	.A(n23813),
	.B(n23815));
   NOR3xp33_ASAP7_75t_SL U21272 (.Y(n23845),
	.A(n25627),
	.B(n25632),
	.C(n25631));
   NAND3xp33_ASAP7_75t_SRAM U21273 (.Y(n25639),
	.A(n23811),
	.B(n23810),
	.C(n23809));
   NAND3xp33_ASAP7_75t_R U21274 (.Y(n25634),
	.A(n23794),
	.B(n23793),
	.C(n25901));
   NAND3xp33_ASAP7_75t_SL U21275 (.Y(n24064),
	.A(n20590),
	.B(n22226),
	.C(n25442));
   NAND3xp33_ASAP7_75t_L U21276 (.Y(n24065),
	.A(n20582),
	.B(n20581),
	.C(n20580));
   NAND2xp33_ASAP7_75t_SRAM U21277 (.Y(n20581),
	.A(FE_OCPN27729_n24362),
	.B(FE_OCPN28386_n17899));
   NAND2xp33_ASAP7_75t_L U21278 (.Y(n20582),
	.A(n20578),
	.B(n20577));
   NAND2xp33_ASAP7_75t_SRAM U21279 (.Y(n20570),
	.A(n20567),
	.B(n20566));
   NOR2xp33_ASAP7_75t_SRAM U21280 (.Y(n20568),
	.A(FE_OCPN27729_n24362),
	.B(n24381));
   OAI21xp33_ASAP7_75t_SRAM U21282 (.Y(n24053),
	.A1(n20555),
	.A2(n20554),
	.B(n23609));
   NAND2xp33_ASAP7_75t_SRAM U21283 (.Y(n16630),
	.A(n19766),
	.B(n19641));
   NOR3xp33_ASAP7_75t_SL U21284 (.Y(n16665),
	.A(n16664),
	.B(n24458),
	.C(n24894));
   NAND3xp33_ASAP7_75t_SL U21285 (.Y(n16664),
	.A(n16662),
	.B(n19644),
	.C(n16661));
   NAND2xp5_ASAP7_75t_L U21286 (.Y(n16662),
	.A(n16660),
	.B(n16659));
   NAND3xp33_ASAP7_75t_SL U21287 (.Y(n16667),
	.A(n23140),
	.B(n19782),
	.C(n16652));
   NAND3xp33_ASAP7_75t_L U21288 (.Y(n16668),
	.A(n16639),
	.B(n19647),
	.C(n16638));
   OAI22xp33_ASAP7_75t_SRAM U21289 (.Y(n16639),
	.A1(n23980),
	.A2(n23119),
	.B1(n19630),
	.B2(n23119));
   NAND2xp33_ASAP7_75t_SL U21290 (.Y(n16635),
	.A(n16580),
	.B(n16579));
   NOR2xp33_ASAP7_75t_L U21291 (.Y(n16579),
	.A(n23996),
	.B(n16578));
   NAND2xp33_ASAP7_75t_SRAM U21292 (.Y(n16578),
	.A(n23120),
	.B(n23028));
   NOR2x1p5_ASAP7_75t_L U21293 (.Y(n23148),
	.A(FE_OFN26161_sa10_4),
	.B(n16581));
   NOR2xp33_ASAP7_75t_SRAM U21295 (.Y(n16613),
	.A(FE_OCPN28040_n19766),
	.B(n21906));
   NAND2xp33_ASAP7_75t_L U21296 (.Y(n16615),
	.A(n16611),
	.B(n16612));
   NOR2xp33_ASAP7_75t_R U21297 (.Y(n16611),
	.A(n23980),
	.B(n21906));
   NOR2xp33_ASAP7_75t_SL U21298 (.Y(n23438),
	.A(n21740),
	.B(n21058));
   OA21x2_ASAP7_75t_L U21299 (.Y(n21076),
	.A1(n21073),
	.A2(n21072),
	.B(n21742));
   NOR2xp33_ASAP7_75t_SRAM U21300 (.Y(n21066),
	.A(FE_OCPN27675_n17986),
	.B(FE_OCPN29314_n));
   NOR3xp33_ASAP7_75t_SL U21302 (.Y(n21065),
	.A(n21062),
	.B(n21754),
	.C(n24440));
   NOR2xp33_ASAP7_75t_R U21303 (.Y(n21063),
	.A(FE_OCPN7584_n23447),
	.B(n21735));
   NOR3xp33_ASAP7_75t_SL U21304 (.Y(n21298),
	.A(n21013),
	.B(n21043),
	.C(FE_OCPN27918_n21042));
   OAI21xp5_ASAP7_75t_L U21305 (.Y(n21013),
	.A1(FE_OCPN27998_n18019),
	.A2(FE_OFN28677_n17998),
	.B(n21046));
   NAND3x1_ASAP7_75t_SL U21306 (.Y(n21754),
	.A(n21026),
	.B(n21025),
	.C(n21024));
   NOR3xp33_ASAP7_75t_SL U21307 (.Y(n21025),
	.A(n21509),
	.B(n18008),
	.C(n21023));
   NAND3xp33_ASAP7_75t_L U21308 (.Y(n23464),
	.A(n23458),
	.B(n23463),
	.C(n23462));
   NOR3xp33_ASAP7_75t_SL U21309 (.Y(n23463),
	.A(n23461),
	.B(n23460),
	.C(n23459));
   NOR3xp33_ASAP7_75t_SRAM U21311 (.Y(n23452),
	.A(FE_OCPN5072_n23451),
	.B(n23450),
	.C(n23449));
   NOR3xp33_ASAP7_75t_SL U21312 (.Y(n23453),
	.A(n23448),
	.B(n23447),
	.C(n23446));
   OAI21xp33_ASAP7_75t_SRAM U21313 (.Y(n23446),
	.A1(FE_OCPN27733_n17996),
	.A2(FE_OFN28677_n17998),
	.B(n23444));
   NAND2xp33_ASAP7_75t_SRAM U21314 (.Y(n23437),
	.A(n23433),
	.B(n23435));
   NAND2xp33_ASAP7_75t_SRAM U21315 (.Y(n23436),
	.A(n17992),
	.B(n23435));
   NOR2xp33_ASAP7_75t_SRAM U21316 (.Y(n23425),
	.A(FE_OCPN27675_n17986),
	.B(FE_OFN27133_n21725));
   OAI21xp33_ASAP7_75t_SRAM U21317 (.Y(n23422),
	.A1(FE_OFN28677_n17998),
	.A2(FE_OCPN29283_n23439),
	.B(FE_OCPN28297_n23417));
   NAND2xp33_ASAP7_75t_SRAM U21318 (.Y(n23421),
	.A(n23419),
	.B(n23418));
   NAND2xp33_ASAP7_75t_SL U21319 (.Y(n21749),
	.A(n21745),
	.B(n21744));
   NAND2xp5_ASAP7_75t_L U21320 (.Y(n21744),
	.A(n21743),
	.B(n21742));
   NAND2xp5_ASAP7_75t_L U21321 (.Y(n21745),
	.A(n21739),
	.B(n21742));
   NOR3xp33_ASAP7_75t_SRAM U21322 (.Y(n21748),
	.A(n23443),
	.B(n21747),
	.C(n21746));
   NOR3xp33_ASAP7_75t_SRAM U21323 (.Y(n21736),
	.A(n21735),
	.B(FE_OCPN28431_n21734),
	.C(n21733));
   NOR3xp33_ASAP7_75t_L U21324 (.Y(n21757),
	.A(n21756),
	.B(FE_OFN29175_n21755),
	.C(n21754));
   NOR3xp33_ASAP7_75t_SRAM U21325 (.Y(n21758),
	.A(n21753),
	.B(n21752),
	.C(n21751));
   NAND3xp33_ASAP7_75t_L U21326 (.Y(n23459),
	.A(n21719),
	.B(n21718),
	.C(n24241));
   OAI21xp5_ASAP7_75t_SL U21327 (.Y(n23448),
	.A1(FE_OFN28886_FE_OCPN27675_n17986),
	.A2(FE_OCPN29283_n23439),
	.B(n21717));
   NOR3xp33_ASAP7_75t_SL U21328 (.Y(n21717),
	.A(n21716),
	.B(n21729),
	.C(n21715));
   NAND3xp33_ASAP7_75t_SL U21329 (.Y(n21716),
	.A(n23419),
	.B(n23418),
	.C(n21714));
   NOR2x1_ASAP7_75t_L U21330 (.Y(n21707),
	.A(n18875),
	.B(FE_OFN28949_n18011));
   NOR2x1_ASAP7_75t_L U21331 (.Y(n21711),
	.A(FE_OCPN27611_n23426),
	.B(n21296));
   NOR3xp33_ASAP7_75t_SL U21332 (.Y(n26457),
	.A(n20388),
	.B(n20387),
	.C(n22194));
   NOR3x1_ASAP7_75t_SL U21333 (.Y(n25069),
	.A(n20416),
	.B(n26461),
	.C(n26460));
   NAND3xp33_ASAP7_75t_SL U21334 (.Y(n20416),
	.A(n26459),
	.B(n20414),
	.C(FE_OCPN28305_n26451));
   NAND2xp33_ASAP7_75t_L U21335 (.Y(n20414),
	.A(n20413),
	.B(n20412));
   NAND2xp33_ASAP7_75t_SRAM U21336 (.Y(n20413),
	.A(n20408),
	.B(n20410));
   AND3x1_ASAP7_75t_SL U21337 (.Y(n20381),
	.A(n25065),
	.B(n25062),
	.C(n25060));
   NAND3xp33_ASAP7_75t_R U21338 (.Y(n20086),
	.A(n20863),
	.B(n20072),
	.C(n20071));
   NAND3x1_ASAP7_75t_SL U21340 (.Y(n20047),
	.A(n16407),
	.B(n16406),
	.C(n16405));
   NAND2xp5_ASAP7_75t_L U21341 (.Y(n16403),
	.A(n16402),
	.B(n16401));
   NAND2xp5_ASAP7_75t_L U21342 (.Y(n16404),
	.A(n16400),
	.B(n16401));
   OAI21xp5_ASAP7_75t_L U21343 (.Y(n20049),
	.A1(n20853),
	.A2(FE_OCPN28008_n16290),
	.B(n16350));
   NAND2xp33_ASAP7_75t_R U21344 (.Y(n20063),
	.A(n20058),
	.B(n21975));
   NAND2xp33_ASAP7_75t_SRAM U21345 (.Y(n20062),
	.A(n20061),
	.B(n21975));
   NAND3xp33_ASAP7_75t_SL U21346 (.Y(n26399),
	.A(FE_OFN29016_n16512),
	.B(FE_OCPN27444_n20064),
	.C(FE_OCPN29483_FE_OFN26014_sa31_3));
   NOR3xp33_ASAP7_75t_L U21347 (.Y(n26406),
	.A(n18066),
	.B(FE_OCPN27316_n25849),
	.C(n20043));
   NAND2xp5_ASAP7_75t_SL U21348 (.Y(n26409),
	.A(n18083),
	.B(n16500));
   NOR3xp33_ASAP7_75t_SL U21349 (.Y(n16500),
	.A(n21928),
	.B(n16499),
	.C(n16498));
   NAND2xp33_ASAP7_75t_R U21351 (.Y(n20349),
	.A(n20348),
	.B(n20347));
   NAND2xp5_ASAP7_75t_SL U21352 (.Y(n20350),
	.A(n20343),
	.B(n20342));
   NAND2xp33_ASAP7_75t_R U21353 (.Y(n20347),
	.A(n22681),
	.B(n20346));
   NAND2xp33_ASAP7_75t_L U21354 (.Y(n22688),
	.A(n20324),
	.B(n20323));
   NAND2xp5_ASAP7_75t_R U21355 (.Y(n20321),
	.A(n20320),
	.B(n20319));
   NAND2xp5_ASAP7_75t_L U21356 (.Y(n16704),
	.A(n16700),
	.B(n16701));
   NAND2xp5_ASAP7_75t_L U21357 (.Y(n16703),
	.A(n16702),
	.B(n16701));
   OAI21xp5_ASAP7_75t_SL U21358 (.Y(n16731),
	.A1(n16860),
	.A2(n16739),
	.B(n26770));
   NOR3x1_ASAP7_75t_SL U21359 (.Y(n24296),
	.A(n16676),
	.B(FE_OFN26055_n),
	.C(n16847));
   NOR2x1p5_ASAP7_75t_L U21360 (.Y(n24297),
	.A(FE_OCPN29391_FE_OFN29162_sa33_2),
	.B(n16953));
   NAND3xp33_ASAP7_75t_L U21361 (.Y(n24299),
	.A(n16737),
	.B(n16674),
	.C(n16846));
   NOR2xp33_ASAP7_75t_L U21362 (.Y(n16674),
	.A(n18431),
	.B(n16723));
   NOR2xp33_ASAP7_75t_SL U21364 (.Y(n24010),
	.A(n20102),
	.B(n20101));
   NOR2xp33_ASAP7_75t_SL U21365 (.Y(n18922),
	.A(n17115),
	.B(n20526));
   NOR2x1_ASAP7_75t_L U21366 (.Y(n22095),
	.A(n17765),
	.B(FE_OCPN29545_n22529));
   NOR3x1_ASAP7_75t_SL U21367 (.Y(n22105),
	.A(n26968),
	.B(n20168),
	.C(n25530));
   INVxp33_ASAP7_75t_L U21368 (.Y(n17785),
	.A(n17784));
   NOR3xp33_ASAP7_75t_L U21369 (.Y(n17786),
	.A(n17783),
	.B(n22894),
	.C(n22532));
   A2O1A1Ixp33_ASAP7_75t_SL U21370 (.Y(n17818),
	.A1(n17817),
	.A2(n17816),
	.B(n27140),
	.C(FE_OCPN27773_n22070));
   NOR3xp33_ASAP7_75t_L U21371 (.Y(n17817),
	.A(FE_OCPN28196_n22547),
	.B(n20995),
	.C(n20138));
   NOR3xp33_ASAP7_75t_SL U21372 (.Y(n17816),
	.A(n17814),
	.B(n20957),
	.C(n21001));
   NOR3xp33_ASAP7_75t_L U21374 (.Y(n17778),
	.A(n22899),
	.B(n20186),
	.C(n20995));
   NAND3xp33_ASAP7_75t_SL U21375 (.Y(n25212),
	.A(n20955),
	.B(n22069),
	.C(FE_OCPN27773_n22070));
   NOR3x1_ASAP7_75t_SL U21376 (.Y(n25524),
	.A(n17771),
	.B(FE_OFN28665_FE_OCPN27566),
	.C(FE_OFN29184_n17744));
   NOR2x1_ASAP7_75t_R U21377 (.Y(n25523),
	.A(n20195),
	.B(n17780));
   NOR3xp33_ASAP7_75t_R U21379 (.Y(n19957),
	.A(n19955),
	.B(n19954),
	.C(n19953));
   NAND2xp33_ASAP7_75t_SRAM U21380 (.Y(n19955),
	.A(FE_OFN28965_n24869),
	.B(n19951));
   NAND3xp33_ASAP7_75t_SL U21381 (.Y(n19959),
	.A(n24648),
	.B(n19949),
	.C(n20114));
   NAND2xp5_ASAP7_75t_L U21382 (.Y(n19949),
	.A(n19948),
	.B(n19947));
   NAND2xp33_ASAP7_75t_R U21383 (.Y(n19947),
	.A(n19946),
	.B(n19945));
   NAND2xp33_ASAP7_75t_R U21384 (.Y(n19948),
	.A(n19944),
	.B(n19945));
   NAND2x1_ASAP7_75t_SL U21386 (.Y(n19936),
	.A(n18338),
	.B(n22403));
   NAND2xp5_ASAP7_75t_SL U21387 (.Y(n19934),
	.A(n19938),
	.B(n18847));
   NAND2xp33_ASAP7_75t_L U21388 (.Y(n21289),
	.A(n21288),
	.B(n21287));
   NAND2xp33_ASAP7_75t_R U21389 (.Y(n21287),
	.A(n21286),
	.B(n21285));
   NAND2xp33_ASAP7_75t_R U21390 (.Y(n21288),
	.A(n21283),
	.B(n21285));
   NOR2xp33_ASAP7_75t_SRAM U21391 (.Y(n21286),
	.A(FE_OFN28614_n21715),
	.B(n21284));
   NAND2xp5_ASAP7_75t_L U21392 (.Y(n21316),
	.A(n21307),
	.B(n21306));
   NAND2xp5_ASAP7_75t_L U21393 (.Y(n21307),
	.A(n21303),
	.B(n24245));
   NOR3xp33_ASAP7_75t_SL U21394 (.Y(n21523),
	.A(n21294),
	.B(n23412),
	.C(n21293));
   OAI21xp33_ASAP7_75t_L U21395 (.Y(n21293),
	.A1(FE_OFN29109_n),
	.A2(n21292),
	.B(n23419));
   NAND2xp33_ASAP7_75t_R U21396 (.Y(n21315),
	.A(n21314),
	.B(n21313));
   NAND2xp33_ASAP7_75t_SRAM U21397 (.Y(n21313),
	.A(n21312),
	.B(n21311));
   NAND2xp33_ASAP7_75t_SRAM U21398 (.Y(n21314),
	.A(n21309),
	.B(n21311));
   NOR3x1_ASAP7_75t_L U21400 (.Y(n21334),
	.A(n21037),
	.B(n21520),
	.C(n21279));
   NAND3xp33_ASAP7_75t_SL U21401 (.Y(n21037),
	.A(FE_OFN28635_n21034),
	.B(n21064),
	.C(n21033));
   NAND2xp5_ASAP7_75t_L U21402 (.Y(n21033),
	.A(n21032),
	.B(n21031));
   NAND2xp5_ASAP7_75t_SL U21403 (.Y(n21333),
	.A(n21331),
	.B(n21330));
   NAND2xp33_ASAP7_75t_L U21404 (.Y(n21330),
	.A(n21329),
	.B(n21328));
   NAND2xp33_ASAP7_75t_SL U21405 (.Y(n21331),
	.A(n21326),
	.B(n21328));
   NOR2xp33_ASAP7_75t_SRAM U21406 (.Y(n21329),
	.A(n21327),
	.B(FE_OCPN27628_n23455));
   NOR3xp33_ASAP7_75t_R U21407 (.Y(n21332),
	.A(n21284),
	.B(n21513),
	.C(n21074));
   O2A1O1Ixp33_ASAP7_75t_L U21408 (.Y(n21270),
	.A1(n21269),
	.A2(n21738),
	.B(FE_OCPN27617_n18016),
	.C(n21268));
   NAND2xp33_ASAP7_75t_L U21409 (.Y(n21271),
	.A(FE_OCPN27617_n18016),
	.B(FE_OFN28589_n21048));
   NOR2xp33_ASAP7_75t_SL U21410 (.Y(n23426),
	.A(FE_OCPN27675_n17986),
	.B(FE_OCPN27998_n18019));
   NAND2x1_ASAP7_75t_SL U21411 (.Y(n21731),
	.A(n18861),
	.B(n21718));
   OAI21xp5_ASAP7_75t_L U21412 (.Y(n21038),
	.A1(FE_OFN27189_n),
	.A2(n21292),
	.B(n19449));
   OAI21xp33_ASAP7_75t_SRAM U21413 (.Y(n24244),
	.A1(n21706),
	.A2(FE_OCPN28184_n18020),
	.B(n21060));
   NAND2xp5_ASAP7_75t_L U21414 (.Y(n21510),
	.A(FE_PSN8306_FE_OFN28689_sa03_5),
	.B(n18874));
   NOR3xp33_ASAP7_75t_SRAM U21415 (.Y(n18905),
	.A(n21735),
	.B(n21752),
	.C(n18904));
   NOR3xp33_ASAP7_75t_SL U21416 (.Y(n18906),
	.A(n18903),
	.B(n18008),
	.C(n18902));
   OAI22xp33_ASAP7_75t_SRAM U21417 (.Y(n18903),
	.A1(n21706),
	.A2(FE_OCPN27948_FE_OFN26173_n21511),
	.B1(FE_OFN27133_n21725),
	.B2(FE_OCPN27948_FE_OFN26173_n21511));
   NAND3xp33_ASAP7_75t_L U21418 (.Y(n18908),
	.A(n19445),
	.B(n21714),
	.C(n21750));
   NAND2xp33_ASAP7_75t_L U21419 (.Y(n18886),
	.A(n18885),
	.B(n18884));
   NAND2xp33_ASAP7_75t_R U21420 (.Y(n18884),
	.A(n18883),
	.B(n18882));
   NAND2xp33_ASAP7_75t_R U21421 (.Y(n18885),
	.A(n18881),
	.B(n18882));
   NOR3xp33_ASAP7_75t_SL U21422 (.Y(n18043),
	.A(n18042),
	.B(FE_OCPN7618_n21027),
	.C(n21015));
   NOR3xp33_ASAP7_75t_SL U21423 (.Y(n18044),
	.A(n18869),
	.B(n23441),
	.C(n21735));
   NAND3xp33_ASAP7_75t_SL U21425 (.Y(n23942),
	.A(n18862),
	.B(n18001),
	.C(n18889));
   NAND2xp33_ASAP7_75t_L U21426 (.Y(n18000),
	.A(n17994),
	.B(n21047));
   NOR3xp33_ASAP7_75t_SL U21427 (.Y(n22066),
	.A(n22064),
	.B(n22561),
	.C(n22063));
   NAND3xp33_ASAP7_75t_SL U21428 (.Y(n22910),
	.A(n22898),
	.B(n22897),
	.C(n22896));
   OAI222xp33_ASAP7_75t_L U21429 (.Y(n22909),
	.A1(n22908),
	.A2(n27140),
	.B1(n22907),
	.B2(n27140),
	.C1(n22906),
	.C2(n27140));
   NOR3xp33_ASAP7_75t_L U21430 (.Y(n22907),
	.A(n22905),
	.B(n25296),
	.C(n22904));
   NOR3xp33_ASAP7_75t_R U21431 (.Y(n22908),
	.A(n22901),
	.B(n22900),
	.C(n22899));
   NAND2xp33_ASAP7_75t_SRAM U21432 (.Y(n22905),
	.A(n22903),
	.B(n22902));
   NAND2xp33_ASAP7_75t_SL U21433 (.Y(n22886),
	.A(n22880),
	.B(n22883));
   NOR2x1_ASAP7_75t_L U21435 (.Y(n23992),
	.A(n24460),
	.B(n21890));
   NAND2xp33_ASAP7_75t_SRAM U21437 (.Y(n23026),
	.A(FE_OFN28916_sa10_4),
	.B(FE_OFN16377_n23998));
   NAND2xp33_ASAP7_75t_SRAM U21438 (.Y(n23025),
	.A(n23024),
	.B(FE_OFN16377_n23998));
   OAI21x1_ASAP7_75t_SL U21439 (.Y(n23999),
	.A1(FE_OCPN27636_sa10_4),
	.A2(n16646),
	.B(n23120));
   NAND2x1_ASAP7_75t_L U21440 (.Y(n23997),
	.A(n23127),
	.B(n19771));
   NAND3xp33_ASAP7_75t_SL U21441 (.Y(n21185),
	.A(n21176),
	.B(n21175),
	.C(n21174));
   NAND2xp5_ASAP7_75t_L U21442 (.Y(n21174),
	.A(n21173),
	.B(n21172));
   NOR3xp33_ASAP7_75t_SL U21443 (.Y(n21176),
	.A(n21165),
	.B(n21164),
	.C(n21163));
   NAND2xp5_ASAP7_75t_R U21444 (.Y(n21172),
	.A(n21171),
	.B(n21170));
   NAND2xp33_ASAP7_75t_L U21446 (.Y(n21153),
	.A(n19812),
	.B(n19811));
   NAND2xp5_ASAP7_75t_R U21447 (.Y(n21159),
	.A(n18655),
	.B(n19835));
   NOR2xp33_ASAP7_75t_L U21448 (.Y(n18655),
	.A(n24348),
	.B(n18654));
   NAND2xp33_ASAP7_75t_L U21449 (.Y(n18654),
	.A(n18653),
	.B(n18652));
   NAND2xp33_ASAP7_75t_SRAM U21451 (.Y(n21156),
	.A(n17254),
	.B(FE_PSN8282_n21154));
   OAI21xp5_ASAP7_75t_SL U21452 (.Y(n24348),
	.A1(FE_OCPN27951_n19098),
	.A2(FE_OFN29062_n18651),
	.B(n18650));
   NOR2xp33_ASAP7_75t_L U21453 (.Y(n18650),
	.A(n21439),
	.B(n18746));
   NAND3x1_ASAP7_75t_L U21455 (.Y(n21462),
	.A(FE_OCPN28021_n21445),
	.B(FE_OCPN27500_n19834),
	.C(FE_OFN29172_sa00_4));
   NAND2xp33_ASAP7_75t_SRAM U21457 (.Y(n21486),
	.A(n21485),
	.B(n21484));
   NAND2xp33_ASAP7_75t_SRAM U21459 (.Y(n21485),
	.A(n21480),
	.B(n21482));
   NAND3xp33_ASAP7_75t_L U21460 (.Y(n21490),
	.A(FE_OCPN28167_n21472),
	.B(n21471),
	.C(FE_OFN16306_n27041));
   NAND3xp33_ASAP7_75t_L U21461 (.Y(n24476),
	.A(n21476),
	.B(n21458),
	.C(FE_OCPN5199_n21457));
   NOR3x1_ASAP7_75t_SL U21463 (.Y(n19598),
	.A(n18736),
	.B(n21147),
	.C(n17297));
   NAND2xp5_ASAP7_75t_SL U21464 (.Y(n18736),
	.A(n21167),
	.B(n19615));
   NAND2x1_ASAP7_75t_L U21466 (.Y(n19602),
	.A(FE_OCPN28021_n21445),
	.B(n21479));
   NOR2xp33_ASAP7_75t_L U21467 (.Y(n21181),
	.A(n19839),
	.B(FE_OFN28958_n17261));
   NOR2xp33_ASAP7_75t_L U21468 (.Y(n18629),
	.A(n19593),
	.B(FE_OCPN27588_n19824));
   NAND2xp5_ASAP7_75t_L U21469 (.Y(n19840),
	.A(n21167),
	.B(n17272));
   INVxp67_ASAP7_75t_L U21470 (.Y(n17241),
	.A(n17239));
   INVxp67_ASAP7_75t_R U21471 (.Y(n19574),
	.A(n24097));
   NAND3xp33_ASAP7_75t_SL U21472 (.Y(n24099),
	.A(FE_OCPN27679_n18631),
	.B(n17245),
	.C(FE_PSN8275_FE_OCPN27818_n17267));
   NOR2x1_ASAP7_75t_L U21473 (.Y(n24086),
	.A(FE_OCPN29415_n17237),
	.B(FE_OCPN27968_n21154));
   A2O1A1Ixp33_ASAP7_75t_SL U21474 (.Y(n24103),
	.A1(n17309),
	.A2(n17308),
	.B(n21493),
	.C(n17307));
   NOR3xp33_ASAP7_75t_SL U21475 (.Y(n17308),
	.A(n17295),
	.B(n19145),
	.C(n19846));
   NOR3xp33_ASAP7_75t_L U21476 (.Y(n25555),
	.A(n18288),
	.B(n17128),
	.C(n25220));
   NAND2xp33_ASAP7_75t_L U21477 (.Y(n25554),
	.A(n17094),
	.B(n17093));
   NAND2xp33_ASAP7_75t_R U21478 (.Y(n17093),
	.A(n17092),
	.B(n20499));
   NAND2xp33_ASAP7_75t_R U21479 (.Y(n17094),
	.A(n17090),
	.B(n20499));
   NAND3xp33_ASAP7_75t_L U21480 (.Y(n25539),
	.A(n18924),
	.B(n25872),
	.C(n17102));
   NOR3xp33_ASAP7_75t_R U21481 (.Y(n25541),
	.A(n20523),
	.B(n19435),
	.C(n19434));
   NAND2x1p5_ASAP7_75t_L U21483 (.Y(n22902),
	.A(FE_OCPN29469_n17747),
	.B(FE_OCPN27771_n19275));
   NOR3xp33_ASAP7_75t_L U21484 (.Y(n22107),
	.A(n20995),
	.B(n20952),
	.C(FE_OFN28924_n25912));
   NAND3xp33_ASAP7_75t_SL U21485 (.Y(n20954),
	.A(n17761),
	.B(n22888),
	.C(FE_OFN27202_n));
   NAND2x1_ASAP7_75t_L U21486 (.Y(n20955),
	.A(FE_OCPN29469_n17747),
	.B(n17757));
   NAND3xp33_ASAP7_75t_L U21487 (.Y(n20957),
	.A(n19280),
	.B(FE_OCPN28303_n20961),
	.C(n20174));
   NAND2xp5_ASAP7_75t_R U21488 (.Y(n22534),
	.A(FE_OCPN27570_n17791),
	.B(FE_OFN108_n26971));
   NOR3xp33_ASAP7_75t_L U21490 (.Y(n20990),
	.A(n20989),
	.B(FE_OCPN27972_n20988),
	.C(n20987));
   NOR3xp33_ASAP7_75t_L U21491 (.Y(n20991),
	.A(n25298),
	.B(n22894),
	.C(n22532));
   NAND3xp33_ASAP7_75t_L U21492 (.Y(n20989),
	.A(n20986),
	.B(n22891),
	.C(n22067));
   NAND3x1_ASAP7_75t_SL U21493 (.Y(n21000),
	.A(n20999),
	.B(n20998),
	.C(n20997));
   NAND3xp33_ASAP7_75t_SL U21494 (.Y(n22547),
	.A(n17788),
	.B(n19255),
	.C(n20214));
   NOR2xp33_ASAP7_75t_SL U21495 (.Y(n17788),
	.A(n20952),
	.B(n20186));
   NAND3xp33_ASAP7_75t_R U21496 (.Y(n22109),
	.A(n20983),
	.B(n22065),
	.C(n22084));
   NOR3xp33_ASAP7_75t_L U21497 (.Y(n20983),
	.A(n25531),
	.B(n20982),
	.C(n20981));
   NOR2x1_ASAP7_75t_L U21498 (.Y(n20190),
	.A(n25297),
	.B(n25296));
   NAND2xp5_ASAP7_75t_SL U21499 (.Y(n25301),
	.A(n19245),
	.B(n19244));
   NAND2xp33_ASAP7_75t_SL U21500 (.Y(n19244),
	.A(n19243),
	.B(n19242));
   NAND2xp33_ASAP7_75t_SL U21501 (.Y(n19245),
	.A(n19241),
	.B(n19242));
   OAI22xp33_ASAP7_75t_L U21502 (.Y(n17774),
	.A1(FE_OFN25998_n17781),
	.A2(n20132),
	.B1(FE_OFN108_n26971),
	.B2(n20132));
   NAND3xp33_ASAP7_75t_R U21503 (.Y(n25309),
	.A(n22085),
	.B(n20992),
	.C(n22878));
   NAND3xp33_ASAP7_75t_SRAM U21504 (.Y(n25310),
	.A(n20955),
	.B(n20954),
	.C(n20202));
   NOR2xp33_ASAP7_75t_L U21505 (.Y(n22058),
	.A(n20194),
	.B(n22872));
   OAI22xp33_ASAP7_75t_SRAM U21506 (.Y(n22059),
	.A1(FE_OCPN27771_n19275),
	.A2(n22533),
	.B1(FE_OCPN29469_n17747),
	.B2(n22533));
   NAND2xp33_ASAP7_75t_SRAM U21508 (.Y(n26969),
	.A(n22074),
	.B(n22073));
   NAND2xp33_ASAP7_75t_L U21509 (.Y(n26967),
	.A(n22076),
	.B(n22075));
   NAND2xp33_ASAP7_75t_L U21510 (.Y(n22082),
	.A(n22079),
	.B(n22078));
   NOR3xp33_ASAP7_75t_R U21512 (.Y(n18282),
	.A(FE_OCPN29541_n25870),
	.B(n18276),
	.C(n18275));
   NOR3xp33_ASAP7_75t_R U21513 (.Y(n18280),
	.A(n18279),
	.B(n20490),
	.C(n20529));
   NOR3xp33_ASAP7_75t_SL U21514 (.Y(n18281),
	.A(n25220),
	.B(FE_OFN28559_n18278),
	.C(n18277));
   NOR3xp33_ASAP7_75t_SRAM U21516 (.Y(n18290),
	.A(n18289),
	.B(n25996),
	.C(n18288));
   NAND2xp33_ASAP7_75t_SRAM U21517 (.Y(n18258),
	.A(n18257),
	.B(n25872));
   OAI21xp33_ASAP7_75t_L U21518 (.Y(n18273),
	.A1(FE_OFN28491_sa13_3),
	.A2(n17033),
	.B(n18241));
   NAND2xp33_ASAP7_75t_SRAM U21519 (.Y(n18252),
	.A(n18248),
	.B(n18249));
   NAND3x1_ASAP7_75t_SL U21520 (.Y(n25287),
	.A(n17138),
	.B(FE_OCPN29569_n18947),
	.C(n19431));
   NAND2xp5_ASAP7_75t_SL U21521 (.Y(n17138),
	.A(n17137),
	.B(n17136));
   NAND2xp33_ASAP7_75t_SL U21522 (.Y(n17136),
	.A(n17135),
	.B(n17134));
   NAND2xp33_ASAP7_75t_SL U21523 (.Y(n17137),
	.A(n17133),
	.B(n17134));
   NAND3xp33_ASAP7_75t_SL U21524 (.Y(n20492),
	.A(FE_OCPN27902_n20514),
	.B(FE_OCPN28137_n17170),
	.C(FE_OCPN29351_FE_OFN26116_sa13_1));
   NAND3xp33_ASAP7_75t_SL U21525 (.Y(n20495),
	.A(n25995),
	.B(FE_OFN26572_n19405),
	.C(n17130));
   NOR3xp33_ASAP7_75t_SL U21526 (.Y(n17130),
	.A(n18277),
	.B(n17129),
	.C(n17128));
   NOR3xp33_ASAP7_75t_SRAM U21527 (.Y(n20504),
	.A(n20503),
	.B(n20502),
	.C(n20501));
   NOR2xp33_ASAP7_75t_R U21528 (.Y(n20520),
	.A(n20507),
	.B(n20506));
   NAND2xp5_ASAP7_75t_SL U21529 (.Y(n20519),
	.A(n20518),
	.B(n20517));
   NAND2xp33_ASAP7_75t_SRAM U21530 (.Y(n20517),
	.A(n20516),
	.B(n20515));
   NAND2xp33_ASAP7_75t_SL U21531 (.Y(n20518),
	.A(n20512),
	.B(n20515));
   NOR3xp33_ASAP7_75t_SL U21532 (.Y(n20531),
	.A(n18265),
	.B(FE_OCPN29525_n18947),
	.C(n18264));
   NAND3xp33_ASAP7_75t_SL U21534 (.Y(n18265),
	.A(n18262),
	.B(n18261),
	.C(n18260));
   NOR3xp33_ASAP7_75t_L U21535 (.Y(n20533),
	.A(n20530),
	.B(n20529),
	.C(n20528));
   NOR2xp33_ASAP7_75t_L U21537 (.Y(n21026),
	.A(n18879),
	.B(n21297));
   NOR3xp33_ASAP7_75t_SL U21538 (.Y(n19484),
	.A(n19482),
	.B(n19481),
	.C(n18902));
   NOR2xp33_ASAP7_75t_SL U21539 (.Y(n19483),
	.A(n21707),
	.B(n19475));
   NOR3xp33_ASAP7_75t_SL U21540 (.Y(n19494),
	.A(n19491),
	.B(n19490),
	.C(n23420));
   NAND2x1_ASAP7_75t_L U21541 (.Y(n21292),
	.A(n18045),
	.B(FE_OCPN27285_n18011));
   NOR3xp33_ASAP7_75t_SRAM U21542 (.Y(n19493),
	.A(n21278),
	.B(n19492),
	.C(n21023));
   NOR3xp33_ASAP7_75t_L U21544 (.Y(n24241),
	.A(n21505),
	.B(n18008),
	.C(n21504));
   NOR2x1_ASAP7_75t_SL U21545 (.Y(n24243),
	.A(FE_OFN29122_n),
	.B(n19450));
   NAND3xp33_ASAP7_75t_SL U21546 (.Y(n24249),
	.A(n21282),
	.B(n21281),
	.C(n21280));
   OAI22xp33_ASAP7_75t_R U21547 (.Y(n21506),
	.A1(FE_OFN28589_n21048),
	.A2(n19478),
	.B1(n21295),
	.B2(n19478));
   NOR3xp33_ASAP7_75t_SL U21548 (.Y(n19688),
	.A(n23038),
	.B(n19791),
	.C(n19686));
   NAND3x1_ASAP7_75t_SL U21549 (.Y(n23144),
	.A(n23048),
	.B(n23028),
	.C(n19660));
   NAND3xp33_ASAP7_75t_SL U21550 (.Y(n19691),
	.A(n19676),
	.B(n19667),
	.C(n24000));
   NOR3xp33_ASAP7_75t_SRAM U21551 (.Y(n19676),
	.A(FE_OFN28923_n21873),
	.B(n21894),
	.C(n21906));
   NOR3x1_ASAP7_75t_L U21552 (.Y(n23955),
	.A(n17202),
	.B(n21893),
	.C(n19679));
   NAND2xp5_ASAP7_75t_L U21553 (.Y(n17202),
	.A(n17200),
	.B(n24896));
   NAND3x1_ASAP7_75t_SL U21554 (.Y(n23958),
	.A(n19637),
	.B(n19636),
	.C(n19635));
   NAND2xp5_ASAP7_75t_L U21555 (.Y(n19636),
	.A(n19634),
	.B(n19633));
   NAND2xp33_ASAP7_75t_R U21556 (.Y(n19634),
	.A(n19629),
	.B(FE_OCPN27906_n23131));
   OAI21xp33_ASAP7_75t_SRAM U21557 (.Y(n24459),
	.A1(n23982),
	.A2(n17191),
	.B(n17187));
   NOR3xp33_ASAP7_75t_SL U21558 (.Y(n24461),
	.A(n19625),
	.B(n19663),
	.C(n17190));
   NAND2x1_ASAP7_75t_SL U21559 (.Y(n24458),
	.A(n16663),
	.B(n19769));
   NAND2xp5_ASAP7_75t_SL U21560 (.Y(n24901),
	.A(n17228),
	.B(n16555));
   NOR3xp33_ASAP7_75t_L U21561 (.Y(n16555),
	.A(n16554),
	.B(n17221),
	.C(n16553));
   NAND2xp33_ASAP7_75t_L U21562 (.Y(n16553),
	.A(n16580),
	.B(n16618));
   NOR2xp33_ASAP7_75t_L U21563 (.Y(n17228),
	.A(n19671),
	.B(n16620));
   NAND2xp33_ASAP7_75t_L U21564 (.Y(n17218),
	.A(n19781),
	.B(n19668));
   NAND2xp5_ASAP7_75t_L U21565 (.Y(n21904),
	.A(n17217),
	.B(n19770));
   OAI21xp33_ASAP7_75t_L U21566 (.Y(n17214),
	.A1(n17213),
	.A2(n17212),
	.B(n17211));
   NOR2xp33_ASAP7_75t_SRAM U21567 (.Y(n17211),
	.A(FE_OFN59_sa10_7),
	.B(FE_OFN131_sa10_6));
   NAND2xp33_ASAP7_75t_L U21568 (.Y(n17213),
	.A(n24967),
	.B(n23955));
   NAND3xp33_ASAP7_75t_R U21569 (.Y(n17212),
	.A(n17210),
	.B(n17209),
	.C(n21896));
   NAND2xp33_ASAP7_75t_R U21570 (.Y(n17198),
	.A(n19781),
	.B(n17197));
   NOR3xp33_ASAP7_75t_L U21571 (.Y(n17229),
	.A(n17227),
	.B(FE_OFN29154_n19753),
	.C(n23998));
   NAND2xp33_ASAP7_75t_SRAM U21572 (.Y(n17227),
	.A(n19635),
	.B(n17222));
   NOR3x1_ASAP7_75t_SL U21573 (.Y(n21882),
	.A(n21875),
	.B(n23133),
	.C(n19765));
   NOR2xp33_ASAP7_75t_SRAM U21575 (.Y(n21913),
	.A(FE_OCPN28358_n21899),
	.B(n23044));
   NAND2xp33_ASAP7_75t_SL U21576 (.Y(n21911),
	.A(n21910),
	.B(n21909));
   NOR3xp33_ASAP7_75t_SL U21577 (.Y(n21912),
	.A(n23958),
	.B(n21901),
	.C(n21900));
   NAND3x1_ASAP7_75t_SL U21578 (.Y(n23998),
	.A(n17226),
	.B(n17225),
	.C(n24461));
   NOR3xp33_ASAP7_75t_SL U21579 (.Y(n17225),
	.A(n17224),
	.B(n23132),
	.C(n21906));
   NAND2xp33_ASAP7_75t_L U21580 (.Y(n17224),
	.A(n19767),
	.B(n19768));
   NAND3xp33_ASAP7_75t_R U21581 (.Y(n21915),
	.A(n21898),
	.B(n21897),
	.C(n21896));
   NAND2xp33_ASAP7_75t_SRAM U21582 (.Y(n21887),
	.A(n21886),
	.B(n21885));
   NOR2xp33_ASAP7_75t_SL U21583 (.Y(n21872),
	.A(n16533),
	.B(n21902));
   NAND2xp33_ASAP7_75t_SL U21585 (.Y(n21874),
	.A(n24949),
	.B(n24951));
   NAND2xp33_ASAP7_75t_SRAM U21586 (.Y(n24727),
	.A(n23129),
	.B(n23128));
   NAND3xp33_ASAP7_75t_SRAM U21587 (.Y(n23126),
	.A(n23980),
	.B(FE_OCPN28323_FE_OFN16427_sa10_3),
	.C(n19756));
   NOR3xp33_ASAP7_75t_SL U21588 (.Y(n23125),
	.A(n16634),
	.B(n23133),
	.C(n16633));
   NOR2xp33_ASAP7_75t_SRAM U21591 (.Y(n23155),
	.A(n24958),
	.B(n23141));
   NAND2xp33_ASAP7_75t_L U21592 (.Y(n23153),
	.A(n23152),
	.B(n23151));
   NOR3xp33_ASAP7_75t_SL U21593 (.Y(n23154),
	.A(n23145),
	.B(n23144),
	.C(n23143));
   NAND3xp33_ASAP7_75t_R U21594 (.Y(n24731),
	.A(FE_OFN16291_n23142),
	.B(n23140),
	.C(n23955));
   NAND3xp33_ASAP7_75t_L U21595 (.Y(n24732),
	.A(n23136),
	.B(FE_OFN28946_n23135),
	.C(n23134));
   NAND2xp5_ASAP7_75t_SL U21596 (.Y(n24742),
	.A(n16589),
	.B(n16642));
   NAND3xp33_ASAP7_75t_SRAM U21597 (.Y(n24735),
	.A(n23121),
	.B(n23120),
	.C(n24669));
   NOR3x1_ASAP7_75t_R U21598 (.Y(n24734),
	.A(n16648),
	.B(FE_OFN26160_sa10_4),
	.C(FE_OCPN29498_n16581));
   NAND3xp33_ASAP7_75t_SL U21599 (.Y(n24733),
	.A(n19776),
	.B(n19775),
	.C(n23134));
   NOR3xp33_ASAP7_75t_L U21600 (.Y(n19776),
	.A(n19773),
	.B(n19772),
	.C(n24976));
   NOR2x1_ASAP7_75t_L U21601 (.Y(n23119),
	.A(FE_OCPN29424_FE_OFN26039_sa10_2),
	.B(n16616));
   NAND2xp5_ASAP7_75t_SL U21602 (.Y(n17219),
	.A(FE_OFN130_sa10_5),
	.B(n19661));
   NOR2xp33_ASAP7_75t_SL U21603 (.Y(n19653),
	.A(n21872),
	.B(n21899));
   NAND2xp33_ASAP7_75t_L U21604 (.Y(n21885),
	.A(n16542),
	.B(n19641));
   NOR2x1p5_ASAP7_75t_SL U21605 (.Y(n19791),
	.A(n16648),
	.B(FE_OFN28910_n16534));
   NOR3x1_ASAP7_75t_SL U21607 (.Y(n24969),
	.A(n16599),
	.B(FE_OFN28923_n21873),
	.C(n24894));
   NAND3x1_ASAP7_75t_SL U21608 (.Y(n16599),
	.A(n16593),
	.B(n19687),
	.C(n23993));
   OAI21xp33_ASAP7_75t_SRAM U21609 (.Y(n16593),
	.A1(FE_OCPN27900_n23949),
	.A2(n23948),
	.B(FE_OFN26161_sa10_4));
   NAND2xp5_ASAP7_75t_SL U21611 (.Y(n16618),
	.A(FE_OCPN28157_n16534),
	.B(n24944));
   NOR3xp33_ASAP7_75t_R U21612 (.Y(n19128),
	.A(n19118),
	.B(n26100),
	.C(n19117));
   NAND2xp5_ASAP7_75t_R U21613 (.Y(n19127),
	.A(n19126),
	.B(n19125));
   NAND2xp33_ASAP7_75t_L U21614 (.Y(n19125),
	.A(n19124),
	.B(n19123));
   NAND2xp33_ASAP7_75t_L U21615 (.Y(n19126),
	.A(n19120),
	.B(n19123));
   NOR3xp33_ASAP7_75t_SRAM U21617 (.Y(n19152),
	.A(n19151),
	.B(n19150),
	.C(n17297));
   NOR2xp33_ASAP7_75t_SRAM U21618 (.Y(n19151),
	.A(FE_OFN26651_n19573),
	.B(FE_OCPN29464_n));
   NAND3xp33_ASAP7_75t_SL U21619 (.Y(n19156),
	.A(n19141),
	.B(n19140),
	.C(n19584));
   NOR3xp33_ASAP7_75t_SRAM U21620 (.Y(n19140),
	.A(n19138),
	.B(n26100),
	.C(n26099));
   NAND2xp33_ASAP7_75t_SRAM U21622 (.Y(n19137),
	.A(FE_OCPN29346_n12998),
	.B(n19609));
   NAND3xp33_ASAP7_75t_L U21624 (.Y(n19596),
	.A(n21473),
	.B(n18742),
	.C(n17302));
   NAND3xp33_ASAP7_75t_L U21625 (.Y(n19105),
	.A(n19104),
	.B(n19103),
	.C(n21177));
   O2A1O1Ixp33_ASAP7_75t_L U21626 (.Y(n19103),
	.A1(FE_OCPN27818_n17267),
	.A2(FE_OFN28514_sa00_1),
	.B(n19122),
	.C(n21491));
   NAND3xp33_ASAP7_75t_SL U21627 (.Y(n24344),
	.A(n19093),
	.B(n19092),
	.C(n19860));
   NOR2xp33_ASAP7_75t_SRAM U21628 (.Y(n19093),
	.A(FE_OFN25980_n19087),
	.B(n19150));
   NAND2xp33_ASAP7_75t_SRAM U21629 (.Y(n19109),
	.A(n19108),
	.B(n19107));
   NOR2x1_ASAP7_75t_L U21630 (.Y(n17653),
	.A(n22623),
	.B(n17647));
   INVx1_ASAP7_75t_L U21631 (.Y(n17647),
	.A(n18496));
   NAND2xp5_ASAP7_75t_L U21633 (.Y(n18396),
	.A(n18395),
	.B(n18394));
   NOR3xp33_ASAP7_75t_L U21634 (.Y(n18395),
	.A(n18387),
	.B(n21608),
	.C(n18508));
   NOR3xp33_ASAP7_75t_SL U21635 (.Y(n18394),
	.A(n24128),
	.B(n19075),
	.C(n18393));
   NOR2xp33_ASAP7_75t_SL U21636 (.Y(n24795),
	.A(n20450),
	.B(n18476));
   NAND3xp33_ASAP7_75t_SL U21637 (.Y(n18476),
	.A(n20467),
	.B(n18475),
	.C(n24759));
   NAND2xp5_ASAP7_75t_L U21638 (.Y(n26024),
	.A(n22167),
	.B(n22166));
   NAND2xp5_ASAP7_75t_L U21640 (.Y(n22129),
	.A(n22123),
	.B(n22126));
   NAND2xp33_ASAP7_75t_L U21641 (.Y(n22128),
	.A(n22127),
	.B(n22126));
   NOR2xp33_ASAP7_75t_L U21642 (.Y(n22127),
	.A(FE_OFN28610_n22125),
	.B(n22124));
   OAI21xp33_ASAP7_75t_SL U21643 (.Y(n22635),
	.A1(FE_OFN25901_n22133),
	.A2(FE_OCPN27428_n26027),
	.B(n22132));
   NOR3x1_ASAP7_75t_L U21644 (.Y(n22617),
	.A(n18494),
	.B(n21601),
	.C(n18493));
   NAND2xp5_ASAP7_75t_L U21645 (.Y(n18493),
	.A(n18492),
	.B(n18491));
   NOR3xp33_ASAP7_75t_R U21646 (.Y(n20477),
	.A(n22640),
	.B(n20450),
	.C(n22613));
   NAND2xp33_ASAP7_75t_L U21647 (.Y(n20485),
	.A(n22654),
	.B(n20483));
   NOR2xp33_ASAP7_75t_L U21648 (.Y(n20478),
	.A(n17645),
	.B(n20439));
   NOR3x1_ASAP7_75t_L U21650 (.Y(n18384),
	.A(n18383),
	.B(n22139),
	.C(n18382));
   NOR3xp33_ASAP7_75t_SRAM U21651 (.Y(n18382),
	.A(n20429),
	.B(FE_OCPN29413_sa30_5),
	.C(n18381));
   NAND2xp5_ASAP7_75t_L U21652 (.Y(n18456),
	.A(n20427),
	.B(n18478));
   NAND3xp33_ASAP7_75t_SL U21653 (.Y(n20433),
	.A(n17613),
	.B(n19063),
	.C(n22625));
   NAND3xp33_ASAP7_75t_L U21654 (.Y(n22619),
	.A(n20432),
	.B(n22132),
	.C(n20431));
   OAI21xp33_ASAP7_75t_SRAM U21655 (.Y(n20430),
	.A1(n20429),
	.A2(FE_PSN8272_n20428),
	.B(n20427));
   NAND2xp33_ASAP7_75t_SRAM U21656 (.Y(n20426),
	.A(n20420),
	.B(n20423));
   NOR3xp33_ASAP7_75t_SRAM U21657 (.Y(n17481),
	.A(n19198),
	.B(FE_OCPN27496_n21820),
	.C(n17462));
   NOR3xp33_ASAP7_75t_SRAM U21658 (.Y(n17479),
	.A(n23281),
	.B(n21823),
	.C(n19194));
   NAND2x1_ASAP7_75t_SL U21659 (.Y(n22508),
	.A(n17488),
	.B(n17487));
   NAND2xp5_ASAP7_75t_SL U21660 (.Y(n17488),
	.A(n17484),
	.B(FE_OFN26031_n22499));
   NAND2xp5_ASAP7_75t_SL U21661 (.Y(n17487),
	.A(n17486),
	.B(FE_OFN26031_n22499));
   NOR2xp33_ASAP7_75t_L U21662 (.Y(n17505),
	.A(n17493),
	.B(n17492));
   NOR3xp33_ASAP7_75t_L U21663 (.Y(n17515),
	.A(n17513),
	.B(n24079),
	.C(n21385));
   OAI21xp33_ASAP7_75t_SRAM U21664 (.Y(n17514),
	.A1(FE_OFN29061_n22505),
	.A2(n19162),
	.B(FE_OCPN5021_n17446));
   NAND3xp33_ASAP7_75t_R U21665 (.Y(n17493),
	.A(FE_OCPN28417_n21396),
	.B(n24548),
	.C(n23260));
   NAND2xp33_ASAP7_75t_SRAM U21666 (.Y(n17455),
	.A(n17502),
	.B(n21362));
   NAND2xp33_ASAP7_75t_SRAM U21668 (.Y(n17449),
	.A(n23269),
	.B(n23391));
   NOR3xp33_ASAP7_75t_SL U21669 (.Y(n19825),
	.A(n17273),
	.B(n19088),
	.C(n24086));
   NAND2xp33_ASAP7_75t_R U21672 (.Y(n19827),
	.A(n19823),
	.B(n19822));
   NAND2xp33_ASAP7_75t_SRAM U21673 (.Y(n19823),
	.A(n19820),
	.B(n19819));
   NAND3xp33_ASAP7_75t_L U21674 (.Y(n19856),
	.A(n21450),
	.B(n19843),
	.C(n19842));
   NOR3xp33_ASAP7_75t_SRAM U21675 (.Y(n19843),
	.A(n19840),
	.B(n26100),
	.C(n21150));
   NAND2xp5_ASAP7_75t_SL U21678 (.Y(n25256),
	.A(n21445),
	.B(n17263));
   NOR2xp33_ASAP7_75t_SL U21679 (.Y(n17263),
	.A(FE_OCPN27338_n19149),
	.B(n17262));
   NAND3xp33_ASAP7_75t_SL U21680 (.Y(n26103),
	.A(FE_OCPN29542_n21151),
	.B(n21154),
	.C(FE_OCPN29396_n19149));
   NAND3xp33_ASAP7_75t_SL U21681 (.Y(n26106),
	.A(n18636),
	.B(n18635),
	.C(n21162));
   NOR3xp33_ASAP7_75t_SRAM U21682 (.Y(n18636),
	.A(n19106),
	.B(n21147),
	.C(n19845));
   NOR3xp33_ASAP7_75t_R U21684 (.Y(n21862),
	.A(n21861),
	.B(FE_OCPN28082_n21860),
	.C(n24561));
   NAND2xp33_ASAP7_75t_SRAM U21685 (.Y(n21861),
	.A(n21859),
	.B(n21858));
   NAND3xp33_ASAP7_75t_SRAM U21686 (.Y(n21865),
	.A(n22484),
	.B(n21846),
	.C(FE_OCPN29416_n22516));
   NAND3xp33_ASAP7_75t_R U21687 (.Y(n17508),
	.A(FE_OCPN27730_n17464),
	.B(FE_OCPN28038_n23252),
	.C(FE_OFN28915_FE_OCPN27241_sa11_1));
   NAND2xp5_ASAP7_75t_SL U21688 (.Y(n17456),
	.A(n23250),
	.B(n23259));
   NAND2xp33_ASAP7_75t_L U21689 (.Y(n24710),
	.A(n21343),
	.B(n21342));
   NAND2xp33_ASAP7_75t_L U21690 (.Y(n21346),
	.A(n23370),
	.B(n21345));
   NOR3xp33_ASAP7_75t_SL U21692 (.Y(n21387),
	.A(n21386),
	.B(n21385),
	.C(n21842));
   OAI21xp5_ASAP7_75t_SL U21693 (.Y(n26084),
	.A1(FE_OCPN28006_n17454),
	.A2(FE_OCPN27313_n21845),
	.B(n21364));
   NOR2x1_ASAP7_75t_SL U21694 (.Y(n21364),
	.A(n23383),
	.B(n21363));
   NAND2xp33_ASAP7_75t_L U21695 (.Y(n24547),
	.A(n22483),
	.B(n22482));
   NAND2xp33_ASAP7_75t_R U21696 (.Y(n22483),
	.A(n22481),
	.B(n22480));
   INVxp67_ASAP7_75t_R U21697 (.Y(n22484),
	.A(n24546));
   NAND3xp33_ASAP7_75t_SRAM U21698 (.Y(n24548),
	.A(FE_OCPN28321_n21341),
	.B(n19171),
	.C(FE_OFN94_sa11_5));
   NAND2xp5_ASAP7_75t_SL U21699 (.Y(n23254),
	.A(n17444),
	.B(FE_OCPN27414_n23359));
   NOR3x1_ASAP7_75t_SL U21701 (.Y(n22515),
	.A(n22513),
	.B(FE_OFN114_n22512),
	.C(n22511));
   NAND3x1_ASAP7_75t_SL U21702 (.Y(n22513),
	.A(n22510),
	.B(n22509),
	.C(n22508));
   NAND3xp33_ASAP7_75t_L U21703 (.Y(n22518),
	.A(FE_OCPN29554_n22507),
	.B(n22506),
	.C(n23371));
   OAI22xp33_ASAP7_75t_SRAM U21704 (.Y(n22506),
	.A1(FE_OFN29061_n22505),
	.A2(n22504),
	.B1(FE_OCPN5021_n17446),
	.B2(n22504));
   NAND3xp33_ASAP7_75t_L U21705 (.Y(n22519),
	.A(n21857),
	.B(n22503),
	.C(n24559));
   NAND3xp33_ASAP7_75t_SL U21706 (.Y(n22499),
	.A(n17483),
	.B(n17482),
	.C(n21425));
   NAND2xp33_ASAP7_75t_SRAM U21707 (.Y(n22494),
	.A(n22493),
	.B(n22492));
   NAND2xp33_ASAP7_75t_R U21708 (.Y(n22493),
	.A(n22491),
	.B(FE_OFN16391_n22490));
   NAND3xp33_ASAP7_75t_SL U21709 (.Y(n21431),
	.A(n23282),
	.B(n21424),
	.C(n23275));
   NOR3xp33_ASAP7_75t_SL U21711 (.Y(n21429),
	.A(n21427),
	.B(n21426),
	.C(n24079));
   NAND2xp33_ASAP7_75t_R U21712 (.Y(n21409),
	.A(n21405),
	.B(n21404));
   NAND2xp33_ASAP7_75t_R U21713 (.Y(n21408),
	.A(n21407),
	.B(n21404));
   NAND2xp5_ASAP7_75t_L U21714 (.Y(n21403),
	.A(n17467),
	.B(n17466));
   NAND2xp33_ASAP7_75t_SRAM U21715 (.Y(n17466),
	.A(n17465),
	.B(FE_OCPN27730_n17464));
   NAND2xp33_ASAP7_75t_SRAM U21716 (.Y(n17467),
	.A(FE_OCPN27903_n19223),
	.B(FE_OCPN27730_n17464));
   NAND2xp33_ASAP7_75t_L U21717 (.Y(n23274),
	.A(n26064),
	.B(n23249));
   NOR3x1_ASAP7_75t_SL U21718 (.Y(n23404),
	.A(n23384),
	.B(n23383),
	.C(n23382));
   NAND2xp33_ASAP7_75t_SRAM U21719 (.Y(n23382),
	.A(n23381),
	.B(n23380));
   NAND3xp33_ASAP7_75t_SL U21720 (.Y(n23384),
	.A(n23379),
	.B(n23378),
	.C(n23377));
   OAI21xp5_ASAP7_75t_SL U21721 (.Y(n23403),
	.A1(n23402),
	.A2(n23401),
	.B(n23400));
   NAND3xp33_ASAP7_75t_SL U21722 (.Y(n23401),
	.A(n23399),
	.B(n23398),
	.C(FE_OCPN29422_n23397));
   NOR3xp33_ASAP7_75t_SL U21723 (.Y(n23398),
	.A(n23396),
	.B(n23395),
	.C(n23394));
   NOR2xp67_ASAP7_75t_SL U21724 (.Y(n23399),
	.A(n24544),
	.B(n23388));
   NOR2xp67_ASAP7_75t_SL U21725 (.Y(n23405),
	.A(n24551),
	.B(n23373));
   NOR3xp33_ASAP7_75t_SL U21726 (.Y(n23369),
	.A(n21853),
	.B(n22498),
	.C(n21852));
   OAI21xp33_ASAP7_75t_SRAM U21727 (.Y(n21852),
	.A1(FE_OCPN28447_n23392),
	.A2(FE_OCPN29378_n23266),
	.B(n21851));
   NOR2xp67_ASAP7_75t_L U21728 (.Y(n23387),
	.A(FE_OCPN27496_n21820),
	.B(n19163));
   NAND2x1p5_ASAP7_75t_SL U21729 (.Y(n26064),
	.A(FE_OFN29054_n17453),
	.B(FE_OCPN29513_n17447));
   NOR2xp33_ASAP7_75t_SL U21730 (.Y(n23365),
	.A(n23273),
	.B(n21406));
   NAND2xp33_ASAP7_75t_SL U21731 (.Y(n23363),
	.A(n23358),
	.B(n23360));
   NAND2xp33_ASAP7_75t_R U21732 (.Y(n23362),
	.A(n23361),
	.B(n23360));
   NAND2xp5_ASAP7_75t_SL U21733 (.Y(n23366),
	.A(n17508),
	.B(n23391));
   OAI21xp33_ASAP7_75t_SRAM U21734 (.Y(n24802),
	.A1(FE_OCPN8207_n18497),
	.A2(n18467),
	.B(FE_OCPN28049_sa30_0));
   NOR3xp33_ASAP7_75t_L U21735 (.Y(n24779),
	.A(n18352),
	.B(FE_OCPN29431_sa30_3),
	.C(FE_OCPN27971_n21627));
   NAND2xp5_ASAP7_75t_SL U21736 (.Y(n19058),
	.A(n18492),
	.B(n18466));
   OAI22xp5_ASAP7_75t_L U21737 (.Y(n18466),
	.A1(FE_OFN28610_n22125),
	.A2(n17616),
	.B1(n18465),
	.B2(n17616));
   NAND3x1_ASAP7_75t_SL U21739 (.Y(n24798),
	.A(n18486),
	.B(FE_OCPN28241_n22142),
	.C(n18485));
   OAI22xp33_ASAP7_75t_R U21740 (.Y(n18486),
	.A1(FE_OCPN29467_n25102),
	.A2(n18484),
	.B1(n18483),
	.B2(n18484));
   NAND2xp33_ASAP7_75t_L U21741 (.Y(n18484),
	.A(n21596),
	.B(n22621));
   NAND3xp33_ASAP7_75t_SL U21742 (.Y(n24797),
	.A(n22617),
	.B(n18496),
	.C(n25115));
   NOR3xp33_ASAP7_75t_SRAM U21743 (.Y(n18511),
	.A(n24761),
	.B(n18510),
	.C(n24762));
   INVxp33_ASAP7_75t_SRAM U21745 (.Y(n26022),
	.A(n24795));
   NAND2xp5_ASAP7_75t_L U21746 (.Y(n21601),
	.A(n18490),
	.B(n18489));
   NAND2xp33_ASAP7_75t_R U21747 (.Y(n21602),
	.A(n22151),
	.B(n22643));
   NOR2xp33_ASAP7_75t_L U21749 (.Y(n21611),
	.A(FE_OFN29094_n21607),
	.B(n21606));
   NAND2xp5_ASAP7_75t_L U21750 (.Y(n21584),
	.A(FE_OFN28896_sa30_2),
	.B(n25083));
   NAND2x1_ASAP7_75t_L U21751 (.Y(n25086),
	.A(n20443),
	.B(n18463));
   NAND2xp33_ASAP7_75t_L U21752 (.Y(n20443),
	.A(n20442),
	.B(n20441));
   NAND3x1_ASAP7_75t_SL U21754 (.Y(n25087),
	.A(n20468),
	.B(n20467),
	.C(n20466));
   NAND2xp33_ASAP7_75t_L U21755 (.Y(n20464),
	.A(n20463),
	.B(n20462));
   NAND3xp33_ASAP7_75t_SL U21756 (.Y(n25118),
	.A(n17640),
	.B(n22130),
	.C(n17639));
   NOR2xp33_ASAP7_75t_L U21757 (.Y(n17639),
	.A(n18458),
	.B(n17638));
   NOR2x1p5_ASAP7_75t_L U21758 (.Y(n25113),
	.A(n18359),
	.B(n20481));
   NAND3x1_ASAP7_75t_SL U21759 (.Y(n25107),
	.A(n19072),
	.B(n18501),
	.C(n17663));
   NAND2xp5_ASAP7_75t_SL U21760 (.Y(n17663),
	.A(n17662),
	.B(n17661));
   NAND2xp5_ASAP7_75t_SL U21761 (.Y(n17661),
	.A(n17660),
	.B(n17659));
   NAND3x1_ASAP7_75t_SL U21762 (.Y(n25104),
	.A(n17606),
	.B(FE_OCPN28057_n17603),
	.C(FE_OFN28896_sa30_2));
   NAND3xp33_ASAP7_75t_L U21763 (.Y(n25103),
	.A(FE_OCPN28378_n22632),
	.B(n22125),
	.C(n18463));
   NOR3xp33_ASAP7_75t_SL U21765 (.Y(n18607),
	.A(n18601),
	.B(n21676),
	.C(FE_OFN28650_n23802));
   NAND3xp33_ASAP7_75t_R U21766 (.Y(n18601),
	.A(n25903),
	.B(FE_OCPN5110_n23721),
	.C(n18598));
   NOR2xp33_ASAP7_75t_R U21767 (.Y(n18598),
	.A(n21648),
	.B(FE_OCPN28017_n18548));
   NAND3x1_ASAP7_75t_SL U21768 (.Y(n23798),
	.A(n18569),
	.B(n20633),
	.C(n18568));
   OAI21xp5_ASAP7_75t_L U21769 (.Y(n18568),
	.A1(n18529),
	.A2(n18567),
	.B(FE_OFN28869_FE_OCPN27715_n23875));
   NOR3x1_ASAP7_75t_SL U21770 (.Y(n18569),
	.A(n18566),
	.B(n18565),
	.C(n21654));
   NAND2xp5_ASAP7_75t_SL U21771 (.Y(n18565),
	.A(n23809),
	.B(n23811));
   NAND3xp33_ASAP7_75t_SL U21772 (.Y(n18609),
	.A(n25637),
	.B(n18581),
	.C(n21200));
   NAND2xp5_ASAP7_75t_SL U21773 (.Y(n18581),
	.A(n18578),
	.B(n18577));
   NAND2xp33_ASAP7_75t_L U21774 (.Y(n18577),
	.A(n18576),
	.B(n18575));
   NAND2xp33_ASAP7_75t_R U21775 (.Y(n18578),
	.A(n18574),
	.B(n18575));
   NAND3xp33_ASAP7_75t_SL U21776 (.Y(n18563),
	.A(n25635),
	.B(n18560),
	.C(n23687));
   NAND2xp33_ASAP7_75t_L U21777 (.Y(n20633),
	.A(n18540),
	.B(n20617));
   NOR2x1p5_ASAP7_75t_SL U21778 (.Y(n23698),
	.A(FE_OFN28815_n18523),
	.B(n21639));
   NAND2xp33_ASAP7_75t_SRAM U21780 (.Y(n18539),
	.A(n21691),
	.B(n18605));
   NAND2xp5_ASAP7_75t_L U21782 (.Y(n18567),
	.A(n21664),
	.B(n23678));
   NOR2xp33_ASAP7_75t_SL U21785 (.Y(n23196),
	.A(n23194),
	.B(n23193));
   NAND2xp33_ASAP7_75t_SRAM U21786 (.Y(n23181),
	.A(n23177),
	.B(n23178));
   NAND2x1_ASAP7_75t_L U21787 (.Y(n23200),
	.A(n22307),
	.B(n22306));
   NOR2x1_ASAP7_75t_L U21788 (.Y(n22306),
	.A(n22305),
	.B(n22304));
   NOR2x1p5_ASAP7_75t_SL U21789 (.Y(n23169),
	.A(n21772),
	.B(n18186));
   NOR2xp33_ASAP7_75t_SL U21790 (.Y(n23170),
	.A(FE_OFN28980_n18169),
	.B(n23303));
   NOR2xp67_ASAP7_75t_L U21791 (.Y(n23168),
	.A(n23160),
	.B(n18178));
   OAI22xp33_ASAP7_75t_L U21792 (.Y(n23190),
	.A1(n23336),
	.A2(n23161),
	.B1(FE_OFN25952_n22312),
	.B2(n23161));
   NAND2xp5_ASAP7_75t_L U21794 (.Y(n20776),
	.A(n20771),
	.B(n20770));
   NAND2xp33_ASAP7_75t_L U21795 (.Y(n20770),
	.A(n20769),
	.B(n20768));
   NAND2xp33_ASAP7_75t_L U21796 (.Y(n20771),
	.A(n20767),
	.B(n20768));
   NAND3xp33_ASAP7_75t_SL U21797 (.Y(n20778),
	.A(n21119),
	.B(n20773),
	.C(n20744));
   NAND2xp33_ASAP7_75t_L U21798 (.Y(n20744),
	.A(n20743),
	.B(n20742));
   NAND2xp33_ASAP7_75t_R U21799 (.Y(n20742),
	.A(n20741),
	.B(n20740));
   NAND2xp33_ASAP7_75t_R U21800 (.Y(n20743),
	.A(n20738),
	.B(n20740));
   NAND2x1_ASAP7_75t_SL U21801 (.Y(n22304),
	.A(n22862),
	.B(n20725));
   NOR3xp33_ASAP7_75t_SL U21802 (.Y(n20725),
	.A(n20724),
	.B(n22827),
	.C(n20749));
   NAND3xp33_ASAP7_75t_SL U21803 (.Y(n20724),
	.A(n21126),
	.B(n21103),
	.C(n21787));
   NAND2xp33_ASAP7_75t_R U21805 (.Y(n20718),
	.A(n20717),
	.B(FE_OFN28647_n21764));
   NAND2xp33_ASAP7_75t_R U21806 (.Y(n20719),
	.A(n20715),
	.B(FE_OFN28647_n21764));
   NOR2x1_ASAP7_75t_L U21807 (.Y(n20702),
	.A(n21130),
	.B(FE_OCPN5182_n21090));
   NAND2xp5_ASAP7_75t_SL U21808 (.Y(n20729),
	.A(FE_OFN55_sa22_5),
	.B(FE_OFN26133_sa22_3));
   NOR2xp33_ASAP7_75t_L U21809 (.Y(n21096),
	.A(n22838),
	.B(n21802));
   NOR2xp33_ASAP7_75t_SL U21810 (.Y(n21094),
	.A(n22278),
	.B(n20746));
   NOR3xp33_ASAP7_75t_R U21812 (.Y(n21137),
	.A(n21136),
	.B(n22321),
	.C(n22825));
   NOR3xp33_ASAP7_75t_SL U21813 (.Y(n21138),
	.A(n21134),
	.B(n21764),
	.C(n23194));
   NAND3xp33_ASAP7_75t_SL U21814 (.Y(n21140),
	.A(n21116),
	.B(n22802),
	.C(n22852));
   NAND3xp33_ASAP7_75t_L U21815 (.Y(n21141),
	.A(n21113),
	.B(n21112),
	.C(n21111));
   NAND2xp33_ASAP7_75t_L U21816 (.Y(n21112),
	.A(n21110),
	.B(n21109));
   NAND2xp33_ASAP7_75t_R U21818 (.Y(n21109),
	.A(n23299),
	.B(n21108));
   NAND2x1p5_ASAP7_75t_L U21819 (.Y(n21124),
	.A(n22795),
	.B(n23336));
   NOR2x1p5_ASAP7_75t_SL U21820 (.Y(n21122),
	.A(FE_OFN25987_n23322),
	.B(n21772));
   NAND3x1_ASAP7_75t_L U21821 (.Y(n23312),
	.A(FE_OFN28680_n),
	.B(n20739),
	.C(FE_OCPN27750_n22293));
   NAND2xp5_ASAP7_75t_SL U21822 (.Y(n22824),
	.A(n22820),
	.B(n22819));
   NAND2xp5_ASAP7_75t_L U21823 (.Y(n22823),
	.A(n22822),
	.B(n22819));
   NAND2xp5_ASAP7_75t_L U21824 (.Y(n22833),
	.A(n22832),
	.B(n22831));
   NAND2xp33_ASAP7_75t_R U21825 (.Y(n22832),
	.A(n22826),
	.B(n22829));
   NAND2xp33_ASAP7_75t_R U21826 (.Y(n22831),
	.A(n22830),
	.B(n22829));
   NAND3xp33_ASAP7_75t_SL U21828 (.Y(n22864),
	.A(n22853),
	.B(n23172),
	.C(n22852));
   NAND2xp33_ASAP7_75t_SL U21829 (.Y(n22853),
	.A(n23183),
	.B(n22851));
   NOR3xp33_ASAP7_75t_SRAM U21831 (.Y(n22860),
	.A(n23162),
	.B(FE_OFN28505_n23296),
	.C(n22859));
   NOR3xp33_ASAP7_75t_SL U21832 (.Y(n22861),
	.A(n22858),
	.B(FE_OFN25941_n22857),
	.C(n22856));
   NAND3xp33_ASAP7_75t_SL U21833 (.Y(n22865),
	.A(n23195),
	.B(n22849),
	.C(n22848));
   NAND2xp33_ASAP7_75t_L U21834 (.Y(n22849),
	.A(n22847),
	.B(n22846));
   NAND2xp33_ASAP7_75t_R U21835 (.Y(n22846),
	.A(n22845),
	.B(n23176));
   NAND2xp33_ASAP7_75t_R U21836 (.Y(n22847),
	.A(n22844),
	.B(n23176));
   NAND2xp5_ASAP7_75t_L U21837 (.Y(n23331),
	.A(n22817),
	.B(n22816));
   NAND2xp5_ASAP7_75t_L U21838 (.Y(n22816),
	.A(n22815),
	.B(n22814));
   NAND2xp5_ASAP7_75t_SL U21839 (.Y(n22802),
	.A(FE_OFN26141_n23307),
	.B(n22828));
   INVxp67_ASAP7_75t_R U21840 (.Y(n23185),
	.A(n18214));
   NAND2xp5_ASAP7_75t_L U21841 (.Y(n22801),
	.A(FE_OFN25952_n22312),
	.B(FE_OCPN27721_n23336));
   NOR2xp33_ASAP7_75t_L U21842 (.Y(n21775),
	.A(n22827),
	.B(FE_OFN28505_n23296));
   NOR2xp33_ASAP7_75t_L U21843 (.Y(n22800),
	.A(n20706),
	.B(n22825));
   NOR2x1_ASAP7_75t_SL U21844 (.Y(n22285),
	.A(n18190),
	.B(n24692));
   OAI21xp33_ASAP7_75t_L U21845 (.Y(n26870),
	.A1(n18186),
	.A2(n21772),
	.B(FE_OCPN28016_n21124));
   NOR2x1p5_ASAP7_75t_SL U21846 (.Y(n26872),
	.A(n22827),
	.B(n18188));
   NAND3x1_ASAP7_75t_SL U21847 (.Y(n18188),
	.A(n23311),
	.B(n21119),
	.C(n21801));
   NAND3x1_ASAP7_75t_SL U21848 (.Y(n26876),
	.A(n21111),
	.B(n18194),
	.C(n18197));
   NOR3xp33_ASAP7_75t_SL U21849 (.Y(n18194),
	.A(n18193),
	.B(n23161),
	.C(n22319));
   NAND3xp33_ASAP7_75t_L U21851 (.Y(n21234),
	.A(n18540),
	.B(n18529),
	.C(FE_OFN29131_FE_OCPN27371_sa20_2));
   NOR2x1_ASAP7_75t_L U21852 (.Y(n23777),
	.A(n23864),
	.B(n25632));
   NAND2xp5_ASAP7_75t_SRAM U21853 (.Y(n21235),
	.A(FE_OFN28986_n18597),
	.B(n20685));
   NOR3xp33_ASAP7_75t_L U21855 (.Y(n21259),
	.A(n21257),
	.B(n21256),
	.C(n23799));
   OAI21xp33_ASAP7_75t_SRAM U21856 (.Y(n21257),
	.A1(n18530),
	.A2(n23677),
	.B(n21254));
   NAND3xp33_ASAP7_75t_L U21857 (.Y(n21261),
	.A(n21252),
	.B(n21251),
	.C(n21250));
   NAND2xp33_ASAP7_75t_L U21858 (.Y(n21251),
	.A(n21245),
	.B(n21244));
   NAND2xp33_ASAP7_75t_L U21859 (.Y(n21250),
	.A(n21249),
	.B(n21248));
   NOR3xp33_ASAP7_75t_SRAM U21860 (.Y(n21252),
	.A(n21241),
	.B(n23863),
	.C(n23835));
   NAND3xp33_ASAP7_75t_L U21861 (.Y(n21237),
	.A(n21222),
	.B(n23803),
	.C(n21636));
   NAND2xp5_ASAP7_75t_R U21862 (.Y(n21222),
	.A(n21214),
	.B(n21213));
   NAND2xp33_ASAP7_75t_L U21863 (.Y(n21213),
	.A(n21212),
	.B(n23832));
   O2A1O1Ixp5_ASAP7_75t_SL U21864 (.Y(n25901),
	.A1(FE_OFN28986_n18597),
	.A2(n20617),
	.B(FE_OCPN27896_n18583),
	.C(n23814));
   O2A1O1Ixp33_ASAP7_75t_L U21865 (.Y(n25903),
	.A1(FE_OFN29076_n18540),
	.A2(FE_OFN28868_FE_OCPN27715_n23875),
	.B(FE_OFN28986_n18597),
	.C(n21682));
   NAND2x1_ASAP7_75t_L U21866 (.Y(n25189),
	.A(FE_OCPN27896_n18583),
	.B(n21669));
   NAND3xp33_ASAP7_75t_SL U21867 (.Y(n21698),
	.A(FE_PSN8329_n21638),
	.B(n21239),
	.C(n21238));
   NOR3xp33_ASAP7_75t_SRAM U21869 (.Y(n21695),
	.A(n21674),
	.B(n23835),
	.C(n21673));
   NAND2xp5_ASAP7_75t_L U21870 (.Y(n21694),
	.A(n21689),
	.B(n21688));
   NAND2xp33_ASAP7_75t_L U21871 (.Y(n21689),
	.A(n21685),
	.B(n21686));
   NOR3xp33_ASAP7_75t_R U21872 (.Y(n21671),
	.A(n21666),
	.B(n23831),
	.C(FE_OFN28607_n23884));
   O2A1O1Ixp33_ASAP7_75t_SRAM U21873 (.Y(n21670),
	.A1(n21669),
	.A2(n20617),
	.B(FE_OCPN27715_n23875),
	.C(n21668));
   NAND3xp33_ASAP7_75t_SL U21874 (.Y(n21647),
	.A(n20631),
	.B(n20630),
	.C(n20629));
   NAND2xp5_ASAP7_75t_SL U21875 (.Y(n20631),
	.A(n20622),
	.B(n20621));
   NAND2xp5_ASAP7_75t_SL U21876 (.Y(n20630),
	.A(n20628),
	.B(n20627));
   NAND2xp33_ASAP7_75t_L U21877 (.Y(n21661),
	.A(n21660),
	.B(n21659));
   NOR2xp33_ASAP7_75t_SRAM U21878 (.Y(n21660),
	.A(FE_OFN28868_FE_OCPN27715_n23875),
	.B(n21658));
   NAND2xp33_ASAP7_75t_L U21879 (.Y(n21662),
	.A(n21657),
	.B(n21659));
   NAND2x2_ASAP7_75t_SL U21880 (.Y(n23711),
	.A(FE_OFN29251_n18536),
	.B(n18521));
   NAND2xp5_ASAP7_75t_SL U21881 (.Y(n18587),
	.A(n18584),
	.B(FE_OCPN27531_n21643));
   NAND2xp5_ASAP7_75t_SL U21882 (.Y(n18586),
	.A(n18585),
	.B(FE_OCPN27531_n21643));
   NOR2xp67_ASAP7_75t_SL U21883 (.Y(n18584),
	.A(n18583),
	.B(n23830));
   NAND3xp33_ASAP7_75t_SL U21884 (.Y(n23733),
	.A(n23718),
	.B(n23717),
	.C(n23779));
   NOR3xp33_ASAP7_75t_SL U21886 (.Y(n23730),
	.A(n23723),
	.B(n23745),
	.C(n26900));
   NAND3xp33_ASAP7_75t_SRAM U21887 (.Y(n23734),
	.A(n23716),
	.B(n23715),
	.C(n23714));
   NAND3xp33_ASAP7_75t_L U21888 (.Y(n23713),
	.A(n25899),
	.B(n23709),
	.C(n23720));
   NOR3xp33_ASAP7_75t_SL U21889 (.Y(n18548),
	.A(n20670),
	.B(FE_OFN28791_n),
	.C(n18571));
   NAND2x2_ASAP7_75t_SL U21890 (.Y(n18530),
	.A(FE_OFN29131_FE_OCPN27371_sa20_2),
	.B(n18529));
   NOR3xp33_ASAP7_75t_R U21892 (.Y(n23868),
	.A(n23865),
	.B(n23864),
	.C(n23863));
   NAND2xp5_ASAP7_75t_SL U21893 (.Y(n23891),
	.A(n23887),
	.B(n23886));
   NOR3xp33_ASAP7_75t_SL U21894 (.Y(n23886),
	.A(n23885),
	.B(n23884),
	.C(n23883));
   NAND2xp5_ASAP7_75t_L U21895 (.Y(n23895),
	.A(n23878),
	.B(n23877));
   NAND2xp5_ASAP7_75t_L U21896 (.Y(n23877),
	.A(n23876),
	.B(n23873));
   NAND2xp33_ASAP7_75t_SL U21897 (.Y(n23878),
	.A(n23874),
	.B(n23873));
   NOR3xp33_ASAP7_75t_R U21898 (.Y(n23894),
	.A(FE_OFN28650_n23802),
	.B(n23880),
	.C(FE_PSN8332_n23879));
   AND3x1_ASAP7_75t_SRAM U21899 (.Y(n23857),
	.A(n25635),
	.B(FE_OFN28477_n23853),
	.C(n23852));
   NOR3xp33_ASAP7_75t_R U21900 (.Y(n18439),
	.A(n18431),
	.B(n18430),
	.C(FE_OCPN28078_n24296));
   NAND3xp33_ASAP7_75t_SL U21901 (.Y(n24298),
	.A(n16675),
	.B(n16680),
	.C(n16679));
   NOR3xp33_ASAP7_75t_R U21902 (.Y(n16680),
	.A(n16678),
	.B(FE_OCPN28141_n),
	.C(FE_OFN28918_n16949));
   NAND2xp33_ASAP7_75t_SRAM U21903 (.Y(n18411),
	.A(n18407),
	.B(n18408));
   NAND2xp33_ASAP7_75t_SRAM U21904 (.Y(n18410),
	.A(n18409),
	.B(n18408));
   OAI22xp33_ASAP7_75t_SRAM U21905 (.Y(n18404),
	.A1(FE_OFN29164_sa33_2),
	.A2(FE_OFN27090_n23558),
	.B1(FE_OFN28592_n16427),
	.B2(FE_OFN27090_n23558));
   NOR3xp33_ASAP7_75t_SL U21907 (.Y(n17438),
	.A(n17425),
	.B(n17424),
	.C(FE_OCPN29577_n24298));
   NOR3xp33_ASAP7_75t_SRAM U21908 (.Y(n17437),
	.A(FE_OCPN7595_n17426),
	.B(n18107),
	.C(n23538));
   AND2x2_ASAP7_75t_R U21909 (.Y(n17421),
	.A(n17420),
	.B(n26120));
   NAND2xp33_ASAP7_75t_SRAM U21910 (.Y(n17403),
	.A(n17397),
	.B(FE_OFN28935_n18104));
   NAND2xp5_ASAP7_75t_SL U21911 (.Y(n16935),
	.A(n26358),
	.B(n16917));
   NAND2xp5_ASAP7_75t_SL U21912 (.Y(n16917),
	.A(n16916),
	.B(n16915));
   NAND2xp33_ASAP7_75t_SL U21913 (.Y(n16916),
	.A(n16954),
	.B(n16914));
   NAND2xp33_ASAP7_75t_L U21914 (.Y(n16915),
	.A(n16956),
	.B(n16914));
   NOR3xp33_ASAP7_75t_R U21915 (.Y(n16933),
	.A(n16932),
	.B(n16931),
	.C(n16930));
   NAND2xp33_ASAP7_75t_SRAM U21916 (.Y(n16932),
	.A(n23533),
	.B(n17432));
   OAI21xp33_ASAP7_75t_SRAM U21917 (.Y(n16934),
	.A1(n16417),
	.A2(n16929),
	.B(n16928));
   NOR3xp33_ASAP7_75t_SL U21918 (.Y(n16967),
	.A(n16950),
	.B(FE_OFN28918_n16949),
	.C(n16948));
   NAND2xp33_ASAP7_75t_L U21919 (.Y(n16944),
	.A(n16943),
	.B(n16942));
   OAI21xp33_ASAP7_75t_L U21920 (.Y(n16966),
	.A1(n16965),
	.A2(n16964),
	.B(n24610));
   NAND3xp33_ASAP7_75t_L U21921 (.Y(n16964),
	.A(n16963),
	.B(n16962),
	.C(n23529));
   NAND2xp33_ASAP7_75t_L U21922 (.Y(n16963),
	.A(n16958),
	.B(n16957));
   NOR3xp33_ASAP7_75t_L U21923 (.Y(n16962),
	.A(n16961),
	.B(n16960),
	.C(n24485));
   NOR3xp33_ASAP7_75t_SL U21924 (.Y(n18108),
	.A(n16947),
	.B(FE_OFN28679_sa33_5),
	.C(FE_OFN25938_sa33_3));
   NOR3x1_ASAP7_75t_SL U21925 (.Y(n18105),
	.A(n17431),
	.B(n18143),
	.C(n17430));
   NAND3xp33_ASAP7_75t_L U21927 (.Y(n18150),
	.A(n23546),
	.B(n18418),
	.C(n18149));
   NAND3xp33_ASAP7_75t_L U21928 (.Y(n18151),
	.A(n18441),
	.B(n18148),
	.C(n18147));
   NAND3xp33_ASAP7_75t_SL U21929 (.Y(n18126),
	.A(n18125),
	.B(n18124),
	.C(n18123));
   NAND2xp33_ASAP7_75t_R U21930 (.Y(n18122),
	.A(n18119),
	.B(n18118));
   NAND2xp33_ASAP7_75t_R U21931 (.Y(n18118),
	.A(n18117),
	.B(n18116));
   NAND2xp33_ASAP7_75t_R U21932 (.Y(n18119),
	.A(n18115),
	.B(n18116));
   NAND2xp33_ASAP7_75t_SRAM U21933 (.Y(n18137),
	.A(n18134),
	.B(n18133));
   NOR3xp33_ASAP7_75t_SL U21934 (.Y(n23547),
	.A(n23545),
	.B(n23544),
	.C(n23543));
   NOR3xp33_ASAP7_75t_L U21935 (.Y(n23561),
	.A(n23559),
	.B(n23558),
	.C(n23557));
   OAI21xp33_ASAP7_75t_R U21936 (.Y(n23559),
	.A1(n23556),
	.A2(FE_OFN29208_n16436),
	.B(n23555));
   NOR3xp33_ASAP7_75t_R U21937 (.Y(n23555),
	.A(n23554),
	.B(n23553),
	.C(n23552));
   OR3x1_ASAP7_75t_L U21938 (.Y(n23534),
	.A(n18132),
	.B(n18426),
	.C(n18131));
   NAND2xp5_ASAP7_75t_L U21939 (.Y(n18132),
	.A(n18129),
	.B(n18128));
   NOR2x1_ASAP7_75t_SL U21941 (.Y(n23558),
	.A(n16429),
	.B(FE_OFN26545_n16447));
   NOR3x1_ASAP7_75t_R U21942 (.Y(n23530),
	.A(n16436),
	.B(FE_OFN28679_sa33_5),
	.C(n16676));
   NOR2x1_ASAP7_75t_L U21943 (.Y(n23552),
	.A(n16473),
	.B(n16874));
   NAND2xp5_ASAP7_75t_SL U21944 (.Y(n18406),
	.A(FE_OFN28592_n16427),
	.B(FE_OFN29101_n16418));
   NOR2x1_ASAP7_75t_R U21945 (.Y(n17408),
	.A(n23553),
	.B(n16833));
   NAND2xp5_ASAP7_75t_SRAM U21946 (.Y(n16833),
	.A(n16832),
	.B(n16880));
   NAND2xp5_ASAP7_75t_SL U21947 (.Y(n17404),
	.A(n16865),
	.B(n16864));
   NOR3xp33_ASAP7_75t_L U21948 (.Y(n16865),
	.A(n16856),
	.B(n18420),
	.C(FE_OCPN28141_n));
   NAND2xp5_ASAP7_75t_L U21949 (.Y(n16856),
	.A(n18140),
	.B(n18130));
   INVx1_ASAP7_75t_SL U21950 (.Y(n25006),
	.A(n25007));
   NAND3x1_ASAP7_75t_SL U21952 (.Y(n26568),
	.A(n22051),
	.B(n19007),
	.C(n22967));
   NAND3xp33_ASAP7_75t_R U21953 (.Y(n26569),
	.A(n20916),
	.B(n22007),
	.C(n19020));
   NAND3xp33_ASAP7_75t_SL U21954 (.Y(n19025),
	.A(n19024),
	.B(n19023),
	.C(n22978));
   NOR3xp33_ASAP7_75t_SL U21955 (.Y(n19023),
	.A(n19022),
	.B(n19021),
	.C(n26559));
   NAND3xp33_ASAP7_75t_L U21956 (.Y(n26550),
	.A(n19014),
	.B(n20238),
	.C(n20237));
   NOR3xp33_ASAP7_75t_SL U21957 (.Y(n22942),
	.A(n22933),
	.B(n26659),
	.C(n24769));
   NAND3x1_ASAP7_75t_SL U21959 (.Y(n22941),
	.A(FE_OCPN27986_n18970),
	.B(FE_OFN28752_n),
	.C(FE_OCPN29374_FE_OFN29191_sa23_2));
   NAND2xp33_ASAP7_75t_R U21960 (.Y(n22940),
	.A(n22939),
	.B(n22938));
   NAND2xp33_ASAP7_75t_SRAM U21961 (.Y(n22938),
	.A(n22937),
	.B(n22936));
   NOR3xp33_ASAP7_75t_L U21963 (.Y(n22958),
	.A(n22956),
	.B(n24765),
	.C(n22955));
   NAND2xp33_ASAP7_75t_L U21964 (.Y(n22922),
	.A(n22928),
	.B(n20922));
   NAND2xp33_ASAP7_75t_SRAM U21965 (.Y(n22919),
	.A(n22918),
	.B(FE_OFN16250_n26165));
   NAND2xp33_ASAP7_75t_SRAM U21966 (.Y(n22920),
	.A(n22916),
	.B(FE_OFN16250_n26165));
   NOR2xp33_ASAP7_75t_SRAM U21967 (.Y(n22916),
	.A(FE_OFN29026_n20911),
	.B(n22998));
   NAND2xp33_ASAP7_75t_SRAM U21968 (.Y(n24775),
	.A(FE_OCPN27986_n18970),
	.B(FE_OFN28787_n19000));
   NOR2x1_ASAP7_75t_L U21969 (.Y(n20234),
	.A(n22973),
	.B(n19314));
   NAND2xp5_ASAP7_75t_L U21970 (.Y(n19314),
	.A(n20941),
	.B(n20930));
   NAND2xp33_ASAP7_75t_SRAM U21971 (.Y(n22038),
	.A(FE_OFN29189_sa23_0),
	.B(n19000));
   NOR3xp33_ASAP7_75t_SL U21973 (.Y(n20279),
	.A(n20271),
	.B(n20270),
	.C(n20269));
   NAND2xp5_ASAP7_75t_L U21974 (.Y(n20278),
	.A(n20277),
	.B(n20276));
   NAND3xp33_ASAP7_75t_SL U21975 (.Y(n20281),
	.A(n20254),
	.B(n20253),
	.C(n24041));
   NOR3xp33_ASAP7_75t_SL U21976 (.Y(n20253),
	.A(n20248),
	.B(n23473),
	.C(n22031));
   NAND2xp33_ASAP7_75t_SRAM U21977 (.Y(n20239),
	.A(n20238),
	.B(n22046));
   NAND3x1_ASAP7_75t_SL U21978 (.Y(n22923),
	.A(n26152),
	.B(n19334),
	.C(n26151));
   NOR3xp33_ASAP7_75t_SL U21979 (.Y(n19334),
	.A(n19331),
	.B(FE_OFN26542_n26155),
	.C(n26154));
   OAI21xp33_ASAP7_75t_SRAM U21980 (.Y(n22003),
	.A1(FE_OCPN28363_n22979),
	.A2(n22980),
	.B(n19329));
   NAND2xp5_ASAP7_75t_L U21981 (.Y(n22006),
	.A(n26660),
	.B(FE_OCPN29480_n20913));
   NAND3xp33_ASAP7_75t_R U21982 (.Y(n22007),
	.A(FE_OCPN27627_sa23_1),
	.B(n18971),
	.C(n19313));
   NAND3xp33_ASAP7_75t_SL U21983 (.Y(n22013),
	.A(n20267),
	.B(n20266),
	.C(n22039));
   NAND2xp5_ASAP7_75t_SL U21984 (.Y(n20266),
	.A(n20264),
	.B(n20263));
   NAND2xp5_ASAP7_75t_L U21985 (.Y(n20263),
	.A(n20262),
	.B(n20261));
   NAND2x1_ASAP7_75t_SL U21986 (.Y(n23514),
	.A(n22012),
	.B(n22011));
   NAND2xp5_ASAP7_75t_L U21988 (.Y(n22002),
	.A(n22046),
	.B(n26160));
   NAND2x1_ASAP7_75t_L U21989 (.Y(n25717),
	.A(FE_OCPN28112_n26664),
	.B(n26660));
   NAND2xp33_ASAP7_75t_SRAM U21990 (.Y(n25716),
	.A(FE_OFN29026_n20911),
	.B(FE_OCPN27727_n22964));
   NAND3xp33_ASAP7_75t_SL U21992 (.Y(n19006),
	.A(n23511),
	.B(n20238),
	.C(n19343));
   NAND3x1_ASAP7_75t_SL U21993 (.Y(n23515),
	.A(n22984),
	.B(n22983),
	.C(n22982));
   NAND3xp33_ASAP7_75t_SL U21994 (.Y(n23006),
	.A(n22994),
	.B(n23501),
	.C(n23517));
   NOR3xp33_ASAP7_75t_R U21996 (.Y(n22974),
	.A(n22973),
	.B(n22972),
	.C(n26148));
   NAND2xp5_ASAP7_75t_SL U21997 (.Y(n22976),
	.A(n19344),
	.B(n20250));
   NAND2xp5_ASAP7_75t_R U21998 (.Y(n22605),
	.A(FE_OCPN27887_n17331),
	.B(n17382));
   NAND2x1_ASAP7_75t_SL U21999 (.Y(n20367),
	.A(FE_OFN27152_n17315),
	.B(n27007));
   NOR2x1_ASAP7_75t_L U22000 (.Y(n21557),
	.A(n22592),
	.B(n18669));
   NAND2xp33_ASAP7_75t_L U22001 (.Y(n18669),
	.A(n22421),
	.B(n21540));
   NOR3xp33_ASAP7_75t_SL U22003 (.Y(n18728),
	.A(n18725),
	.B(n21560),
	.C(n18724));
   NAND2xp33_ASAP7_75t_L U22005 (.Y(n18715),
	.A(n24389),
	.B(n24390));
   NAND2xp5_ASAP7_75t_L U22006 (.Y(n23112),
	.A(n23111),
	.B(n23110));
   NAND2xp33_ASAP7_75t_SL U22007 (.Y(n23110),
	.A(n23109),
	.B(n23108));
   NOR2xp33_ASAP7_75t_L U22008 (.Y(n23109),
	.A(FE_OFN16208_n23101),
	.B(n23106));
   NOR3xp33_ASAP7_75t_SRAM U22009 (.Y(n23084),
	.A(n23083),
	.B(FE_OCPN28397_n23082),
	.C(n27012));
   NOR3xp33_ASAP7_75t_SRAM U22010 (.Y(n23085),
	.A(n23081),
	.B(n23092),
	.C(n23080));
   NAND2xp33_ASAP7_75t_L U22011 (.Y(n23081),
	.A(n23074),
	.B(FE_OFN28558_n23073));
   NAND2xp5_ASAP7_75t_L U22012 (.Y(n23096),
	.A(n23091),
	.B(n23090));
   NAND2xp5_ASAP7_75t_R U22013 (.Y(n23090),
	.A(n23089),
	.B(n23088));
   NAND2xp5_ASAP7_75t_R U22014 (.Y(n23091),
	.A(n23086),
	.B(n23088));
   NAND2xp5_ASAP7_75t_R U22015 (.Y(n23069),
	.A(FE_OCPN29309_n26452),
	.B(n18677));
   NOR3x1_ASAP7_75t_L U22016 (.Y(n25057),
	.A(n20366),
	.B(n22436),
	.C(n20365));
   NAND2xp33_ASAP7_75t_L U22017 (.Y(n23068),
	.A(n23067),
	.B(n23066));
   NAND2xp33_ASAP7_75t_R U22018 (.Y(n23066),
	.A(n23065),
	.B(n23064));
   NAND2xp33_ASAP7_75t_R U22019 (.Y(n23067),
	.A(n23061),
	.B(n23064));
   NOR3xp33_ASAP7_75t_SL U22020 (.Y(n24221),
	.A(n17379),
	.B(n17383),
	.C(n18666));
   NAND3xp33_ASAP7_75t_SL U22021 (.Y(n24227),
	.A(n22182),
	.B(n22589),
	.C(n21554));
   NAND2xp33_ASAP7_75t_L U22022 (.Y(n24228),
	.A(n22432),
	.B(n17380));
   NOR3x1_ASAP7_75t_L U22023 (.Y(n24222),
	.A(n17371),
	.B(n23087),
	.C(FE_OFN78_n22457));
   NOR3xp33_ASAP7_75t_SL U22024 (.Y(n24220),
	.A(n17333),
	.B(n27006),
	.C(n18717));
   NOR2x1_ASAP7_75t_SL U22025 (.Y(n22584),
	.A(n18693),
	.B(n22450));
   NOR3x1_ASAP7_75t_SL U22026 (.Y(n22585),
	.A(n18684),
	.B(FE_OFN28736_FE_OCPN28216_sa01_5),
	.C(n18693));
   NOR3xp33_ASAP7_75t_SRAM U22027 (.Y(n27002),
	.A(n22583),
	.B(n22582),
	.C(n23092));
   NAND2x1p5_ASAP7_75t_SL U22029 (.Y(n27012),
	.A(n21535),
	.B(n22458));
   NAND2xp5_ASAP7_75t_L U22030 (.Y(n27011),
	.A(n22415),
	.B(FE_OCPN5188_n22414));
   NAND2xp33_ASAP7_75t_R U22031 (.Y(n22578),
	.A(n22576),
	.B(n27008));
   NAND2xp33_ASAP7_75t_R U22032 (.Y(n22445),
	.A(n22444),
	.B(n22443));
   NAND2xp33_ASAP7_75t_SRAM U22033 (.Y(n22443),
	.A(n22442),
	.B(FE_OFN27064_n22438));
   NOR3x1_ASAP7_75t_SL U22034 (.Y(n22456),
	.A(n18712),
	.B(n20401),
	.C(n18711));
   NOR3xp33_ASAP7_75t_SRAM U22035 (.Y(n18711),
	.A(FE_OCPN29406_n18710),
	.B(FE_OCPN29429_FE_OFN16141_sa01_3),
	.C(FE_OCPN28217_sa01_5));
   NAND2xp5_ASAP7_75t_L U22036 (.Y(n18705),
	.A(n18703),
	.B(n18702));
   NOR3xp33_ASAP7_75t_SRAM U22037 (.Y(n22455),
	.A(n22452),
	.B(n26461),
	.C(n22451));
   OAI21xp33_ASAP7_75t_SRAM U22038 (.Y(n22452),
	.A1(FE_OCPN28000_n22450),
	.A2(n23107),
	.B(n22449));
   NOR3xp33_ASAP7_75t_SL U22039 (.Y(n22474),
	.A(n22583),
	.B(n23099),
	.C(n23062));
   NOR3xp33_ASAP7_75t_L U22040 (.Y(n22473),
	.A(n22472),
	.B(n23083),
	.C(n22471));
   NAND3xp33_ASAP7_75t_L U22041 (.Y(n22472),
	.A(n23097),
	.B(n27008),
	.C(n22467));
   NAND2xp33_ASAP7_75t_L U22043 (.Y(n22427),
	.A(n22423),
	.B(n22424));
   NAND2xp33_ASAP7_75t_R U22044 (.Y(n22426),
	.A(n22425),
	.B(n22424));
   NAND2xp33_ASAP7_75t_SRAM U22045 (.Y(n22419),
	.A(n22418),
	.B(n22417));
   NAND2xp33_ASAP7_75t_SRAM U22046 (.Y(n19542),
	.A(n22778),
	.B(n23235));
   NAND3xp33_ASAP7_75t_SRAM U22047 (.Y(n19537),
	.A(n23608),
	.B(n19520),
	.C(n22244));
   NAND3xp33_ASAP7_75t_SL U22048 (.Y(n23572),
	.A(n19536),
	.B(n23613),
	.C(FE_OCPN8224_n22773));
   NOR3xp33_ASAP7_75t_L U22049 (.Y(n19536),
	.A(n22760),
	.B(n20596),
	.C(n22743));
   NAND3x1_ASAP7_75t_L U22050 (.Y(n22247),
	.A(n17977),
	.B(n17919),
	.C(n17918));
   NOR3xp33_ASAP7_75t_L U22051 (.Y(n17919),
	.A(n17917),
	.B(n24370),
	.C(n20562));
   NAND3xp33_ASAP7_75t_L U22052 (.Y(n17917),
	.A(n22722),
	.B(n20595),
	.C(n24592));
   NOR2xp33_ASAP7_75t_L U22054 (.Y(n19565),
	.A(n20584),
	.B(n19563));
   NOR3xp33_ASAP7_75t_L U22055 (.Y(n19564),
	.A(n23224),
	.B(n22750),
	.C(n23581));
   NAND3xp33_ASAP7_75t_L U22056 (.Y(n19563),
	.A(n20791),
	.B(n20819),
	.C(n24586));
   NOR2xp33_ASAP7_75t_SRAM U22057 (.Y(n19506),
	.A(FE_OFN29075_n22745),
	.B(FE_OFN28654_n22751));
   NAND3xp33_ASAP7_75t_SRAM U22058 (.Y(n20792),
	.A(n20814),
	.B(n24056),
	.C(n20542));
   OAI21xp33_ASAP7_75t_SRAM U22059 (.Y(n19515),
	.A1(n19510),
	.A2(n19509),
	.B(n24592));
   NAND2xp33_ASAP7_75t_R U22060 (.Y(n19508),
	.A(n19504),
	.B(n19505));
   NOR2xp33_ASAP7_75t_SRAM U22061 (.Y(n19504),
	.A(n24362),
	.B(FE_OFN28654_n22751));
   NOR2xp33_ASAP7_75t_L U22062 (.Y(n22752),
	.A(FE_OFN26158_n22224),
	.B(n17935));
   INVxp33_ASAP7_75t_L U22063 (.Y(n17935),
	.A(n24362));
   OAI21xp33_ASAP7_75t_L U22066 (.Y(n17979),
	.A1(n24051),
	.A2(n17978),
	.B(n25682));
   NAND3xp33_ASAP7_75t_L U22067 (.Y(n17978),
	.A(n17977),
	.B(n17976),
	.C(n22261));
   NOR3xp33_ASAP7_75t_R U22068 (.Y(n17976),
	.A(n17975),
	.B(n22235),
	.C(n17974));
   NAND2xp33_ASAP7_75t_SL U22069 (.Y(n17974),
	.A(n22251),
	.B(n22228));
   NOR3xp33_ASAP7_75t_SL U22070 (.Y(n17980),
	.A(n17956),
	.B(n24055),
	.C(n17955));
   NAND3xp33_ASAP7_75t_L U22071 (.Y(n17956),
	.A(n22728),
	.B(n20828),
	.C(n22253));
   NOR2xp33_ASAP7_75t_SL U22072 (.Y(n17938),
	.A(n22247),
	.B(n17934));
   NAND3xp33_ASAP7_75t_L U22073 (.Y(n17934),
	.A(n22786),
	.B(n22720),
	.C(n19534));
   NAND2xp5_ASAP7_75t_L U22074 (.Y(n25737),
	.A(n20550),
	.B(n17907));
   NOR2xp33_ASAP7_75t_L U22075 (.Y(n17907),
	.A(n23214),
	.B(n23602));
   NAND2xp5_ASAP7_75t_SL U22076 (.Y(n23616),
	.A(n17904),
	.B(n17903));
   NAND2xp33_ASAP7_75t_R U22077 (.Y(n17904),
	.A(n17902),
	.B(n17901));
   INVxp33_ASAP7_75t_SRAM U22078 (.Y(n22740),
	.A(n22739));
   NAND2xp33_ASAP7_75t_L U22079 (.Y(n22741),
	.A(n22738),
	.B(n22737));
   NAND2xp33_ASAP7_75t_SRAM U22080 (.Y(n22738),
	.A(n22736),
	.B(n22735));
   NAND2xp33_ASAP7_75t_L U22083 (.Y(n22787),
	.A(n22785),
	.B(n22784));
   NAND2xp33_ASAP7_75t_R U22084 (.Y(n22784),
	.A(n22783),
	.B(n22782));
   NAND2xp33_ASAP7_75t_SL U22085 (.Y(n22785),
	.A(n22780),
	.B(n22782));
   NAND2xp33_ASAP7_75t_SL U22086 (.Y(n22790),
	.A(n23598),
	.B(n22256));
   NAND3xp33_ASAP7_75t_SL U22087 (.Y(n22789),
	.A(n22764),
	.B(n22763),
	.C(n22762));
   NOR3xp33_ASAP7_75t_SRAM U22088 (.Y(n22763),
	.A(n22761),
	.B(FE_OFN28475_n23573),
	.C(n22760));
   NAND3x1_ASAP7_75t_SL U22089 (.Y(n23237),
	.A(n22755),
	.B(n22754),
	.C(n23611));
   NAND2xp5_ASAP7_75t_SL U22090 (.Y(n22755),
	.A(n22748),
	.B(n22747));
   NOR3xp33_ASAP7_75t_SL U22091 (.Y(n22754),
	.A(n25740),
	.B(FE_OFN28723_n22750),
	.C(n23602));
   NAND2xp33_ASAP7_75t_SL U22092 (.Y(n22747),
	.A(n22746),
	.B(n20814));
   NOR2xp67_ASAP7_75t_L U22093 (.Y(n22718),
	.A(FE_OFN26158_n22224),
	.B(n22223));
   NAND2xp5_ASAP7_75t_SL U22094 (.Y(n22719),
	.A(n19541),
	.B(n19540));
   NOR2xp67_ASAP7_75t_SL U22095 (.Y(n19541),
	.A(n22781),
	.B(n20540));
   NOR3x1_ASAP7_75t_SL U22096 (.Y(n24370),
	.A(FE_OFN27145_n23216),
	.B(FE_OFN28882_FE_OCPN27356_sa12_0),
	.C(n17952));
   NAND2xp33_ASAP7_75t_R U22097 (.Y(n22756),
	.A(n23242),
	.B(n22725));
   NAND2xp5_ASAP7_75t_SL U22098 (.Y(n22720),
	.A(n17929),
	.B(FE_OFN26589_sa12_1));
   NAND2xp33_ASAP7_75t_SL U22099 (.Y(n17929),
	.A(n17927),
	.B(n17926));
   NOR2xp33_ASAP7_75t_L U22100 (.Y(n17927),
	.A(FE_OCPN29511_n22226),
	.B(n23573));
   INVxp67_ASAP7_75t_L U22101 (.Y(n17926),
	.A(n17925));
   NAND2x1_ASAP7_75t_SL U22102 (.Y(n23235),
	.A(FE_OCPN5137_n23600),
	.B(n24367));
   NOR3x1_ASAP7_75t_L U22103 (.Y(n22726),
	.A(n19502),
	.B(FE_OCPN29494_sa12_4),
	.C(n17949));
   NAND2xp33_ASAP7_75t_SRAM U22104 (.Y(n22234),
	.A(FE_OFN25907_sa12_2),
	.B(n22233));
   NAND3xp33_ASAP7_75t_L U22105 (.Y(n22262),
	.A(n22261),
	.B(n22260),
	.C(n23240));
   NOR3xp33_ASAP7_75t_L U22106 (.Y(n22260),
	.A(n22257),
	.B(n23588),
	.C(n22790));
   NAND3xp33_ASAP7_75t_SRAM U22107 (.Y(n22257),
	.A(n22252),
	.B(n22251),
	.C(n22250));
   NAND2xp33_ASAP7_75t_L U22108 (.Y(n22241),
	.A(n22762),
	.B(n22764));
   NAND2xp5_ASAP7_75t_R U22109 (.Y(n22242),
	.A(n20602),
	.B(n20812));
   NAND3xp33_ASAP7_75t_R U22110 (.Y(n22229),
	.A(n22228),
	.B(n23612),
	.C(n22227));
   NAND3xp33_ASAP7_75t_L U22111 (.Y(n22230),
	.A(FE_OCPN28309_n22779),
	.B(n22226),
	.C(n22225));
   NOR2xp33_ASAP7_75t_L U22112 (.Y(n24591),
	.A(n22751),
	.B(n22765));
   NAND3x1_ASAP7_75t_SL U22113 (.Y(n24589),
	.A(n23595),
	.B(n20809),
	.C(n22758));
   NOR3xp33_ASAP7_75t_SL U22114 (.Y(n20809),
	.A(n22719),
	.B(n22233),
	.C(FE_OFN26556_n23236));
   NAND3xp33_ASAP7_75t_SL U22115 (.Y(n23585),
	.A(n17948),
	.B(n17947),
	.C(n22250));
   NOR3xp33_ASAP7_75t_R U22116 (.Y(n17948),
	.A(n22774),
	.B(n20596),
	.C(FE_OFN28567_n19514));
   NAND2xp5_ASAP7_75t_L U22117 (.Y(n17947),
	.A(n17944),
	.B(n17943));
   NAND2xp33_ASAP7_75t_SL U22118 (.Y(n17943),
	.A(n17942),
	.B(n17941));
   NOR2x1_ASAP7_75t_L U22119 (.Y(n23584),
	.A(n22752),
	.B(n24370));
   NOR2xp33_ASAP7_75t_SRAM U22120 (.Y(n23575),
	.A(n24364),
	.B(n24363));
   NOR2xp33_ASAP7_75t_R U22122 (.Y(n23577),
	.A(FE_OCPN27729_n24362),
	.B(n24363));
   NOR3xp33_ASAP7_75t_SL U22123 (.Y(n24365),
	.A(n23574),
	.B(FE_OFN28475_n23573),
	.C(n23572));
   NAND3xp33_ASAP7_75t_SL U22124 (.Y(n20826),
	.A(n20819),
	.B(n20818),
	.C(n20817));
   NOR3xp33_ASAP7_75t_L U22125 (.Y(n20818),
	.A(n20816),
	.B(n23225),
	.C(n24368));
   NOR2x1p5_ASAP7_75t_SL U22126 (.Y(n25439),
	.A(FE_OCPN29492_sa12_4),
	.B(n17921));
   NAND3x1_ASAP7_75t_SL U22127 (.Y(n26599),
	.A(FE_OCPN28309_n22779),
	.B(n20558),
	.C(n20789));
   NAND2x1_ASAP7_75t_SL U22128 (.Y(n25438),
	.A(n22228),
	.B(n22778));
   NOR3xp33_ASAP7_75t_SL U22129 (.Y(n27101),
	.A(n25283),
	.B(n25282),
	.C(n25281));
   NAND3xp33_ASAP7_75t_L U22130 (.Y(n25283),
	.A(n25280),
	.B(n25279),
	.C(n25880));
   NOR2x1_ASAP7_75t_SL U22131 (.Y(n19924),
	.A(n18846),
	.B(n22368));
   NAND2xp5_ASAP7_75t_R U22132 (.Y(n18317),
	.A(n18316),
	.B(n24646));
   NAND2xp33_ASAP7_75t_L U22133 (.Y(n18318),
	.A(n18315),
	.B(n24646));
   NAND3xp33_ASAP7_75t_SL U22135 (.Y(n17598),
	.A(n20093),
	.B(n22386),
	.C(n17579));
   NOR2xp33_ASAP7_75t_SL U22136 (.Y(n17596),
	.A(n20112),
	.B(n17595));
   NOR3xp33_ASAP7_75t_SL U22137 (.Y(n23898),
	.A(n17562),
	.B(FE_OFN16232_n17691),
	.C(n20106));
   NAND3xp33_ASAP7_75t_L U22138 (.Y(n17562),
	.A(n19956),
	.B(n24853),
	.C(n24645));
   NAND3x1_ASAP7_75t_SL U22139 (.Y(n19720),
	.A(FE_OCPN29449_n17521),
	.B(FE_OCPN28434_n17546),
	.C(FE_OCPN29421_FE_OFN16128_sa32_2));
   NAND2xp33_ASAP7_75t_R U22140 (.Y(n18812),
	.A(n18810),
	.B(n18809));
   NAND2xp33_ASAP7_75t_R U22141 (.Y(n18809),
	.A(n18808),
	.B(n18807));
   NAND2xp33_ASAP7_75t_SRAM U22142 (.Y(n18810),
	.A(n18806),
	.B(n18807));
   NOR2xp33_ASAP7_75t_SL U22144 (.Y(n18823),
	.A(n18822),
	.B(n18821));
   OAI21xp33_ASAP7_75t_SRAM U22145 (.Y(n18822),
	.A1(n18818),
	.A2(FE_OCPN27882_n18829),
	.B(n25025));
   NAND2xp33_ASAP7_75t_R U22147 (.Y(n18849),
	.A(n18845),
	.B(n18848));
   NOR3xp33_ASAP7_75t_SL U22148 (.Y(n18850),
	.A(n22387),
	.B(n24991),
	.C(n22398));
   NAND3xp33_ASAP7_75t_L U22149 (.Y(n18853),
	.A(n18835),
	.B(n18834),
	.C(n18833));
   NOR3xp33_ASAP7_75t_SL U22151 (.Y(n18835),
	.A(n18831),
	.B(n18830),
	.C(n19919));
   NAND3xp33_ASAP7_75t_SL U22153 (.Y(n19935),
	.A(n18801),
	.B(n18800),
	.C(n18824));
   NAND2xp33_ASAP7_75t_SRAM U22155 (.Y(n18792),
	.A(n24856),
	.B(n18790));
   NOR2xp67_ASAP7_75t_L U22156 (.Y(n22367),
	.A(FE_OCPN29348_n17592),
	.B(n17700));
   NAND2xp33_ASAP7_75t_L U22157 (.Y(n22366),
	.A(FE_OFN16231_n17691),
	.B(n18330));
   NOR3x1_ASAP7_75t_L U22158 (.Y(n22368),
	.A(FE_OCPN29348_n17592),
	.B(FE_OCPN29459_n),
	.C(FE_OCPN29323_n19721));
   NOR3x1_ASAP7_75t_R U22159 (.Y(n22369),
	.A(FE_OCPN29348_n17592),
	.B(FE_OCPN29459_n),
	.C(FE_OCPN27882_n18829));
   NAND2xp5_ASAP7_75t_L U22160 (.Y(n22372),
	.A(n17527),
	.B(n17546));
   NOR3xp33_ASAP7_75t_SRAM U22161 (.Y(n22402),
	.A(n22400),
	.B(n22399),
	.C(n22398));
   NAND3xp33_ASAP7_75t_L U22162 (.Y(n22407),
	.A(n22391),
	.B(n22390),
	.C(n22389));
   NOR2xp33_ASAP7_75t_L U22163 (.Y(n22391),
	.A(n22388),
	.B(n22387));
   NAND2xp33_ASAP7_75t_SRAM U22165 (.Y(n22394),
	.A(FE_OCPN29449_n17521),
	.B(n22392));
   NAND3x1_ASAP7_75t_SL U22166 (.Y(n22380),
	.A(n17697),
	.B(n18309),
	.C(n17696));
   NOR2xp67_ASAP7_75t_SL U22167 (.Y(n17696),
	.A(n17695),
	.B(n17694));
   NAND2xp5_ASAP7_75t_L U22168 (.Y(n17695),
	.A(n17711),
	.B(n20117));
   NAND2xp33_ASAP7_75t_L U22169 (.Y(n22381),
	.A(n18839),
	.B(n22397));
   NAND2xp33_ASAP7_75t_L U22170 (.Y(n22385),
	.A(n18300),
	.B(n18299));
   OAI21xp33_ASAP7_75t_SL U22171 (.Y(n22383),
	.A1(FE_OFN69_sa32_4),
	.A2(n18320),
	.B(n19917));
   NAND2xp33_ASAP7_75t_SRAM U22172 (.Y(n16756),
	.A(n16752),
	.B(n16753));
   NAND2xp33_ASAP7_75t_L U22175 (.Y(n16822),
	.A(n16821),
	.B(n16820));
   NOR3xp33_ASAP7_75t_L U22176 (.Y(n16823),
	.A(n16816),
	.B(n20334),
	.C(n17857));
   NAND2xp33_ASAP7_75t_R U22177 (.Y(n16820),
	.A(n16819),
	.B(n23662));
   NAND3xp33_ASAP7_75t_SL U22178 (.Y(n16825),
	.A(n16805),
	.B(n16804),
	.C(n22339));
   O2A1O1Ixp33_ASAP7_75t_L U22179 (.Y(n16805),
	.A1(n16808),
	.A2(FE_OFN29023_n16750),
	.B(FE_OFN28778_FE_OCPN28352_n16748),
	.C(n24254));
   NAND2xp5_ASAP7_75t_L U22180 (.Y(n16804),
	.A(n16797),
	.B(n16796));
   NAND2xp5_ASAP7_75t_R U22181 (.Y(n16797),
	.A(n16794),
	.B(n16795));
   NAND3xp33_ASAP7_75t_SL U22182 (.Y(n16787),
	.A(n16782),
	.B(n23656),
	.C(n23654));
   NAND3xp33_ASAP7_75t_SRAM U22183 (.Y(n16788),
	.A(n20332),
	.B(n20009),
	.C(n23668));
   NAND2xp5_ASAP7_75t_L U22185 (.Y(n17887),
	.A(FE_OCPN29265_FE_OFN28698_sa21_1),
	.B(n17886));
   NOR2xp33_ASAP7_75t_SL U22186 (.Y(n17888),
	.A(n25589),
	.B(n17883));
   NAND2xp33_ASAP7_75t_L U22187 (.Y(n17886),
	.A(n17885),
	.B(n17884));
   NAND3xp33_ASAP7_75t_SL U22188 (.Y(n17890),
	.A(n17884),
	.B(n17859),
	.C(n24281));
   NAND3xp33_ASAP7_75t_R U22190 (.Y(n17891),
	.A(n17853),
	.B(n17852),
	.C(n17851));
   NAND2xp33_ASAP7_75t_R U22191 (.Y(n17851),
	.A(n17850),
	.B(n17849));
   NAND2xp5_ASAP7_75t_L U22192 (.Y(n22335),
	.A(n17841),
	.B(n20299));
   NAND2xp33_ASAP7_75t_R U22193 (.Y(n17837),
	.A(n17834),
	.B(n20323));
   NAND2xp33_ASAP7_75t_SRAM U22194 (.Y(n17836),
	.A(n17835),
	.B(n20323));
   NAND2x1p5_ASAP7_75t_L U22195 (.Y(n20011),
	.A(n16791),
	.B(FE_OCPN27774_n25351));
   NAND2xp5_ASAP7_75t_SL U22197 (.Y(n25581),
	.A(n22669),
	.B(n22340));
   NAND2xp5_ASAP7_75t_R U22198 (.Y(n25579),
	.A(n20312),
	.B(n19973));
   NAND3xp33_ASAP7_75t_L U22199 (.Y(n25582),
	.A(n20002),
	.B(n22657),
	.C(n22670));
   NAND2xp5_ASAP7_75t_R U22200 (.Y(n24279),
	.A(n20326),
	.B(n20299));
   NOR3x1_ASAP7_75t_SL U22201 (.Y(n22339),
	.A(n16803),
	.B(FE_OCPN5079_n20287),
	.C(n23651));
   NAND3xp33_ASAP7_75t_SL U22202 (.Y(n16803),
	.A(n22354),
	.B(n19867),
	.C(n20003));
   NAND3xp33_ASAP7_75t_L U22203 (.Y(n22359),
	.A(n22358),
	.B(n22357),
	.C(n22356));
   NOR2xp33_ASAP7_75t_L U22204 (.Y(n22358),
	.A(n22349),
	.B(n25579));
   NOR3xp33_ASAP7_75t_R U22205 (.Y(n22357),
	.A(n23658),
	.B(n23652),
	.C(n22355));
   NOR3xp33_ASAP7_75t_SL U22207 (.Y(n22347),
	.A(n22345),
	.B(n22344),
	.C(n25577));
   NAND2xp33_ASAP7_75t_R U22208 (.Y(n22345),
	.A(n23654),
	.B(n22343));
   NOR2xp67_ASAP7_75t_SL U22209 (.Y(n22363),
	.A(n20314),
	.B(n20313));
   NAND3xp33_ASAP7_75t_SL U22210 (.Y(n20313),
	.A(n22661),
	.B(n20312),
	.C(n20311));
   NAND2xp5_ASAP7_75t_SL U22211 (.Y(n20311),
	.A(n20310),
	.B(n20309));
   NAND2xp33_ASAP7_75t_SL U22212 (.Y(n20309),
	.A(n20308),
	.B(n20307));
   NAND2xp5_ASAP7_75t_L U22213 (.Y(n23638),
	.A(n22340),
	.B(n22667));
   NAND3xp33_ASAP7_75t_SL U22214 (.Y(n22692),
	.A(n22356),
	.B(n19895),
	.C(n19894));
   NOR3xp33_ASAP7_75t_SL U22215 (.Y(n19895),
	.A(n19893),
	.B(n19892),
	.C(FE_OFN27179_n20327));
   NAND2xp33_ASAP7_75t_SRAM U22216 (.Y(n22334),
	.A(n22346),
	.B(n22333));
   NAND2xp5_ASAP7_75t_L U22217 (.Y(n24278),
	.A(n20315),
	.B(n22340));
   NOR2x1p5_ASAP7_75t_SL U22218 (.Y(n22330),
	.A(FE_OFN28823_n17860),
	.B(FE_OFN28820_n));
   NAND2xp5_ASAP7_75t_L U22220 (.Y(n23666),
	.A(n23665),
	.B(n23664));
   NOR3x1_ASAP7_75t_L U22221 (.Y(n23667),
	.A(n23659),
	.B(n23658),
	.C(n23657));
   NAND2xp33_ASAP7_75t_SRAM U22222 (.Y(n23664),
	.A(n23663),
	.B(n23662));
   NAND3xp33_ASAP7_75t_L U22223 (.Y(n23670),
	.A(n23655),
	.B(n23656),
	.C(n23654));
   NAND3xp33_ASAP7_75t_L U22224 (.Y(n23671),
	.A(n22687),
	.B(n22686),
	.C(n22685));
   NAND2xp33_ASAP7_75t_L U22225 (.Y(n22685),
	.A(n22684),
	.B(n22683));
   NAND2xp33_ASAP7_75t_L U22226 (.Y(n23648),
	.A(n23642),
	.B(n23645));
   NAND2xp5_ASAP7_75t_L U22227 (.Y(n24843),
	.A(n25007),
	.B(n24841));
   NAND2xp33_ASAP7_75t_L U22228 (.Y(n24833),
	.A(n26836),
	.B(FE_OFN26058_w3_1));
   NAND3xp33_ASAP7_75t_SL U22229 (.Y(n21995),
	.A(n21994),
	.B(n21993),
	.C(n21992));
   OAI22xp33_ASAP7_75t_SRAM U22230 (.Y(n21994),
	.A1(n21989),
	.A2(n21988),
	.B1(n21987),
	.B2(n21988));
   NOR3xp33_ASAP7_75t_SL U22231 (.Y(n21993),
	.A(n24180),
	.B(n21991),
	.C(n21990));
   NOR3xp33_ASAP7_75t_L U22233 (.Y(n21985),
	.A(n21983),
	.B(n21982),
	.C(n27072));
   OAI21xp33_ASAP7_75t_R U22234 (.Y(n21983),
	.A1(FE_OCPN7597_n21981),
	.A2(FE_OFN29117_n),
	.B(n21979));
   NOR3xp33_ASAP7_75t_SL U22236 (.Y(n21963),
	.A(n21939),
	.B(FE_OFN28719_n20025),
	.C(n21980));
   NAND2xp5_ASAP7_75t_SL U22237 (.Y(n21962),
	.A(n21932),
	.B(n16335));
   NOR2x1_ASAP7_75t_L U22239 (.Y(n21968),
	.A(n20074),
	.B(FE_OCPN28334_n16497));
   NOR2x1_ASAP7_75t_L U22240 (.Y(n21922),
	.A(FE_OCPN27697_n16309),
	.B(n21980));
   NOR3xp33_ASAP7_75t_SL U22241 (.Y(n21921),
	.A(n16497),
	.B(FE_OCPN29482_FE_OFN26014_sa31_3),
	.C(n16340));
   NAND2xp5_ASAP7_75t_SL U22242 (.Y(n25325),
	.A(n21925),
	.B(n21924));
   NAND3xp33_ASAP7_75t_SL U22243 (.Y(n21930),
	.A(n20875),
	.B(n20874),
	.C(n20873));
   NAND2xp5_ASAP7_75t_SL U22244 (.Y(n20875),
	.A(n20872),
	.B(n20871));
   NAND2xp33_ASAP7_75t_SL U22245 (.Y(n20871),
	.A(n20870),
	.B(FE_OFN26569_n20866));
   NAND2xp33_ASAP7_75t_L U22246 (.Y(n20872),
	.A(n20867),
	.B(FE_OFN26569_n20866));
   NAND2xp33_ASAP7_75t_L U22247 (.Y(n21929),
	.A(n16406),
	.B(n18069));
   NOR3xp33_ASAP7_75t_SL U22248 (.Y(n21953),
	.A(n21943),
	.B(n21942),
	.C(n21941));
   OAI21xp33_ASAP7_75t_SRAM U22249 (.Y(n21941),
	.A1(n21940),
	.A2(n21939),
	.B(n21938));
   NAND2x1_ASAP7_75t_SL U22251 (.Y(n20890),
	.A(n20889),
	.B(n20888));
   NAND2xp5_ASAP7_75t_SL U22252 (.Y(n20888),
	.A(n20887),
	.B(n20884));
   NAND2xp5_ASAP7_75t_SL U22253 (.Y(n20889),
	.A(n20885),
	.B(n20884));
   NAND3xp33_ASAP7_75t_L U22254 (.Y(n20892),
	.A(n20865),
	.B(n20864),
	.C(n20863));
   NAND2xp5_ASAP7_75t_L U22255 (.Y(n20864),
	.A(n20862),
	.B(n20861));
   NAND2xp33_ASAP7_75t_L U22256 (.Y(n20861),
	.A(n20860),
	.B(n20859));
   NAND2xp33_ASAP7_75t_L U22257 (.Y(n20862),
	.A(n20857),
	.B(n20859));
   NAND2xp33_ASAP7_75t_L U22258 (.Y(n26297),
	.A(n16346),
	.B(n16385));
   NOR3xp33_ASAP7_75t_L U22259 (.Y(n16346),
	.A(n16361),
	.B(n18072),
	.C(n16372));
   NAND2xp33_ASAP7_75t_SRAM U22260 (.Y(n20848),
	.A(n20847),
	.B(n21932));
   NAND3xp33_ASAP7_75t_SL U22261 (.Y(n20893),
	.A(n16513),
	.B(n20034),
	.C(n16359));
   NAND3xp33_ASAP7_75t_SL U22262 (.Y(n20851),
	.A(n16407),
	.B(n20052),
	.C(n16311));
   NOR3xp33_ASAP7_75t_SL U22263 (.Y(n16311),
	.A(n16310),
	.B(n25848),
	.C(n18085));
   NAND2xp33_ASAP7_75t_L U22264 (.Y(n21974),
	.A(n20836),
	.B(n20835));
   NOR3xp33_ASAP7_75t_SL U22265 (.Y(n25849),
	.A(n16321),
	.B(FE_OFN28669_sa31_5),
	.C(n20854));
   NOR3x1_ASAP7_75t_SL U22267 (.Y(n26006),
	.A(n20047),
	.B(FE_OFN26550_n16331),
	.C(n20070));
   NAND3xp33_ASAP7_75t_R U22268 (.Y(n26008),
	.A(n20849),
	.B(n18082),
	.C(n16396));
   NOR3x1_ASAP7_75t_L U22269 (.Y(n26007),
	.A(n16297),
	.B(n21977),
	.C(n21962));
   NAND2xp33_ASAP7_75t_L U22270 (.Y(n16297),
	.A(n25322),
	.B(n26399));
   NAND3xp33_ASAP7_75t_L U22272 (.Y(n26303),
	.A(n18078),
	.B(n16339),
	.C(n16338));
   NAND3xp33_ASAP7_75t_SL U22273 (.Y(n26304),
	.A(n16333),
	.B(n16332),
	.C(n16503));
   NOR3xp33_ASAP7_75t_L U22274 (.Y(n16333),
	.A(n25318),
	.B(n20059),
	.C(n18062));
   NOR3xp33_ASAP7_75t_SL U22275 (.Y(n16332),
	.A(n16328),
	.B(n20876),
	.C(n20850));
   OAI21xp5_ASAP7_75t_SL U22276 (.Y(n25825),
	.A1(n25823),
	.A2(n27168),
	.B(n25822));
   NAND2xp33_ASAP7_75t_SRAM U22277 (.Y(n25821),
	.A(n25816),
	.B(n25815));
   A2O1A1Ixp33_ASAP7_75t_SL U22278 (.Y(n24598),
	.A1(FE_OFN16169_n26567),
	.A2(n24812),
	.B(n24596),
	.C(n24595));
   NAND2xp33_ASAP7_75t_SL U22279 (.Y(n24596),
	.A(FE_OFN27169_n26683),
	.B(n24608));
   O2A1O1Ixp33_ASAP7_75t_SL U22281 (.Y(n25770),
	.A1(FE_OCPN28346_n24051),
	.A2(n24050),
	.B(n26139),
	.C(n24049));
   NAND2xp33_ASAP7_75t_SRAM U22283 (.Y(n24060),
	.A(n24059),
	.B(n24058));
   NOR3xp33_ASAP7_75t_L U22284 (.Y(n24061),
	.A(n24053),
	.B(n24052),
	.C(n24381));
   A2O1A1Ixp33_ASAP7_75t_L U22285 (.Y(n24069),
	.A1(n26679),
	.A2(n26678),
	.B(n24067),
	.C(n24066));
   NAND2xp5_ASAP7_75t_L U22286 (.Y(n24067),
	.A(n26673),
	.B(n24073));
   NOR2x1_ASAP7_75t_L U22287 (.Y(n24034),
	.A(n25494),
	.B(FE_OCPN27753_n26685));
   NAND2x1p5_ASAP7_75t_L U22288 (.Y(n22661),
	.A(FE_OCPN27631_n16774),
	.B(n16757));
   NAND3x1_ASAP7_75t_SL U22289 (.Y(n22663),
	.A(n16783),
	.B(FE_OFN25989_sa21_4),
	.C(FE_OFN28678_sa21_3));
   NAND3xp33_ASAP7_75t_L U22290 (.Y(n24254),
	.A(n20312),
	.B(n23625),
	.C(n20315));
   NAND2x1_ASAP7_75t_SL U22291 (.Y(n22662),
	.A(FE_OCPN27328_sa21_2),
	.B(n16747));
   NAND2xp5_ASAP7_75t_R U22292 (.Y(n26817),
	.A(FE_OFN16271_n26814),
	.B(n26838));
   OAI222xp33_ASAP7_75t_L U22293 (.Y(n25494),
	.A1(n24032),
	.A2(n26687),
	.B1(n24031),
	.B2(n26687),
	.C1(n24030),
	.C2(n26687));
   NAND2xp33_ASAP7_75t_SRAM U22294 (.Y(n24017),
	.A(n24013),
	.B(sa21_7_));
   NAND2xp33_ASAP7_75t_L U22295 (.Y(n24016),
	.A(n24015),
	.B(sa21_7_));
   NAND2xp33_ASAP7_75t_R U22296 (.Y(n24656),
	.A(n24903),
	.B(FE_OFN7_w3_22));
   NAND3xp33_ASAP7_75t_SRAM U22297 (.Y(n24649),
	.A(FE_OFN28533_n24995),
	.B(n24648),
	.C(FE_OCPN7596_n24647));
   A2O1A1Ixp33_ASAP7_75t_R U22298 (.Y(n25508),
	.A1(n26407),
	.A2(n25510),
	.B(FE_OCPN29444_n25507),
	.C(FE_OCPN27770_n26049));
   O2A1O1Ixp5_ASAP7_75t_SL U22299 (.Y(n24877),
	.A1(n24875),
	.A2(n24874),
	.B(n25367),
	.C(n25363));
   NAND2xp33_ASAP7_75t_SRAM U22300 (.Y(n24873),
	.A(n24860),
	.B(n24859));
   NAND3x1_ASAP7_75t_SL U22301 (.Y(n24891),
	.A(n16812),
	.B(n16811),
	.C(n16810));
   NAND2xp33_ASAP7_75t_SRAM U22302 (.Y(n16811),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(FE_OFN29023_n16750));
   NOR3x1_ASAP7_75t_SL U22303 (.Y(n16812),
	.A(n17854),
	.B(n20314),
	.C(n16809));
   NAND2xp33_ASAP7_75t_SRAM U22305 (.Y(n27046),
	.A(n27038),
	.B(FE_OFN163_sa00_7));
   NAND2xp33_ASAP7_75t_SRAM U22306 (.Y(n27045),
	.A(n27044),
	.B(FE_OFN163_sa00_7));
   NAND2xp33_ASAP7_75t_L U22307 (.Y(n27051),
	.A(FE_OFN29224_FE_OCPN28074_n27049),
	.B(FE_OFN133_n24306));
   A2O1A1Ixp33_ASAP7_75t_SL U22308 (.Y(n27050),
	.A1(n27117),
	.A2(n27052),
	.B(FE_OFN29142_n27049),
	.C(n24306));
   O2A1O1Ixp5_ASAP7_75t_SL U22310 (.Y(n25193),
	.A1(n25191),
	.A2(n25190),
	.B(n27207),
	.C(n25832));
   NAND3xp33_ASAP7_75t_SRAM U22311 (.Y(n25190),
	.A(n25189),
	.B(FE_OFN29096_n25188),
	.C(FE_OCPN28366_n25329));
   NAND2xp33_ASAP7_75t_L U22312 (.Y(n25836),
	.A(n25833),
	.B(n25841));
   NOR2x1_ASAP7_75t_SL U22313 (.Y(n25565),
	.A(n25564),
	.B(n25563));
   NAND2xp33_ASAP7_75t_L U22315 (.Y(n27075),
	.A(sa31_7_),
	.B(FE_OFN25970_n));
   NAND2xp33_ASAP7_75t_R U22317 (.Y(n25404),
	.A(n25396),
	.B(FE_OFN175_sa12_6));
   NOR2xp33_ASAP7_75t_SRAM U22318 (.Y(n25396),
	.A(n25395),
	.B(FE_OFN165_sa12_7));
   NAND2x1_ASAP7_75t_SL U22320 (.Y(n24324),
	.A(n16952),
	.B(n18133));
   NAND2xp5_ASAP7_75t_SL U22321 (.Y(n24326),
	.A(n16851),
	.B(FE_OFN28995_n16850));
   NAND3xp33_ASAP7_75t_SL U22322 (.Y(n24325),
	.A(n18120),
	.B(n16869),
	.C(n16868));
   NOR2xp33_ASAP7_75t_L U22323 (.Y(n16869),
	.A(n16882),
	.B(n17415));
   NOR3x1_ASAP7_75t_SL U22324 (.Y(n24328),
	.A(n16874),
	.B(FE_OFN29164_sa33_2),
	.C(FE_OCPN27539_n16875));
   NOR2xp33_ASAP7_75t_SRAM U22325 (.Y(n24327),
	.A(FE_OFN29164_sa33_2),
	.B(FE_OFN25960_n));
   O2A1O1Ixp5_ASAP7_75t_SL U22326 (.Y(n24480),
	.A1(FE_OFN28553_n25599),
	.A2(n24477),
	.B(FE_OFN16170_n26637),
	.C(n26535));
   NAND2xp33_ASAP7_75t_R U22328 (.Y(n26670),
	.A(n26668),
	.B(n26667));
   NAND2xp33_ASAP7_75t_SRAM U22329 (.Y(n26667),
	.A(n26666),
	.B(n26665));
   NAND2xp33_ASAP7_75t_SRAM U22330 (.Y(n26668),
	.A(n26662),
	.B(n26665));
   NAND2xp5_ASAP7_75t_SL U22332 (.Y(n26677),
	.A(n26673),
	.B(FE_OFN86_n26674));
   NAND2xp5_ASAP7_75t_SL U22334 (.Y(n26530),
	.A(FE_OCPN29390_n26528),
	.B(FE_OFN25927_n26527));
   A2O1A1Ixp33_ASAP7_75t_SL U22335 (.Y(n14084),
	.A1(n14082),
	.A2(n14081),
	.B(n15704),
	.C(n14080));
   NAND2xp33_ASAP7_75t_L U22336 (.Y(n14081),
	.A(n14040),
	.B(n14039));
   NAND3xp33_ASAP7_75t_L U22338 (.Y(n14087),
	.A(n14028),
	.B(n14027),
	.C(n14026));
   OAI22xp33_ASAP7_75t_SRAM U22339 (.Y(n14026),
	.A1(FE_OFN16426_w3_20),
	.A2(n14025),
	.B1(n14369),
	.B2(n14025));
   NAND2xp33_ASAP7_75t_L U22340 (.Y(n14027),
	.A(n14024),
	.B(n14023));
   O2A1O1Ixp5_ASAP7_75t_SL U22342 (.Y(n15770),
	.A1(n15259),
	.A2(n14605),
	.B(n14604),
	.C(n14603));
   A2O1A1Ixp33_ASAP7_75t_SL U22344 (.Y(n14245),
	.A1(n14243),
	.A2(n14242),
	.B(FE_OFN28682_n15888),
	.C(n14241));
   NAND2xp33_ASAP7_75t_L U22345 (.Y(n14243),
	.A(n14201),
	.B(n14200));
   NAND2xp33_ASAP7_75t_L U22346 (.Y(n14242),
	.A(n14208),
	.B(n14207));
   O2A1O1Ixp5_ASAP7_75t_SL U22347 (.Y(n13861),
	.A1(n13860),
	.A2(n13859),
	.B(n16042),
	.C(n13858));
   OAI21xp33_ASAP7_75t_SRAM U22348 (.Y(n13860),
	.A1(n13815),
	.A2(FE_OFN28856_n15450),
	.B(n14640));
   A2O1A1Ixp33_ASAP7_75t_L U22349 (.Y(n13858),
	.A1(n13857),
	.A2(n13856),
	.B(n15969),
	.C(n13855));
   OAI21xp33_ASAP7_75t_L U22350 (.Y(n13859),
	.A1(n14959),
	.A2(n16016),
	.B(n13825));
   NAND2xp33_ASAP7_75t_L U22351 (.Y(n13813),
	.A(n13810),
	.B(n13809));
   NAND2xp33_ASAP7_75t_R U22352 (.Y(n13809),
	.A(n13808),
	.B(n13807));
   NOR3xp33_ASAP7_75t_SRAM U22353 (.Y(n13811),
	.A(FE_OFN26007_n16010),
	.B(FE_OFN26003_n15992),
	.C(n14695));
   NAND3xp33_ASAP7_75t_SRAM U22354 (.Y(n13803),
	.A(n13802),
	.B(n13801),
	.C(n13800));
   INVxp67_ASAP7_75t_SL U22355 (.Y(n13862),
	.A(n13861));
   NAND2xp5_ASAP7_75t_SL U22357 (.Y(n14178),
	.A(n14177),
	.B(n14176));
   NAND2xp33_ASAP7_75t_SL U22358 (.Y(n14177),
	.A(n14172),
	.B(n14174));
   NAND2xp5_ASAP7_75t_L U22359 (.Y(n14176),
	.A(n14175),
	.B(n14174));
   NOR2xp33_ASAP7_75t_L U22360 (.Y(n14172),
	.A(n14157),
	.B(n14173));
   NAND2xp5_ASAP7_75t_L U22361 (.Y(n14110),
	.A(n14106),
	.B(n14105));
   NAND2xp33_ASAP7_75t_L U22362 (.Y(n14105),
	.A(n14104),
	.B(n14103));
   NAND2xp5_ASAP7_75t_R U22363 (.Y(n14106),
	.A(n14101),
	.B(n14103));
   NOR2xp33_ASAP7_75t_SRAM U22364 (.Y(n14104),
	.A(FE_OCPN29520_n24755),
	.B(n14102));
   NAND2xp33_ASAP7_75t_SRAM U22365 (.Y(n14111),
	.A(n14097),
	.B(n14096));
   NAND2xp33_ASAP7_75t_SRAM U22366 (.Y(n14096),
	.A(n14095),
	.B(n14094));
   NAND2xp33_ASAP7_75t_SRAM U22367 (.Y(n14097),
	.A(n14093),
	.B(n14094));
   NAND2xp33_ASAP7_75t_SRAM U22368 (.Y(n14108),
	.A(n14907),
	.B(n14107));
   NAND2xp33_ASAP7_75t_SRAM U22369 (.Y(n14107),
	.A(n14912),
	.B(n14919));
   OAI222xp33_ASAP7_75t_R U22372 (.Y(n14817),
	.A1(FE_PSN8276_FE_OFN28712_n),
	.A2(n14768),
	.B1(n14767),
	.B2(n14768),
	.C1(FE_OFN28628_n15667),
	.C2(n14768));
   NAND2xp5_ASAP7_75t_SL U22373 (.Y(n14816),
	.A(n14788),
	.B(n14787));
   NOR3xp33_ASAP7_75t_L U22374 (.Y(n14763),
	.A(n14762),
	.B(n15281),
	.C(n15682));
   NAND3xp33_ASAP7_75t_R U22375 (.Y(n14762),
	.A(n14761),
	.B(n14760),
	.C(n14759));
   O2A1O1Ixp33_ASAP7_75t_SL U22376 (.Y(n13329),
	.A1(n13287),
	.A2(n13328),
	.B(n15271),
	.C(n13327));
   OAI21xp33_ASAP7_75t_R U22377 (.Y(n13328),
	.A1(FE_OFN26104_n13659),
	.A2(n13428),
	.B(n13299));
   A2O1A1Ixp33_ASAP7_75t_L U22378 (.Y(n13327),
	.A1(n13326),
	.A2(n13325),
	.B(n13689),
	.C(n13324));
   NAND2xp5_ASAP7_75t_SL U22379 (.Y(n13285),
	.A(n13284),
	.B(n13283));
   NAND2xp33_ASAP7_75t_L U22380 (.Y(n13284),
	.A(n13279),
	.B(n13281));
   NAND2xp33_ASAP7_75t_L U22381 (.Y(n13283),
	.A(n13282),
	.B(n13281));
   NOR2xp33_ASAP7_75t_SRAM U22382 (.Y(n13279),
	.A(n14515),
	.B(n13280));
   INVxp33_ASAP7_75t_L U22383 (.Y(n14491),
	.A(n13650));
   NAND2xp5_ASAP7_75t_SL U22385 (.Y(n13793),
	.A(n13765),
	.B(n13764));
   NAND3xp33_ASAP7_75t_R U22386 (.Y(n13790),
	.A(n13774),
	.B(n13773),
	.C(n14872));
   A2O1A1Ixp33_ASAP7_75t_SL U22387 (.Y(n13933),
	.A1(n13931),
	.A2(n13930),
	.B(n13901),
	.C(n13929));
   NAND2xp33_ASAP7_75t_R U22388 (.Y(n13930),
	.A(n13900),
	.B(n13899));
   NOR3xp33_ASAP7_75t_SRAM U22389 (.Y(n13931),
	.A(n13894),
	.B(n15507),
	.C(n13893));
   OAI21xp5_ASAP7_75t_SL U22390 (.Y(n13936),
	.A1(n13888),
	.A2(FE_OFN27074_n13868),
	.B(n13887));
   OAI22xp33_ASAP7_75t_SRAM U22391 (.Y(n13888),
	.A1(FE_OFN5_w3_22),
	.A2(n15341),
	.B1(FE_OFN28623_n13874),
	.B2(n15341));
   NAND2xp5_ASAP7_75t_L U22392 (.Y(n13887),
	.A(n13886),
	.B(n13885));
   NAND2xp33_ASAP7_75t_R U22393 (.Y(n13885),
	.A(n13884),
	.B(n13883));
   INVxp67_ASAP7_75t_SL U22394 (.Y(n13932),
	.A(n13933));
   NAND2xp33_ASAP7_75t_L U22395 (.Y(n14620),
	.A(n14619),
	.B(n14618));
   NAND2xp33_ASAP7_75t_L U22396 (.Y(n14619),
	.A(n14613),
	.B(n14616));
   NOR2xp33_ASAP7_75t_SRAM U22397 (.Y(n14613),
	.A(FE_OFN29017_n15921),
	.B(n14614));
   NAND2xp33_ASAP7_75t_SRAM U22398 (.Y(n14608),
	.A(n15934),
	.B(n14607));
   A2O1A1Ixp33_ASAP7_75t_SL U22399 (.Y(n14658),
	.A1(n14656),
	.A2(n14655),
	.B(n16023),
	.C(n14654));
   O2A1O1Ixp33_ASAP7_75t_SRAM U22400 (.Y(n14655),
	.A1(n14940),
	.A2(n14626),
	.B(FE_OCPN28407_FE_OFN16433_w3_11),
	.C(n14625));
   O2A1O1Ixp5_ASAP7_75t_L U22401 (.Y(n14654),
	.A1(n14716),
	.A2(n14653),
	.B(n14971),
	.C(n14652));
   A2O1A1Ixp33_ASAP7_75t_SL U22402 (.Y(n15360),
	.A1(n15358),
	.A2(n15357),
	.B(n13901),
	.C(n15356));
   NAND2xp33_ASAP7_75t_R U22403 (.Y(n15357),
	.A(n15318),
	.B(n15317));
   NAND2xp33_ASAP7_75t_L U22404 (.Y(n15358),
	.A(n15311),
	.B(n15310));
   NAND3xp33_ASAP7_75t_SL U22405 (.Y(n15363),
	.A(n15293),
	.B(n15292),
	.C(n15291));
   OAI22xp33_ASAP7_75t_SRAM U22406 (.Y(n15291),
	.A1(n15290),
	.A2(n15661),
	.B1(n15744),
	.B2(n15661));
   NAND2xp33_ASAP7_75t_SRAM U22407 (.Y(n15293),
	.A(n15279),
	.B(n15278));
   NAND2xp33_ASAP7_75t_L U22408 (.Y(n15292),
	.A(n15289),
	.B(n15288));
   INVxp67_ASAP7_75t_SL U22409 (.Y(n15359),
	.A(n15360));
   NAND3xp33_ASAP7_75t_SL U22410 (.Y(n13406),
	.A(n13404),
	.B(n13403),
	.C(n13402));
   NAND2xp33_ASAP7_75t_SL U22411 (.Y(n13404),
	.A(n13368),
	.B(n13367));
   NAND2xp33_ASAP7_75t_SL U22412 (.Y(n13402),
	.A(n13401),
	.B(n13400));
   A2O1A1Ixp33_ASAP7_75t_SL U22415 (.Y(n15052),
	.A1(n15051),
	.A2(n15050),
	.B(FE_OFN28682_n15888),
	.C(n15049));
   NAND3xp33_ASAP7_75t_SL U22416 (.Y(n15054),
	.A(n15018),
	.B(n15017),
	.C(n15016));
   NAND2xp33_ASAP7_75t_L U22417 (.Y(n14995),
	.A(n14984),
	.B(n14983));
   NAND2xp33_ASAP7_75t_R U22418 (.Y(n14983),
	.A(n14982),
	.B(n14981));
   NAND2xp33_ASAP7_75t_R U22419 (.Y(n14984),
	.A(n14979),
	.B(n14981));
   NAND2xp33_ASAP7_75t_L U22420 (.Y(n14994),
	.A(n14993),
	.B(n14992));
   NAND2xp33_ASAP7_75t_SRAM U22421 (.Y(n14992),
	.A(n14991),
	.B(n14990));
   NAND2xp33_ASAP7_75t_SRAM U22422 (.Y(n14993),
	.A(n14987),
	.B(n14990));
   NAND2xp5_ASAP7_75t_L U22424 (.Y(n15394),
	.A(n15393),
	.B(n15392));
   NAND2xp33_ASAP7_75t_L U22425 (.Y(n15392),
	.A(n15391),
	.B(n15390));
   NAND2xp33_ASAP7_75t_L U22426 (.Y(n15393),
	.A(n15388),
	.B(n15390));
   NOR2xp33_ASAP7_75t_SRAM U22427 (.Y(n15391),
	.A(n16000),
	.B(n15389));
   OAI21xp33_ASAP7_75t_SRAM U22428 (.Y(n15396),
	.A1(n15378),
	.A2(n15377),
	.B(n15956));
   NOR2xp33_ASAP7_75t_SRAM U22429 (.Y(n15378),
	.A(n15374),
	.B(FE_OFN26007_n16010));
   NAND2xp33_ASAP7_75t_L U22430 (.Y(n15463),
	.A(n15421),
	.B(n15420));
   NAND2xp33_ASAP7_75t_L U22431 (.Y(n15464),
	.A(n15406),
	.B(n15405));
   NAND2xp5_ASAP7_75t_L U22433 (.Y(n14262),
	.A(n14261),
	.B(n14260));
   NAND2xp33_ASAP7_75t_SRAM U22434 (.Y(n14261),
	.A(n14253),
	.B(n15349));
   NAND3xp33_ASAP7_75t_SL U22435 (.Y(n14323),
	.A(n14322),
	.B(n14321),
	.C(n14320));
   NAND2xp33_ASAP7_75t_SL U22436 (.Y(n14322),
	.A(n14275),
	.B(n14274));
   A2O1A1Ixp33_ASAP7_75t_L U22437 (.Y(n14321),
	.A1(FE_OFN27066_n13869),
	.A2(n15527),
	.B(n14285),
	.C(n15757));
   NAND2xp5_ASAP7_75t_SL U22438 (.Y(n15652),
	.A(n15651),
	.B(n15650));
   NAND2xp5_ASAP7_75t_L U22439 (.Y(n15650),
	.A(n15649),
	.B(n15648));
   INVx1_ASAP7_75t_SL U22440 (.Y(n15648),
	.A(n15623));
   NOR3xp33_ASAP7_75t_R U22441 (.Y(n15584),
	.A(n15574),
	.B(n15573),
	.C(n15572));
   NOR2xp33_ASAP7_75t_SRAM U22442 (.Y(n15572),
	.A(n15571),
	.B(n15570));
   NOR2xp33_ASAP7_75t_SRAM U22443 (.Y(n15573),
	.A(n15568),
	.B(n15813));
   NAND2xp33_ASAP7_75t_SRAM U22444 (.Y(n15583),
	.A(n15582),
	.B(n15581));
   NAND2xp33_ASAP7_75t_SRAM U22445 (.Y(n15581),
	.A(n15580),
	.B(n15579));
   NAND2xp33_ASAP7_75t_SRAM U22446 (.Y(n15582),
	.A(n15576),
	.B(n15579));
   NAND2xp5_ASAP7_75t_L U22448 (.Y(n15557),
	.A(n15556),
	.B(n15555));
   NAND2xp33_ASAP7_75t_SL U22449 (.Y(n15558),
	.A(n15533),
	.B(n15555));
   NOR2xp33_ASAP7_75t_SL U22450 (.Y(n15556),
	.A(n15554),
	.B(n15553));
   NOR3xp33_ASAP7_75t_L U22451 (.Y(n15563),
	.A(n15490),
	.B(n15489),
	.C(n15488));
   NOR2xp33_ASAP7_75t_SRAM U22452 (.Y(n15488),
	.A(n15487),
	.B(n15486));
   NAND3xp33_ASAP7_75t_L U22453 (.Y(n15490),
	.A(n15483),
	.B(n15482),
	.C(n15481));
   OAI22xp33_ASAP7_75t_L U22455 (.Y(n15091),
	.A1(n15780),
	.A2(n15078),
	.B1(n15834),
	.B2(n15078));
   O2A1O1Ixp33_ASAP7_75t_SL U22456 (.Y(n15072),
	.A1(n15835),
	.A2(n15577),
	.B(n15635),
	.C(n15071));
   OAI21xp33_ASAP7_75t_L U22457 (.Y(n15071),
	.A1(n13725),
	.A2(n15070),
	.B(n15069));
   NAND2xp33_ASAP7_75t_R U22458 (.Y(n15069),
	.A(n15068),
	.B(n15067));
   INVxp33_ASAP7_75t_SRAM U22459 (.Y(n15070),
	.A(n15589));
   NOR2x1_ASAP7_75t_L U22461 (.Y(n16042),
	.A(w3_10_),
	.B(FE_OFN25961_w3_8));
   O2A1O1Ixp5_ASAP7_75t_SL U22462 (.Y(n14738),
	.A1(n14737),
	.A2(n14736),
	.B(n14971),
	.C(n14735));
   NAND3xp33_ASAP7_75t_SL U22463 (.Y(n14736),
	.A(n14693),
	.B(n14692),
	.C(n14691));
   A2O1A1Ixp33_ASAP7_75t_SL U22464 (.Y(n14735),
	.A1(n14734),
	.A2(n14733),
	.B(n16023),
	.C(n14732));
   NAND2xp33_ASAP7_75t_R U22465 (.Y(n14678),
	.A(n14676),
	.B(n14675));
   NAND2xp33_ASAP7_75t_R U22466 (.Y(n14675),
	.A(n14674),
	.B(n14673));
   NAND2xp33_ASAP7_75t_R U22467 (.Y(n14676),
	.A(n14671),
	.B(n14673));
   O2A1O1Ixp5_ASAP7_75t_SRAM U22468 (.Y(n14679),
	.A1(n13804),
	.A2(n14667),
	.B(FE_OFN29017_n15921),
	.C(n14666));
   INVxp67_ASAP7_75t_SL U22469 (.Y(n14739),
	.A(n14738));
   NAND2xp5_ASAP7_75t_L U22470 (.Y(n15767),
	.A(n15678),
	.B(n15677));
   NAND2xp33_ASAP7_75t_L U22471 (.Y(n15678),
	.A(n15672),
	.B(n15675));
   NAND2xp33_ASAP7_75t_L U22472 (.Y(n15677),
	.A(n15676),
	.B(n15675));
   NOR2xp33_ASAP7_75t_SRAM U22473 (.Y(n15672),
	.A(n15664),
	.B(n15673));
   A2O1A1Ixp33_ASAP7_75t_SL U22474 (.Y(n15761),
	.A1(n15760),
	.A2(n15759),
	.B(n15758),
	.C(n15757));
   NAND2xp33_ASAP7_75t_SRAM U22475 (.Y(n15759),
	.A(n15480),
	.B(n15738));
   NAND2xp33_ASAP7_75t_R U22476 (.Y(n13719),
	.A(n13712),
	.B(n13711));
   NAND2xp33_ASAP7_75t_SRAM U22477 (.Y(n13711),
	.A(n14566),
	.B(n13710));
   NAND2xp33_ASAP7_75t_SRAM U22478 (.Y(n13712),
	.A(n13709),
	.B(n13710));
   NOR3xp33_ASAP7_75t_SRAM U22480 (.Y(n13716),
	.A(FE_OFN26104_n13659),
	.B(FE_OFN28603_n14534),
	.C(n15155));
   NOR2xp33_ASAP7_75t_SRAM U22481 (.Y(n13714),
	.A(FE_OCPN29571_n26355),
	.B(n13713));
   OAI21xp33_ASAP7_75t_SRAM U22482 (.Y(n13715),
	.A1(n15145),
	.A2(FE_OFN27209_w3_30),
	.B(FE_OFN28817_n));
   NAND2xp5_ASAP7_75t_SL U22483 (.Y(n13704),
	.A(n13698),
	.B(n13701));
   NOR2xp33_ASAP7_75t_SL U22484 (.Y(n13698),
	.A(n15246),
	.B(n13699));
   NAND2xp33_ASAP7_75t_SRAM U22485 (.Y(n13707),
	.A(n13645),
	.B(n13644));
   NAND2xp33_ASAP7_75t_SRAM U22486 (.Y(n13645),
	.A(n13641),
	.B(n13640));
   NAND2xp33_ASAP7_75t_SRAM U22487 (.Y(n13706),
	.A(n13654),
	.B(n13653));
   NAND2xp33_ASAP7_75t_SRAM U22488 (.Y(n13653),
	.A(n13652),
	.B(n13651));
   NAND2xp33_ASAP7_75t_SRAM U22489 (.Y(n13654),
	.A(n13709),
	.B(n13651));
   A2O1A1Ixp33_ASAP7_75t_L U22490 (.Y(n26795),
	.A1(FE_OCPN29586_n26857),
	.A2(n26793),
	.B(n26792),
	.C(n26791));
   A2O1A1Ixp33_ASAP7_75t_R U22491 (.Y(n26791),
	.A1(n26793),
	.A2(FE_OCPN29586_n26857),
	.B(n26787),
	.C(n26789));
   OAI21xp5_ASAP7_75t_L U22492 (.Y(n26794),
	.A1(FE_OFN28482_ld_r),
	.A2(FE_OCPN29381_n26796),
	.B(n26795));
   OAI21xp5_ASAP7_75t_SL U22493 (.Y(n25771),
	.A1(FE_OFN16213_ld_r),
	.A2(n26713),
	.B(n25772));
   A2O1A1Ixp33_ASAP7_75t_SL U22494 (.Y(n25772),
	.A1(FE_OCPN28023_n25770),
	.A2(FE_OCPN27815_n25769),
	.B(FE_OCPN27421_n25768),
	.C(n25767));
   NAND3xp33_ASAP7_75t_SL U22495 (.Y(n25767),
	.A(FE_OCPN27815_n25769),
	.B(FE_OCPN28023_n25770),
	.C(n25768));
   A2O1A1Ixp33_ASAP7_75t_SL U22496 (.Y(n26214),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(n26212),
	.C(n26211));
   NAND2xp5_ASAP7_75t_L U22497 (.Y(n26212),
	.A(FE_OFN25939_n26275),
	.B(n26210));
   A2O1A1Ixp33_ASAP7_75t_SL U22498 (.Y(n26211),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(FE_OFN27123_n26275),
	.C(w1_17_));
   OAI21xp5_ASAP7_75t_SL U22499 (.Y(n26432),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OCPN27525_n26434),
	.B(n26433));
   NOR2xp33_ASAP7_75t_R U22500 (.Y(n26430),
	.A(FE_OFN16265_n26527),
	.B(FE_OCPN28024_n26427));
   O2A1O1Ixp33_ASAP7_75t_L U22501 (.Y(n26429),
	.A1(FE_OFN16180_n26542),
	.A2(n26431),
	.B(FE_OCPN27637_n26428),
	.C(FE_OFN25927_n26527));
   OAI21xp5_ASAP7_75t_SL U22502 (.Y(n25779),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27787_n26728),
	.B(n25780));
   A2O1A1Ixp33_ASAP7_75t_SL U22503 (.Y(n25780),
	.A1(FE_OCPN27991_n26336),
	.A2(FE_OCPN28110_n),
	.B(n25778),
	.C(n25777));
   NAND3xp33_ASAP7_75t_SL U22504 (.Y(n25777),
	.A(FE_OCPN28110_n),
	.B(FE_OCPN27991_n26336),
	.C(n25778));
   A2O1A1Ixp33_ASAP7_75t_SRAM U22505 (.Y(n26284),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(n26280),
	.C(n26279));
   NAND2xp33_ASAP7_75t_SRAM U22506 (.Y(n26280),
	.A(FE_OFN28990_n26276),
	.B(FE_OFN25939_n26275));
   XNOR2xp5_ASAP7_75t_SL U22507 (.Y(n16206),
	.A(w2_30_),
	.B(n16197));
   FAx1_ASAP7_75t_SL U22508 (.SN(n25758),
	.A(n25756),
	.B(FE_OCPN27322_n25755),
	.CI(n25754));
   A2O1A1Ixp33_ASAP7_75t_SL U22509 (.Y(n25756),
	.A1(n26249),
	.A2(n25736),
	.B(n25735),
	.C(n25734));
   NAND2xp5_ASAP7_75t_L U22510 (.Y(n25735),
	.A(FE_OFN28904_n25733),
	.B(n25732));
   A2O1A1Ixp33_ASAP7_75t_SL U22511 (.Y(n24638),
	.A1(n24636),
	.A2(n24635),
	.B(n24719),
	.C(n24634));
   NAND3xp33_ASAP7_75t_SL U22512 (.Y(n24634),
	.A(n24635),
	.B(n24636),
	.C(n24719));
   O2A1O1Ixp33_ASAP7_75t_L U22513 (.Y(n24635),
	.A1(n24624),
	.A2(n24623),
	.B(n26770),
	.C(n24622));
   NAND2x1_ASAP7_75t_SL U22514 (.Y(n26391),
	.A(n26388),
	.B(n26764));
   A2O1A1Ixp33_ASAP7_75t_SL U22515 (.Y(n26261),
	.A1(n26139),
	.A2(n26138),
	.B(n25075),
	.C(n25074));
   NAND2xp5_ASAP7_75t_R U22516 (.Y(n25075),
	.A(n26134),
	.B(n25072));
   A2O1A1Ixp33_ASAP7_75t_L U22518 (.Y(n25014),
	.A1(n26857),
	.A2(n19640),
	.B(n25013),
	.C(n25012));
   NAND2xp33_ASAP7_75t_R U22519 (.Y(n25013),
	.A(FE_OCPN27664_w3_25),
	.B(n25010));
   OAI22xp33_ASAP7_75t_SRAM U22520 (.Y(n25015),
	.A1(text_in_r_25_),
	.A2(FE_OFN28490_ld_r),
	.B1(FE_OCPN27659_w3_25),
	.B2(FE_OFN28490_ld_r));
   NAND2xp33_ASAP7_75t_L U22522 (.Y(n26855),
	.A(n26852),
	.B(n26850));
   OAI21xp5_ASAP7_75t_SL U22523 (.Y(n26413),
	.A1(FE_OFN1_ld_r),
	.A2(FE_OCPN7625_n26501),
	.B(n26414));
   NAND2xp5_ASAP7_75t_SL U22524 (.Y(n26928),
	.A(n26927),
	.B(n26929));
   A2O1A1Ixp33_ASAP7_75t_SL U22526 (.Y(n26653),
	.A1(n26651),
	.A2(FE_OCPN29471_n24175),
	.B(n26649),
	.C(n26648));
   O2A1O1Ixp33_ASAP7_75t_SRAM U22527 (.Y(n26471),
	.A1(n27004),
	.A2(n26702),
	.B(n26469),
	.C(n26468));
   NOR2xp33_ASAP7_75t_SRAM U22528 (.Y(n26469),
	.A(n26466),
	.B(n26697));
   O2A1O1Ixp33_ASAP7_75t_SRAM U22529 (.Y(n26468),
	.A1(n27004),
	.A2(n26702),
	.B(n26699),
	.C(n26467));
   OAI22xp5_ASAP7_75t_SL U22530 (.Y(n16249),
	.A1(w2_16_),
	.A2(n16125),
	.B1(n16250),
	.B2(n16125));
   NAND3xp33_ASAP7_75t_SL U22531 (.Y(n26114),
	.A(FE_OFN28484_ld_r),
	.B(n26116),
	.C(n26784));
   A2O1A1Ixp33_ASAP7_75t_SL U22532 (.Y(n26844),
	.A1(n22405),
	.A2(FE_OCPN27940_n26842),
	.B(n26841),
	.C(n26840));
   NAND2xp5_ASAP7_75t_SL U22533 (.Y(n26841),
	.A(FE_OCPN27234_n26837),
	.B(n26836));
   A2O1A1Ixp33_ASAP7_75t_L U22534 (.Y(n26840),
	.A1(FE_OCPN27940_n26842),
	.A2(n22405),
	.B(n26839),
	.C(n26838));
   OAI21xp5_ASAP7_75t_SL U22535 (.Y(n24466),
	.A1(FE_OFN28482_ld_r),
	.A2(n24468),
	.B(n24467));
   NOR2xp33_ASAP7_75t_L U22536 (.Y(n27166),
	.A(n27178),
	.B(FE_OFN26650_n27164));
   O2A1O1Ixp5_ASAP7_75t_L U22537 (.Y(n27165),
	.A1(n27168),
	.A2(n27167),
	.B(n27163),
	.C(FE_OFN105_n27178));
   NOR2x1p5_ASAP7_75t_SL U22538 (.Y(n27209),
	.A(n25311),
	.B(FE_OCPN29287_n27210));
   NAND2xp33_ASAP7_75t_SL U22539 (.Y(n27205),
	.A(n27201),
	.B(n27200));
   NAND2xp33_ASAP7_75t_SRAM U22540 (.Y(n27214),
	.A(w2_18_),
	.B(n27211));
   NOR3xp33_ASAP7_75t_SL U22541 (.Y(n26233),
	.A(FE_OCPN27451_n26236),
	.B(n26234),
	.C(n26235));
   NOR3xp33_ASAP7_75t_L U22542 (.Y(n26266),
	.A(n26268),
	.B(n26638),
	.C(n26267));
   NOR3xp33_ASAP7_75t_SL U22543 (.Y(n26269),
	.A(n26270),
	.B(FE_OFN2_ld_r),
	.C(FE_OFN26024_n26115));
   NOR3xp33_ASAP7_75t_SL U22547 (.Y(n17710),
	.A(n17709),
	.B(n20102),
	.C(n19729));
   OAI222xp33_ASAP7_75t_SRAM U22548 (.Y(n17719),
	.A1(n17718),
	.A2(n26346),
	.B1(n20094),
	.B2(n26346),
	.C1(n17717),
	.C2(n26346));
   NAND3xp33_ASAP7_75t_R U22549 (.Y(n25368),
	.A(n24648),
	.B(n17688),
	.C(FE_OCPN7596_n24647));
   NOR2xp33_ASAP7_75t_SRAM U22550 (.Y(n17687),
	.A(n17560),
	.B(FE_OFN27138_n24012));
   NOR3xp33_ASAP7_75t_SRAM U22551 (.Y(n17053),
	.A(FE_OCPN7612_n25229),
	.B(n27186),
	.C(n17052));
   OAI222xp33_ASAP7_75t_SRAM U22552 (.Y(n17052),
	.A1(n25223),
	.A2(n26959),
	.B1(n17051),
	.B2(n26959),
	.C1(n17050),
	.C2(n26959));
   NOR3x1_ASAP7_75t_SL U22554 (.Y(n25228),
	.A(n17149),
	.B(n19379),
	.C(n17043));
   NAND2xp33_ASAP7_75t_SRAM U22555 (.Y(n16999),
	.A(n25290),
	.B(n16995));
   INVxp33_ASAP7_75t_SRAM U22558 (.Y(n25895),
	.A(w2_28_));
   INVxp33_ASAP7_75t_SRAM U22563 (.Y(n26615),
	.A(w2_7_));
   NOR3xp33_ASAP7_75t_L U22565 (.Y(n21041),
	.A(n21040),
	.B(n21754),
	.C(n23461));
   NAND3xp33_ASAP7_75t_SRAM U22566 (.Y(n21040),
	.A(n21726),
	.B(n21271),
	.C(n21014));
   A2O1A1Ixp33_ASAP7_75t_SL U22567 (.Y(n26245),
	.A1(n23525),
	.A2(n23524),
	.B(n26710),
	.C(n23523));
   NOR3xp33_ASAP7_75t_L U22568 (.Y(n23525),
	.A(n23486),
	.B(n23485),
	.C(n23484));
   NAND2xp5_ASAP7_75t_L U22569 (.Y(n23524),
	.A(n23495),
	.B(n23494));
   NAND3x1_ASAP7_75t_SL U22571 (.Y(n26248),
	.A(n23482),
	.B(n23481),
	.C(n23480));
   NOR2xp33_ASAP7_75t_L U22572 (.Y(n23481),
	.A(n23479),
	.B(n23478));
   NAND3xp33_ASAP7_75t_SL U22573 (.Y(n23478),
	.A(n23477),
	.B(n23476),
	.C(n23475));
   NAND3xp33_ASAP7_75t_SL U22577 (.Y(n16733),
	.A(n16706),
	.B(n16736),
	.C(n16737));
   NAND2xp5_ASAP7_75t_L U22578 (.Y(n16706),
	.A(n16704),
	.B(n16703));
   O2A1O1Ixp5_ASAP7_75t_SRAM U22580 (.Y(n16740),
	.A1(n16860),
	.A2(n16739),
	.B(n26770),
	.C(n16738));
   OAI222xp33_ASAP7_75t_SL U22581 (.Y(n16738),
	.A1(n16737),
	.A2(n23548),
	.B1(n16736),
	.B2(n23548),
	.C1(n16735),
	.C2(n23548));
   OAI21xp5_ASAP7_75t_L U22582 (.Y(n25077),
	.A1(n17672),
	.A2(n26687),
	.B(n17671));
   O2A1O1Ixp5_ASAP7_75t_SRAM U22583 (.Y(n17671),
	.A1(n24134),
	.A2(n24133),
	.B(FE_OFN16163_n26584),
	.C(n25762));
   NAND2xp33_ASAP7_75t_L U22584 (.Y(n25080),
	.A(n24137),
	.B(n24136));
   INVxp33_ASAP7_75t_SRAM U22586 (.Y(n26656),
	.A(w2_21_));
   A2O1A1Ixp33_ASAP7_75t_SL U22587 (.Y(n24927),
	.A1(n22403),
	.A2(n20124),
	.B(n26346),
	.C(n20123));
   NOR2x1_ASAP7_75t_L U22588 (.Y(n20124),
	.A(n24992),
	.B(n20110));
   NOR2xp33_ASAP7_75t_SL U22589 (.Y(n20123),
	.A(n20122),
	.B(n20121));
   NOR3xp33_ASAP7_75t_SRAM U22591 (.Y(n18964),
	.A(n18963),
	.B(n26003),
	.C(FE_OCPN5051_n25883));
   NOR2x1_ASAP7_75t_L U22592 (.Y(n25882),
	.A(n17021),
	.B(n17098));
   NAND2xp5_ASAP7_75t_SL U22593 (.Y(n17098),
	.A(n24165),
	.B(n19385));
   INVxp33_ASAP7_75t_SRAM U22596 (.Y(n26919),
	.A(w2_26_));
   INVxp33_ASAP7_75t_SRAM U22597 (.Y(n26240),
	.A(w2_29_));
   A2O1A1Ixp33_ASAP7_75t_SL U22598 (.Y(n26223),
	.A1(n18786),
	.A2(n18785),
	.B(n21493),
	.C(n18784));
   NOR3xp33_ASAP7_75t_SRAM U22599 (.Y(n18785),
	.A(n18754),
	.B(FE_OFN28783_n26099),
	.C(n18753));
   INVxp33_ASAP7_75t_R U22600 (.Y(n18786),
	.A(FE_PSN8274_n21164));
   INVxp33_ASAP7_75t_SRAM U22603 (.Y(n26760),
	.A(w2_24_));
   NOR3xp33_ASAP7_75t_SRAM U22605 (.Y(n19440),
	.A(n19439),
	.B(FE_OCPN8245_n25295),
	.C(n25291));
   NOR3xp33_ASAP7_75t_SRAM U22606 (.Y(n19417),
	.A(n19415),
	.B(n25282),
	.C(n25281));
   NOR2x1_ASAP7_75t_L U22607 (.Y(n25286),
	.A(FE_OCPN28189_n20491),
	.B(n19405));
   NAND2xp33_ASAP7_75t_SRAM U22608 (.Y(n19407),
	.A(n19403),
	.B(n19402));
   NAND2xp33_ASAP7_75t_SRAM U22609 (.Y(n19403),
	.A(n19400),
	.B(FE_OFN27147_n25284));
   NAND2xp33_ASAP7_75t_SRAM U22610 (.Y(n19402),
	.A(n19401),
	.B(FE_OFN27147_n25284));
   INVxp33_ASAP7_75t_SRAM U22620 (.Y(n18515),
	.A(w1_0_));
   OAI222xp33_ASAP7_75t_SRAM U22621 (.Y(n21616),
	.A1(FE_OCPN28169_n25121),
	.A2(n26926),
	.B1(n21600),
	.B2(n26926),
	.C1(FE_OFN28540_n21599),
	.C2(n26926));
   NOR2xp33_ASAP7_75t_SRAM U22623 (.Y(n21631),
	.A(n25116),
	.B(n21630));
   NOR3xp33_ASAP7_75t_L U22629 (.Y(n21811),
	.A(n21784),
	.B(n22309),
	.C(n21783));
   NAND3xp33_ASAP7_75t_SL U22630 (.Y(n26531),
	.A(n21768),
	.B(n21781),
	.C(n22280));
   NOR3xp33_ASAP7_75t_L U22631 (.Y(n21768),
	.A(n21767),
	.B(n21766),
	.C(n23194));
   OAI21xp33_ASAP7_75t_SRAM U22632 (.Y(n21767),
	.A1(n18166),
	.A2(FE_OFN16450_n23315),
	.B(n21765));
   INVxp33_ASAP7_75t_SRAM U22634 (.Y(n27173),
	.A(w2_8_));
   O2A1O1Ixp33_ASAP7_75t_L U22636 (.Y(n23893),
	.A1(n23892),
	.A2(n23891),
	.B(n26323),
	.C(n23890));
   NOR2x1_ASAP7_75t_SL U22637 (.Y(n26052),
	.A(FE_OCPN5132_n23890),
	.B(n23889));
   A2O1A1Ixp33_ASAP7_75t_SL U22638 (.Y(n23889),
	.A1(n23895),
	.A2(n23894),
	.B(n26517),
	.C(n23888));
   OAI21xp33_ASAP7_75t_L U22639 (.Y(n23888),
	.A1(n23892),
	.A2(n23891),
	.B(n26323));
   O2A1O1Ixp5_ASAP7_75t_SRAM U22645 (.Y(n25592),
	.A1(n25577),
	.A2(n25576),
	.B(n25575),
	.C(FE_OCPN5115_n25574));
   A2O1A1Ixp33_ASAP7_75t_L U22646 (.Y(n25008),
	.A1(n26857),
	.A2(n26793),
	.B(n26787),
	.C(n25007));
   NAND2xp33_ASAP7_75t_L U22647 (.Y(n25009),
	.A(FE_OCPN27435_n26790),
	.B(n25006));
   INVxp33_ASAP7_75t_SRAM U22648 (.Y(n26041),
	.A(w1_10_));
   INVxp33_ASAP7_75t_SRAM U22649 (.Y(n26932),
	.A(w1_8_));
   NOR3xp33_ASAP7_75t_R U22650 (.Y(n22055),
	.A(n22032),
	.B(n26659),
	.C(n22031));
   INVxp33_ASAP7_75t_SRAM U22652 (.Y(n26287),
	.A(w1_26_));
   INVxp33_ASAP7_75t_SRAM U22654 (.Y(n26474),
	.A(w1_29_));
   INVxp33_ASAP7_75t_SRAM U22655 (.Y(n26611),
	.A(w1_24_));
   INVxp33_ASAP7_75t_SRAM U22656 (.Y(n25184),
	.A(w1_27_));
   NOR3xp33_ASAP7_75t_R U22660 (.Y(n23622),
	.A(n23586),
	.B(FE_OFN26140_n23585),
	.C(n24368));
   NAND3xp33_ASAP7_75t_SRAM U22661 (.Y(n23586),
	.A(n24375),
	.B(n23617),
	.C(n23584));
   INVxp33_ASAP7_75t_L U22662 (.Y(n25451),
	.A(n25452));
   NAND2xp5_ASAP7_75t_SL U22663 (.Y(n25455),
	.A(n24365),
	.B(n23580));
   NAND2xp33_ASAP7_75t_SL U22664 (.Y(n23580),
	.A(n23579),
	.B(n23578));
   NAND2xp33_ASAP7_75t_L U22665 (.Y(n23578),
	.A(n23577),
	.B(n23576));
   NAND2xp33_ASAP7_75t_L U22666 (.Y(n23579),
	.A(n23575),
	.B(n23576));
   INVxp33_ASAP7_75t_SRAM U22668 (.Y(n27106),
	.A(w2_25_));
   INVxp33_ASAP7_75t_L U22669 (.Y(n24286),
	.A(n24996));
   NAND3x1_ASAP7_75t_SL U22670 (.Y(n24289),
	.A(n17550),
	.B(n24988),
	.C(n17549));
   OAI22xp33_ASAP7_75t_SRAM U22671 (.Y(n17549),
	.A1(FE_OCPN28434_n17546),
	.A2(n24991),
	.B1(n17548),
	.B2(n24991));
   NOR3xp33_ASAP7_75t_SRAM U22672 (.Y(n17550),
	.A(n24992),
	.B(FE_OFN27138_n24012),
	.C(n24998));
   A2O1A1Ixp33_ASAP7_75t_SL U22673 (.Y(n25002),
	.A1(n22363),
	.A2(n22362),
	.B(n25585),
	.C(n22361));
   NOR3xp33_ASAP7_75t_L U22674 (.Y(n22362),
	.A(n22342),
	.B(n22341),
	.C(n23638));
   NAND3xp33_ASAP7_75t_R U22675 (.Y(n22342),
	.A(n23650),
	.B(n23640),
	.C(n22339));
   INVxp33_ASAP7_75t_SRAM U22678 (.Y(n21961),
	.A(n27168));
   INVxp33_ASAP7_75t_SRAM U22681 (.Y(n26424),
	.A(w2_30_));
   NOR3xp33_ASAP7_75t_L U22684 (.Y(n24490),
	.A(FE_OCPN29481_n26537),
	.B(n24491),
	.C(n25610));
   INVxp33_ASAP7_75t_SRAM U22686 (.Y(n25490),
	.A(w1_30_));
   INVxp33_ASAP7_75t_SRAM U22687 (.Y(n26448),
	.A(w1_31_));
   INVxp33_ASAP7_75t_SRAM U22688 (.Y(n25499),
	.A(w1_14_));
   OAI21xp5_ASAP7_75t_SL U22689 (.Y(n25497),
	.A1(n24424),
	.A2(n24420),
	.B(n24423));
   A2O1A1Ixp33_ASAP7_75t_SL U22690 (.Y(n24423),
	.A1(FE_OFN16164_n25081),
	.A2(n24422),
	.B(n24421),
	.C(n24420));
   NAND2xp5_ASAP7_75t_SL U22691 (.Y(n24424),
	.A(n24417),
	.B(n24416));
   NAND3xp33_ASAP7_75t_L U22692 (.Y(n26048),
	.A(n25506),
	.B(FE_OCPN5086_n26050),
	.C(n27074));
   NOR3xp33_ASAP7_75t_L U22693 (.Y(n26058),
	.A(n26059),
	.B(FE_OFN1_ld_r),
	.C(FE_OCPN29397_n26502));
   INVxp33_ASAP7_75t_SRAM U22694 (.Y(n26061),
	.A(w2_31_));
   INVxp33_ASAP7_75t_SRAM U22695 (.Y(n25516),
	.A(w2_6_));
   OAI21xp5_ASAP7_75t_SL U22696 (.Y(n25244),
	.A1(FE_OFN1_ld_r),
	.A2(FE_OCPN28138_n26654),
	.B(n25245));
   NOR2xp33_ASAP7_75t_R U22697 (.Y(n25243),
	.A(FE_OCPN27770_n26049),
	.B(FE_OFN28528_n25241));
   NAND2xp5_ASAP7_75t_SL U22699 (.Y(n25195),
	.A(FE_OCPN29443_n25507),
	.B(n25192));
   A2O1A1Ixp33_ASAP7_75t_SL U22700 (.Y(n25194),
	.A1(n26407),
	.A2(n25510),
	.B(FE_OCPN8218_n25507),
	.C(n25193));
   INVxp33_ASAP7_75t_SRAM U22702 (.Y(n25841),
	.A(w2_22_));
   INVxp33_ASAP7_75t_SRAM U22703 (.Y(n24236),
	.A(w1_6_));
   INVxp33_ASAP7_75t_SRAM U22704 (.Y(n25411),
	.A(w1_15_));
   NAND2xp33_ASAP7_75t_L U22705 (.Y(n25406),
	.A(n25404),
	.B(n25403));
   NAND2xp33_ASAP7_75t_R U22706 (.Y(n25403),
	.A(n25402),
	.B(FE_OFN175_sa12_6));
   NOR3xp33_ASAP7_75t_SL U22707 (.Y(n25408),
	.A(n25409),
	.B(FE_OFN16213_ld_r),
	.C(FE_OCPN27519_n25407));
   NAND3xp33_ASAP7_75t_SL U22709 (.Y(n26622),
	.A(n26623),
	.B(n26625),
	.C(n26624));
   A2O1A1Ixp33_ASAP7_75t_SL U22710 (.Y(n26623),
	.A1(n26621),
	.A2(FE_OCPN5133_n26620),
	.B(n26619),
	.C(n26618));
   NAND3xp33_ASAP7_75t_SRAM U22711 (.Y(n26624),
	.A(sa31_6_),
	.B(FE_OFN16334_n25823),
	.C(sa31_7_));
   INVxp33_ASAP7_75t_SRAM U22712 (.Y(n26692),
	.A(w1_7_));
   A2O1A1Ixp33_ASAP7_75t_SL U22714 (.Y(n16143),
	.A1(w2_31_),
	.A2(FE_OFN22_n16125),
	.B(n16131),
	.C(n16130));
   OAI21xp33_ASAP7_75t_SL U22715 (.Y(n16130),
	.A1(ld),
	.A2(w2_31_),
	.B(n16131));
   OAI22xp5_ASAP7_75t_SL U22716 (.Y(n16150),
	.A1(n26692),
	.A2(FE_OFN25891_n15770),
	.B1(n15771),
	.B2(w1_7_));
   A2O1A1Ixp33_ASAP7_75t_SL U22717 (.Y(n14974),
	.A1(n14971),
	.A2(n13865),
	.B(n13864),
	.C(n13863));
   NAND2xp33_ASAP7_75t_L U22718 (.Y(n13864),
	.A(n13861),
	.B(n27064));
   A2O1A1Ixp33_ASAP7_75t_L U22719 (.Y(n13863),
	.A1(n14971),
	.A2(n13865),
	.B(n13862),
	.C(w0_23_));
   NAND3xp33_ASAP7_75t_R U22720 (.Y(n13865),
	.A(n13814),
	.B(n13813),
	.C(n13812));
   AOI22xp5_ASAP7_75t_SL U22721 (.Y(n16069),
	.A1(w1_23_),
	.A2(n14974),
	.B1(n14973),
	.B2(n24608));
   INVxp67_ASAP7_75t_SL U22722 (.Y(n14973),
	.A(n14974));
   OAI21xp5_ASAP7_75t_L U22723 (.Y(n16114),
	.A1(n16069),
	.A2(n27195),
	.B(n16068));
   O2A1O1Ixp33_ASAP7_75t_L U22725 (.Y(n14404),
	.A1(n15704),
	.A2(n14406),
	.B(n14403),
	.C(n26645));
   NOR2xp33_ASAP7_75t_SL U22726 (.Y(n14405),
	.A(w0_30_),
	.B(n14402));
   XNOR2x1_ASAP7_75t_SL U22727 (.Y(n16197),
	.A(w1_30_),
	.B(n15904));
   A2O1A1Ixp33_ASAP7_75t_SL U22728 (.Y(n16117),
	.A1(n15896),
	.A2(n15895),
	.B(n15894),
	.C(n15893));
   NAND2xp5_ASAP7_75t_L U22729 (.Y(n15894),
	.A(n15891),
	.B(n26095));
   NAND3xp33_ASAP7_75t_SL U22730 (.Y(n15895),
	.A(n15807),
	.B(n15806),
	.C(n15805));
   A2O1A1Ixp33_ASAP7_75t_SL U22731 (.Y(n14823),
	.A1(n15757),
	.A2(n14822),
	.B(n14821),
	.C(n14820));
   NAND2xp5_ASAP7_75t_SL U22732 (.Y(n14821),
	.A(w0_29_),
	.B(n14818));
   A2O1A1Ixp33_ASAP7_75t_SL U22733 (.Y(n14820),
	.A1(n14822),
	.A2(n15757),
	.B(n14819),
	.C(n26385));
   XNOR2x1_ASAP7_75t_SL U22734 (.Y(n16186),
	.A(w1_29_),
	.B(n16119));
   A2O1A1Ixp33_ASAP7_75t_SL U22735 (.Y(n16189),
	.A1(w2_29_),
	.A2(FE_OFN22_n16125),
	.B(n16186),
	.C(n16185));
   OAI21xp5_ASAP7_75t_SL U22736 (.Y(n16185),
	.A1(ld),
	.A2(w2_29_),
	.B(n16186));
   A2O1A1Ixp33_ASAP7_75t_SL U22737 (.Y(n14826),
	.A1(n14971),
	.A2(n14002),
	.B(n14001),
	.C(n14000));
   NAND2xp5_ASAP7_75t_L U22738 (.Y(n14001),
	.A(n13998),
	.B(n24358));
   NAND3xp33_ASAP7_75t_R U22739 (.Y(n14002),
	.A(n13948),
	.B(n13947),
	.C(n13946));
   AOI22x1_ASAP7_75t_SL U22740 (.Y(n16103),
	.A1(w1_21_),
	.A2(FE_OFN16300_n14826),
	.B1(FE_OFN28531_FE_OFN56_n14826),
	.B2(n24435));
   OAI21x1_ASAP7_75t_SL U22742 (.Y(n16110),
	.A1(n16103),
	.A2(n26656),
	.B(n16102));
   XNOR2x1_ASAP7_75t_SL U22744 (.Y(n16106),
	.A(w1_28_),
	.B(n15906));
   A2O1A1Ixp33_ASAP7_75t_SL U22745 (.Y(n16113),
	.A1(w2_28_),
	.A2(FE_OFN22_n16125),
	.B(n16106),
	.C(n16105));
   OAI21xp5_ASAP7_75t_SL U22746 (.Y(n16105),
	.A1(ld),
	.A2(w2_28_),
	.B(n16106));
   A2O1A1Ixp33_ASAP7_75t_SL U22747 (.Y(n14664),
	.A1(n13634),
	.A2(n13633),
	.B(n13632),
	.C(n13631));
   NAND2xp5_ASAP7_75t_L U22748 (.Y(n13632),
	.A(n13629),
	.B(n25802));
   A2O1A1Ixp33_ASAP7_75t_SL U22750 (.Y(n14892),
	.A1(FE_OFN16411_n15884),
	.A2(n14894),
	.B(n14891),
	.C(w0_12_));
   NAND2xp33_ASAP7_75t_SL U22751 (.Y(n14879),
	.A(n14878),
	.B(n14877));
   A2O1A1Ixp33_ASAP7_75t_L U22752 (.Y(n14659),
	.A1(n16042),
	.A2(n14661),
	.B(n14658),
	.C(w0_20_));
   NAND2xp5_ASAP7_75t_R U22753 (.Y(n14660),
	.A(n14657),
	.B(n26884));
   NAND2xp33_ASAP7_75t_L U22754 (.Y(n14661),
	.A(n14621),
	.B(n14620));
   AOI22xp5_ASAP7_75t_SL U22755 (.Y(n16213),
	.A1(w1_20_),
	.A2(n16045),
	.B1(n16044),
	.B2(n26698));
   INVx1_ASAP7_75t_SL U22756 (.Y(n16044),
	.A(n16045));
   XNOR2x2_ASAP7_75t_SL U22757 (.Y(n16135),
	.A(u0_rcon_27_),
	.B(n15364));
   A2O1A1Ixp33_ASAP7_75t_SL U22758 (.Y(n15364),
	.A1(n15757),
	.A2(n15363),
	.B(n15362),
	.C(n15361));
   NAND2xp5_ASAP7_75t_SL U22759 (.Y(n15362),
	.A(w0_27_),
	.B(n15359));
   A2O1A1Ixp33_ASAP7_75t_SL U22760 (.Y(n15361),
	.A1(n15363),
	.A2(n15757),
	.B(n15360),
	.C(n24721));
   A2O1A1Ixp33_ASAP7_75t_L U22764 (.Y(n15467),
	.A1(n16042),
	.A2(n15469),
	.B(n15466),
	.C(w0_18_));
   NAND2xp5_ASAP7_75t_SL U22765 (.Y(n15468),
	.A(n15465),
	.B(n24118));
   NAND3xp33_ASAP7_75t_L U22766 (.Y(n15469),
	.A(n15396),
	.B(n15395),
	.C(n15394));
   XNOR2x2_ASAP7_75t_SL U22767 (.Y(n16065),
	.A(u0_rcon_26_),
	.B(n14328));
   O2A1O1Ixp5_ASAP7_75t_SL U22768 (.Y(n14328),
	.A1(n15704),
	.A2(n14327),
	.B(n14326),
	.C(n14325));
   NOR2xp33_ASAP7_75t_L U22769 (.Y(n14326),
	.A(w0_26_),
	.B(n14323));
   O2A1O1Ixp33_ASAP7_75t_SL U22770 (.Y(n14325),
	.A1(n15704),
	.A2(n14327),
	.B(n14324),
	.C(n26396));
   XNOR2x1_ASAP7_75t_SL U22771 (.Y(n16158),
	.A(w1_26_),
	.B(n16065));
   A2O1A1Ixp33_ASAP7_75t_L U22772 (.Y(n16162),
	.A1(w2_26_),
	.A2(FE_OFN22_n16125),
	.B(n16158),
	.C(n16157));
   OAI21xp5_ASAP7_75t_SL U22773 (.Y(n16157),
	.A1(ld),
	.A2(w2_26_),
	.B(n16158));
   A2O1A1Ixp33_ASAP7_75t_SL U22774 (.Y(n14011),
	.A1(n13595),
	.A2(n13479),
	.B(n13478),
	.C(n13477));
   NAND2xp5_ASAP7_75t_L U22775 (.Y(n13478),
	.A(n13475),
	.B(n25265));
   NAND3xp33_ASAP7_75t_L U22776 (.Y(n13479),
	.A(n13425),
	.B(n13424),
	.C(n13423));
   NAND2xp33_ASAP7_75t_R U22777 (.Y(n14970),
	.A(n14902),
	.B(n15457));
   INVxp67_ASAP7_75t_SL U22779 (.Y(n16062),
	.A(n16063));
   OAI21xp5_ASAP7_75t_L U22780 (.Y(n16191),
	.A1(n16175),
	.A2(n26512),
	.B(n16174));
   XNOR2x2_ASAP7_75t_SL U22782 (.Y(n16163),
	.A(u0_rcon_24_),
	.B(n15564));
   O2A1O1Ixp33_ASAP7_75t_SL U22783 (.Y(n15564),
	.A1(n15704),
	.A2(n15563),
	.B(n15562),
	.C(n15561));
   O2A1O1Ixp33_ASAP7_75t_SL U22784 (.Y(n15561),
	.A1(n15704),
	.A2(n15563),
	.B(n15560),
	.C(n26436));
   NOR2xp33_ASAP7_75t_SL U22785 (.Y(n15562),
	.A(w0_24_),
	.B(n15559));
   A2O1A1Ixp33_ASAP7_75t_SL U22786 (.Y(n14091),
	.A1(n15263),
	.A2(n13548),
	.B(n13547),
	.C(n13546));
   NAND2xp33_ASAP7_75t_R U22787 (.Y(n13547),
	.A(n13544),
	.B(n26772));
   NAND3xp33_ASAP7_75t_L U22788 (.Y(n13548),
	.A(n13498),
	.B(n13497),
	.C(n13496));
   AOI22xp5_ASAP7_75t_SL U22789 (.Y(n16194),
	.A1(w1_13_),
	.A2(FE_OCPN29581_n16097),
	.B1(n16096),
	.B2(n25774));
   OAI21xp5_ASAP7_75t_SL U22790 (.Y(n16240),
	.A1(n16194),
	.A2(n26416),
	.B(n16193));
   NAND2xp33_ASAP7_75t_SL U22792 (.Y(n14741),
	.A(n14738),
	.B(n25975));
   A2O1A1Ixp33_ASAP7_75t_SL U22793 (.Y(n14740),
	.A1(n16042),
	.A2(n14742),
	.B(n14739),
	.C(w0_17_));
   NAND3xp33_ASAP7_75t_SL U22794 (.Y(n14742),
	.A(n14679),
	.B(n14678),
	.C(n14677));
   O2A1O1Ixp5_ASAP7_75t_SL U22795 (.Y(n15768),
	.A1(n13901),
	.A2(n15767),
	.B(n15766),
	.C(n15765));
   NOR2xp33_ASAP7_75t_L U22796 (.Y(n15766),
	.A(w0_25_),
	.B(n15763));
   O2A1O1Ixp33_ASAP7_75t_SL U22797 (.Y(n15765),
	.A1(n13901),
	.A2(n15767),
	.B(n15764),
	.C(n24575));
   XNOR2x1_ASAP7_75t_SL U22798 (.Y(n16237),
	.A(w1_25_),
	.B(n16138));
   A2O1A1Ixp33_ASAP7_75t_L U22799 (.Y(n16263),
	.A1(w2_25_),
	.A2(FE_OFN22_n16125),
	.B(n16237),
	.C(n16236));
   OAI21xp5_ASAP7_75t_SL U22800 (.Y(n16236),
	.A1(ld),
	.A2(w2_25_),
	.B(n16237));
   AOI22xp5_ASAP7_75t_SL U22801 (.Y(n16199),
	.A1(w1_9_),
	.A2(FE_OCPN29468_n15919),
	.B1(n15918),
	.B2(n24821));
   OAI22xp5_ASAP7_75t_SL U22802 (.Y(n16248),
	.A1(n25729),
	.A2(n16076),
	.B1(n16075),
	.B2(w1_16_));
   OAI21xp5_ASAP7_75t_SL U22803 (.Y(n16273),
	.A1(w2_6_),
	.A2(n16184),
	.B(n16183));
   NOR2xp33_ASAP7_75t_SRAM U22805 (.Y(n16275),
	.A(key_6_),
	.B(FE_OFN22_n16125));
   INVxp33_ASAP7_75t_SRAM U22806 (.Y(n16287),
	.A(u0_r0_rcnt_3_));
   INVxp33_ASAP7_75t_SRAM U22807 (.Y(n13269),
	.A(u0_r0_rcnt_1_));
   NOR2xp33_ASAP7_75t_SRAM U22808 (.Y(n16285),
	.A(n13269),
	.B(n16286));
   O2A1O1Ixp5_ASAP7_75t_L U22809 (.Y(n440),
	.A1(w1_3_),
	.A2(text_in_r_67_),
	.B(n26593),
	.C(n26592));
   O2A1O1Ixp5_ASAP7_75t_SL U22810 (.Y(n26592),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(FE_OCPN27519_n25407),
	.B(n26591),
	.C(n26590));
   A2O1A1Ixp33_ASAP7_75t_SL U22811 (.Y(n340),
	.A1(n26800),
	.A2(n26799),
	.B(FE_OFN25881_w3_24),
	.C(n26797));
   A2O1A1Ixp33_ASAP7_75t_L U22812 (.Y(n26800),
	.A1(FE_OCPN29381_n26796),
	.A2(FE_OFN28490_ld_r),
	.B(n26795),
	.C(n26794));
   NAND2xp33_ASAP7_75t_SRAM U22813 (.Y(n26799),
	.A(FE_OFN28482_ld_r),
	.B(text_in_r_24_));
   A2O1A1Ixp33_ASAP7_75t_SL U22814 (.Y(n478),
	.A1(n25776),
	.A2(n25775),
	.B(n25774),
	.C(n25773));
   NAND3xp33_ASAP7_75t_SL U22815 (.Y(n25773),
	.A(n25774),
	.B(n25776),
	.C(n25775));
   A2O1A1Ixp33_ASAP7_75t_SL U22816 (.Y(n25776),
	.A1(n26713),
	.A2(FE_OFN28487_ld_r),
	.B(n25772),
	.C(n25771));
   NAND2xp33_ASAP7_75t_SRAM U22817 (.Y(n25775),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_77_));
   OAI21xp33_ASAP7_75t_SRAM U22818 (.Y(n24532),
	.A1(text_in_r_98_),
	.A2(n24531),
	.B(n24530));
   OAI21xp5_ASAP7_75t_SL U22819 (.Y(n24533),
	.A1(n24535),
	.A2(n24534),
	.B(FE_OFN28484_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22820 (.Y(n24530),
	.A1(text_in_r_98_),
	.A2(FE_OFN28484_ld_r),
	.B1(n24531),
	.B2(FE_OFN28484_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22821 (.Y(n23938),
	.A1(text_in_r_2_),
	.A2(n23937),
	.B(n23936));
   OAI21xp33_ASAP7_75t_SL U22822 (.Y(n23939),
	.A1(n23940),
	.A2(n25423),
	.B(FE_OFN28489_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22823 (.Y(n23936),
	.A1(text_in_r_2_),
	.A2(FE_OFN28489_ld_r),
	.B1(n23937),
	.B2(FE_OFN28489_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22824 (.Y(n26019),
	.A1(text_in_r_44_),
	.A2(n26018),
	.B(n26017));
   A2O1A1Ixp33_ASAP7_75t_SL U22825 (.Y(n329),
	.A1(n26921),
	.A2(n26920),
	.B(n26919),
	.C(n26918));
   NAND2xp33_ASAP7_75t_SRAM U22826 (.Y(n26920),
	.A(FE_OFN1_ld_r),
	.B(text_in_r_58_));
   O2A1O1Ixp33_ASAP7_75t_SL U22827 (.Y(n26896),
	.A1(FE_OFN2_ld_r),
	.A2(n26895),
	.B(n26894),
	.C(n26893));
   NOR2x1_ASAP7_75t_SL U22828 (.Y(n26893),
	.A(n26892),
	.B(n26894));
   A2O1A1Ixp33_ASAP7_75t_SL U22829 (.Y(n509),
	.A1(n26613),
	.A2(n26612),
	.B(n26611),
	.C(n26610));
   NAND2xp33_ASAP7_75t_SRAM U22830 (.Y(n26612),
	.A(FE_OFN16213_ld_r),
	.B(text_in_r_88_));
   A2O1A1Ixp33_ASAP7_75t_L U22831 (.Y(n16177),
	.A1(FE_OFN29087_n),
	.A2(FE_OFN28460_ld),
	.B(n16176),
	.C(FE_OCPN29371_n16191));
   NOR2xp33_ASAP7_75t_SRAM U22832 (.Y(n16176),
	.A(key_19_),
	.B(FE_OFN28460_ld));
   OAI21xp5_ASAP7_75t_SL U22833 (.Y(n627),
	.A1(n16172),
	.A2(FE_OFN28674_n),
	.B(n16147));
   NOR2xp33_ASAP7_75t_SRAM U22834 (.Y(n16146),
	.A(key_17_),
	.B(FE_OFN26_n16125));
   OAI21xp33_ASAP7_75t_SRAM U22835 (.Y(n27130),
	.A1(text_in_r_101_),
	.A2(n27129),
	.B(n27128));
   OAI22xp33_ASAP7_75t_SRAM U22836 (.Y(n27128),
	.A1(text_in_r_101_),
	.A2(FE_OFN28484_ld_r),
	.B1(n27129),
	.B2(FE_OFN28484_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22837 (.Y(n23975),
	.A1(text_in_r_18_),
	.A2(FE_OFN16421_n23974),
	.B(n23973));
   OAI21xp5_ASAP7_75t_SL U22838 (.Y(n23976),
	.A1(n23978),
	.A2(n23977),
	.B(FE_OFN28489_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22839 (.Y(n23973),
	.A1(text_in_r_18_),
	.A2(FE_OFN28489_ld_r),
	.B1(FE_OFN16421_n23974),
	.B2(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U22840 (.Y(n424),
	.A1(n26043),
	.A2(n26042),
	.B(n26041),
	.C(n26040));
   NAND3xp33_ASAP7_75t_L U22841 (.Y(n26040),
	.A(n26041),
	.B(n26043),
	.C(n26042));
   NAND2xp33_ASAP7_75t_SRAM U22842 (.Y(n26042),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_74_));
   A2O1A1Ixp33_ASAP7_75t_SL U22843 (.Y(n464),
	.A1(n25784),
	.A2(n25783),
	.B(FE_OFN26163_w3_13),
	.C(n25781));
   NAND2xp33_ASAP7_75t_SRAM U22845 (.Y(n25783),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_13_));
   A2O1A1Ixp33_ASAP7_75t_SL U22846 (.Y(n401),
	.A1(n26289),
	.A2(n26288),
	.B(n26287),
	.C(n26286));
   A2O1A1Ixp33_ASAP7_75t_SL U22847 (.Y(n26289),
	.A1(n26285),
	.A2(FE_OFN28487_ld_r),
	.B(n26284),
	.C(n26283));
   NAND2xp33_ASAP7_75t_SRAM U22848 (.Y(n26288),
	.A(FE_OFN16213_ld_r),
	.B(text_in_r_90_));
   NOR3xp33_ASAP7_75t_SL U22849 (.Y(n26987),
	.A(n26989),
	.B(w2_16_),
	.C(n26988));
   NOR3xp33_ASAP7_75t_SL U22850 (.Y(n26988),
	.A(n27147),
	.B(FE_OFN12_FE_DBTN0_ld_r),
	.C(n26986));
   OAI21xp33_ASAP7_75t_SL U22851 (.Y(n648),
	.A1(n16265),
	.A2(FE_OCPN28408_FE_OFN16433_w3_11),
	.B(n16227));
   NOR2xp33_ASAP7_75t_SRAM U22852 (.Y(n16226),
	.A(key_11_),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SL U22853 (.Y(n650),
	.A1(n16207),
	.A2(n16206),
	.B(n16205));
   NAND2xp33_ASAP7_75t_SRAM U22854 (.Y(n16207),
	.A(FE_OFN28472_ld),
	.B(n24688));
   OAI21xp5_ASAP7_75t_L U22855 (.Y(n16205),
	.A1(FE_OFN21_n16125),
	.A2(FE_OFN27206_w3_30),
	.B(n16204));
   OAI21xp5_ASAP7_75t_SL U22856 (.Y(n16204),
	.A1(key_30_),
	.A2(FE_OFN28472_ld),
	.B(n16203));
   OAI21xp33_ASAP7_75t_SRAM U22857 (.Y(n25571),
	.A1(text_in_r_59_),
	.A2(n25570),
	.B(n25569));
   OAI21xp33_ASAP7_75t_SRAM U22858 (.Y(n24722),
	.A1(text_in_r_123_),
	.A2(n24721),
	.B(n24720));
   OAI21xp33_ASAP7_75t_L U22859 (.Y(n24723),
	.A1(n24724),
	.A2(FE_OCPN29540_FE_OFN25927_n26527),
	.B(FE_OFN28483_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22860 (.Y(n24720),
	.A1(text_in_r_123_),
	.A2(FE_OFN28483_ld_r),
	.B1(n24721),
	.B2(FE_OFN28483_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U22861 (.Y(n15373),
	.A1(FE_OFN28732_n),
	.A2(FE_OFN26_n16125),
	.B(n15372),
	.C(n15916));
   NOR2xp33_ASAP7_75t_SRAM U22862 (.Y(n15372),
	.A(key_1_),
	.B(FE_OFN26_n16125));
   OAI22xp33_ASAP7_75t_SRAM U22863 (.Y(n25760),
	.A1(w1_19_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_83_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U22864 (.Y(n25759),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27884_n26717),
	.B(FE_OCPN5080_n25758),
	.C(n25757));
   NOR2xp33_ASAP7_75t_SL U22865 (.Y(n25757),
	.A(n26714),
	.B(n25758));
   OAI21xp33_ASAP7_75t_SRAM U22866 (.Y(n24436),
	.A1(text_in_r_85_),
	.A2(n24435),
	.B(n24434));
   OAI21xp33_ASAP7_75t_SRAM U22867 (.Y(n25434),
	.A1(text_in_r_11_),
	.A2(FE_OFN28853_FE_OCPN28408),
	.B(n25432));
   OAI21xp33_ASAP7_75t_L U22868 (.Y(n25435),
	.A1(n25436),
	.A2(FE_OCPN27282_n25437),
	.B(FE_OFN28489_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22869 (.Y(n26131),
	.A1(text_in_r_108_),
	.A2(n26130),
	.B(n26129));
   OAI21xp33_ASAP7_75t_SL U22870 (.Y(n26132),
	.A1(n26133),
	.A2(FE_OCPN27321_n26380),
	.B(FE_OFN28483_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U22871 (.Y(n25665),
	.A1(FE_OFN16214_ld_r),
	.A2(n26852),
	.B(n25664),
	.C(n25663));
   OAI21xp33_ASAP7_75t_SRAM U22872 (.Y(n24027),
	.A1(text_in_r_5_),
	.A2(FE_OFN16276_w3_5),
	.B(n24025));
   OAI21xp5_ASAP7_75t_SL U22873 (.Y(n24028),
	.A1(n24029),
	.A2(FE_OCPN27505_n24684),
	.B(FE_OFN28490_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22874 (.Y(n24025),
	.A1(text_in_r_5_),
	.A2(FE_OFN28490_ld_r),
	.B1(FE_OFN16276_w3_5),
	.B2(FE_OFN28490_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U22875 (.Y(n443),
	.A1(FE_OCPN27362_n25679),
	.A2(n25678),
	.B(n25677),
	.C(n25676));
   OAI21xp33_ASAP7_75t_SRAM U22876 (.Y(n25676),
	.A1(text_in_r_27_),
	.A2(FE_OFN26120_n),
	.B(n25674));
   A2O1A1Ixp33_ASAP7_75t_SL U22878 (.Y(n470),
	.A1(n25053),
	.A2(n25052),
	.B(n25051),
	.C(n25050));
   A2O1A1Ixp33_ASAP7_75t_SL U22880 (.Y(n25053),
	.A1(FE_OCPN27292_n25389),
	.A2(FE_OFN28489_ld_r),
	.B(n25049),
	.C(n25048));
   OAI21xp33_ASAP7_75t_SRAM U22881 (.Y(n25896),
	.A1(text_in_r_60_),
	.A2(n25895),
	.B(n25894));
   OAI21xp5_ASAP7_75t_SL U22882 (.Y(n25897),
	.A1(n25898),
	.A2(FE_OCPN29356_n27110),
	.B(FE_OFN16_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22883 (.Y(n26096),
	.A1(text_in_r_107_),
	.A2(n26095),
	.B(n26094));
   OAI21xp33_ASAP7_75t_SL U22885 (.Y(n24120),
	.A1(n24121),
	.A2(FE_OCPN27941_n),
	.B(FE_OFN28484_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22886 (.Y(n24119),
	.A1(text_in_r_114_),
	.A2(n24118),
	.B(n24117));
   O2A1O1Ixp5_ASAP7_75t_SL U22887 (.Y(n24121),
	.A1(FE_OFN28934_n24552),
	.A2(n24112),
	.B(n24111),
	.C(n24110));
   A2O1A1Ixp33_ASAP7_75t_SL U22888 (.Y(n425),
	.A1(FE_OCPN29572_n24468),
	.A2(n24295),
	.B(n24294),
	.C(n24293));
   OAI21xp33_ASAP7_75t_SRAM U22889 (.Y(n24293),
	.A1(text_in_r_9_),
	.A2(FE_OFN27111_n),
	.B(n24291));
   OAI21xp33_ASAP7_75t_SL U22890 (.Y(n24294),
	.A1(n24295),
	.A2(FE_OCPN29572_n24468),
	.B(FE_OFN28489_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22891 (.Y(n25691),
	.A1(text_in_r_75_),
	.A2(n25690),
	.B(n25689));
   OAI21xp33_ASAP7_75t_L U22892 (.Y(n25692),
	.A1(n25693),
	.A2(FE_OCPN7585_FE_OFN25926_n26922),
	.B(FE_OFN28486_ld_r));
   NAND3xp33_ASAP7_75t_SL U22893 (.Y(n25728),
	.A(n25729),
	.B(n25731),
	.C(n25730));
   NAND3xp33_ASAP7_75t_R U22894 (.Y(n25730),
	.A(n25727),
	.B(FE_OFN28486_ld_r),
	.C(FE_OCPN27884_n26717));
   A2O1A1Ixp33_ASAP7_75t_SL U22895 (.Y(n476),
	.A1(n24643),
	.A2(n24642),
	.B(n24641),
	.C(n24640));
   NAND3xp33_ASAP7_75t_SL U22896 (.Y(n24640),
	.A(n24641),
	.B(n24643),
	.C(n24642));
   A2O1A1Ixp33_ASAP7_75t_SL U22897 (.Y(n24643),
	.A1(FE_OCPN29365_n24639),
	.A2(FE_OFN28483_ld_r),
	.B(n24638),
	.C(n24637));
   NAND2xp33_ASAP7_75t_SRAM U22898 (.Y(n24642),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_106_));
   A2O1A1Ixp33_ASAP7_75t_SL U22899 (.Y(n376),
	.A1(n26398),
	.A2(n26397),
	.B(n26396),
	.C(n26395));
   NAND2xp33_ASAP7_75t_SRAM U22901 (.Y(n26397),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_122_));
   O2A1O1Ixp33_ASAP7_75t_SL U22902 (.Y(n26231),
	.A1(FE_OFN2_ld_r),
	.A2(n26895),
	.B(FE_OCPN5043_n26230),
	.C(n26229));
   NOR2xp33_ASAP7_75t_SL U22903 (.Y(n26229),
	.A(n26892),
	.B(n26230));
   A2O1A1Ixp33_ASAP7_75t_SL U22904 (.Y(n481),
	.A1(n26189),
	.A2(n26188),
	.B(n26187),
	.C(n26186));
   OAI21xp33_ASAP7_75t_SRAM U22905 (.Y(n26186),
	.A1(text_in_r_66_),
	.A2(n26185),
	.B(n26184));
   OAI21x1_ASAP7_75t_SL U22906 (.Y(n26187),
	.A1(n26189),
	.A2(n26188),
	.B(FE_OFN14_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22907 (.Y(n24359),
	.A1(text_in_r_117_),
	.A2(n24358),
	.B(n24357));
   OAI21xp5_ASAP7_75t_SL U22908 (.Y(n24360),
	.A1(n24361),
	.A2(FE_OCPN27412_n24491),
	.B(FE_OFN15_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_SL U22909 (.Y(n24823),
	.A1(n24824),
	.A2(FE_OCPN27439_n27030),
	.B(FE_OFN28486_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22910 (.Y(n24413),
	.A1(text_in_r_82_),
	.A2(n24412),
	.B(n24411));
   OAI21xp33_ASAP7_75t_L U22911 (.Y(n24414),
	.A1(n24415),
	.A2(n26285),
	.B(FE_OFN28487_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22912 (.Y(n24150),
	.A1(text_in_r_69_),
	.A2(n24149),
	.B(n24148));
   OAI22xp33_ASAP7_75t_SRAM U22913 (.Y(n24148),
	.A1(text_in_r_69_),
	.A2(FE_OFN28487_ld_r),
	.B1(n24149),
	.B2(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U22914 (.Y(n518),
	.A1(FE_OCPN8212_n26261),
	.A2(n25131),
	.B(n25130),
	.C(n25129));
   OAI21xp33_ASAP7_75t_SRAM U22915 (.Y(n25129),
	.A1(text_in_r_76_),
	.A2(n25128),
	.B(n25127));
   OAI21xp33_ASAP7_75t_SL U22916 (.Y(n25130),
	.A1(n25131),
	.A2(FE_OCPN8212_n26261),
	.B(FE_OFN28486_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22917 (.Y(n25127),
	.A1(text_in_r_76_),
	.A2(FE_OFN28486_ld_r),
	.B1(n25128),
	.B2(FE_OFN28486_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22918 (.Y(n27196),
	.A1(text_in_r_55_),
	.A2(n27195),
	.B(n27194));
   OAI21xp33_ASAP7_75t_SRAM U22919 (.Y(n25185),
	.A1(text_in_r_91_),
	.A2(n25184),
	.B(n25183));
   OAI21xp33_ASAP7_75t_L U22920 (.Y(n25186),
	.A1(n25187),
	.A2(FE_OCPN27560_n25755),
	.B(FE_OFN28487_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U22921 (.Y(n25271),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OFN26024_n26115),
	.B(n25270),
	.C(n25269));
   NOR2x1_ASAP7_75t_L U22922 (.Y(n25269),
	.A(n26781),
	.B(n25270));
   OAI21xp33_ASAP7_75t_SRAM U22923 (.Y(n24321),
	.A1(text_in_r_105_),
	.A2(n24320),
	.B(n24319));
   O2A1O1Ixp33_ASAP7_75t_SL U22925 (.Y(n26208),
	.A1(FE_OFN1_ld_r),
	.A2(n26330),
	.B(FE_OCPN5146_n26207),
	.C(n26206));
   NOR2xp33_ASAP7_75t_SL U22926 (.Y(n26206),
	.A(n26327),
	.B(n26207));
   A2O1A1Ixp33_ASAP7_75t_SL U22927 (.Y(n480),
	.A1(n26418),
	.A2(n26417),
	.B(n26416),
	.C(n26415));
   NAND3xp33_ASAP7_75t_SL U22928 (.Y(n26415),
	.A(n26416),
	.B(n26418),
	.C(n26417));
   NAND2xp33_ASAP7_75t_SRAM U22930 (.Y(n26417),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_45_));
   A2O1A1Ixp33_ASAP7_75t_SL U22931 (.Y(n491),
	.A1(n26658),
	.A2(n26657),
	.B(n26656),
	.C(n26655));
   NAND2xp33_ASAP7_75t_SRAM U22932 (.Y(n26657),
	.A(FE_OFN12_FE_DBTN0_ld_r),
	.B(text_in_r_53_));
   A2O1A1Ixp33_ASAP7_75t_SL U22933 (.Y(n454),
	.A1(n26476),
	.A2(n26475),
	.B(n26474),
	.C(n26473));
   NAND2xp33_ASAP7_75t_SRAM U22934 (.Y(n26475),
	.A(FE_OFN16213_ld_r),
	.B(text_in_r_93_));
   NAND3xp33_ASAP7_75t_SL U22935 (.Y(n26810),
	.A(n26811),
	.B(n26813),
	.C(n26812));
   A2O1A1Ixp33_ASAP7_75t_SL U22936 (.Y(n26813),
	.A1(FE_OCPN27379_n26809),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B(n26808),
	.C(n26807));
   NAND2xp33_ASAP7_75t_SRAM U22937 (.Y(n26812),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_127_));
   OAI21xp33_ASAP7_75t_SL U22938 (.Y(n641),
	.A1(n16078),
	.A2(FE_OFN26073_n),
	.B(n16061));
   NOR2xp33_ASAP7_75t_SRAM U22939 (.Y(n16060),
	.A(key_4_),
	.B(FE_OFN26_n16125));
   O2A1O1Ixp5_ASAP7_75t_SL U22940 (.Y(n344),
	.A1(FE_OFN38_w0_17),
	.A2(text_in_r_113_),
	.B(n25986),
	.C(n25985));
   OAI22xp33_ASAP7_75t_SRAM U22941 (.Y(n25986),
	.A1(FE_OFN38_w0_17),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_113_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U22942 (.Y(n25985),
	.A1(FE_OFN2_ld_r),
	.A2(n26895),
	.B(FE_OCPN5068_n25984),
	.C(n25983));
   NOR3xp33_ASAP7_75t_SL U22943 (.Y(n24455),
	.A(n24457),
	.B(FE_OFN16432_w3_16),
	.C(n24456));
   OAI21xp5_ASAP7_75t_SL U22944 (.Y(n24457),
	.A1(text_in_r_16_),
	.A2(FE_OFN28489_ld_r),
	.B(n24453));
   NOR3xp33_ASAP7_75t_SL U22945 (.Y(n24456),
	.A(n24454),
	.B(FE_OFN16214_ld_r),
	.C(n25390));
   OAI21xp33_ASAP7_75t_L U22946 (.Y(n24577),
	.A1(n24578),
	.A2(FE_OCPN29540_FE_OFN25927_n26527),
	.B(FE_OFN28483_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22947 (.Y(n24574),
	.A1(text_in_r_121_),
	.A2(FE_OFN28483_ld_r),
	.B1(n24575),
	.B2(FE_OFN28483_ld_r));
   NOR3xp33_ASAP7_75t_SL U22949 (.Y(n26117),
	.A(n26119),
	.B(w0_0_),
	.C(n26118));
   NOR3xp33_ASAP7_75t_SL U22950 (.Y(n26118),
	.A(n26116),
	.B(FE_OFN2_ld_r),
	.C(n26784));
   OAI21xp33_ASAP7_75t_SRAM U22951 (.Y(n25347),
	.A1(text_in_r_41_),
	.A2(n25346),
	.B(n25345));
   NAND3xp33_ASAP7_75t_SL U22953 (.Y(n26743),
	.A(n26744),
	.B(n26746),
	.C(n26745));
   NAND2xp33_ASAP7_75t_SRAM U22954 (.Y(n26745),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_104_));
   A2O1A1Ixp33_ASAP7_75t_SL U22955 (.Y(n390),
	.A1(n26849),
	.A2(n26848),
	.B(FE_OFN25961_w3_8),
	.C(n26846));
   NAND2xp33_ASAP7_75t_SRAM U22956 (.Y(n26848),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_8_));
   OAI21xp5_ASAP7_75t_L U22957 (.Y(n25460),
	.A1(n25461),
	.A2(FE_OCPN29382_n26674),
	.B(FE_OFN28487_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22958 (.Y(n25457),
	.A1(text_in_r_89_),
	.A2(FE_OFN28487_ld_r),
	.B1(FE_OFN66_w1_25),
	.B2(FE_OFN28487_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U22959 (.Y(n25393),
	.A1(FE_OFN16214_ld_r),
	.A2(n26732),
	.B(n25392),
	.C(n25391));
   NOR2x1_ASAP7_75t_SL U22960 (.Y(n25391),
	.A(n26729),
	.B(n25392));
   O2A1O1Ixp5_ASAP7_75t_SL U22961 (.Y(n25943),
	.A1(FE_OFN1_ld_r),
	.A2(n26330),
	.B(n25942),
	.C(n25941));
   NOR2x1_ASAP7_75t_SL U22962 (.Y(n25941),
	.A(n26327),
	.B(n25942));
   NAND2xp33_ASAP7_75t_SRAM U22964 (.Y(n27174),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_40_));
   OAI21xp33_ASAP7_75t_SRAM U22965 (.Y(n24985),
	.A1(text_in_r_28_),
	.A2(FE_OFN28571_w3_28),
	.B(n24983));
   OAI21xp5_ASAP7_75t_L U22966 (.Y(n24986),
	.A1(n24987),
	.A2(FE_OCPN27787_n26728),
	.B(FE_OFN28490_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22967 (.Y(n24983),
	.A1(text_in_r_28_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(FE_OFN28571_w3_28),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   O2A1O1Ixp5_ASAP7_75t_L U22968 (.Y(n27148),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(n27147),
	.B(n27146),
	.C(n27145));
   NOR2x1_ASAP7_75t_L U22969 (.Y(n27145),
	.A(n27144),
	.B(n27146));
   OAI21xp33_ASAP7_75t_SRAM U22970 (.Y(n26143),
	.A1(text_in_r_92_),
	.A2(n26142),
	.B(n26141));
   OAI22xp33_ASAP7_75t_SRAM U22971 (.Y(n26141),
	.A1(text_in_r_92_),
	.A2(FE_OFN28487_ld_r),
	.B1(n26142),
	.B2(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U22972 (.Y(n444),
	.A1(n26343),
	.A2(n26342),
	.B(FE_OCPN29428_FE_OFN27131_w3_29),
	.C(n26340));
   NAND3xp33_ASAP7_75t_SL U22973 (.Y(n26340),
	.A(FE_OCPN29428_FE_OFN27131_w3_29),
	.B(n26343),
	.C(n26342));
   OAI21xp33_ASAP7_75t_SL U22974 (.Y(n25618),
	.A1(n25620),
	.A2(n25619),
	.B(FE_OFN15_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U22975 (.Y(n25617),
	.A1(text_in_r_118_),
	.A2(n25616),
	.B(n25615));
   AOI22xp33_ASAP7_75t_SRAM U22976 (.Y(n25619),
	.A1(FE_OCPN27447_n26638),
	.A2(n25616),
	.B1(w0_22_),
	.B2(n26639));
   A2O1A1Ixp33_ASAP7_75t_L U22977 (.Y(n447),
	.A1(n26953),
	.A2(n26952),
	.B(n26951),
	.C(n26950));
   NAND3xp33_ASAP7_75t_L U22978 (.Y(n26950),
	.A(n26951),
	.B(n26953),
	.C(n26952));
   NAND2xp33_ASAP7_75t_SRAM U22979 (.Y(n26952),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_42_));
   OAI21xp5_ASAP7_75t_SL U22980 (.Y(n25707),
	.A1(text_in_r_64_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B(n25703));
   NOR3xp33_ASAP7_75t_SL U22981 (.Y(n25706),
	.A(FE_OCPN27519_n25407),
	.B(FE_OFN12_FE_DBTN0_ld_r),
	.C(n25704));
   A2O1A1Ixp33_ASAP7_75t_SL U22982 (.Y(n449),
	.A1(n27223),
	.A2(n27222),
	.B(n27221),
	.C(n27220));
   OAI21xp33_ASAP7_75t_SRAM U22983 (.Y(n27220),
	.A1(text_in_r_50_),
	.A2(n27219),
	.B(n27218));
   OAI21x1_ASAP7_75t_SL U22984 (.Y(n27221),
	.A1(n27223),
	.A2(n27222),
	.B(FE_OFN16215_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22985 (.Y(n27218),
	.A1(text_in_r_50_),
	.A2(FE_OFN16215_ld_r),
	.B1(n27219),
	.B2(FE_OFN16215_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U22986 (.Y(n452),
	.A1(FE_OCPN28122_n27157),
	.A2(n26378),
	.B(n26377),
	.C(n26376));
   OAI21xp33_ASAP7_75t_SRAM U22987 (.Y(n26376),
	.A1(text_in_r_124_),
	.A2(n26375),
	.B(n26374));
   OAI21xp5_ASAP7_75t_SL U22988 (.Y(n26377),
	.A1(n26378),
	.A2(FE_OCPN28122_n27157),
	.B(FE_OFN28483_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22989 (.Y(n26524),
	.A1(w2_19_),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B1(text_in_r_51_),
	.B2(FE_OFN16_FE_DBTN0_ld_r));
   O2A1O1Ixp5_ASAP7_75t_L U22990 (.Y(n26523),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(n27147),
	.B(n26522),
	.C(n26521));
   NOR2xp67_ASAP7_75t_SL U22991 (.Y(n26521),
	.A(n27144),
	.B(n26522));
   O2A1O1Ixp5_ASAP7_75t_SL U22992 (.Y(n459),
	.A1(FE_OCPN8254_w3_3),
	.A2(text_in_r_3_),
	.B(n25156),
	.C(n25155));
   O2A1O1Ixp33_ASAP7_75t_SL U22993 (.Y(n25155),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27476_n26852),
	.B(n25154),
	.C(n25153));
   OAI21xp33_ASAP7_75t_SRAM U22994 (.Y(n26964),
	.A1(text_in_r_43_),
	.A2(n26963),
	.B(n26962));
   OAI21xp33_ASAP7_75t_L U22995 (.Y(n26965),
	.A1(n26966),
	.A2(n27176),
	.B(FE_OFN16215_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22996 (.Y(n27036),
	.A1(w1_1_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_65_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U22999 (.Y(n26332),
	.A1(w2_3_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_35_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL U23000 (.Y(n26328),
	.A(n26327),
	.B(n26329));
   A2O1A1Ixp33_ASAP7_75t_SL U23001 (.Y(n472),
	.A1(n26242),
	.A2(n26241),
	.B(n26240),
	.C(n26239));
   NAND3xp33_ASAP7_75t_SL U23002 (.Y(n26239),
	.A(n26240),
	.B(n26242),
	.C(n26241));
   A2O1A1Ixp33_ASAP7_75t_SL U23003 (.Y(n26242),
	.A1(FE_OCPN28138_n26654),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B(n26238),
	.C(n26237));
   NAND2xp33_ASAP7_75t_SRAM U23004 (.Y(n26241),
	.A(FE_OFN1_ld_r),
	.B(text_in_r_61_));
   OAI21xp33_ASAP7_75t_SRAM U23005 (.Y(n24201),
	.A1(text_in_r_37_),
	.A2(n24200),
	.B(n24199));
   OAI21xp33_ASAP7_75t_L U23006 (.Y(n24202),
	.A1(n24204),
	.A2(n24203),
	.B(FE_OFN14_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U23007 (.Y(n24199),
	.A1(text_in_r_37_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(n24200),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U23008 (.Y(n26506),
	.A1(w2_20_),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B1(text_in_r_52_),
	.B2(FE_OFN16_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL U23009 (.Y(n26503),
	.A(n27144),
	.B(n26504));
   OAI22xp33_ASAP7_75t_SRAM U23010 (.Y(n25814),
	.A1(w0_4_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_100_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   NOR2x1_ASAP7_75t_SL U23011 (.Y(n25811),
	.A(n26781),
	.B(n25812));
   OAI22xp33_ASAP7_75t_SRAM U23012 (.Y(n26719),
	.A1(w1_20_),
	.A2(FE_OFN28486_ld_r),
	.B1(text_in_r_84_),
	.B2(FE_OFN28486_ld_r));
   O2A1O1Ixp33_ASAP7_75t_L U23013 (.Y(n26718),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27884_n26717),
	.B(FE_OCPN5022_n26716),
	.C(n26715));
   NOR2x1_ASAP7_75t_SL U23014 (.Y(n26715),
	.A(n26714),
	.B(FE_OCPN5022_n26716));
   NAND3xp33_ASAP7_75t_SL U23015 (.Y(n25373),
	.A(FE_OFN26640_w3_14),
	.B(n25376),
	.C(n25375));
   NAND2xp33_ASAP7_75t_SRAM U23016 (.Y(n25375),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_14_));
   A2O1A1Ixp33_ASAP7_75t_SL U23017 (.Y(n504),
	.A1(n26274),
	.A2(n26273),
	.B(n26272),
	.C(n26271));
   NAND3xp33_ASAP7_75t_SL U23018 (.Y(n26271),
	.A(n26272),
	.B(n26274),
	.C(n26273));
   NAND2xp5_ASAP7_75t_L U23019 (.Y(n26273),
	.A(n26781),
	.B(n26270));
   NOR2xp33_ASAP7_75t_SRAM U23021 (.Y(n15911),
	.A(key_3_),
	.B(FE_OFN26_n16125));
   A2O1A1Ixp33_ASAP7_75t_SL U23023 (.Y(n16142),
	.A1(FE_OFN28470_ld),
	.A2(FE_OCPN29571_n26355),
	.B(n16141),
	.C(FE_OFN25904_n16143));
   NOR2xp33_ASAP7_75t_SRAM U23024 (.Y(n16141),
	.A(key_31_),
	.B(FE_OFN28470_ld));
   OAI21xp33_ASAP7_75t_SRAM U23025 (.Y(n930),
	.A1(ld),
	.A2(n13010),
	.B(rst));
   NAND2xp33_ASAP7_75t_SRAM U23026 (.Y(n19240),
	.A(n26803),
	.B(n27064));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23027 (.Y(n272),
	.A1(n25575),
	.A2(n25475),
	.B(n20021),
	.C(n20020));
   NAND2xp33_ASAP7_75t_SRAM U23028 (.Y(n20021),
	.A(n25471),
	.B(FE_OFN26129_w3_15));
   NAND2xp33_ASAP7_75t_SRAM U23029 (.Y(n18103),
	.A(n26625),
	.B(n25516));
   NAND2xp33_ASAP7_75t_SRAM U23030 (.Y(n23245),
	.A(FE_OCPN29457_n25722),
	.B(n24608));
   NAND2xp33_ASAP7_75t_SRAM U23031 (.Y(n19085),
	.A(n26686),
	.B(n24236));
   NAND2xp33_ASAP7_75t_SRAM U23032 (.Y(n23295),
	.A(n27057),
	.B(n25616));
   NAND2xp33_ASAP7_75t_SRAM U23033 (.Y(n22656),
	.A(n24416),
	.B(n24149));
   NAND2xp33_ASAP7_75t_SRAM U23034 (.Y(n23354),
	.A(FE_OFN29224_FE_OCPN28074_n27049),
	.B(n24495));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23035 (.Y(n280),
	.A1(n23571),
	.A2(FE_OFN16275_n26536),
	.B(n16489),
	.C(n16488));
   NAND2xp33_ASAP7_75t_SRAM U23036 (.Y(n23790),
	.A(FE_OCPN29448_n27189),
	.B(n25247));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23037 (.Y(n283),
	.A1(n26915),
	.A2(n17057),
	.B(n17056),
	.C(n17055));
   NAND2xp33_ASAP7_75t_R U23038 (.Y(n17056),
	.A(n17053),
	.B(n25841));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23039 (.Y(n17055),
	.A1(n26915),
	.A2(n17057),
	.B(n17054),
	.C(w2_22_));
   NAND2xp33_ASAP7_75t_SRAM U23040 (.Y(n17057),
	.A(n25228),
	.B(n17000));
   NAND2xp33_ASAP7_75t_SRAM U23041 (.Y(n19287),
	.A(n25833),
	.B(n26424));
   NAND2xp33_ASAP7_75t_SRAM U23042 (.Y(n19752),
	.A(n25361),
	.B(FE_OFN16276_w3_5));
   NAND2xp33_ASAP7_75t_SRAM U23043 (.Y(n20951),
	.A(n24602),
	.B(n25499));
   NAND2xp33_ASAP7_75t_SRAM U23044 (.Y(n19357),
	.A(n19354),
	.B(n25774));
   NAND2xp33_ASAP7_75t_SRAM U23046 (.Y(n20185),
	.A(FE_OFN25911_n26491),
	.B(n25895));
   NAND2xp33_ASAP7_75t_SRAM U23047 (.Y(n22575),
	.A(FE_OFN104_n27179),
	.B(n26061));
   NAND2xp33_ASAP7_75t_SRAM U23048 (.Y(n22328),
	.A(n26364),
	.B(n26130));
   NAND2xp33_ASAP7_75t_SRAM U23049 (.Y(n19810),
	.A(n19808),
	.B(FE_OFN7_w3_22));
   INVxp33_ASAP7_75t_SRAM U23050 (.Y(n19808),
	.A(n24899));
   NAND2xp33_ASAP7_75t_SRAM U23051 (.Y(n20701),
	.A(FE_OFN28616_n26191),
	.B(n26018));
   NAND2xp33_ASAP7_75t_SRAM U23052 (.Y(n22221),
	.A(n25167),
	.B(n26448));
   NAND2xp33_ASAP7_75t_SRAM U23053 (.Y(n21580),
	.A(n26673),
	.B(n25490));
   NAND2xp33_ASAP7_75t_SRAM U23054 (.Y(n19623),
	.A(FE_OFN29024_n),
	.B(n26375));
   NAND2xp33_ASAP7_75t_SRAM U23055 (.Y(n18665),
	.A(n25251),
	.B(n26811));
   NAND2xp33_ASAP7_75t_SRAM U23056 (.Y(n23850),
	.A(n23848),
	.B(n26951));
   NAND2xp33_ASAP7_75t_R U23058 (.Y(n20611),
	.A(n20608),
	.B(n24435));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23059 (.Y(n299),
	.A1(n26942),
	.A2(n16531),
	.B(n16530),
	.C(n16529));
   NAND2xp33_ASAP7_75t_SRAM U23060 (.Y(n16531),
	.A(n25337),
	.B(n16492));
   NAND2xp33_ASAP7_75t_SRAM U23061 (.Y(n16672),
	.A(n26850),
	.B(FE_OCPN29502_w3_23));
   NAND2xp33_ASAP7_75t_SRAM U23062 (.Y(n23471),
	.A(n24903),
	.B(FE_OFN27209_w3_30));
   NAND2xp33_ASAP7_75t_SRAM U23063 (.Y(n21763),
	.A(FE_OCPN7599_n26721),
	.B(FE_OFN28571_w3_28));
   NAND2xp33_ASAP7_75t_SRAM U23064 (.Y(n20419),
	.A(FE_OCPN29527_n24138),
	.B(n26142));
   NAND2xp33_ASAP7_75t_SRAM U23065 (.Y(n20091),
	.A(FE_OCPN29443_n25507),
	.B(n24200));
   NAND2xp33_ASAP7_75t_SRAM U23066 (.Y(n20357),
	.A(n20355),
	.B(FE_OFN26163_w3_13));
   INVxp33_ASAP7_75t_L U23067 (.Y(n20355),
	.A(FE_OCPN29342_n25357));
   A2O1A1Ixp33_ASAP7_75t_SL U23068 (.Y(n308),
	.A1(n23571),
	.A2(n16746),
	.B(n16745),
	.C(n16744));
   NAND2xp33_ASAP7_75t_SRAM U23069 (.Y(n16745),
	.A(FE_OCPN7656_n24301),
	.B(n26544));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23070 (.Y(n16744),
	.A1(n23571),
	.A2(n16746),
	.B(n16743),
	.C(w0_7_));
   NAND3xp33_ASAP7_75t_SRAM U23071 (.Y(n16746),
	.A(n16683),
	.B(n16682),
	.C(n16681));
   NAND2xp33_ASAP7_75t_SRAM U23072 (.Y(n19396),
	.A(n19393),
	.B(n27195));
   NAND2xp33_ASAP7_75t_SRAM U23073 (.Y(n17183),
	.A(n17180),
	.B(n26656));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23075 (.Y(n313),
	.A1(n26915),
	.A2(n18968),
	.B(n18967),
	.C(n18966));
   NAND2xp33_ASAP7_75t_R U23076 (.Y(n18967),
	.A(n18964),
	.B(FE_OFN70_w2_20));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23077 (.Y(n18966),
	.A1(n26915),
	.A2(n18968),
	.B(n18965),
	.C(w2_20_));
   NAND3xp33_ASAP7_75t_SRAM U23078 (.Y(n18968),
	.A(n25882),
	.B(n18920),
	.C(n25880));
   NAND2xp33_ASAP7_75t_SRAM U23079 (.Y(n17823),
	.A(n27211),
	.B(n26919));
   NAND2xp33_ASAP7_75t_SRAM U23080 (.Y(n19964),
	.A(n24826),
	.B(FE_OCPN29501_FE_OFN28662_w3_7));
   NAND2xp33_ASAP7_75t_SRAM U23081 (.Y(n21339),
	.A(FE_OFN16322_n25946),
	.B(FE_OCPN29428_FE_OFN27131_w3_29));
   NAND2xp33_ASAP7_75t_SRAM U23083 (.Y(n18060),
	.A(FE_OCPN28089_n23913),
	.B(n24470));
   NAND2xp33_ASAP7_75t_SRAM U23084 (.Y(n22915),
	.A(FE_OCPN29470_n24175),
	.B(n26240));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23085 (.Y(n320),
	.A1(n24974),
	.A2(n23058),
	.B(n23057),
	.C(n23056));
   NAND2xp33_ASAP7_75t_SRAM U23086 (.Y(n23057),
	.A(n23054),
	.B(n25961));
   NAND2xp33_ASAP7_75t_SRAM U23087 (.Y(n21191),
	.A(n26631),
	.B(n26385));
   NAND2xp33_ASAP7_75t_SRAM U23088 (.Y(n21498),
	.A(n21496),
	.B(n26645));
   NAND2xp33_ASAP7_75t_SRAM U23090 (.Y(n17313),
	.A(FE_OFN164_n24529),
	.B(n26396));
   NAND2xp33_ASAP7_75t_SRAM U23091 (.Y(n17112),
	.A(n17109),
	.B(n26512));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23092 (.Y(n17111),
	.A1(n26915),
	.A2(n17113),
	.B(n17110),
	.C(w2_19_));
   NAND2xp33_ASAP7_75t_SRAM U23093 (.Y(n21011),
	.A(n21009),
	.B(n25570));
   INVxp33_ASAP7_75t_SRAM U23094 (.Y(n21009),
	.A(FE_OCPN7610_n25861));
   NAND2xp33_ASAP7_75t_R U23095 (.Y(n20221),
	.A(n20218),
	.B(n27106));
   NAND2xp33_ASAP7_75t_SRAM U23096 (.Y(n20222),
	.A(n25504),
	.B(n20193));
   NAND2xp33_ASAP7_75t_SRAM U23097 (.Y(n22120),
	.A(n22118),
	.B(n26760));
   NAND2xp33_ASAP7_75t_SRAM U23098 (.Y(n22121),
	.A(n25915),
	.B(n22072));
   NAND2xp33_ASAP7_75t_SRAM U23099 (.Y(n18297),
	.A(FE_OFN26558_n26911),
	.B(n27219));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23100 (.Y(n331),
	.A1(n26915),
	.A2(n19444),
	.B(n19443),
	.C(n19442));
   NAND2xp33_ASAP7_75t_SRAM U23101 (.Y(n19443),
	.A(n19440),
	.B(n27135));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23102 (.Y(n19442),
	.A1(n26915),
	.A2(n19444),
	.B(n19441),
	.C(w2_17_));
   NAND3xp33_ASAP7_75t_SRAM U23103 (.Y(n19444),
	.A(n19407),
	.B(n19406),
	.C(n25286));
   NAND2xp33_ASAP7_75t_SRAM U23104 (.Y(n20539),
	.A(FE_OCPN27541_n26748),
	.B(n20537));
   INVxp33_ASAP7_75t_SRAM U23105 (.Y(n20537),
	.A(w2_16_));
   NAND2xp33_ASAP7_75t_SRAM U23106 (.Y(n19500),
	.A(n19498),
	.B(FE_OFN25881_w3_24));
   NAND2xp33_ASAP7_75t_SRAM U23107 (.Y(n21533),
	.A(n24841),
	.B(FE_OCPN27659_w3_25));
   NAND2xp33_ASAP7_75t_SRAM U23108 (.Y(n19696),
	.A(n25010),
	.B(FE_OFN28674_n));
   NAND2xp33_ASAP7_75t_SRAM U23109 (.Y(n17234),
	.A(n25041),
	.B(FE_OFN16421_n23974));
   INVxp33_ASAP7_75t_SRAM U23110 (.Y(n21918),
	.A(FE_OFN16432_w3_16));
   NAND2xp33_ASAP7_75t_SRAM U23111 (.Y(n23159),
	.A(n24935),
	.B(FE_OFN28713_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23112 (.Y(n343),
	.A1(n24974),
	.A2(n16607),
	.B(n16606),
	.C(n16605));
   NAND2xp33_ASAP7_75t_SRAM U23113 (.Y(n16606),
	.A(n16603),
	.B(FE_OFN29087_n));
   NAND2xp33_ASAP7_75t_SRAM U23114 (.Y(n19160),
	.A(n24522),
	.B(n24575));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23115 (.Y(n346),
	.A1(n25081),
	.A2(n18403),
	.B(n18402),
	.C(n18401));
   NAND2xp33_ASAP7_75t_SRAM U23116 (.Y(n18402),
	.A(n18400),
	.B(n26692));
   NAND2xp33_ASAP7_75t_SRAM U23117 (.Y(n22174),
	.A(n26580),
	.B(n26185));
   NAND2xp33_ASAP7_75t_SRAM U23118 (.Y(n20489),
	.A(n26179),
	.B(n26991));
   NAND2xp33_ASAP7_75t_SRAM U23119 (.Y(n17520),
	.A(FE_OCPN29503_n24627),
	.B(n24118));
   NAND2xp33_ASAP7_75t_SRAM U23120 (.Y(n19862),
	.A(n24540),
	.B(n26436));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23122 (.Y(n354),
	.A1(n27062),
	.A2(n21391),
	.B(n21390),
	.C(n21389));
   NAND2xp33_ASAP7_75t_SRAM U23123 (.Y(n21390),
	.A(n24714),
	.B(n26221));
   NAND2xp33_ASAP7_75t_R U23124 (.Y(n21391),
	.A(n26071),
	.B(n21348));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23125 (.Y(n356),
	.A1(n27062),
	.A2(FE_OFN171_n26739),
	.B(n22524),
	.C(n22523));
   NAND2xp33_ASAP7_75t_SRAM U23126 (.Y(n22524),
	.A(n26736),
	.B(n26486));
   NAND2xp33_ASAP7_75t_SRAM U23128 (.Y(n21437),
	.A(n26368),
	.B(n26884));
   NAND2xp33_ASAP7_75t_SRAM U23129 (.Y(n23411),
	.A(FE_OFN27075_n23409),
	.B(n24358));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23130 (.Y(n360),
	.A1(n25081),
	.A2(n18520),
	.B(n18519),
	.C(n18518));
   NAND2xp33_ASAP7_75t_R U23131 (.Y(n18519),
	.A(n18516),
	.B(n18515));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23132 (.Y(n361),
	.A1(n26584),
	.A2(n21635),
	.B(n21634),
	.C(n21633));
   NAND2xp33_ASAP7_75t_SRAM U23133 (.Y(n21634),
	.A(n21617),
	.B(n26578));
   A2O1A1Ixp33_ASAP7_75t_R U23134 (.Y(n21633),
	.A1(n26584),
	.A2(n21635),
	.B(n21632),
	.C(w1_3_));
   NOR3xp33_ASAP7_75t_SRAM U23135 (.Y(n21617),
	.A(n21630),
	.B(n21616),
	.C(n25116));
   NAND2xp33_ASAP7_75t_SRAM U23136 (.Y(n18613),
	.A(FE_OFN26019_n26319),
	.B(n26963));
   NAND2xp33_ASAP7_75t_SRAM U23137 (.Y(n23205),
	.A(FE_OFN16263_n25976),
	.B(n24320));
   NAND2xp33_ASAP7_75t_SRAM U23138 (.Y(n20783),
	.A(FE_OFN29011_n27113),
	.B(n27160));
   NAND2xp33_ASAP7_75t_SRAM U23139 (.Y(n21146),
	.A(n21144),
	.B(n24641));
   NAND2xp33_ASAP7_75t_SRAM U23140 (.Y(n22870),
	.A(n26477),
	.B(n26744));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23141 (.Y(n368),
	.A1(n26878),
	.A2(n18240),
	.B(n18239),
	.C(n18238));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23142 (.Y(n18238),
	.A1(n26878),
	.A2(n18240),
	.B(n18237),
	.C(w0_11_));
   NAND2xp33_ASAP7_75t_SRAM U23143 (.Y(n18239),
	.A(n18236),
	.B(n26095));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23144 (.Y(n371),
	.A1(n26323),
	.A2(n21267),
	.B(n21266),
	.C(n21265));
   NAND2xp33_ASAP7_75t_SRAM U23145 (.Y(n21266),
	.A(n21264),
	.B(n27173));
   NAND2xp33_ASAP7_75t_SRAM U23146 (.Y(n21704),
	.A(FE_OFN16324_n25832),
	.B(n26416));
   NAND2xp33_ASAP7_75t_SRAM U23148 (.Y(n23738),
	.A(n27201),
	.B(n25346));
   NAND2xp33_ASAP7_75t_SRAM U23149 (.Y(n18451),
	.A(n26764),
	.B(n24531));
   NAND2xp33_ASAP7_75t_SRAM U23150 (.Y(n17443),
	.A(FE_OFN27172_n17441),
	.B(n25265));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23151 (.Y(n379),
	.A1(n23571),
	.A2(n16974),
	.B(n16973),
	.C(n16972));
   NAND2xp33_ASAP7_75t_SRAM U23152 (.Y(n16973),
	.A(FE_OCPN27637_n26428),
	.B(n16971));
   INVxp33_ASAP7_75t_SRAM U23153 (.Y(n16971),
	.A(w0_0_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23154 (.Y(n380),
	.A1(n23571),
	.A2(FE_OFN28546_n26091),
	.B(n18157),
	.C(n18156));
   NAND2xp33_ASAP7_75t_SRAM U23155 (.Y(n18157),
	.A(n26088),
	.B(n26772));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23156 (.Y(n381),
	.A1(n23571),
	.A2(n23570),
	.B(n23569),
	.C(n23568));
   NAND2xp33_ASAP7_75t_SRAM U23157 (.Y(n23569),
	.A(n26124),
	.B(n25802));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23158 (.Y(n382),
	.A1(n24610),
	.A2(n16907),
	.B(n16906),
	.C(n16905));
   NAND2xp33_ASAP7_75t_SRAM U23159 (.Y(n16906),
	.A(n16903),
	.B(n27129));
   NAND2xp33_ASAP7_75t_SRAM U23160 (.Y(n16907),
	.A(n16849),
	.B(n24336));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23161 (.Y(n384),
	.A1(n26249),
	.A2(n19032),
	.B(n19031),
	.C(n19030));
   NAND2xp33_ASAP7_75t_SRAM U23162 (.Y(n19031),
	.A(n19029),
	.B(n25690));
   NAND3xp33_ASAP7_75t_SRAM U23163 (.Y(n19032),
	.A(n18979),
	.B(FE_OFN27165_n),
	.C(n18978));
   NAND2xp33_ASAP7_75t_SRAM U23164 (.Y(n22963),
	.A(FE_OFN28904_n25733),
	.B(n26041));
   NAND2xp33_ASAP7_75t_SRAM U23165 (.Y(n20285),
	.A(n25698),
	.B(n26932));
   NAND2xp33_ASAP7_75t_SRAM U23167 (.Y(n23010),
	.A(FE_OFN27169_n26683),
	.B(n25411));
   INVxp33_ASAP7_75t_SRAM U23168 (.Y(n18731),
	.A(FE_OCPN7598_n25174));
   NAND2xp33_ASAP7_75t_SRAM U23169 (.Y(n23118),
	.A(FE_OFN25939_n26275),
	.B(FE_OFN66_w1_25));
   NAND2xp33_ASAP7_75t_SRAM U23170 (.Y(n17396),
	.A(n24122),
	.B(n26474));
   NAND2xp33_ASAP7_75t_SRAM U23171 (.Y(n22612),
	.A(FE_OFN29143_n25444),
	.B(n26611));
   NAND2xp33_ASAP7_75t_SRAM U23172 (.Y(n22479),
	.A(FE_OFN28525_n25751),
	.B(n25184));
   NAND2xp33_ASAP7_75t_SRAM U23173 (.Y(n19571),
	.A(n25179),
	.B(n25732));
   NAND2xp33_ASAP7_75t_SRAM U23174 (.Y(n17984),
	.A(FE_OFN16292_n25175),
	.B(n24412));
   NAND2xp33_ASAP7_75t_SRAM U23175 (.Y(n22794),
	.A(n26134),
	.B(n26698));
   NAND2xp33_ASAP7_75t_SRAM U23176 (.Y(n22268),
	.A(n24210),
	.B(n24073));
   NAND2xp33_ASAP7_75t_SRAM U23177 (.Y(n20830),
	.A(n20822),
	.B(n25729));
   NOR2xp33_ASAP7_75t_SRAM U23178 (.Y(n20822),
	.A(n20821),
	.B(n26597));
   OAI21xp33_ASAP7_75t_SRAM U23179 (.Y(n27107),
	.A1(text_in_r_57_),
	.A2(n27106),
	.B(n27105));
   NAND2xp33_ASAP7_75t_SRAM U23180 (.Y(n18348),
	.A(FE_OFN29020_n25146),
	.B(n23937));
   NAND2xp33_ASAP7_75t_SRAM U23182 (.Y(n18857),
	.A(n26836),
	.B(n25596));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23183 (.Y(n415),
	.A1(n25367),
	.A2(FE_OFN16189_n25672),
	.B(n22412),
	.C(n22411));
   NAND2xp33_ASAP7_75t_SRAM U23184 (.Y(n22412),
	.A(n25669),
	.B(FE_OFN25886_w3_3));
   NAND2xp33_ASAP7_75t_SRAM U23186 (.Y(n16830),
	.A(n16828),
	.B(FE_OFN28853_FE_OCPN28408));
   INVxp33_ASAP7_75t_SRAM U23187 (.Y(n16828),
	.A(FE_OCPN29262_n24750));
   NAND2xp33_ASAP7_75t_SRAM U23188 (.Y(n17896),
	.A(n23965),
	.B(n25051));
   NAND2xp33_ASAP7_75t_SRAM U23189 (.Y(n19906),
	.A(n25378),
	.B(FE_OFN25961_w3_8));
   NAND2xp33_ASAP7_75t_SRAM U23190 (.Y(n23676),
	.A(FE_OFN28504_n25956),
	.B(FE_OCPN29520_n24755));
   O2A1O1Ixp5_ASAP7_75t_SL U23191 (.Y(n24850),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27476_n26852),
	.B(n24849),
	.C(n24848));
   NOR2x1_ASAP7_75t_SL U23192 (.Y(n24848),
	.A(n25152),
	.B(n24849));
   NAND2xp33_ASAP7_75t_SRAM U23193 (.Y(n22001),
	.A(n26936),
	.B(n25931));
   NAND2xp33_ASAP7_75t_SRAM U23194 (.Y(n21959),
	.A(n27163),
	.B(n21957));
   INVxp33_ASAP7_75t_SRAM U23195 (.Y(n21957),
	.A(w2_0_));
   NAND2xp33_ASAP7_75t_SRAM U23196 (.Y(n20898),
	.A(n26197),
	.B(n26310));
   NAND2xp33_ASAP7_75t_SRAM U23197 (.Y(n16414),
	.A(n16411),
	.B(n26202));
   NAND2xp33_ASAP7_75t_SRAM U23198 (.Y(n16355),
	.A(n26902),
	.B(n25648));
   NAND3xp33_ASAP7_75t_SL U23199 (.Y(n24687),
	.A(FE_OFN27209_w3_30),
	.B(n24690),
	.C(n24689));
   A2O1A1Ixp33_ASAP7_75t_SL U23200 (.Y(n24690),
	.A1(FE_OCPN27375_n26860),
	.A2(FE_OFN28490_ld_r),
	.B(n24686),
	.C(n24685));
   NAND2xp33_ASAP7_75t_SRAM U23201 (.Y(n24689),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_30_));
   NAND2xp33_ASAP7_75t_SL U23202 (.Y(n26356),
	.A(n26729),
	.B(n26353));
   A2O1A1Ixp33_ASAP7_75t_SL U23203 (.Y(n485),
	.A1(n26647),
	.A2(n26646),
	.B(n26645),
	.C(n26644));
   NAND3xp33_ASAP7_75t_SL U23204 (.Y(n26644),
	.A(n26645),
	.B(n26647),
	.C(n26646));
   NAND2xp33_ASAP7_75t_SRAM U23205 (.Y(n26646),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_126_));
   OAI21xp33_ASAP7_75t_SRAM U23206 (.Y(n24607),
	.A1(text_in_r_87_),
	.A2(n24608),
	.B(FE_OFN12_FE_DBTN0_ld_r));
   NAND2xp5_ASAP7_75t_SL U23207 (.Y(n24604),
	.A(n24603),
	.B(n24605));
   A2O1A1Ixp33_ASAP7_75t_SL U23208 (.Y(n488),
	.A1(n24497),
	.A2(n24496),
	.B(n24495),
	.C(n24494));
   A2O1A1Ixp33_ASAP7_75t_SL U23209 (.Y(n24497),
	.A1(FE_OCPN27379_n26809),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B(n24493),
	.C(n24492));
   NAND2xp33_ASAP7_75t_SRAM U23210 (.Y(n24496),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_110_));
   OAI21xp33_ASAP7_75t_SRAM U23211 (.Y(n24074),
	.A1(text_in_r_86_),
	.A2(n24073),
	.B(n24072));
   OAI22xp33_ASAP7_75t_SRAM U23212 (.Y(n24072),
	.A1(text_in_r_86_),
	.A2(FE_OFN28486_ld_r),
	.B1(n24073),
	.B2(FE_OFN28486_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U23213 (.Y(n490),
	.A1(n25492),
	.A2(n25491),
	.B(n25490),
	.C(n25489));
   NAND3xp33_ASAP7_75t_SL U23214 (.Y(n25489),
	.A(n25490),
	.B(n25492),
	.C(n25491));
   NAND2xp33_ASAP7_75t_SRAM U23215 (.Y(n25491),
	.A(FE_OFN16213_ld_r),
	.B(text_in_r_94_));
   A2O1A1Ixp33_ASAP7_75t_L U23216 (.Y(n493),
	.A1(n26450),
	.A2(n26449),
	.B(n26448),
	.C(n26447));
   NAND2xp5_ASAP7_75t_L U23217 (.Y(n26449),
	.A(n26446),
	.B(n26445));
   A2O1A1Ixp33_ASAP7_75t_SL U23218 (.Y(n495),
	.A1(n26835),
	.A2(n26834),
	.B(n26833),
	.C(n26832));
   OAI21xp5_ASAP7_75t_SL U23219 (.Y(n26833),
	.A1(n26835),
	.A2(n26834),
	.B(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SRAM U23220 (.Y(n26834),
	.A1(n26829),
	.A2(n26828),
	.B(n26827),
	.C(n26826));
   A2O1A1Ixp33_ASAP7_75t_L U23221 (.Y(n501),
	.A1(n26063),
	.A2(n26062),
	.B(n26061),
	.C(n26060));
   NAND3xp33_ASAP7_75t_SL U23222 (.Y(n26060),
	.A(n26061),
	.B(n26063),
	.C(n26062));
   NAND3xp33_ASAP7_75t_R U23223 (.Y(n26062),
	.A(n26059),
	.B(FE_OFN16215_ld_r),
	.C(FE_OCPN29397_n26502));
   A2O1A1Ixp33_ASAP7_75t_SL U23224 (.Y(n502),
	.A1(FE_OCPN27375_n26860),
	.A2(n24666),
	.B(n24665),
	.C(n24664));
   OAI21xp33_ASAP7_75t_SRAM U23225 (.Y(n24664),
	.A1(text_in_r_22_),
	.A2(FE_OFN7_w3_22),
	.B(n24662));
   OAI21xp5_ASAP7_75t_L U23226 (.Y(n24665),
	.A1(n24666),
	.A2(FE_OCPN27375_n26860),
	.B(FE_OFN28489_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U23227 (.Y(n25517),
	.A1(text_in_r_38_),
	.A2(n25516),
	.B(n25515));
   OAI21xp5_ASAP7_75t_SL U23228 (.Y(n25518),
	.A1(n25520),
	.A2(n25519),
	.B(FE_OFN14_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U23229 (.Y(n24914),
	.A1(text_in_r_6_),
	.A2(n24913),
	.B(n24912));
   OAI21xp33_ASAP7_75t_SRAM U23230 (.Y(n27065),
	.A1(text_in_r_119_),
	.A2(n27064),
	.B(n27063));
   NAND2xp33_ASAP7_75t_SRAM U23231 (.Y(n25248),
	.A(FE_OFN13_FE_DBTN0_ld_r),
	.B(text_in_r_46_));
   OAI21xp33_ASAP7_75t_SRAM U23232 (.Y(n25842),
	.A1(text_in_r_54_),
	.A2(n25841),
	.B(n25840));
   OAI21xp33_ASAP7_75t_SL U23233 (.Y(n25843),
	.A1(n25845),
	.A2(n25844),
	.B(FE_OFN16_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_L U23234 (.Y(n24238),
	.A1(n24240),
	.A2(n24239),
	.B(FE_OFN14_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U23235 (.Y(n24235),
	.A1(text_in_r_70_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(n24236),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U23236 (.Y(n516),
	.A1(n27087),
	.A2(n27086),
	.B(n27085),
	.C(n27084));
   NAND3xp33_ASAP7_75t_SL U23237 (.Y(n27084),
	.A(n27085),
	.B(n27087),
	.C(n27086));
   NAND2xp33_ASAP7_75t_SRAM U23238 (.Y(n27086),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_47_));
   A2O1A1Ixp33_ASAP7_75t_SL U23239 (.Y(n520),
	.A1(n25413),
	.A2(n25412),
	.B(n25411),
	.C(n25410));
   NAND3xp33_ASAP7_75t_SL U23240 (.Y(n25410),
	.A(n25411),
	.B(n25413),
	.C(n25412));
   NAND2xp5_ASAP7_75t_R U23241 (.Y(n25412),
	.A(n27031),
	.B(n25409));
   OAI21xp5_ASAP7_75t_L U23242 (.Y(n24508),
	.A1(n24509),
	.A2(FE_OCPN27379_n26809),
	.B(FE_OFN15_FE_DBTN0_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U23243 (.Y(n24507),
	.A1(text_in_r_102_),
	.A2(n24506),
	.B(n24505));
   A2O1A1Ixp33_ASAP7_75t_SL U23244 (.Y(n522),
	.A1(n25481),
	.A2(n25480),
	.B(n25479),
	.C(n25478));
   OAI21xp33_ASAP7_75t_SRAM U23245 (.Y(n25478),
	.A1(text_in_r_7_),
	.A2(FE_OCPN29501_FE_OFN28662_w3_7),
	.B(n25476));
   OAI22xp33_ASAP7_75t_SRAM U23246 (.Y(n26629),
	.A1(w2_7_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_39_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_L U23247 (.Y(n26628),
	.A1(FE_OFN12_FE_DBTN0_ld_r),
	.A2(n27147),
	.B(n26627),
	.C(n26626));
   NOR2x1_ASAP7_75t_SL U23248 (.Y(n26626),
	.A(n27144),
	.B(n26627));
   OAI21xp33_ASAP7_75t_SRAM U23249 (.Y(n26693),
	.A1(text_in_r_71_),
	.A2(n26692),
	.B(n26691));
   A2O1A1Ixp33_ASAP7_75t_SL U23251 (.Y(n525),
	.A1(n26548),
	.A2(n26547),
	.B(n26546),
	.C(n26545));
   OAI21xp33_ASAP7_75t_SRAM U23252 (.Y(n26545),
	.A1(text_in_r_103_),
	.A2(n26544),
	.B(n26543));
   OAI21xp5_ASAP7_75t_SL U23253 (.Y(n26546),
	.A1(n26548),
	.A2(n26547),
	.B(FE_OFN28484_ld_r));
   OAI21xp33_ASAP7_75t_SRAM U23254 (.Y(n527),
	.A1(key_127_),
	.A2(FE_OFN28468_ld),
	.B(n14089));
   NAND2xp33_ASAP7_75t_SRAM U23255 (.Y(n16057),
	.A(n16056),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23257 (.Y(n14606),
	.A(FE_OFN25891_n15770),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23258 (.Y(n15772),
	.A(n16150),
	.B(FE_OFN28463_ld));
   NAND2xp33_ASAP7_75t_SRAM U23259 (.Y(n14249),
	.A(FE_OCPN28327_n15899),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23260 (.Y(n15900),
	.A(n16127),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23261 (.Y(n13866),
	.A(n14974),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23262 (.Y(n14975),
	.A(FE_OCPN8267_n16069),
	.B(FE_OFN28462_ld));
   NAND2xp33_ASAP7_75t_SRAM U23264 (.Y(n14409),
	.A(n14408),
	.B(FE_OFN28467_ld));
   NAND2xp33_ASAP7_75t_R U23266 (.Y(n15905),
	.A(n16197),
	.B(FE_OFN28472_ld));
   NAND2xp33_ASAP7_75t_SRAM U23268 (.Y(n16054),
	.A(n16182),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23269 (.Y(n15897),
	.A(FE_OFN16405_n16117),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23270 (.Y(n16118),
	.A(n16225),
	.B(FE_OFN28464_ld));
   NAND2xp33_ASAP7_75t_SRAM U23271 (.Y(n14184),
	.A(n15774),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23272 (.Y(n15775),
	.A(n16134),
	.B(FE_OFN27_n16125));
   OAI22xp33_ASAP7_75t_SL U23273 (.Y(n550),
	.A1(ld),
	.A2(FE_OFN28538_n16166),
	.B1(key_54_),
	.B2(FE_OFN28538_n16166));
   NAND2xp33_ASAP7_75t_SRAM U23274 (.Y(n14824),
	.A(n16119),
	.B(FE_OFN28468_ld));
   NAND2xp33_ASAP7_75t_R U23275 (.Y(n16121),
	.A(n16120),
	.B(FE_OFN22_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23277 (.Y(n554),
	.A1(key_101_),
	.A2(FE_OFN28472_ld),
	.B(n13334));
   NAND2xp33_ASAP7_75t_SRAM U23278 (.Y(n13334),
	.A(n14004),
	.B(FE_OFN28472_ld));
   NAND2xp33_ASAP7_75t_SRAM U23279 (.Y(n14006),
	.A(n15367),
	.B(FE_OFN28462_ld));
   OAI21xp33_ASAP7_75t_SRAM U23280 (.Y(n557),
	.A1(key_110_),
	.A2(FE_OFN26_n16125),
	.B(n13799));
   NAND2xp33_ASAP7_75t_SRAM U23281 (.Y(n14746),
	.A(n16091),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23282 (.Y(n14003),
	.A(FE_OFN16300_n14826),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23283 (.Y(n14827),
	.A(n16103),
	.B(FE_OFN27_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23285 (.Y(n13938),
	.A(n15906),
	.B(FE_OFN28461_ld));
   NAND2xp33_ASAP7_75t_R U23286 (.Y(n15908),
	.A(n15907),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23288 (.Y(n13635),
	.A(FE_OFN16274_n14664),
	.B(FE_OFN28472_ld));
   NAND2xp33_ASAP7_75t_SRAM U23289 (.Y(n14665),
	.A(n16059),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23290 (.Y(n569),
	.A1(key_108_),
	.A2(FE_OFN28460_ld),
	.B(n14895));
   NAND2xp33_ASAP7_75t_SRAM U23291 (.Y(n14895),
	.A(FE_OFN25929_n16073),
	.B(FE_OFN28460_ld));
   NAND2xp33_ASAP7_75t_SRAM U23292 (.Y(n16074),
	.A(n16179),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23293 (.Y(n572),
	.A1(key_116_),
	.A2(FE_OFN25_n16125),
	.B(n14662));
   NAND2xp33_ASAP7_75t_SRAM U23294 (.Y(n14662),
	.A(n16045),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23295 (.Y(n16046),
	.A(n16213),
	.B(FE_OFN27_n16125));
   INVxp67_ASAP7_75t_L U23296 (.Y(n16214),
	.A(n16231));
   NAND2xp33_ASAP7_75t_SRAM U23297 (.Y(n15365),
	.A(n16135),
	.B(FE_OFN28461_ld));
   NAND2xp33_ASAP7_75t_SRAM U23298 (.Y(n16137),
	.A(n16136),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23300 (.Y(n13410),
	.A(n14007),
	.B(FE_OFN28471_ld));
   NAND2xp33_ASAP7_75t_SRAM U23302 (.Y(n15060),
	.A(n16088),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23303 (.Y(n16089),
	.A(n16219),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23305 (.Y(n15470),
	.A(FE_PSN8277_n16099),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23306 (.Y(n16101),
	.A(n16243),
	.B(FE_OFN27_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23307 (.Y(n14329),
	.A(n16065),
	.B(FE_OFN28468_ld));
   NAND2xp33_ASAP7_75t_R U23308 (.Y(n16067),
	.A(n16066),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23310 (.Y(n13480),
	.A(FE_OFN16240_n14011),
	.B(FE_OFN28471_ld));
   NAND2xp33_ASAP7_75t_SRAM U23311 (.Y(n14012),
	.A(n15371),
	.B(FE_OFN28463_ld));
   NAND2xp33_ASAP7_75t_SRAM U23312 (.Y(n15657),
	.A(FE_OCPN28186_n16123),
	.B(FE_OFN26_n16125));
   OAI21xp33_ASAP7_75t_L U23313 (.Y(n594),
	.A1(key_72_),
	.A2(FE_OFN25_n16125),
	.B(n16124));
   NAND2xp33_ASAP7_75t_SRAM U23314 (.Y(n14972),
	.A(FE_OCPN8223_n16063),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23315 (.Y(n16064),
	.A(n16175),
	.B(FE_OFN27_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23316 (.Y(n599),
	.A1(key_120_),
	.A2(FE_OFN28468_ld),
	.B(n15565));
   NAND2xp33_ASAP7_75t_SRAM U23317 (.Y(n15565),
	.A(n16163),
	.B(FE_OFN28468_ld));
   NAND2xp33_ASAP7_75t_R U23318 (.Y(n16165),
	.A(n16164),
	.B(FE_OFN19_n16125));
   OAI22xp5_ASAP7_75t_SL U23320 (.Y(n601),
	.A1(ld),
	.A2(FE_OFN25882_n16262),
	.B1(key_56_),
	.B2(FE_OFN25882_n16262));
   NAND2xp33_ASAP7_75t_SRAM U23321 (.Y(n13549),
	.A(n14090),
	.B(FE_OFN28471_ld));
   NAND2xp33_ASAP7_75t_R U23322 (.Y(n14092),
	.A(n15910),
	.B(FE_OFN28463_ld));
   NAND2xp33_ASAP7_75t_SRAM U23324 (.Y(n15143),
	.A(FE_OCPN29581_n16097),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SL U23325 (.Y(n16098),
	.A(n16194),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23327 (.Y(n16049),
	.A(FE_OCPN8248_n16145),
	.B(FE_OFN28462_ld));
   NAND2xp33_ASAP7_75t_SRAM U23328 (.Y(n15769),
	.A(n16138),
	.B(FE_OFN28468_ld));
   NAND2xp33_ASAP7_75t_SRAM U23329 (.Y(n16140),
	.A(n16139),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U23331 (.Y(n13724),
	.A(FE_OFN25971_n14472),
	.B(FE_OFN28472_ld));
   INVx1_ASAP7_75t_SL U23333 (.Y(n16083),
	.A(n16086));
   OAI21xp33_ASAP7_75t_SRAM U23334 (.Y(n617),
	.A1(key_105_),
	.A2(FE_OFN28460_ld),
	.B(n14471));
   NAND2xp33_ASAP7_75t_SRAM U23335 (.Y(n14471),
	.A(FE_OCPN29468_n15919),
	.B(FE_OFN28460_ld));
   NAND2xp33_ASAP7_75t_SRAM U23336 (.Y(n15920),
	.A(n16199),
	.B(FE_OFN28462_ld));
   NAND2xp33_ASAP7_75t_SRAM U23337 (.Y(n16043),
	.A(n16076),
	.B(FE_OFN28462_ld));
   NAND2xp33_ASAP7_75t_R U23338 (.Y(n16077),
	.A(FE_OFN26549_n16248),
	.B(FE_OFN28462_ld));
   A2O1A1Ixp33_ASAP7_75t_SL U23339 (.Y(n16085),
	.A1(n25596),
	.A2(FE_OFN26139_n16125),
	.B(n16084),
	.C(n16086));
   NOR2xp33_ASAP7_75t_SRAM U23340 (.Y(n16084),
	.A(key_0_),
	.B(FE_OFN26139_n16125));
   OAI21xp33_ASAP7_75t_SL U23341 (.Y(n630),
	.A1(FE_OFN16370_n16261),
	.A2(FE_OFN16159_w3_24),
	.B(n16260));
   NOR2xp33_ASAP7_75t_SRAM U23342 (.Y(n16259),
	.A(key_24_),
	.B(FE_OFN28470_ld));
   OAI21xp33_ASAP7_75t_SL U23343 (.Y(n632),
	.A1(n16271),
	.A2(FE_OFN25961_w3_8),
	.B(n16270));
   NOR2xp33_ASAP7_75t_SRAM U23344 (.Y(n16269),
	.A(key_8_),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SL U23345 (.Y(n644),
	.A1(n16094),
	.A2(FE_PSN8297_FE_OFN8_w3_14),
	.B(n16093));
   NOR2xp33_ASAP7_75t_SRAM U23346 (.Y(n16092),
	.A(key_14_),
	.B(FE_OFN25_n16125));
   NAND2xp5_ASAP7_75t_SL U23347 (.Y(n647),
	.A(n16171),
	.B(n16170));
   NAND2xp5_ASAP7_75t_SL U23348 (.Y(n16170),
	.A(FE_PSN8299_FE_OFN4_w3_22),
	.B(FE_OFN28538_n16166));
   NOR2xp33_ASAP7_75t_SRAM U23349 (.Y(n16167),
	.A(ld),
	.B(FE_PSN8299_FE_OFN4_w3_22));
   OAI21xp33_ASAP7_75t_L U23350 (.Y(n16279),
	.A1(n16275),
	.A2(n16274),
	.B(n16273));
   NOR2xp33_ASAP7_75t_SRAM U23351 (.Y(n16274),
	.A(FE_OFN21_n16125),
	.B(FE_OFN28699_w3_6));
   NAND2xp33_ASAP7_75t_SRAM U23352 (.Y(n659),
	.A(n16282),
	.B(n13273));
   OAI22xp33_ASAP7_75t_SRAM U23353 (.Y(n662),
	.A1(u0_r0_rcnt_2_),
	.A2(ld),
	.B1(n16285),
	.B2(ld));
   NAND2xp33_ASAP7_75t_SRAM U23354 (.Y(n663),
	.A(n13271),
	.B(FE_OFN28461_ld));
   NAND2xp33_ASAP7_75t_SRAM U23355 (.Y(n666),
	.A(FE_OFN28461_ld),
	.B(n16286));
   NAND2xp33_ASAP7_75t_SRAM U23356 (.Y(n13258),
	.A(n13257),
	.B(FE_OFN28469_ld));
   NAND2xp33_ASAP7_75t_SRAM U23357 (.Y(n13256),
	.A(n13255),
	.B(FE_OFN28470_ld));
   NAND2xp33_ASAP7_75t_SRAM U23358 (.Y(n13238),
	.A(FE_OFN28470_ld),
	.B(n13237));
   INVxp33_ASAP7_75t_SRAM U23359 (.Y(n13237),
	.A(text_in_r_2_));
   OAI21xp33_ASAP7_75t_SRAM U23360 (.Y(n673),
	.A1(text_in_3_),
	.A2(FE_OFN28470_ld),
	.B(n13158));
   NAND2xp33_ASAP7_75t_SRAM U23361 (.Y(n13158),
	.A(n13157),
	.B(FE_OFN28470_ld));
   INVxp33_ASAP7_75t_SRAM U23362 (.Y(n13157),
	.A(text_in_r_3_));
   OAI21xp33_ASAP7_75t_SRAM U23363 (.Y(n675),
	.A1(text_in_4_),
	.A2(FE_OFN28470_ld),
	.B(n13160));
   NAND2xp33_ASAP7_75t_SRAM U23364 (.Y(n13160),
	.A(n13159),
	.B(FE_OFN28470_ld));
   OAI21xp33_ASAP7_75t_SRAM U23365 (.Y(n677),
	.A1(text_in_5_),
	.A2(FE_OFN28470_ld),
	.B(n13230));
   NAND2xp33_ASAP7_75t_SRAM U23366 (.Y(n13230),
	.A(FE_OFN28470_ld),
	.B(n13229));
   INVxp33_ASAP7_75t_SRAM U23367 (.Y(n13229),
	.A(text_in_r_5_));
   OAI21xp33_ASAP7_75t_SRAM U23368 (.Y(n679),
	.A1(text_in_6_),
	.A2(FE_OFN28469_ld),
	.B(n13232));
   OAI21xp33_ASAP7_75t_SRAM U23369 (.Y(n681),
	.A1(text_in_7_),
	.A2(FE_OFN26139_n16125),
	.B(n13228));
   NAND2xp33_ASAP7_75t_SRAM U23370 (.Y(n13228),
	.A(FE_OFN26139_n16125),
	.B(n13227));
   OAI21xp33_ASAP7_75t_SRAM U23371 (.Y(n683),
	.A1(text_in_8_),
	.A2(FE_OFN28457_ld),
	.B(n13162));
   NAND2xp33_ASAP7_75t_SRAM U23372 (.Y(n13162),
	.A(n13161),
	.B(FE_OFN28457_ld));
   INVxp33_ASAP7_75t_SRAM U23373 (.Y(n13161),
	.A(text_in_r_8_));
   NAND2xp33_ASAP7_75t_SRAM U23374 (.Y(n13150),
	.A(FE_OFN28457_ld),
	.B(n13149));
   INVxp33_ASAP7_75t_SRAM U23375 (.Y(n13149),
	.A(text_in_r_9_));
   NAND2xp33_ASAP7_75t_SRAM U23376 (.Y(n13156),
	.A(n13155),
	.B(FE_OFN28457_ld));
   NAND2xp33_ASAP7_75t_SRAM U23377 (.Y(n13152),
	.A(FE_OFN28457_ld),
	.B(n13151));
   INVxp33_ASAP7_75t_SRAM U23378 (.Y(n13151),
	.A(text_in_r_11_));
   NAND2xp33_ASAP7_75t_SRAM U23379 (.Y(n13146),
	.A(FE_OFN28457_ld),
	.B(n13145));
   NAND2xp33_ASAP7_75t_SRAM U23380 (.Y(n13154),
	.A(FE_OFN28457_ld),
	.B(n13153));
   INVxp33_ASAP7_75t_SRAM U23381 (.Y(n13153),
	.A(text_in_r_14_));
   NAND2xp33_ASAP7_75t_SRAM U23382 (.Y(n13148),
	.A(FE_OFN28457_ld),
	.B(n13147));
   INVxp33_ASAP7_75t_SRAM U23383 (.Y(n13147),
	.A(text_in_r_15_));
   OAI21xp33_ASAP7_75t_SRAM U23384 (.Y(n699),
	.A1(text_in_16_),
	.A2(FE_OFN26139_n16125),
	.B(n13234));
   NAND2xp33_ASAP7_75t_SRAM U23385 (.Y(n13234),
	.A(n13233),
	.B(FE_OFN26139_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23386 (.Y(n701),
	.A1(text_in_17_),
	.A2(FE_OFN26139_n16125),
	.B(n13242));
   NAND2xp33_ASAP7_75t_SRAM U23387 (.Y(n13242),
	.A(n13241),
	.B(FE_OFN26139_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23388 (.Y(n703),
	.A1(text_in_18_),
	.A2(FE_OFN28469_ld),
	.B(n13070));
   NAND2xp33_ASAP7_75t_SRAM U23389 (.Y(n13070),
	.A(FE_OFN28469_ld),
	.B(n13069));
   INVxp33_ASAP7_75t_SRAM U23390 (.Y(n13069),
	.A(text_in_r_18_));
   OAI21xp33_ASAP7_75t_SRAM U23391 (.Y(n705),
	.A1(text_in_19_),
	.A2(FE_OFN28470_ld),
	.B(n13224));
   NAND2xp33_ASAP7_75t_SRAM U23392 (.Y(n13224),
	.A(n13223),
	.B(FE_OFN28470_ld));
   OAI21xp33_ASAP7_75t_SRAM U23393 (.Y(n707),
	.A1(text_in_20_),
	.A2(FE_OFN26139_n16125),
	.B(n13200));
   OAI21xp33_ASAP7_75t_SRAM U23394 (.Y(n709),
	.A1(text_in_21_),
	.A2(FE_OFN28457_ld),
	.B(n13044));
   NAND2xp33_ASAP7_75t_SRAM U23395 (.Y(n13044),
	.A(FE_OFN28457_ld),
	.B(n13043));
   OAI21xp33_ASAP7_75t_SRAM U23396 (.Y(n711),
	.A1(text_in_22_),
	.A2(FE_OFN28470_ld),
	.B(n13046));
   NAND2xp33_ASAP7_75t_SRAM U23397 (.Y(n13046),
	.A(FE_OFN28470_ld),
	.B(n13045));
   INVxp33_ASAP7_75t_SRAM U23398 (.Y(n13045),
	.A(text_in_r_22_));
   OAI21xp33_ASAP7_75t_SRAM U23399 (.Y(n713),
	.A1(text_in_23_),
	.A2(FE_OFN26139_n16125),
	.B(n13038));
   NAND2xp33_ASAP7_75t_SRAM U23400 (.Y(n13038),
	.A(FE_OFN26139_n16125),
	.B(n13037));
   INVxp33_ASAP7_75t_SRAM U23401 (.Y(n13037),
	.A(text_in_r_23_));
   OAI21xp33_ASAP7_75t_SRAM U23402 (.Y(n715),
	.A1(text_in_24_),
	.A2(FE_OFN28469_ld),
	.B(n13184));
   NAND2xp33_ASAP7_75t_SRAM U23403 (.Y(n13184),
	.A(n13183),
	.B(FE_OFN28469_ld));
   OAI21xp33_ASAP7_75t_SRAM U23404 (.Y(n717),
	.A1(text_in_25_),
	.A2(FE_OFN28469_ld),
	.B(n13036));
   NAND2xp33_ASAP7_75t_SRAM U23405 (.Y(n13036),
	.A(FE_OFN28469_ld),
	.B(n13035));
   INVxp33_ASAP7_75t_SRAM U23406 (.Y(n13035),
	.A(text_in_r_25_));
   OAI21xp33_ASAP7_75t_SRAM U23407 (.Y(n719),
	.A1(text_in_26_),
	.A2(FE_OFN28469_ld),
	.B(n13192));
   NAND2xp33_ASAP7_75t_SRAM U23408 (.Y(n13192),
	.A(n13191),
	.B(FE_OFN28469_ld));
   OAI21xp33_ASAP7_75t_SRAM U23409 (.Y(n721),
	.A1(text_in_27_),
	.A2(FE_OFN28470_ld),
	.B(n13042));
   NAND2xp33_ASAP7_75t_SRAM U23410 (.Y(n13042),
	.A(FE_OFN28470_ld),
	.B(n13041));
   INVxp33_ASAP7_75t_SRAM U23411 (.Y(n13039),
	.A(text_in_r_28_));
   OAI21xp33_ASAP7_75t_SRAM U23412 (.Y(n725),
	.A1(text_in_29_),
	.A2(FE_OFN28469_ld),
	.B(n13186));
   NAND2xp33_ASAP7_75t_SRAM U23413 (.Y(n13186),
	.A(n13185),
	.B(FE_OFN28469_ld));
   INVxp33_ASAP7_75t_SRAM U23414 (.Y(n13185),
	.A(text_in_r_29_));
   OAI21xp33_ASAP7_75t_SRAM U23415 (.Y(n727),
	.A1(text_in_30_),
	.A2(FE_OFN28470_ld),
	.B(n13064));
   NAND2xp33_ASAP7_75t_SRAM U23416 (.Y(n13064),
	.A(FE_OFN28470_ld),
	.B(n13063));
   INVxp33_ASAP7_75t_SRAM U23417 (.Y(n13063),
	.A(text_in_r_30_));
   OAI21xp33_ASAP7_75t_SRAM U23418 (.Y(n729),
	.A1(text_in_31_),
	.A2(FE_OFN28469_ld),
	.B(n13066));
   NAND2xp33_ASAP7_75t_SRAM U23419 (.Y(n13066),
	.A(FE_OFN28469_ld),
	.B(n13065));
   INVxp33_ASAP7_75t_SRAM U23420 (.Y(n13065),
	.A(text_in_r_31_));
   OAI21xp33_ASAP7_75t_SRAM U23421 (.Y(n731),
	.A1(text_in_32_),
	.A2(FE_OFN22_n16125),
	.B(n13196));
   NAND2xp33_ASAP7_75t_SRAM U23422 (.Y(n13196),
	.A(n13195),
	.B(FE_OFN22_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23423 (.Y(n733),
	.A1(text_in_33_),
	.A2(FE_OFN22_n16125),
	.B(n13218));
   NAND2xp33_ASAP7_75t_SRAM U23424 (.Y(n13218),
	.A(n13217),
	.B(FE_OFN22_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23425 (.Y(n735),
	.A1(text_in_34_),
	.A2(FE_OFN22_n16125),
	.B(n13068));
   NAND2xp33_ASAP7_75t_SRAM U23426 (.Y(n13068),
	.A(FE_OFN22_n16125),
	.B(n13067));
   OAI21xp33_ASAP7_75t_SRAM U23427 (.Y(n737),
	.A1(text_in_35_),
	.A2(FE_OFN22_n16125),
	.B(n13208));
   OAI21xp33_ASAP7_75t_SRAM U23428 (.Y(n739),
	.A1(text_in_36_),
	.A2(FE_OFN22_n16125),
	.B(n13240));
   NAND2xp33_ASAP7_75t_SRAM U23429 (.Y(n13240),
	.A(n13239),
	.B(FE_OFN22_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23430 (.Y(n741),
	.A1(text_in_37_),
	.A2(FE_OFN19_n16125),
	.B(n13048));
   NAND2xp33_ASAP7_75t_SRAM U23431 (.Y(n13048),
	.A(FE_OFN19_n16125),
	.B(n13047));
   INVxp33_ASAP7_75t_SRAM U23432 (.Y(n13047),
	.A(text_in_r_37_));
   OAI21xp33_ASAP7_75t_SRAM U23433 (.Y(n743),
	.A1(text_in_38_),
	.A2(FE_OFN22_n16125),
	.B(n13050));
   NAND2xp33_ASAP7_75t_SRAM U23434 (.Y(n13050),
	.A(FE_OFN22_n16125),
	.B(n13049));
   OAI21xp33_ASAP7_75t_SRAM U23435 (.Y(n745),
	.A1(text_in_39_),
	.A2(FE_OFN28458_ld),
	.B(n13052));
   NAND2xp33_ASAP7_75t_SRAM U23436 (.Y(n13052),
	.A(FE_OFN28458_ld),
	.B(n13051));
   OAI21xp33_ASAP7_75t_SRAM U23437 (.Y(n747),
	.A1(text_in_40_),
	.A2(FE_OFN19_n16125),
	.B(n13262));
   NAND2xp33_ASAP7_75t_SRAM U23438 (.Y(n13262),
	.A(n13261),
	.B(FE_OFN19_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23439 (.Y(n749),
	.A1(text_in_41_),
	.A2(FE_OFN22_n16125),
	.B(n13054));
   NAND2xp33_ASAP7_75t_SRAM U23440 (.Y(n13054),
	.A(FE_OFN22_n16125),
	.B(n13053));
   INVxp33_ASAP7_75t_SRAM U23441 (.Y(n13053),
	.A(text_in_r_41_));
   OAI21xp33_ASAP7_75t_SRAM U23442 (.Y(n751),
	.A1(text_in_42_),
	.A2(FE_OFN19_n16125),
	.B(n13264));
   NAND2xp33_ASAP7_75t_SRAM U23443 (.Y(n13264),
	.A(n13263),
	.B(FE_OFN19_n16125));
   INVxp33_ASAP7_75t_SRAM U23444 (.Y(n13055),
	.A(text_in_r_43_));
   OAI21xp33_ASAP7_75t_SRAM U23445 (.Y(n755),
	.A1(text_in_44_),
	.A2(FE_OFN22_n16125),
	.B(n13058));
   NAND2xp33_ASAP7_75t_SRAM U23446 (.Y(n13058),
	.A(FE_OFN22_n16125),
	.B(n13057));
   INVxp33_ASAP7_75t_SRAM U23447 (.Y(n13057),
	.A(text_in_r_44_));
   OAI21xp33_ASAP7_75t_SRAM U23448 (.Y(n757),
	.A1(text_in_45_),
	.A2(FE_OFN19_n16125),
	.B(n13194));
   NAND2xp33_ASAP7_75t_SRAM U23449 (.Y(n13194),
	.A(n13193),
	.B(FE_OFN19_n16125));
   INVxp33_ASAP7_75t_SRAM U23450 (.Y(n13193),
	.A(text_in_r_45_));
   OAI21xp33_ASAP7_75t_SRAM U23451 (.Y(n759),
	.A1(text_in_46_),
	.A2(FE_OFN22_n16125),
	.B(n13060));
   NAND2xp33_ASAP7_75t_SRAM U23452 (.Y(n13060),
	.A(FE_OFN22_n16125),
	.B(n13059));
   INVxp33_ASAP7_75t_SRAM U23453 (.Y(n13059),
	.A(text_in_r_46_));
   OAI21xp33_ASAP7_75t_SRAM U23454 (.Y(n761),
	.A1(text_in_47_),
	.A2(FE_OFN22_n16125),
	.B(n13188));
   NAND2xp33_ASAP7_75t_SRAM U23455 (.Y(n13188),
	.A(n13187),
	.B(FE_OFN22_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23456 (.Y(n763),
	.A1(text_in_48_),
	.A2(FE_OFN28458_ld),
	.B(n13206));
   NAND2xp33_ASAP7_75t_SRAM U23457 (.Y(n13206),
	.A(n13205),
	.B(FE_OFN28458_ld));
   OAI21xp33_ASAP7_75t_SRAM U23458 (.Y(n765),
	.A1(text_in_49_),
	.A2(FE_OFN28458_ld),
	.B(n13226));
   NAND2xp33_ASAP7_75t_SRAM U23459 (.Y(n13226),
	.A(n13225),
	.B(FE_OFN28458_ld));
   OAI21xp33_ASAP7_75t_SRAM U23460 (.Y(n767),
	.A1(text_in_50_),
	.A2(FE_OFN28459_ld),
	.B(n13062));
   OAI21xp33_ASAP7_75t_SRAM U23461 (.Y(n769),
	.A1(text_in_51_),
	.A2(FE_OFN28458_ld),
	.B(n13222));
   NAND2xp33_ASAP7_75t_SRAM U23462 (.Y(n13222),
	.A(n13221),
	.B(FE_OFN28458_ld));
   INVxp33_ASAP7_75t_SRAM U23463 (.Y(n13221),
	.A(text_in_r_51_));
   OAI21xp33_ASAP7_75t_SRAM U23464 (.Y(n771),
	.A1(text_in_52_),
	.A2(FE_OFN28458_ld),
	.B(n13210));
   NAND2xp33_ASAP7_75t_SRAM U23465 (.Y(n13210),
	.A(n13209),
	.B(FE_OFN28458_ld));
   OAI21xp33_ASAP7_75t_SRAM U23466 (.Y(n773),
	.A1(text_in_53_),
	.A2(FE_OFN28458_ld),
	.B(n13190));
   NAND2xp33_ASAP7_75t_SRAM U23467 (.Y(n13190),
	.A(n13189),
	.B(FE_OFN28458_ld));
   OAI21xp33_ASAP7_75t_SRAM U23468 (.Y(n775),
	.A1(text_in_54_),
	.A2(FE_OFN28458_ld),
	.B(n13072));
   NAND2xp33_ASAP7_75t_SRAM U23469 (.Y(n13072),
	.A(FE_OFN28459_ld),
	.B(n13071));
   OAI21xp33_ASAP7_75t_SRAM U23470 (.Y(n777),
	.A1(text_in_55_),
	.A2(FE_OFN19_n16125),
	.B(n13074));
   NAND2xp33_ASAP7_75t_SRAM U23471 (.Y(n13074),
	.A(FE_OFN19_n16125),
	.B(n13073));
   OAI21xp33_ASAP7_75t_SRAM U23472 (.Y(n779),
	.A1(text_in_56_),
	.A2(FE_OFN28459_ld),
	.B(n13212));
   NAND2xp33_ASAP7_75t_SRAM U23473 (.Y(n13212),
	.A(n13211),
	.B(FE_OFN28459_ld));
   OAI21xp33_ASAP7_75t_SRAM U23474 (.Y(n781),
	.A1(text_in_57_),
	.A2(FE_OFN28459_ld),
	.B(n13076));
   NAND2xp33_ASAP7_75t_SRAM U23475 (.Y(n13076),
	.A(FE_OFN28459_ld),
	.B(n13075));
   INVxp33_ASAP7_75t_SRAM U23476 (.Y(n13075),
	.A(text_in_r_57_));
   INVxp33_ASAP7_75t_SRAM U23477 (.Y(n13077),
	.A(text_in_r_58_));
   OAI21xp33_ASAP7_75t_SRAM U23478 (.Y(n785),
	.A1(text_in_59_),
	.A2(FE_OFN28459_ld),
	.B(n13080));
   NAND2xp33_ASAP7_75t_SRAM U23479 (.Y(n13080),
	.A(FE_OFN28459_ld),
	.B(n13079));
   INVxp33_ASAP7_75t_SRAM U23480 (.Y(n13079),
	.A(text_in_r_59_));
   OAI21xp33_ASAP7_75t_SRAM U23481 (.Y(n787),
	.A1(text_in_60_),
	.A2(FE_OFN28459_ld),
	.B(n13082));
   NAND2xp33_ASAP7_75t_SRAM U23482 (.Y(n13082),
	.A(FE_OFN28459_ld),
	.B(n13081));
   INVxp33_ASAP7_75t_SRAM U23483 (.Y(n13081),
	.A(text_in_r_60_));
   OAI21xp33_ASAP7_75t_SRAM U23484 (.Y(n789),
	.A1(text_in_61_),
	.A2(FE_OFN28459_ld),
	.B(n13182));
   NAND2xp33_ASAP7_75t_SRAM U23485 (.Y(n13182),
	.A(n13181),
	.B(FE_OFN28459_ld));
   OAI21xp33_ASAP7_75t_SRAM U23486 (.Y(n791),
	.A1(text_in_62_),
	.A2(FE_OFN28459_ld),
	.B(n13174));
   NAND2xp33_ASAP7_75t_SRAM U23487 (.Y(n13174),
	.A(n13173),
	.B(FE_OFN28459_ld));
   INVxp33_ASAP7_75t_SRAM U23488 (.Y(n13173),
	.A(text_in_r_62_));
   OAI21xp33_ASAP7_75t_SRAM U23489 (.Y(n793),
	.A1(text_in_63_),
	.A2(FE_OFN28459_ld),
	.B(n13084));
   NAND2xp33_ASAP7_75t_SRAM U23490 (.Y(n13084),
	.A(FE_OFN28459_ld),
	.B(n13083));
   INVxp33_ASAP7_75t_SRAM U23491 (.Y(n13083),
	.A(text_in_r_63_));
   OAI21xp33_ASAP7_75t_SRAM U23492 (.Y(n795),
	.A1(text_in_64_),
	.A2(FE_OFN28462_ld),
	.B(n13214));
   NAND2xp33_ASAP7_75t_SRAM U23493 (.Y(n13214),
	.A(n13213),
	.B(FE_OFN28462_ld));
   INVxp33_ASAP7_75t_SRAM U23494 (.Y(n13213),
	.A(text_in_r_64_));
   OAI21xp33_ASAP7_75t_SRAM U23495 (.Y(n797),
	.A1(text_in_65_),
	.A2(FE_OFN28463_ld),
	.B(n13202));
   OAI21xp33_ASAP7_75t_SRAM U23496 (.Y(n799),
	.A1(text_in_66_),
	.A2(FE_OFN25_n16125),
	.B(n13086));
   NAND2xp33_ASAP7_75t_SRAM U23497 (.Y(n13086),
	.A(FE_OFN25_n16125),
	.B(n13085));
   OAI21xp33_ASAP7_75t_SRAM U23498 (.Y(n801),
	.A1(text_in_67_),
	.A2(FE_OFN28463_ld),
	.B(n13088));
   NAND2xp33_ASAP7_75t_SRAM U23499 (.Y(n13088),
	.A(FE_OFN28463_ld),
	.B(n13087));
   INVxp33_ASAP7_75t_SRAM U23500 (.Y(n13087),
	.A(text_in_r_67_));
   OAI21xp33_ASAP7_75t_SRAM U23501 (.Y(n803),
	.A1(text_in_68_),
	.A2(FE_OFN25_n16125),
	.B(n13254));
   NAND2xp33_ASAP7_75t_SRAM U23502 (.Y(n13254),
	.A(n13253),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23503 (.Y(n805),
	.A1(text_in_69_),
	.A2(FE_OFN27_n16125),
	.B(n13090));
   NAND2xp33_ASAP7_75t_SRAM U23504 (.Y(n13090),
	.A(FE_OFN27_n16125),
	.B(n13089));
   INVxp33_ASAP7_75t_SRAM U23505 (.Y(n13089),
	.A(text_in_r_69_));
   OAI21xp33_ASAP7_75t_SRAM U23506 (.Y(n807),
	.A1(text_in_70_),
	.A2(FE_OFN28463_ld),
	.B(n13092));
   NAND2xp33_ASAP7_75t_SRAM U23507 (.Y(n13092),
	.A(FE_OFN28463_ld),
	.B(n13091));
   INVxp33_ASAP7_75t_SRAM U23508 (.Y(n13091),
	.A(text_in_r_70_));
   OAI21xp33_ASAP7_75t_SRAM U23509 (.Y(n809),
	.A1(text_in_71_),
	.A2(FE_OFN28463_ld),
	.B(n13094));
   NAND2xp33_ASAP7_75t_SRAM U23510 (.Y(n13094),
	.A(FE_OFN28463_ld),
	.B(n13093));
   INVxp33_ASAP7_75t_SRAM U23511 (.Y(n13093),
	.A(text_in_r_71_));
   OAI21xp33_ASAP7_75t_SRAM U23512 (.Y(n811),
	.A1(text_in_72_),
	.A2(FE_OFN28457_ld),
	.B(n13096));
   NAND2xp33_ASAP7_75t_SRAM U23513 (.Y(n13096),
	.A(FE_OFN28457_ld),
	.B(n13095));
   INVxp33_ASAP7_75t_SRAM U23514 (.Y(n13097),
	.A(text_in_r_73_));
   OAI21xp33_ASAP7_75t_SRAM U23515 (.Y(n815),
	.A1(text_in_74_),
	.A2(FE_OFN28457_ld),
	.B(n13102));
   NAND2xp33_ASAP7_75t_SRAM U23516 (.Y(n13102),
	.A(FE_OFN28457_ld),
	.B(n13101));
   OAI21xp33_ASAP7_75t_SRAM U23517 (.Y(n817),
	.A1(text_in_75_),
	.A2(FE_OFN28457_ld),
	.B(n13104));
   NAND2xp33_ASAP7_75t_SRAM U23518 (.Y(n13104),
	.A(FE_OFN28457_ld),
	.B(n13103));
   OAI21xp33_ASAP7_75t_SRAM U23519 (.Y(n819),
	.A1(text_in_76_),
	.A2(FE_OFN28464_ld),
	.B(n13106));
   NAND2xp33_ASAP7_75t_SRAM U23520 (.Y(n13106),
	.A(FE_OFN28464_ld),
	.B(n13105));
   INVxp33_ASAP7_75t_SRAM U23521 (.Y(n13105),
	.A(text_in_r_76_));
   OAI21xp33_ASAP7_75t_SRAM U23522 (.Y(n821),
	.A1(text_in_77_),
	.A2(FE_OFN28457_ld),
	.B(n13108));
   NAND2xp33_ASAP7_75t_SRAM U23523 (.Y(n13108),
	.A(FE_OFN28457_ld),
	.B(n13107));
   INVxp33_ASAP7_75t_SRAM U23524 (.Y(n13107),
	.A(text_in_r_77_));
   OAI21xp33_ASAP7_75t_SRAM U23525 (.Y(n823),
	.A1(text_in_78_),
	.A2(FE_OFN28457_ld),
	.B(n13176));
   NAND2xp33_ASAP7_75t_SRAM U23526 (.Y(n13176),
	.A(n13175),
	.B(FE_OFN28457_ld));
   OAI21xp33_ASAP7_75t_SRAM U23527 (.Y(n825),
	.A1(text_in_79_),
	.A2(FE_OFN28464_ld),
	.B(n13114));
   NAND2xp33_ASAP7_75t_SRAM U23528 (.Y(n13114),
	.A(FE_OFN28464_ld),
	.B(n13113));
   INVxp33_ASAP7_75t_SRAM U23529 (.Y(n13113),
	.A(text_in_r_79_));
   OAI21xp33_ASAP7_75t_SRAM U23530 (.Y(n827),
	.A1(text_in_80_),
	.A2(FE_OFN28464_ld),
	.B(n13178));
   OAI21xp33_ASAP7_75t_SRAM U23531 (.Y(n829),
	.A1(text_in_81_),
	.A2(FE_OFN27_n16125),
	.B(n13126));
   NAND2xp33_ASAP7_75t_SRAM U23532 (.Y(n13126),
	.A(FE_OFN27_n16125),
	.B(n13125));
   INVxp33_ASAP7_75t_SRAM U23533 (.Y(n13125),
	.A(text_in_r_81_));
   OAI21xp33_ASAP7_75t_SRAM U23534 (.Y(n831),
	.A1(text_in_82_),
	.A2(FE_OFN27_n16125),
	.B(n13110));
   NAND2xp33_ASAP7_75t_SRAM U23535 (.Y(n13110),
	.A(FE_OFN27_n16125),
	.B(n13109));
   INVxp33_ASAP7_75t_SRAM U23536 (.Y(n13109),
	.A(text_in_r_82_));
   OAI21xp33_ASAP7_75t_SRAM U23537 (.Y(n833),
	.A1(text_in_83_),
	.A2(FE_OFN28464_ld),
	.B(n13216));
   NAND2xp33_ASAP7_75t_SRAM U23538 (.Y(n13216),
	.A(n13215),
	.B(FE_OFN28464_ld));
   OAI21xp33_ASAP7_75t_SRAM U23539 (.Y(n835),
	.A1(text_in_84_),
	.A2(FE_OFN28464_ld),
	.B(n13124));
   NAND2xp33_ASAP7_75t_SRAM U23540 (.Y(n13124),
	.A(FE_OFN28464_ld),
	.B(n13123));
   OAI21xp33_ASAP7_75t_SRAM U23541 (.Y(n837),
	.A1(text_in_85_),
	.A2(FE_OFN27_n16125),
	.B(n13136));
   NAND2xp33_ASAP7_75t_SRAM U23542 (.Y(n13136),
	.A(FE_OFN27_n16125),
	.B(n13135));
   INVxp33_ASAP7_75t_SRAM U23543 (.Y(n13135),
	.A(text_in_r_85_));
   OAI21xp33_ASAP7_75t_SRAM U23544 (.Y(n839),
	.A1(text_in_86_),
	.A2(FE_OFN28464_ld),
	.B(n13138));
   NAND2xp33_ASAP7_75t_SRAM U23545 (.Y(n13138),
	.A(FE_OFN28464_ld),
	.B(n13137));
   INVxp33_ASAP7_75t_SRAM U23546 (.Y(n13137),
	.A(text_in_r_86_));
   OAI21xp33_ASAP7_75t_SRAM U23547 (.Y(n841),
	.A1(text_in_87_),
	.A2(FE_OFN27_n16125),
	.B(n13128));
   NAND2xp33_ASAP7_75t_SRAM U23548 (.Y(n13128),
	.A(FE_OFN27_n16125),
	.B(n13127));
   INVxp33_ASAP7_75t_SRAM U23549 (.Y(n13127),
	.A(text_in_r_87_));
   OAI21xp33_ASAP7_75t_SRAM U23550 (.Y(n845),
	.A1(text_in_89_),
	.A2(FE_OFN27_n16125),
	.B(n13018));
   NAND2xp33_ASAP7_75t_SRAM U23551 (.Y(n13018),
	.A(FE_OFN27_n16125),
	.B(n13017));
   OAI21xp33_ASAP7_75t_SRAM U23552 (.Y(n847),
	.A1(text_in_90_),
	.A2(FE_OFN27_n16125),
	.B(n13022));
   NAND2xp33_ASAP7_75t_SRAM U23553 (.Y(n13022),
	.A(FE_OFN27_n16125),
	.B(n13021));
   OAI21xp33_ASAP7_75t_SRAM U23554 (.Y(n849),
	.A1(text_in_91_),
	.A2(FE_OFN27_n16125),
	.B(n13030));
   NAND2xp33_ASAP7_75t_SRAM U23555 (.Y(n13030),
	.A(FE_OFN27_n16125),
	.B(n13029));
   OAI21xp33_ASAP7_75t_SRAM U23556 (.Y(n851),
	.A1(text_in_92_),
	.A2(FE_OFN27_n16125),
	.B(n13100));
   NAND2xp33_ASAP7_75t_SRAM U23557 (.Y(n13100),
	.A(FE_OFN27_n16125),
	.B(n13099));
   INVxp33_ASAP7_75t_SRAM U23558 (.Y(n13099),
	.A(text_in_r_92_));
   OAI21xp33_ASAP7_75t_SRAM U23559 (.Y(n853),
	.A1(text_in_93_),
	.A2(FE_OFN27_n16125),
	.B(n13204));
   NAND2xp33_ASAP7_75t_SRAM U23560 (.Y(n13204),
	.A(n13203),
	.B(FE_OFN27_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23561 (.Y(n855),
	.A1(text_in_94_),
	.A2(FE_OFN27_n16125),
	.B(n13120));
   NAND2xp33_ASAP7_75t_SRAM U23562 (.Y(n13120),
	.A(FE_OFN27_n16125),
	.B(n13119));
   OAI21xp33_ASAP7_75t_SRAM U23563 (.Y(n857),
	.A1(text_in_95_),
	.A2(FE_OFN28457_ld),
	.B(n13180));
   OAI21xp33_ASAP7_75t_SRAM U23564 (.Y(n859),
	.A1(text_in_96_),
	.A2(FE_OFN28471_ld),
	.B(n13248));
   NAND2xp33_ASAP7_75t_SRAM U23565 (.Y(n13248),
	.A(n13247),
	.B(FE_OFN28471_ld));
   OAI21xp33_ASAP7_75t_SRAM U23566 (.Y(n861),
	.A1(text_in_97_),
	.A2(FE_OFN28471_ld),
	.B(n13250));
   NAND2xp33_ASAP7_75t_SRAM U23567 (.Y(n13250),
	.A(n13249),
	.B(FE_OFN28471_ld));
   OAI21xp33_ASAP7_75t_SRAM U23568 (.Y(n863),
	.A1(text_in_98_),
	.A2(FE_OFN28471_ld),
	.B(n13172));
   NAND2xp33_ASAP7_75t_SRAM U23569 (.Y(n13172),
	.A(FE_OFN28471_ld),
	.B(n13171));
   INVxp33_ASAP7_75t_SRAM U23570 (.Y(n13171),
	.A(text_in_r_98_));
   OAI21xp33_ASAP7_75t_SRAM U23571 (.Y(n865),
	.A1(text_in_99_),
	.A2(FE_OFN28471_ld),
	.B(n13164));
   NAND2xp33_ASAP7_75t_SRAM U23572 (.Y(n13164),
	.A(FE_OFN28471_ld),
	.B(n13163));
   INVxp33_ASAP7_75t_SRAM U23573 (.Y(n13163),
	.A(text_in_r_99_));
   OAI21xp33_ASAP7_75t_SRAM U23574 (.Y(n867),
	.A1(text_in_100_),
	.A2(FE_OFN28471_ld),
	.B(n13252));
   NAND2xp33_ASAP7_75t_SRAM U23575 (.Y(n13252),
	.A(n13251),
	.B(FE_OFN28471_ld));
   OAI21xp33_ASAP7_75t_SRAM U23576 (.Y(n869),
	.A1(text_in_101_),
	.A2(FE_OFN28471_ld),
	.B(n13170));
   NAND2xp33_ASAP7_75t_SRAM U23577 (.Y(n13170),
	.A(FE_OFN28471_ld),
	.B(n13169));
   OAI21xp33_ASAP7_75t_SRAM U23578 (.Y(n871),
	.A1(text_in_102_),
	.A2(FE_OFN28471_ld),
	.B(n13166));
   NAND2xp33_ASAP7_75t_SRAM U23579 (.Y(n13166),
	.A(FE_OFN28471_ld),
	.B(n13165));
   INVxp33_ASAP7_75t_SRAM U23580 (.Y(n13165),
	.A(text_in_r_102_));
   INVxp33_ASAP7_75t_SRAM U23581 (.Y(n13111),
	.A(text_in_r_103_));
   OAI21xp33_ASAP7_75t_SRAM U23582 (.Y(n875),
	.A1(text_in_104_),
	.A2(FE_OFN20_n16125),
	.B(n13116));
   NAND2xp33_ASAP7_75t_SRAM U23583 (.Y(n13116),
	.A(FE_OFN20_n16125),
	.B(n13115));
   OAI21xp33_ASAP7_75t_SRAM U23584 (.Y(n877),
	.A1(text_in_105_),
	.A2(FE_OFN28460_ld),
	.B(n13012));
   NAND2xp33_ASAP7_75t_SRAM U23585 (.Y(n13012),
	.A(FE_OFN28460_ld),
	.B(n13011));
   OAI21xp33_ASAP7_75t_SRAM U23586 (.Y(n879),
	.A1(text_in_106_),
	.A2(FE_OFN20_n16125),
	.B(n13028));
   NAND2xp33_ASAP7_75t_SRAM U23587 (.Y(n13028),
	.A(FE_OFN20_n16125),
	.B(n13027));
   OAI21xp33_ASAP7_75t_SRAM U23588 (.Y(n881),
	.A1(text_in_107_),
	.A2(FE_OFN28461_ld),
	.B(n13032));
   NAND2xp33_ASAP7_75t_SRAM U23589 (.Y(n13032),
	.A(FE_OFN28461_ld),
	.B(n13031));
   OAI21xp33_ASAP7_75t_SRAM U23590 (.Y(n883),
	.A1(text_in_108_),
	.A2(FE_OFN28471_ld),
	.B(n13026));
   NAND2xp33_ASAP7_75t_SRAM U23591 (.Y(n13026),
	.A(FE_OFN28471_ld),
	.B(n13025));
   OAI21xp33_ASAP7_75t_SRAM U23592 (.Y(n885),
	.A1(text_in_109_),
	.A2(FE_OFN20_n16125),
	.B(n13246));
   NAND2xp33_ASAP7_75t_SRAM U23593 (.Y(n13246),
	.A(n13245),
	.B(FE_OFN20_n16125));
   OAI21xp33_ASAP7_75t_SRAM U23594 (.Y(n887),
	.A1(text_in_110_),
	.A2(FE_OFN28460_ld),
	.B(n13140));
   OAI21xp33_ASAP7_75t_SRAM U23595 (.Y(n889),
	.A1(text_in_111_),
	.A2(FE_OFN28460_ld),
	.B(n13168));
   NAND2xp33_ASAP7_75t_SRAM U23596 (.Y(n13168),
	.A(FE_OFN28460_ld),
	.B(n13167));
   OAI21xp33_ASAP7_75t_SRAM U23597 (.Y(n891),
	.A1(text_in_112_),
	.A2(FE_OFN28471_ld),
	.B(n13122));
   NAND2xp33_ASAP7_75t_SRAM U23598 (.Y(n13122),
	.A(FE_OFN28471_ld),
	.B(n13121));
   INVxp33_ASAP7_75t_SRAM U23599 (.Y(n13121),
	.A(text_in_r_112_));
   OAI21xp33_ASAP7_75t_SRAM U23600 (.Y(n893),
	.A1(text_in_113_),
	.A2(FE_OFN28472_ld),
	.B(n13244));
   NAND2xp33_ASAP7_75t_SRAM U23601 (.Y(n13244),
	.A(n13243),
	.B(FE_OFN28472_ld));
   OAI21xp33_ASAP7_75t_SRAM U23602 (.Y(n895),
	.A1(text_in_114_),
	.A2(FE_OFN28471_ld),
	.B(n13130));
   NAND2xp33_ASAP7_75t_SRAM U23603 (.Y(n13130),
	.A(FE_OFN28471_ld),
	.B(n13129));
   INVxp33_ASAP7_75t_SRAM U23604 (.Y(n13129),
	.A(text_in_r_114_));
   OAI21xp33_ASAP7_75t_SRAM U23605 (.Y(n897),
	.A1(text_in_115_),
	.A2(FE_OFN28472_ld),
	.B(n13220));
   NAND2xp33_ASAP7_75t_SRAM U23606 (.Y(n13220),
	.A(n13219),
	.B(FE_OFN28472_ld));
   OAI21xp33_ASAP7_75t_SRAM U23607 (.Y(n899),
	.A1(text_in_116_),
	.A2(FE_OFN28472_ld),
	.B(n13198));
   NAND2xp33_ASAP7_75t_SRAM U23608 (.Y(n13198),
	.A(n13197),
	.B(FE_OFN28472_ld));
   OAI21xp33_ASAP7_75t_SRAM U23609 (.Y(n901),
	.A1(text_in_117_),
	.A2(FE_OFN28460_ld),
	.B(n13144));
   NAND2xp33_ASAP7_75t_SRAM U23610 (.Y(n13144),
	.A(FE_OFN28460_ld),
	.B(n13143));
   INVxp33_ASAP7_75t_SRAM U23611 (.Y(n13143),
	.A(text_in_r_117_));
   INVxp33_ASAP7_75t_SRAM U23612 (.Y(n13117),
	.A(text_in_r_118_));
   OAI21xp33_ASAP7_75t_SRAM U23613 (.Y(n905),
	.A1(text_in_119_),
	.A2(FE_OFN28460_ld),
	.B(n13016));
   NAND2xp33_ASAP7_75t_SRAM U23614 (.Y(n13016),
	.A(FE_OFN28460_ld),
	.B(n13015));
   OAI21xp33_ASAP7_75t_SRAM U23615 (.Y(n907),
	.A1(text_in_120_),
	.A2(FE_OFN28467_ld),
	.B(n13260));
   NAND2xp33_ASAP7_75t_SRAM U23616 (.Y(n13260),
	.A(n13259),
	.B(FE_OFN28467_ld));
   OAI21xp33_ASAP7_75t_SRAM U23617 (.Y(n909),
	.A1(text_in_121_),
	.A2(FE_OFN28467_ld),
	.B(n13142));
   NAND2xp33_ASAP7_75t_SRAM U23618 (.Y(n13142),
	.A(FE_OFN28467_ld),
	.B(n13141));
   INVxp33_ASAP7_75t_SRAM U23619 (.Y(n13141),
	.A(text_in_r_121_));
   OAI21xp33_ASAP7_75t_SRAM U23620 (.Y(n911),
	.A1(text_in_122_),
	.A2(FE_OFN28467_ld),
	.B(n13134));
   NAND2xp33_ASAP7_75t_SRAM U23621 (.Y(n13134),
	.A(FE_OFN28467_ld),
	.B(n13133));
   INVxp33_ASAP7_75t_SRAM U23622 (.Y(n13133),
	.A(text_in_r_122_));
   OAI21xp33_ASAP7_75t_SRAM U23623 (.Y(n913),
	.A1(text_in_123_),
	.A2(FE_OFN28467_ld),
	.B(n13014));
   NAND2xp33_ASAP7_75t_SRAM U23624 (.Y(n13014),
	.A(FE_OFN28467_ld),
	.B(n13013));
   OAI21xp33_ASAP7_75t_SRAM U23625 (.Y(n915),
	.A1(text_in_124_),
	.A2(FE_OFN28468_ld),
	.B(n13132));
   NAND2xp33_ASAP7_75t_SRAM U23626 (.Y(n13132),
	.A(FE_OFN28468_ld),
	.B(n13131));
   OAI21xp33_ASAP7_75t_SRAM U23627 (.Y(n917),
	.A1(text_in_125_),
	.A2(FE_OFN28467_ld),
	.B(n13266));
   OAI21xp33_ASAP7_75t_SRAM U23628 (.Y(n919),
	.A1(text_in_126_),
	.A2(FE_OFN28467_ld),
	.B(n13020));
   NAND2xp33_ASAP7_75t_SRAM U23629 (.Y(n13020),
	.A(FE_OFN28467_ld),
	.B(n13019));
   NAND2xp33_ASAP7_75t_SRAM U23630 (.Y(n13034),
	.A(FE_OFN28468_ld),
	.B(n13033));
   INVxp33_ASAP7_75t_SRAM U23631 (.Y(n13033),
	.A(text_in_r_127_));
   OAI21xp33_ASAP7_75t_SRAM U23632 (.Y(n924),
	.A1(ld),
	.A2(n13009),
	.B(rst));
   NAND2xp33_ASAP7_75t_SRAM U23633 (.Y(n926),
	.A(rst),
	.B(n13001));
   OAI21xp33_ASAP7_75t_SRAM U23634 (.Y(n928),
	.A1(ld),
	.A2(n13004),
	.B(rst));
   O2A1O1Ixp5_ASAP7_75t_SL U23635 (.Y(n26422),
	.A1(FE_OFN116_n27187),
	.A2(n27186),
	.B(FE_OCPN7589_n26420),
	.C(n26419));
   NAND2xp5_ASAP7_75t_L U23636 (.Y(n24305),
	.A(FE_OCPN29390_n26528),
	.B(FE_OCPN27333_n25250));
   NAND2xp33_ASAP7_75t_R U23637 (.Y(n25969),
	.A(FE_OCPN29390_n26528),
	.B(n25966));
   OAI21xp5_ASAP7_75t_SL U23639 (.Y(n26642),
	.A1(FE_OFN2_ld_r),
	.A2(FE_OFN16329_n27151),
	.B(n26643));
   NOR2x1_ASAP7_75t_SL U23640 (.Y(n20876),
	.A(n16290),
	.B(n20853));
   A2O1A1Ixp33_ASAP7_75t_SL U23641 (.Y(n26837),
	.A1(n17580),
	.A2(n24830),
	.B(n24276),
	.C(n24275));
   OAI21xp5_ASAP7_75t_SL U23642 (.Y(n24322),
	.A1(n24323),
	.A2(FE_OCPN27310_n26389),
	.B(FE_OFN28483_ld_r));
   NOR2xp33_ASAP7_75t_SL U23644 (.Y(n19119),
	.A(sa00_0_),
	.B(sa00_1_));
   OAI21xp33_ASAP7_75t_SRAM U23645 (.Y(n15574),
	.A1(n15567),
	.A2(n13725),
	.B(n15566));
   OAI21xp5_ASAP7_75t_SL U23647 (.Y(n27082),
	.A1(FE_OFN1_ld_r),
	.A2(n27110),
	.B(n27083));
   OAI21xp5_ASAP7_75t_SL U23648 (.Y(n17750),
	.A1(n17791),
	.A2(FE_OCPN27838_n17747),
	.B(n20142));
   NOR2x1p5_ASAP7_75t_SL U23650 (.Y(n16980),
	.A(FE_OFN28478_sa13_2),
	.B(n19360));
   NOR2x2_ASAP7_75t_SL U23651 (.Y(n17445),
	.A(FE_OFN29137_FE_OCPN27228_sa11_2),
	.B(n17501));
   NOR2x1p5_ASAP7_75t_SL U23652 (.Y(n20617),
	.A(FE_OCPN29430_FE_OFN31_sa20_0),
	.B(n18582));
   NOR2x2_ASAP7_75t_SL U23653 (.Y(n17446),
	.A(FE_OFN28874_FE_OCPN27551_sa11_4),
	.B(n17494));
   NOR2x1_ASAP7_75t_SL U23654 (.Y(n16422),
	.A(FE_OFN29134_sa33_0),
	.B(FE_OFN28727_sa33_1));
   NAND2x1p5_ASAP7_75t_SL U23655 (.Y(n17318),
	.A(FE_OCPN29429_FE_OFN16141_sa01_3),
	.B(n17317));
   NOR2x2_ASAP7_75t_SL U23656 (.Y(n17447),
	.A(FE_OFN28874_FE_OCPN27551_sa11_4),
	.B(n21355));
   NOR2x1p5_ASAP7_75t_SL U23657 (.Y(n18540),
	.A(FE_OCPN27580_n),
	.B(n18602));
   NOR2x1p5_ASAP7_75t_L U23664 (.Y(n18970),
	.A(FE_OFN29189_sa23_0),
	.B(FE_OCPN27627_sa23_1));
   NOR2x1p5_ASAP7_75t_SL U23665 (.Y(n17906),
	.A(FE_OCPN29453_sa12_4),
	.B(FE_OFN73_sa12_5));
   NOR2x1p5_ASAP7_75t_SL U23666 (.Y(n18177),
	.A(FE_OFN16135_sa22_4),
	.B(n21123));
   NOR2x1_ASAP7_75t_SL U23667 (.Y(n16747),
	.A(FE_OFN28698_sa21_1),
	.B(FE_OCPN29418_n));
   NOR2x1p5_ASAP7_75t_SL U23668 (.Y(n17525),
	.A(FE_OFN27148_sa32_3),
	.B(n17679));
   NAND2x1_ASAP7_75t_SL U23669 (.Y(n16290),
	.A(FE_OFN28719_n20025),
	.B(n20028));
   NOR2x1p5_ASAP7_75t_SL U23672 (.Y(n17331),
	.A(FE_OCPN27423_sa01_0),
	.B(FE_OFN28718_sa01_1));
   NOR2x1_ASAP7_75t_SL U23673 (.Y(n16758),
	.A(FE_OCPN27328_sa21_2),
	.B(FE_OCPN27554_n20007));
   NOR2x1p5_ASAP7_75t_SL U23674 (.Y(n16757),
	.A(FE_OCPN27328_sa21_2),
	.B(n17843));
   NAND2x2_ASAP7_75t_SL U23675 (.Y(n16533),
	.A(FE_OFN28751_n),
	.B(n17216));
   NAND2x1p5_ASAP7_75t_L U23676 (.Y(n13890),
	.A(FE_OFN16426_w3_20),
	.B(n15485));
   NAND2x1_ASAP7_75t_SL U23677 (.Y(n14289),
	.A(FE_OFN16426_w3_20),
	.B(n15667));
   NOR2xp33_ASAP7_75t_SL U23679 (.Y(n25213),
	.A(n22872),
	.B(n22095));
   NOR2x1_ASAP7_75t_L U23680 (.Y(n17899),
	.A(FE_OCPN27888_sa12_2),
	.B(FE_OFN29225_sa12_0));
   NOR2x1p5_ASAP7_75t_SL U23681 (.Y(n13804),
	.A(FE_OFN26642_w3_14),
	.B(n15987));
   NOR2xp33_ASAP7_75t_SL U23682 (.Y(n16749),
	.A(n16783),
	.B(n20289));
   NOR2x1_ASAP7_75t_L U23683 (.Y(n17900),
	.A(FE_OCPN27888_sa12_2),
	.B(n17923));
   INVxp67_ASAP7_75t_SL U23686 (.Y(n14354),
	.A(n15719));
   NOR2x1_ASAP7_75t_SL U23687 (.Y(n18527),
	.A(FE_OFN29251_n18536),
	.B(n23689));
   OAI21xp5_ASAP7_75t_L U23688 (.Y(n14579),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OCPN27656_w3_25),
	.B(FE_OFN27207_w3_30));
   NOR2x1p5_ASAP7_75t_L U23689 (.Y(n17329),
	.A(FE_OFN16141_sa01_3),
	.B(n25054));
   NOR2x1_ASAP7_75t_L U23691 (.Y(n18597),
	.A(FE_OFN29250_FE_OCPN27371_sa20_2),
	.B(n23819));
   NOR2x1p5_ASAP7_75t_SL U23695 (.Y(n17321),
	.A(FE_OFN28736_FE_OCPN28216_sa01_5),
	.B(n18684));
   NOR2x1_ASAP7_75t_L U23696 (.Y(n17317),
	.A(FE_OCPN28217_sa01_5),
	.B(n17326));
   NOR2x1p5_ASAP7_75t_SL U23697 (.Y(n17603),
	.A(FE_OCPN28049_sa30_0),
	.B(FE_OFN16247_sa30_1));
   NOR2x2_ASAP7_75t_SL U23699 (.Y(n18161),
	.A(n23308),
	.B(n18169));
   NOR2x1p5_ASAP7_75t_SL U23703 (.Y(n17521),
	.A(FE_OFN28686_FE_OCPN27812),
	.B(FE_OFN26035_n));
   NOR2x1_ASAP7_75t_L U23706 (.Y(n16977),
	.A(FE_OFN16444_sa13_1),
	.B(n16982));
   NOR2x1p5_ASAP7_75t_SL U23707 (.Y(n16748),
	.A(FE_OFN28903_sa21_0),
	.B(n17881));
   NAND2x2_ASAP7_75t_SL U23708 (.Y(n17236),
	.A(FE_OCPN27908_FE_OFN16156_sa00_2),
	.B(FE_OCPN29474_n19119));
   INVx1_ASAP7_75t_SL U23710 (.Y(n14559),
	.A(n14579));
   NAND2xp33_ASAP7_75t_SRAM U23711 (.Y(n14574),
	.A(n14573),
	.B(n14572));
   NAND2xp5_ASAP7_75t_R U23712 (.Y(n14560),
	.A(FE_OFN16206_n15240),
	.B(n14559));
   INVxp67_ASAP7_75t_L U23713 (.Y(n14042),
	.A(n13875));
   NOR2xp33_ASAP7_75t_SL U23714 (.Y(n17803),
	.A(n17761),
	.B(n22533));
   NAND2xp33_ASAP7_75t_R U23715 (.Y(n14548),
	.A(n14544),
	.B(n15224));
   NAND2xp33_ASAP7_75t_L U23716 (.Y(n14122),
	.A(n14117),
	.B(n14119));
   NAND2xp33_ASAP7_75t_R U23717 (.Y(n15330),
	.A(n15329),
	.B(FE_OFN28600_n14289));
   NAND2xp33_ASAP7_75t_SL U23718 (.Y(n13687),
	.A(n13683),
	.B(n13684));
   OAI21xp5_ASAP7_75t_SL U23719 (.Y(n16455),
	.A1(n16418),
	.A2(n16853),
	.B(FE_OFN16430_sa33_3));
   NAND2xp5_ASAP7_75t_L U23721 (.Y(n14380),
	.A(n14379),
	.B(n14378));
   NAND2xp33_ASAP7_75t_SL U23722 (.Y(n14162),
	.A(n14161),
	.B(n14160));
   NAND2xp33_ASAP7_75t_SRAM U23724 (.Y(n13588),
	.A(n14534),
	.B(FE_OFN25966_n13646));
   OAI21xp5_ASAP7_75t_L U23726 (.Y(n14298),
	.A1(n12994),
	.A2(n14398),
	.B(n14297));
   AND2x2_ASAP7_75t_L U23728 (.Y(n26067),
	.A(n26065),
	.B(n26064));
   NOR2xp33_ASAP7_75t_SRAM U23729 (.Y(n21321),
	.A(n21708),
	.B(n21502));
   NAND2xp33_ASAP7_75t_SRAM U23730 (.Y(n14385),
	.A(n14384),
	.B(n14383));
   INVxp33_ASAP7_75t_SRAM U23731 (.Y(n14330),
	.A(n14766));
   NAND2xp33_ASAP7_75t_SRAM U23732 (.Y(n14132),
	.A(n14138),
	.B(n15954));
   NAND2xp33_ASAP7_75t_L U23733 (.Y(n13388),
	.A(n13385),
	.B(n13386));
   NAND2xp33_ASAP7_75t_L U23734 (.Y(n13457),
	.A(n13456),
	.B(n13455));
   NAND2xp33_ASAP7_75t_R U23735 (.Y(n15499),
	.A(n15498),
	.B(n15497));
   OAI22xp33_ASAP7_75t_SRAM U23736 (.Y(n13637),
	.A1(FE_OCPN27656_w3_25),
	.A2(FE_PSN8307_FE_OFN27207_w3_30),
	.B1(FE_OFN26051_w3_27),
	.B2(FE_PSN8307_FE_OFN27207_w3_30));
   NOR2xp33_ASAP7_75t_SRAM U23737 (.Y(n24782),
	.A(n24780),
	.B(n24779));
   NOR2xp33_ASAP7_75t_SL U23738 (.Y(n16656),
	.A(n16542),
	.B(n23133));
   NOR2xp33_ASAP7_75t_L U23740 (.Y(n20686),
	.A(n20685),
	.B(n23792));
   NAND2xp33_ASAP7_75t_SL U23741 (.Y(n20031),
	.A(n20030),
	.B(FE_OFN25972_n20056));
   NAND2xp33_ASAP7_75t_L U23742 (.Y(n14134),
	.A(n14132),
	.B(n14131));
   AND3x1_ASAP7_75t_R U23743 (.Y(n13779),
	.A(n15575),
	.B(n15099),
	.C(n15585));
   NOR2x1_ASAP7_75t_SL U23744 (.Y(n14377),
	.A(FE_OFN6_w3_22),
	.B(FE_OFN26053_n25415));
   NAND2xp5_ASAP7_75t_L U23745 (.Y(n15187),
	.A(FE_OFN28452_w3_29),
	.B(FE_OFN27130_w3_28));
   NAND2xp33_ASAP7_75t_L U23746 (.Y(n15282),
	.A(n15281),
	.B(n15694));
   OR3x1_ASAP7_75t_SRAM U23748 (.Y(n15439),
	.A(n15435),
	.B(n15434),
	.C(FE_OFN28542_n15433));
   NOR3xp33_ASAP7_75t_SRAM U23749 (.Y(n14271),
	.A(FE_OFN28623_n13874),
	.B(FE_OCPN27987_FE_OFN4_w3_22),
	.C(FE_OCPN8264_n13890));
   NAND2xp33_ASAP7_75t_SRAM U23750 (.Y(n14953),
	.A(n14939),
	.B(n14938));
   NOR2xp33_ASAP7_75t_SRAM U23751 (.Y(n15472),
	.A(FE_OFN26535_w3_19),
	.B(FE_OFN28909_w3_23));
   OAI22xp33_ASAP7_75t_SRAM U23752 (.Y(n15617),
	.A1(FE_OFN28721_n),
	.A2(FE_OCPN27978_w3_3),
	.B1(FE_OFN28732_n),
	.B2(FE_OCPN27978_w3_3));
   OR2x2_ASAP7_75t_R U23753 (.Y(n14720),
	.A(n14929),
	.B(n14719));
   NAND2xp33_ASAP7_75t_R U23754 (.Y(n15706),
	.A(FE_OFN26538_w3_19),
	.B(n15719));
   NAND2xp33_ASAP7_75t_L U23755 (.Y(n24783),
	.A(n24782),
	.B(FE_OFN16326_n19058));
   NOR2xp33_ASAP7_75t_SRAM U23756 (.Y(n23953),
	.A(FE_OCPN27900_n23949),
	.B(n23948));
   NAND2xp33_ASAP7_75t_L U23757 (.Y(n24260),
	.A(n24255),
	.B(n24883));
   NOR2xp33_ASAP7_75t_L U23758 (.Y(n17005),
	.A(n16978),
	.B(n24155));
   NAND2xp33_ASAP7_75t_SRAM U23760 (.Y(n18573),
	.A(FE_OFN29140_n18527),
	.B(FE_OFN27083_n));
   NOR2xp33_ASAP7_75t_SL U23761 (.Y(n18554),
	.A(n18526),
	.B(FE_OCPN27532_n21643));
   NAND2xp5_ASAP7_75t_L U23762 (.Y(n17533),
	.A(n17528),
	.B(n17530));
   AND3x2_ASAP7_75t_SL U23764 (.Y(n16461),
	.A(n16459),
	.B(FE_OCPN29561_n23532),
	.C(n16458));
   O2A1O1Ixp33_ASAP7_75t_SRAM U23765 (.Y(n13499),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OFN28859_FE_OCPN27664_w3_25),
	.B(FE_OFN27212_w3_30),
	.C(n15155));
   NAND2xp33_ASAP7_75t_SRAM U23766 (.Y(n15824),
	.A(n15823),
	.B(n15834));
   OAI22xp5_ASAP7_75t_L U23767 (.Y(n15433),
	.A1(FE_OCPN28407_FE_OFN16433_w3_11),
	.A2(FE_OFN26639_w3_14),
	.B1(FE_OCPN29506_FE_OFN16184_w3_9),
	.B2(FE_OFN26639_w3_14));
   NAND2xp33_ASAP7_75t_R U23768 (.Y(n14752),
	.A(n14751),
	.B(n14750));
   NAND2xp33_ASAP7_75t_L U23769 (.Y(n13781),
	.A(n13780),
	.B(n13779));
   NAND2xp33_ASAP7_75t_L U23770 (.Y(n13988),
	.A(n13987),
	.B(n13986));
   NAND2xp5_ASAP7_75t_SL U23771 (.Y(n13926),
	.A(n13923),
	.B(n13922));
   NAND2xp33_ASAP7_75t_SL U23774 (.Y(n14923),
	.A(n14922),
	.B(n14921));
   NAND2xp33_ASAP7_75t_SL U23775 (.Y(n14433),
	.A(n14432),
	.B(n14431));
   NOR3xp33_ASAP7_75t_SL U23776 (.Y(n17029),
	.A(n19374),
	.B(FE_OCPN27589_n25987),
	.C(n18930));
   NAND2xp33_ASAP7_75t_SL U23777 (.Y(n23606),
	.A(n23605),
	.B(n23604));
   NOR2xp33_ASAP7_75t_R U23778 (.Y(n27005),
	.A(n27001),
	.B(n27000));
   NAND2xp33_ASAP7_75t_SRAM U23779 (.Y(n24129),
	.A(n24785),
	.B(n24127));
   NOR2xp33_ASAP7_75t_SL U23780 (.Y(n19230),
	.A(n17444),
	.B(n23402));
   AND3x1_ASAP7_75t_R U23781 (.Y(n23768),
	.A(n23767),
	.B(n23766),
	.C(n23765));
   OAI22xp33_ASAP7_75t_SRAM U23782 (.Y(n19304),
	.A1(FE_OFN29003_n23491),
	.A2(n19301),
	.B1(n19019),
	.B2(n19301));
   NOR2xp33_ASAP7_75t_SRAM U23783 (.Y(n22209),
	.A(FE_OCPN27871_n17317),
	.B(n22597));
   NAND2xp33_ASAP7_75t_SRAM U23784 (.Y(n23801),
	.A(FE_OFN28776_n18532),
	.B(n18540));
   NOR3xp33_ASAP7_75t_SRAM U23785 (.Y(n23500),
	.A(n22971),
	.B(FE_OCPN29441_sa23_4),
	.C(n22951));
   NOR2xp33_ASAP7_75t_L U23786 (.Y(n16685),
	.A(n18415),
	.B(n16684));
   NAND2xp67_ASAP7_75t_SL U23787 (.Y(n17007),
	.A(n17003),
	.B(n17004));
   NOR2xp33_ASAP7_75t_SL U23788 (.Y(n20966),
	.A(FE_OCPN29546_n),
	.B(n20965));
   NAND2xp33_ASAP7_75t_SL U23789 (.Y(n19454),
	.A(n19453),
	.B(n19452));
   NAND2xp33_ASAP7_75t_SRAM U23790 (.Y(n18371),
	.A(n22166),
	.B(n19035));
   NAND2xp5_ASAP7_75t_L U23791 (.Y(n21178),
	.A(FE_OCPN27500_n19834),
	.B(n21154));
   AND3x1_ASAP7_75t_SL U23793 (.Y(n20761),
	.A(n26872),
	.B(n20759),
	.C(n23343));
   OAI22xp33_ASAP7_75t_SRAM U23794 (.Y(n18228),
	.A1(FE_OCPN27722_n23336),
	.A2(n23169),
	.B1(n18159),
	.B2(n23169));
   NOR2xp33_ASAP7_75t_L U23795 (.Y(n21216),
	.A(FE_OFN29081_n18526),
	.B(n21217));
   NAND2xp33_ASAP7_75t_SL U23796 (.Y(n18556),
	.A(n18553),
	.B(n21637));
   NAND2xp33_ASAP7_75t_L U23797 (.Y(n16958),
	.A(n16954),
	.B(n16955));
   NOR2xp33_ASAP7_75t_R U23798 (.Y(n16858),
	.A(FE_OFN28999_n16923),
	.B(n16859));
   OAI21xp33_ASAP7_75t_L U23799 (.Y(n23106),
	.A1(n23107),
	.A2(FE_OCPN29334_n17330),
	.B(n23100));
   NAND2xp33_ASAP7_75t_L U23801 (.Y(n20548),
	.A(n20545),
	.B(n20544));
   NOR3x1_ASAP7_75t_L U23802 (.Y(n19880),
	.A(n19878),
	.B(n19877),
	.C(n19876));
   OAI22xp33_ASAP7_75t_SRAM U23803 (.Y(n16802),
	.A1(FE_OCPN28298_n),
	.A2(n22696),
	.B1(n16757),
	.B2(n22696));
   NAND2xp33_ASAP7_75t_SRAM U23804 (.Y(n20065),
	.A(FE_OCPN27516_n26292),
	.B(FE_OCPN27444_n20064));
   NAND2x1_ASAP7_75t_L U23807 (.Y(n16464),
	.A(n16460),
	.B(n16461));
   AND3x1_ASAP7_75t_SL U23808 (.Y(n17289),
	.A(n21462),
	.B(FE_OCPN27843_n18750),
	.C(n21457));
   OAI21xp33_ASAP7_75t_SL U23809 (.Y(n14400),
	.A1(n15349),
	.A2(n13875),
	.B(n14399));
   INVxp33_ASAP7_75t_L U23810 (.Y(n15163),
	.A(n15160));
   OAI21xp33_ASAP7_75t_R U23811 (.Y(n14694),
	.A1(FE_OFN26639_w3_14),
	.A2(FE_OFN16459_n),
	.B(FE_OCPN29583_n15422));
   NAND2xp33_ASAP7_75t_R U23812 (.Y(n14761),
	.A(n14753),
	.B(n14752));
   NAND2xp5_ASAP7_75t_R U23814 (.Y(n13989),
	.A(n13988),
	.B(FE_OFN27135_n15992));
   NOR2x1p5_ASAP7_75t_SL U23815 (.Y(n14927),
	.A(FE_OFN28884_n),
	.B(n16016));
   OAI22xp33_ASAP7_75t_R U23816 (.Y(n14872),
	.A1(n15636),
	.A2(n15032),
	.B1(n15835),
	.B2(n15032));
   NAND2xp33_ASAP7_75t_R U23818 (.Y(n15000),
	.A(n14999),
	.B(n14998));
   NAND2xp5_ASAP7_75t_R U23819 (.Y(n14274),
	.A(n14273),
	.B(n14272));
   NOR2x1_ASAP7_75t_L U23820 (.Y(n15993),
	.A(FE_OCPN29535_FE_OFN8_w3_14),
	.B(n15414));
   NAND2xp33_ASAP7_75t_L U23821 (.Y(n15078),
	.A(n15077),
	.B(n15076));
   OAI21xp33_ASAP7_75t_R U23822 (.Y(n15923),
	.A1(FE_OFN28883_n),
	.A2(n15447),
	.B(n15446));
   INVxp33_ASAP7_75t_L U23823 (.Y(n13643),
	.A(n14571));
   NAND2xp5_ASAP7_75t_SL U23824 (.Y(n25114),
	.A(n25112),
	.B(n25111));
   NAND2xp33_ASAP7_75t_SRAM U23825 (.Y(n25320),
	.A(FE_PSN8293_n25317),
	.B(n25316));
   NOR2xp33_ASAP7_75t_SL U23826 (.Y(n23842),
	.A(FE_OFN29076_n18540),
	.B(n23840));
   NAND2xp5_ASAP7_75t_L U23827 (.Y(n17388),
	.A(n17326),
	.B(n17387));
   OAI21xp33_ASAP7_75t_SL U23828 (.Y(n26881),
	.A1(n26880),
	.A2(n26879),
	.B(n26878));
   NAND2xp5_ASAP7_75t_L U23829 (.Y(n19233),
	.A(n19232),
	.B(n19231));
   NAND2xp33_ASAP7_75t_SRAM U23830 (.Y(n18097),
	.A(n18094),
	.B(n18093));
   NOR2xp33_ASAP7_75t_L U23832 (.Y(n17497),
	.A(FE_OCPN27730_n17464),
	.B(n19192));
   OAI21xp33_ASAP7_75t_L U23833 (.Y(n23821),
	.A1(FE_OCPN28353_n18534),
	.A2(n20670),
	.B(n23773));
   OAI21xp5_ASAP7_75t_SL U23834 (.Y(n19281),
	.A1(FE_OFN28961_n17744),
	.A2(FE_OCPN27503_n20195),
	.B(n19273));
   NOR2x1_ASAP7_75t_SL U23835 (.Y(n22978),
	.A(n26149),
	.B(n20224));
   NAND2xp33_ASAP7_75t_SRAM U23836 (.Y(n22200),
	.A(n22199),
	.B(n22198));
   OAI21xp33_ASAP7_75t_L U23837 (.Y(n19612),
	.A1(FE_OCPN28270_n17237),
	.A2(FE_OFN26172_n19609),
	.B(n21461));
   NAND2xp33_ASAP7_75t_R U23838 (.Y(n23817),
	.A(n23816),
	.B(n23815));
   NAND2xp33_ASAP7_75t_SL U23839 (.Y(n23506),
	.A(n23505),
	.B(n23502));
   OAI21x1_ASAP7_75t_L U23840 (.Y(n20378),
	.A1(n23107),
	.A2(FE_OCPN28000_n22450),
	.B(n18685));
   NAND2xp33_ASAP7_75t_SRAM U23842 (.Y(n20113),
	.A(n20111),
	.B(n24872));
   NOR2xp33_ASAP7_75t_SRAM U23843 (.Y(n21309),
	.A(n21708),
	.B(n18008));
   NOR2x1_ASAP7_75t_L U23845 (.Y(n22900),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(n20153));
   NOR2xp33_ASAP7_75t_SRAM U23846 (.Y(n17164),
	.A(FE_OCPN29358_n17159),
	.B(n17165));
   NOR2xp33_ASAP7_75t_L U23847 (.Y(n19463),
	.A(FE_OCPN7618_n21027),
	.B(n19462));
   NAND2xp33_ASAP7_75t_SL U23848 (.Y(n21022),
	.A(n21021),
	.B(n21020));
   NOR3xp33_ASAP7_75t_SL U23849 (.Y(n22140),
	.A(n25107),
	.B(n22168),
	.C(n22139));
   NAND2xp5_ASAP7_75t_L U23850 (.Y(n18360),
	.A(n22125),
	.B(FE_OCPN8207_n18497));
   NAND2xp5_ASAP7_75t_L U23851 (.Y(n19851),
	.A(n19850),
	.B(n19849));
   NOR2xp33_ASAP7_75t_R U23853 (.Y(n22501),
	.A(FE_OCPN29378_n23266),
	.B(FE_OCPN28447_n23392));
   NAND2x1_ASAP7_75t_SL U23855 (.Y(n21847),
	.A(n17445),
	.B(FE_OCPN29439_n17447));
   NAND2xp33_ASAP7_75t_R U23856 (.Y(n21622),
	.A(n21621),
	.B(n21620));
   NAND2xp33_ASAP7_75t_L U23858 (.Y(n20731),
	.A(n20728),
	.B(n20727));
   NAND2xp33_ASAP7_75t_SRAM U23859 (.Y(n21136),
	.A(n21135),
	.B(n22802));
   NAND2xp5_ASAP7_75t_L U23860 (.Y(n20722),
	.A(n20721),
	.B(n22318));
   NAND2xp33_ASAP7_75t_L U23862 (.Y(n21214),
	.A(n21210),
	.B(n23832));
   NAND2xp5_ASAP7_75t_L U23863 (.Y(n18547),
	.A(n23856),
	.B(n18540));
   NAND2xp5_ASAP7_75t_SL U23864 (.Y(n16881),
	.A(n16879),
	.B(n16878));
   NAND2xp5_ASAP7_75t_L U23865 (.Y(n16945),
	.A(n16418),
	.B(n16854));
   NOR3xp33_ASAP7_75t_SL U23866 (.Y(n22932),
	.A(n22931),
	.B(n22930),
	.C(n22929));
   AND3x1_ASAP7_75t_R U23868 (.Y(n23108),
	.A(n23104),
	.B(n23103),
	.C(n23102));
   NAND2xp5_ASAP7_75t_SL U23869 (.Y(n17340),
	.A(n17336),
	.B(n17337));
   NAND2xp5_ASAP7_75t_SL U23871 (.Y(n22259),
	.A(n23596),
	.B(n23609));
   NAND2xp33_ASAP7_75t_L U23872 (.Y(n19533),
	.A(n19525),
	.B(n19524));
   NOR2xp33_ASAP7_75t_SRAM U23873 (.Y(n17536),
	.A(n22392),
	.B(n24868));
   NAND2xp33_ASAP7_75t_R U23875 (.Y(n17849),
	.A(n17848),
	.B(n17847));
   OAI21xp5_ASAP7_75t_L U23876 (.Y(n24256),
	.A1(n23633),
	.A2(n16762),
	.B(n22661));
   OAI22xp33_ASAP7_75t_L U23877 (.Y(n21947),
	.A1(FE_OFN27043_n),
	.A2(n21972),
	.B1(n21946),
	.B2(n21972));
   NOR3xp33_ASAP7_75t_SRAM U23878 (.Y(n16395),
	.A(n21939),
	.B(FE_OFN28719_n20025),
	.C(n16394));
   NAND2xp5_ASAP7_75t_L U23879 (.Y(n16328),
	.A(n21986),
	.B(n20052));
   NAND2xp33_ASAP7_75t_SRAM U23880 (.Y(n24059),
	.A(n24054),
	.B(n24056));
   NAND2xp33_ASAP7_75t_R U23881 (.Y(n18648),
	.A(n18644),
	.B(n18645));
   OAI21xp5_ASAP7_75t_SL U23882 (.Y(n22981),
	.A1(FE_OFN28841_n22980),
	.A2(FE_OCPN28363_n22979),
	.B(n22978));
   NAND2xp5_ASAP7_75t_SL U23883 (.Y(n17292),
	.A(n17288),
	.B(n17289));
   INVxp33_ASAP7_75t_SRAM U23884 (.Y(n14495),
	.A(n14493));
   O2A1O1Ixp5_ASAP7_75t_SRAM U23885 (.Y(n14186),
	.A1(n14439),
	.A2(FE_OFN16276_w3_5),
	.B(n14185),
	.C(n15596));
   NAND2xp33_ASAP7_75t_SRAM U23886 (.Y(n13800),
	.A(FE_PSN8271_n15924),
	.B(n14897));
   NAND2xp33_ASAP7_75t_SRAM U23887 (.Y(n15153),
	.A(n15148),
	.B(n15150));
   AND3x1_ASAP7_75t_L U23889 (.Y(n13281),
	.A(n13278),
	.B(n13636),
	.C(n13277));
   NAND2xp33_ASAP7_75t_R U23890 (.Y(n13886),
	.A(n13880),
	.B(n13883));
   INVx1_ASAP7_75t_SL U23891 (.Y(n15356),
	.A(n15355));
   NAND2xp33_ASAP7_75t_L U23892 (.Y(n13368),
	.A(n13362),
	.B(n13365));
   INVx1_ASAP7_75t_L U23893 (.Y(n15390),
	.A(n15387));
   NAND2xp5_ASAP7_75t_SL U23894 (.Y(n13470),
	.A(n13469),
	.B(n13468));
   OAI21xp33_ASAP7_75t_SRAM U23895 (.Y(n14911),
	.A1(n15993),
	.A2(n13805),
	.B(n14903));
   NAND2xp33_ASAP7_75t_SL U23896 (.Y(n13703),
	.A(n13702),
	.B(n13701));
   NAND2x1_ASAP7_75t_L U23897 (.Y(n14417),
	.A(n15835),
	.B(n15834));
   NAND2xp33_ASAP7_75t_R U23900 (.Y(n23594),
	.A(n23589),
	.B(FE_OFN85_n23588));
   NAND2xp5_ASAP7_75t_R U23901 (.Y(n20465),
	.A(n20461),
	.B(n20462));
   NOR3xp33_ASAP7_75t_SRAM U23902 (.Y(n25321),
	.A(n25320),
	.B(n25319),
	.C(n25318));
   NOR3xp33_ASAP7_75t_SRAM U23903 (.Y(n18931),
	.A(n25990),
	.B(FE_OCPN27589_n25987),
	.C(n18930));
   NOR3xp33_ASAP7_75t_SRAM U23904 (.Y(n26167),
	.A(n26166),
	.B(n22917),
	.C(n26164));
   NAND2xp33_ASAP7_75t_L U23905 (.Y(n19195),
	.A(n19186),
	.B(n19185));
   OAI21xp33_ASAP7_75t_SRAM U23906 (.Y(n19977),
	.A1(n22662),
	.A2(FE_OCPN27246_n22663),
	.B(n19972));
   NAND2xp5_ASAP7_75t_L U23907 (.Y(n18505),
	.A(FE_OFN28610_n22125),
	.B(n22157));
   OAI22xp33_ASAP7_75t_L U23908 (.Y(n21375),
	.A1(FE_OFN29054_n17453),
	.A2(FE_OCPN28082_n21860),
	.B1(n17444),
	.B2(FE_OCPN28082_n21860));
   NAND2xp33_ASAP7_75t_R U23910 (.Y(n22701),
	.A(n22700),
	.B(n22699));
   NAND2xp33_ASAP7_75t_L U23911 (.Y(n19953),
	.A(n22372),
	.B(n19741));
   NAND2x1p5_ASAP7_75t_SL U23912 (.Y(n19721),
	.A(FE_OFN28892_n),
	.B(n17565));
   NOR3xp33_ASAP7_75t_SL U23913 (.Y(n23949),
	.A(n16556),
	.B(FE_OFN28751_n),
	.C(n16581));
   NAND2xp33_ASAP7_75t_SL U23914 (.Y(n20615),
	.A(n20614),
	.B(n20693));
   NAND2xp33_ASAP7_75t_L U23916 (.Y(n20682),
	.A(n20681),
	.B(n20680));
   NAND2xp5_ASAP7_75t_SL U23917 (.Y(n16629),
	.A(n16597),
	.B(n16596));
   NOR2x1_ASAP7_75t_SL U23918 (.Y(n21752),
	.A(FE_OFN28886_FE_OCPN27675_n17986),
	.B(FE_OCPN29283_n23439));
   NAND2xp5_ASAP7_75t_SL U23919 (.Y(n23508),
	.A(n23507),
	.B(n23506));
   NAND2xp5_ASAP7_75t_SL U23921 (.Y(n16405),
	.A(n16404),
	.B(n16403));
   NOR2xp33_ASAP7_75t_L U23922 (.Y(n16798),
	.A(FE_OCPN27289_sa21_5),
	.B(n23628));
   INVx1_ASAP7_75t_L U23923 (.Y(n16705),
	.A(FE_OCPN27460_n16913));
   NOR3xp33_ASAP7_75t_SRAM U23924 (.Y(n17605),
	.A(n18503),
	.B(FE_OFN28895_sa30_2),
	.C(n19051));
   NAND2xp5_ASAP7_75t_L U23926 (.Y(n21306),
	.A(n21305),
	.B(n24245));
   O2A1O1Ixp5_ASAP7_75t_SRAM U23927 (.Y(n18876),
	.A1(n21269),
	.A2(n21738),
	.B(FE_OCPN27617_n18016),
	.C(n21752));
   NOR2x1_ASAP7_75t_L U23928 (.Y(n21740),
	.A(FE_OCPN29283_n23439),
	.B(FE_OFN28588_n21048));
   NAND2xp5_ASAP7_75t_SL U23930 (.Y(n21157),
	.A(FE_OFN26146_n18774),
	.B(n19609));
   NAND2xp33_ASAP7_75t_SRAM U23931 (.Y(n18761),
	.A(FE_OCPN29346_n12998),
	.B(FE_OFN28835_n));
   OAI21xp5_ASAP7_75t_L U23932 (.Y(n17307),
	.A1(n18735),
	.A2(n17306),
	.B(n26637));
   NAND2xp5_ASAP7_75t_R U23933 (.Y(n18288),
	.A(n17131),
	.B(n17086));
   NOR2x1p5_ASAP7_75t_SL U23934 (.Y(n20993),
	.A(FE_OFN26077_n),
	.B(FE_OFN16136_sa02_5));
   NOR2xp33_ASAP7_75t_SRAM U23935 (.Y(n17770),
	.A(n20161),
	.B(n20987));
   NAND2xp33_ASAP7_75t_R U23936 (.Y(n22102),
	.A(n22101),
	.B(n22100));
   NOR2x1p5_ASAP7_75t_SL U23938 (.Y(n20529),
	.A(FE_OFN28491_sa13_3),
	.B(n17033));
   OR3x1_ASAP7_75t_R U23939 (.Y(n19482),
	.A(n19480),
	.B(n21301),
	.C(n21728));
   NAND2xp33_ASAP7_75t_SL U23940 (.Y(n21294),
	.A(n21291),
	.B(n21290));
   NOR2x1_ASAP7_75t_L U23941 (.Y(n23430),
	.A(FE_OFN28677_n17998),
	.B(n21725));
   NAND2xp5_ASAP7_75t_L U23943 (.Y(n19633),
	.A(n19632),
	.B(FE_OCPN27906_n23131));
   NOR3xp33_ASAP7_75t_SRAM U23944 (.Y(n16550),
	.A(n23997),
	.B(n19661),
	.C(FE_OFN29159_n21892));
   NAND2xp5_ASAP7_75t_SL U23945 (.Y(n19153),
	.A(n19148),
	.B(n19147));
   NAND2xp5_ASAP7_75t_SL U23946 (.Y(n22642),
	.A(n21613),
	.B(FE_OCPN28241_n22142));
   OAI21xp33_ASAP7_75t_SRAM U23947 (.Y(n23281),
	.A1(FE_OCPN28006_n17454),
	.A2(FE_OFN28996_n17464),
	.B(FE_OCPN28417_n21396));
   NAND2xp5_ASAP7_75t_SL U23948 (.Y(n21384),
	.A(n21381),
	.B(n21380));
   NOR3xp33_ASAP7_75t_SL U23949 (.Y(n23275),
	.A(n21423),
	.B(n21834),
	.C(n21422));
   NOR2x1_ASAP7_75t_SL U23950 (.Y(n21854),
	.A(FE_OFN29170_n17510),
	.B(n21374));
   NAND2xp33_ASAP7_75t_L U23951 (.Y(n18471),
	.A(FE_OCPN29467_n25102),
	.B(n25108));
   NAND2xp33_ASAP7_75t_SL U23953 (.Y(n17662),
	.A(FE_OFN16333_sa30_4),
	.B(n17659));
   NAND2xp5_ASAP7_75t_L U23954 (.Y(n18523),
	.A(FE_OCPN27371_sa20_2),
	.B(n23856));
   NAND2xp5_ASAP7_75t_SL U23955 (.Y(n23164),
	.A(n18216),
	.B(n21135));
   NAND2xp5_ASAP7_75t_R U23956 (.Y(n22834),
	.A(n22824),
	.B(n22823));
   NAND2x2_ASAP7_75t_SL U23957 (.Y(n18178),
	.A(n23308),
	.B(n18199));
   NOR2x1_ASAP7_75t_SL U23959 (.Y(n21193),
	.A(n18530),
	.B(n23677));
   NOR3xp33_ASAP7_75t_SL U23960 (.Y(n21253),
	.A(n23711),
	.B(n18522),
	.C(FE_OCPN7626_n18582));
   NAND2xp33_ASAP7_75t_SRAM U23961 (.Y(n18428),
	.A(n18441),
	.B(n18427));
   NOR2xp33_ASAP7_75t_R U23962 (.Y(n17420),
	.A(n18108),
	.B(n18107));
   NAND2xp5_ASAP7_75t_SL U23963 (.Y(n16864),
	.A(n16863),
	.B(n16862));
   NAND2xp33_ASAP7_75t_SRAM U23965 (.Y(n22939),
	.A(n22934),
	.B(n22936));
   NAND2xp33_ASAP7_75t_L U23966 (.Y(n23111),
	.A(n23105),
	.B(n23108));
   NOR2x1_ASAP7_75t_SL U23967 (.Y(n22582),
	.A(FE_OFN25878_n17329),
	.B(FE_OCPN29406_n18710));
   NAND2xp33_ASAP7_75t_SRAM U23968 (.Y(n22444),
	.A(n22439),
	.B(FE_OFN27064_n22438));
   OAI21xp33_ASAP7_75t_SRAM U23969 (.Y(n19545),
	.A1(n19539),
	.A2(FE_OFN28520_n22753),
	.B(FE_OCPN27368_sa12_3));
   NAND2xp33_ASAP7_75t_R U23970 (.Y(n17955),
	.A(n22261),
	.B(n25399));
   NAND2x1p5_ASAP7_75t_L U23971 (.Y(n22722),
	.A(FE_OCPN28198_n22776),
	.B(n24362));
   NOR2x1p5_ASAP7_75t_L U23972 (.Y(n23600),
	.A(FE_OCPN29485_sa12_3),
	.B(n19509));
   NAND2xp33_ASAP7_75t_SRAM U23973 (.Y(n17556),
	.A(n19941),
	.B(n19720));
   NOR2x1p5_ASAP7_75t_L U23974 (.Y(n19926),
	.A(FE_OCPN29298_n25028),
	.B(FE_OCPN29323_n19721));
   OAI21xp5_ASAP7_75t_SL U23975 (.Y(n18789),
	.A1(FE_OFN26577_n),
	.A2(FE_OCPN27267_n18794),
	.B(n22397));
   NOR3x1_ASAP7_75t_L U23976 (.Y(n19975),
	.A(FE_OCPN27556_n17843),
	.B(FE_OCPN27328_sa21_2),
	.C(n16801));
   NOR2xp33_ASAP7_75t_SRAM U23977 (.Y(n23642),
	.A(FE_OFN16153_n16747),
	.B(n23643));
   INVxp67_ASAP7_75t_L U23978 (.Y(n16397),
	.A(n20050));
   NAND2xp33_ASAP7_75t_SL U23979 (.Y(n18081),
	.A(n18078),
	.B(n20849));
   NAND2xp5_ASAP7_75t_L U23981 (.Y(n16331),
	.A(n20841),
	.B(FE_OFN27043_n));
   NOR2x1_ASAP7_75t_L U23982 (.Y(n20251),
	.A(n22010),
	.B(FE_OCPN27288_n25091));
   NAND2xp33_ASAP7_75t_L U23983 (.Y(n24675),
	.A(n24670),
	.B(FE_OFN131_sa10_6));
   NAND2xp5_ASAP7_75t_SL U23984 (.Y(n19659),
	.A(n19655),
	.B(n19656));
   NAND2xp33_ASAP7_75t_L U23985 (.Y(n18649),
	.A(n18648),
	.B(n18647));
   NOR2xp33_ASAP7_75t_SRAM U23986 (.Y(n17173),
	.A(FE_OCPN27902_n20514),
	.B(n17174));
   OAI22xp33_ASAP7_75t_L U23987 (.Y(n20629),
	.A1(FE_OCPN27606_n23869),
	.A2(n23792),
	.B1(FE_OFN29139_n18527),
	.B2(n23792));
   NAND2xp5_ASAP7_75t_SL U23988 (.Y(n18995),
	.A(n18994),
	.B(n18993));
   NAND2xp33_ASAP7_75t_L U23989 (.Y(n14497),
	.A(n14492),
	.B(n14494));
   NAND2xp33_ASAP7_75t_L U23990 (.Y(n13810),
	.A(n13806),
	.B(n13807));
   NAND2xp33_ASAP7_75t_SRAM U23991 (.Y(n15803),
	.A(n15802),
	.B(n15801));
   NAND2xp33_ASAP7_75t_L U23993 (.Y(n13555),
	.A(n13553),
	.B(n13552));
   NAND2xp33_ASAP7_75t_R U23994 (.Y(n14618),
	.A(n14617),
	.B(n14616));
   OAI22xp5_ASAP7_75t_L U23995 (.Y(n15209),
	.A1(FE_OCPN29350_w3_25),
	.A2(FE_OFN27206_w3_30),
	.B1(FE_OFN26048_w3_27),
	.B2(FE_OFN27206_w3_30));
   OAI21xp33_ASAP7_75t_SRAM U23996 (.Y(n14263),
	.A1(n15478),
	.A2(n15693),
	.B(FE_OFN27074_n13868));
   NAND2xp5_ASAP7_75t_L U23997 (.Y(n15651),
	.A(n15624),
	.B(n15648));
   NAND2xp33_ASAP7_75t_L U23999 (.Y(n13494),
	.A(n13490),
	.B(n13491));
   NAND2xp33_ASAP7_75t_SL U24000 (.Y(n13705),
	.A(n13704),
	.B(n13703));
   NAND2x1_ASAP7_75t_SL U24001 (.Y(n25199),
	.A(FE_OCPN29523_n25544),
	.B(n17031));
   NOR2x1p5_ASAP7_75t_SL U24002 (.Y(n25612),
	.A(n25610),
	.B(FE_OCPN29481_n26537));
   NAND2x1_ASAP7_75t_SL U24005 (.Y(n26009),
	.A(n16525),
	.B(n16378));
   NOR2xp33_ASAP7_75t_SRAM U24007 (.Y(n23313),
	.A(n18177),
	.B(n23314));
   NAND2xp5_ASAP7_75t_L U24008 (.Y(n19993),
	.A(FE_OFN28981_n16767),
	.B(FE_OFN16447_n16749));
   NAND2xp33_ASAP7_75t_L U24009 (.Y(n16448),
	.A(n16427),
	.B(FE_OCPN27555_n16422));
   NOR3xp33_ASAP7_75t_SRAM U24010 (.Y(n17702),
	.A(n17699),
	.B(FE_OCPN28392_n22380),
	.C(n17698));
   NAND2xp33_ASAP7_75t_SRAM U24011 (.Y(n17025),
	.A(n17024),
	.B(n17023));
   NOR3xp33_ASAP7_75t_SRAM U24012 (.Y(n19298),
	.A(n19297),
	.B(n20251),
	.C(FE_OFN27046_n22024));
   NAND2xp5_ASAP7_75t_SL U24013 (.Y(n22891),
	.A(n20170),
	.B(n17757));
   OAI21xp33_ASAP7_75t_SRAM U24014 (.Y(n19778),
	.A1(FE_OFN130_sa10_5),
	.A2(n23951),
	.B(n19777));
   NAND2xp33_ASAP7_75t_L U24015 (.Y(n20651),
	.A(n20650),
	.B(n20649));
   OAI21xp33_ASAP7_75t_SRAM U24016 (.Y(n22192),
	.A1(FE_OFN27152_n17315),
	.A2(n22191),
	.B(n22190));
   NAND2xp5_ASAP7_75t_L U24017 (.Y(n21548),
	.A(FE_OCPN28305_n26451),
	.B(n17373));
   NAND2xp33_ASAP7_75t_SRAM U24018 (.Y(n20569),
	.A(n20568),
	.B(n20566));
   NOR2xp33_ASAP7_75t_L U24019 (.Y(n23415),
	.A(n23413),
	.B(n23412));
   NOR2xp33_ASAP7_75t_R U24020 (.Y(n20382),
	.A(FE_OCPN27988_n26454),
	.B(n20380));
   NAND2x1p5_ASAP7_75t_SL U24021 (.Y(n16801),
	.A(FE_OFN28678_sa21_3),
	.B(n16783));
   NAND2x1p5_ASAP7_75t_SL U24022 (.Y(n18381),
	.A(FE_OCPN29431_sa30_3),
	.B(FE_OFN28901_sa30_4));
   NAND2xp33_ASAP7_75t_L U24024 (.Y(n18256),
	.A(FE_OFN16162_n25869),
	.B(FE_OFN28801_n16978));
   NOR2xp33_ASAP7_75t_SRAM U24026 (.Y(n19913),
	.A(FE_OCPN28268_n19911),
	.B(n19910));
   NAND2x1p5_ASAP7_75t_SL U24027 (.Y(n23981),
	.A(FE_OFN27196_n),
	.B(n19756));
   NAND2xp5_ASAP7_75t_L U24029 (.Y(n25914),
	.A(FE_OCPN29469_n17747),
	.B(FE_OCPN27384_n22888));
   INVxp67_ASAP7_75t_L U24030 (.Y(n18249),
	.A(n19408));
   NAND2xp5_ASAP7_75t_SL U24031 (.Y(n20532),
	.A(n19376),
	.B(FE_OFN26170_n19361));
   NAND2xp5_ASAP7_75t_SL U24032 (.Y(n25995),
	.A(FE_OFN29074_n17170),
	.B(n16983));
   NOR2x1_ASAP7_75t_L U24033 (.Y(n23454),
	.A(n21015),
	.B(n18048));
   OAI21xp33_ASAP7_75t_SRAM U24035 (.Y(n19645),
	.A1(n16533),
	.A2(n23982),
	.B(n19642));
   NOR2xp33_ASAP7_75t_SRAM U24038 (.Y(n20420),
	.A(FE_PSN8335_n17606),
	.B(n20421));
   NAND2x1p5_ASAP7_75t_SL U24039 (.Y(n21374),
	.A(FE_OFN29137_FE_OCPN27228_sa11_2),
	.B(n19206));
   NOR2x1p5_ASAP7_75t_SL U24040 (.Y(n19090),
	.A(FE_OCPN29411_n),
	.B(n21152));
   NAND2xp33_ASAP7_75t_SRAM U24043 (.Y(n21652),
	.A(FE_OCPN27896_n18583),
	.B(FE_OFN28986_n18597));
   NAND2xp5_ASAP7_75t_SL U24044 (.Y(n23892),
	.A(n23777),
	.B(n23776));
   NAND2x1_ASAP7_75t_SL U24045 (.Y(n17418),
	.A(FE_OFN29134_sa33_0),
	.B(n16423));
   NAND2x1p5_ASAP7_75t_R U24047 (.Y(n18446),
	.A(FE_OFN29164_sa33_2),
	.B(n16472));
   NAND2x1_ASAP7_75t_SL U24048 (.Y(n16473),
	.A(FE_OCPN29391_FE_OFN29162_sa33_2),
	.B(n16873));
   NAND2xp33_ASAP7_75t_SL U24049 (.Y(n18983),
	.A(FE_OFN28598_n20933),
	.B(n18981));
   OAI21xp33_ASAP7_75t_SL U24050 (.Y(n22031),
	.A1(FE_OCPN29488_FE_OFN25883_n22945),
	.A2(n20920),
	.B(n20247));
   NOR2x1_ASAP7_75t_SL U24051 (.Y(n20389),
	.A(n18726),
	.B(n21545));
   NAND2x2_ASAP7_75t_SL U24052 (.Y(n18667),
	.A(FE_OFN29254_n),
	.B(n17331));
   NAND2x1p5_ASAP7_75t_L U24055 (.Y(n23617),
	.A(FE_OCPN27429_sa12_3),
	.B(n23208));
   NOR3x1_ASAP7_75t_SL U24056 (.Y(n22773),
	.A(n19535),
	.B(FE_OFN28723_n22750),
	.C(n23602));
   NAND2x1p5_ASAP7_75t_L U24057 (.Y(n18832),
	.A(FE_OFN16463_sa32_0),
	.B(FE_OCPN29304_n17526));
   NOR2xp33_ASAP7_75t_SRAM U24058 (.Y(n24858),
	.A(FE_OCPN28268_n19911),
	.B(n20095));
   NAND2xp5_ASAP7_75t_L U24059 (.Y(n17869),
	.A(FE_OCPN27690_n16757),
	.B(FE_OCPN28299_n));
   NAND2xp33_ASAP7_75t_L U24060 (.Y(n22341),
	.A(n19974),
	.B(n19973));
   NOR2xp33_ASAP7_75t_SRAM U24061 (.Y(n23631),
	.A(FE_OFN28836_FE_OCPN27631_n16774),
	.B(n23632));
   NOR2xp33_ASAP7_75t_L U24063 (.Y(n16316),
	.A(FE_OFN29032_FE_OCPN27728_n21981),
	.B(n20049));
   AND3x1_ASAP7_75t_SRAM U24064 (.Y(n16367),
	.A(n25815),
	.B(n24182),
	.C(n16365));
   NAND2xp5_ASAP7_75t_SL U24065 (.Y(n24906),
	.A(n24903),
	.B(n24902));
   NAND2xp33_ASAP7_75t_SRAM U24066 (.Y(n18996),
	.A(n23511),
	.B(n20238));
   NAND2xp33_ASAP7_75t_L U24067 (.Y(n23488),
	.A(n22975),
	.B(n22974));
   OAI22xp33_ASAP7_75t_SRAM U24068 (.Y(n13814),
	.A1(n15986),
	.A2(n13803),
	.B1(n13949),
	.B2(n13803));
   INVxp67_ASAP7_75t_SL U24069 (.Y(n13998),
	.A(n13999));
   NAND2xp33_ASAP7_75t_L U24070 (.Y(n14843),
	.A(n14842),
	.B(n14841));
   NAND2xp33_ASAP7_75t_L U24071 (.Y(n13347),
	.A(n13342),
	.B(n13341));
   INVxp67_ASAP7_75t_SL U24072 (.Y(n13475),
	.A(n13476));
   AOI21xp5_ASAP7_75t_SL U24073 (.Y(n27155),
	.A1(FE_OFN28483_ld_r),
	.A2(FE_OCPN28122_n27157),
	.B(n27156));
   NAND2xp33_ASAP7_75t_SL U24074 (.Y(n26112),
	.A(n26110),
	.B(n26109));
   O2A1O1Ixp5_ASAP7_75t_SL U24075 (.Y(n24108),
	.A1(n26777),
	.A2(n26776),
	.B(n24106),
	.C(n24105));
   NAND2xp33_ASAP7_75t_SRAM U24076 (.Y(n24380),
	.A(n24366),
	.B(n24365));
   O2A1O1Ixp33_ASAP7_75t_SL U24077 (.Y(n25421),
	.A1(n25420),
	.A2(FE_OFN28561_n25419),
	.B(n25418),
	.C(n25417));
   OAI21x1_ASAP7_75t_SL U24078 (.Y(n23966),
	.A1(n25149),
	.A2(n26346),
	.B(n25146));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24079 (.Y(n26089),
	.A1(FE_OFN16180_n26542),
	.A2(n18158),
	.B(n26088),
	.C(n26095));
   NOR2x1_ASAP7_75t_R U24080 (.Y(n25073),
	.A(n25071),
	.B(n25070));
   NAND2xp33_ASAP7_75t_L U24081 (.Y(n19971),
	.A(n19965),
	.B(FE_OCPN5167_n22336));
   NAND2xp33_ASAP7_75t_R U24082 (.Y(n23212),
	.A(n23207),
	.B(n23209));
   NAND2xp33_ASAP7_75t_SRAM U24083 (.Y(n23261),
	.A(n23260),
	.B(n23259));
   OAI21xp33_ASAP7_75t_SRAM U24084 (.Y(n23304),
	.A1(n23303),
	.A2(FE_OCPN29305_n23302),
	.B(n23301));
   NAND2xp33_ASAP7_75t_SL U24085 (.Y(n22660),
	.A(n17845),
	.B(n19993));
   OAI21xp33_ASAP7_75t_L U24086 (.Y(n23757),
	.A1(n23677),
	.A2(FE_OFN28815_n18523),
	.B(n23755));
   NAND2xp5_ASAP7_75t_L U24087 (.Y(n17684),
	.A(n17680),
	.B(n17681));
   NAND2xp33_ASAP7_75t_SL U24088 (.Y(n20640),
	.A(n20639),
	.B(n20638));
   OAI21xp5_ASAP7_75t_SL U24089 (.Y(n19586),
	.A1(FE_OCPN29292_n18640),
	.A2(n19817),
	.B(n21183));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24090 (.Y(n20605),
	.A1(n24065),
	.A2(n24064),
	.B(n25682),
	.C(n24049));
   NAND2xp5_ASAP7_75t_L U24091 (.Y(n27071),
	.A(n20073),
	.B(n16491));
   OR3x1_ASAP7_75t_SL U24093 (.Y(n23442),
	.A(n23422),
	.B(n23421),
	.C(n23420));
   OAI21xp5_ASAP7_75t_SL U24094 (.Y(n21308),
	.A1(FE_OCPN28184_n18020),
	.A2(n18011),
	.B(n21034));
   NOR2x1_ASAP7_75t_SL U24095 (.Y(n21546),
	.A(n17330),
	.B(FE_OCPN29406_n18710));
   NOR3x1_ASAP7_75t_SL U24096 (.Y(n22350),
	.A(n20302),
	.B(n20301),
	.C(n25580));
   NOR2x1p5_ASAP7_75t_L U24097 (.Y(n25528),
	.A(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(FE_OCPN28303_n20961));
   NAND2xp33_ASAP7_75t_SRAM U24098 (.Y(n23052),
	.A(n23026),
	.B(n23025));
   NOR2x1p5_ASAP7_75t_L U24099 (.Y(n21148),
	.A(n19097),
	.B(FE_OCPN28270_n17237));
   NAND2xp5_ASAP7_75t_L U24100 (.Y(n18735),
	.A(n17296),
	.B(n19572));
   NOR2x1_ASAP7_75t_L U24101 (.Y(n22881),
	.A(n20962),
	.B(n22083));
   NAND2xp33_ASAP7_75t_SRAM U24102 (.Y(n22071),
	.A(FE_OFN28515_n22062),
	.B(n25914));
   NAND2xp33_ASAP7_75t_SL U24103 (.Y(n21876),
	.A(n16536),
	.B(n19669));
   O2A1O1Ixp5_ASAP7_75t_L U24104 (.Y(n19858),
	.A1(n19857),
	.A2(n19856),
	.B(n26637),
	.C(n19855));
   O2A1O1Ixp33_ASAP7_75t_SL U24106 (.Y(n21433),
	.A1(n21432),
	.A2(n21431),
	.B(n26082),
	.C(n21430));
   NAND2xp5_ASAP7_75t_SL U24107 (.Y(n19193),
	.A(n21398),
	.B(n21428));
   NOR2xp33_ASAP7_75t_SRAM U24108 (.Y(n18495),
	.A(n18463),
	.B(n17618));
   O2A1O1Ixp33_ASAP7_75t_L U24109 (.Y(n23201),
	.A1(n23200),
	.A2(n23199),
	.B(n26878),
	.C(n23198));
   NAND2xp33_ASAP7_75t_L U24111 (.Y(n21206),
	.A(n23778),
	.B(n21204));
   NAND2xp33_ASAP7_75t_L U24112 (.Y(n23684),
	.A(n23679),
	.B(n23681));
   NAND2xp5_ASAP7_75t_SL U24113 (.Y(n23543),
	.A(FE_OFN16400_n17404),
	.B(n17406));
   O2A1O1Ixp5_ASAP7_75t_SL U24114 (.Y(n20282),
	.A1(n22923),
	.A2(n20281),
	.B(n26249),
	.C(n20280));
   OAI21xp33_ASAP7_75t_L U24115 (.Y(n17356),
	.A1(FE_OCPN27423_sa01_0),
	.A2(n22175),
	.B(n17373));
   NAND2xp5_ASAP7_75t_L U24116 (.Y(n22238),
	.A(n20598),
	.B(n19513));
   OAI22xp33_ASAP7_75t_SRAM U24117 (.Y(n20821),
	.A1(n20828),
	.A2(n26607),
	.B1(n26594),
	.B2(n26607));
   OAI21x1_ASAP7_75t_SL U24118 (.Y(n26051),
	.A1(n25566),
	.A2(n27102),
	.B(n25565));
   OAI21xp33_ASAP7_75t_R U24119 (.Y(n17831),
	.A1(FE_OCPN29414_n),
	.A2(n23628),
	.B(n23668));
   NAND2xp33_ASAP7_75t_R U24120 (.Y(n23636),
	.A(n23631),
	.B(n23630));
   NOR2x1_ASAP7_75t_L U24121 (.Y(n21982),
	.A(n20074),
	.B(FE_OCPN28008_n16290));
   NAND2xp33_ASAP7_75t_R U24122 (.Y(n24682),
	.A(n24676),
	.B(n24679));
   NAND2xp5_ASAP7_75t_L U24123 (.Y(n24659),
	.A(n24017),
	.B(n24016));
   NAND2xp33_ASAP7_75t_L U24124 (.Y(n24232),
	.A(n24416),
	.B(n24229));
   NAND2xp33_ASAP7_75t_R U24126 (.Y(n25604),
	.A(n25600),
	.B(sa00_6_));
   NAND2xp5_ASAP7_75t_SL U24128 (.Y(n14893),
	.A(n14879),
	.B(n26130));
   NAND2xp5_ASAP7_75t_L U24129 (.Y(n15059),
	.A(n14995),
	.B(n14994));
   O2A1O1Ixp33_ASAP7_75t_SL U24131 (.Y(n27158),
	.A1(FE_OCPN28122_n27157),
	.A2(FE_OFN2_ld_r),
	.B(n27156),
	.C(n27155));
   OAI22xp33_ASAP7_75t_SRAM U24132 (.Y(n27194),
	.A1(text_in_r_55_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(n27195),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL U24133 (.Y(n25983),
	.A(n26892),
	.B(n25984));
   O2A1O1Ixp5_ASAP7_75t_SL U24134 (.Y(n24454),
	.A1(n24837),
	.A2(n24448),
	.B(FE_OCPN28131_n26796),
	.C(n24447));
   OAI21xp5_ASAP7_75t_L U24135 (.Y(n26381),
	.A1(FE_OFN2_ld_r),
	.A2(n26383),
	.B(n26382));
   OAI22xp33_ASAP7_75t_SRAM U24136 (.Y(n24820),
	.A1(text_in_r_73_),
	.A2(FE_OFN28486_ld_r),
	.B1(n24821),
	.B2(FE_OFN28486_ld_r));
   NAND2xp5_ASAP7_75t_L U24137 (.Y(n26366),
	.A(n26364),
	.B(n26361));
   OAI21xp33_ASAP7_75t_SRAM U24138 (.Y(n24024),
	.A1(FE_OFN27138_n24012),
	.A2(n24011),
	.B(n22405));
   OAI21xp5_ASAP7_75t_L U24139 (.Y(n25048),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27292_n25389),
	.B(n25049));
   INVxp33_ASAP7_75t_R U24140 (.Y(n23924),
	.A(n23901));
   NAND2xp5_ASAP7_75t_L U24141 (.Y(n26177),
	.A(n26170),
	.B(n26169));
   OAI21xp5_ASAP7_75t_SL U24142 (.Y(n26608),
	.A1(FE_OFN16213_ld_r),
	.A2(FE_OCPN29382_n26674),
	.B(n26609));
   NOR2xp33_ASAP7_75t_SL U24143 (.Y(n26730),
	.A(n26729),
	.B(n26731));
   XNOR2xp5_ASAP7_75t_SL U24144 (.Y(n16131),
	.A(w1_31_),
	.B(n16055));
   INVx1_ASAP7_75t_SL U24145 (.Y(n24416),
	.A(n24421));
   INVxp33_ASAP7_75t_SRAM U24146 (.Y(n26538),
	.A(FE_OCPN29481_n26537));
   NAND2xp5_ASAP7_75t_R U24147 (.Y(n23887),
	.A(n20641),
	.B(n20640));
   NOR2xp33_ASAP7_75t_SRAM U24148 (.Y(n20553),
	.A(FE_OCPN28346_n24051),
	.B(n20552));
   INVxp67_ASAP7_75t_R U24149 (.Y(n26512),
	.A(w2_19_));
   NOR3xp33_ASAP7_75t_SRAM U24152 (.Y(n21508),
	.A(n21507),
	.B(n24243),
	.C(FE_OFN28922_n24249));
   NOR2xp33_ASAP7_75t_SRAM U24155 (.Y(n19816),
	.A(n26106),
	.B(n19815));
   INVxp33_ASAP7_75t_SRAM U24157 (.Y(n21144),
	.A(n24114));
   NAND2x1_ASAP7_75t_SL U24160 (.Y(n22428),
	.A(n20375),
	.B(n20374));
   OAI21xp5_ASAP7_75t_L U24161 (.Y(n26135),
	.A1(n22792),
	.A2(n26607),
	.B(n22791));
   INVx2_ASAP7_75t_SL U24162 (.Y(n25669),
	.A(n25667));
   O2A1O1Ixp33_ASAP7_75t_SL U24165 (.Y(n25496),
	.A1(FE_OCPN27753_n26685),
	.A2(n25494),
	.B(FE_OFN160_n26440),
	.C(n25493));
   NAND2xp33_ASAP7_75t_SRAM U24167 (.Y(n25474),
	.A(FE_OFN25979_n),
	.B(n25471));
   AOI22x1_ASAP7_75t_SL U24168 (.Y(n16225),
	.A1(w1_11_),
	.A2(FE_OFN16405_n16117),
	.B1(FE_OFN16403_n16117),
	.B2(n25690));
   AOI22x1_ASAP7_75t_SL U24169 (.Y(n15371),
	.A1(w1_1_),
	.A2(FE_OCPN29363_n14011),
	.B1(FE_OFN26020_n14010),
	.B2(n26991));
   INVxp33_ASAP7_75t_SRAM U24170 (.Y(n13145),
	.A(text_in_r_12_));
   INVxp33_ASAP7_75t_SRAM U24171 (.Y(n13041),
	.A(text_in_r_27_));
   INVxp33_ASAP7_75t_SRAM U24172 (.Y(n13261),
	.A(text_in_r_40_));
   INVxp33_ASAP7_75t_SRAM U24173 (.Y(n13071),
	.A(text_in_r_54_));
   INVxp33_ASAP7_75t_SRAM U24174 (.Y(n13253),
	.A(text_in_r_68_));
   INVxp33_ASAP7_75t_SRAM U24175 (.Y(n13177),
	.A(text_in_r_80_));
   INVxp33_ASAP7_75t_SRAM U24176 (.Y(n13119),
	.A(text_in_r_94_));
   INVxp33_ASAP7_75t_SRAM U24177 (.Y(n13025),
	.A(text_in_r_108_));
   INVxp33_ASAP7_75t_SRAM U24178 (.Y(n13259),
	.A(text_in_r_120_));
   NAND2xp33_ASAP7_75t_SRAM U24179 (.Y(n26863),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_15_));
   OAI21x1_ASAP7_75t_SL U24180 (.Y(n16078),
	.A1(n16059),
	.A2(n26202),
	.B(n16058));
   OAI21xp33_ASAP7_75t_SRAM U24181 (.Y(n25017),
	.A1(text_in_r_25_),
	.A2(FE_OCPN27659_w3_25),
	.B(n25015));
   OAI21xp33_ASAP7_75t_SRAM U24182 (.Y(n24576),
	.A1(text_in_r_121_),
	.A2(n24575),
	.B(n24574));
   OAI21xp33_ASAP7_75t_SRAM U24183 (.Y(n25459),
	.A1(text_in_r_89_),
	.A2(FE_OFN66_w1_25),
	.B(n25457));
   OAI21xp33_ASAP7_75t_SRAM U24185 (.Y(n24822),
	.A1(text_in_r_73_),
	.A2(n24821),
	.B(n24820));
   NAND2xp33_ASAP7_75t_SRAM U24186 (.Y(n26342),
	.A(FE_OFN28482_ld_r),
	.B(text_in_r_29_));
   INVxp33_ASAP7_75t_SRAM U24187 (.Y(n25729),
	.A(w1_16_));
   OAI21xp33_ASAP7_75t_SRAM U24188 (.Y(n25649),
	.A1(text_in_r_34_),
	.A2(n25648),
	.B(n25647));
   NAND2xp33_ASAP7_75t_SRAM U24189 (.Y(n25052),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_10_));
   O2A1O1Ixp33_ASAP7_75t_L U24190 (.Y(n24204),
	.A1(FE_OCPN5053_n25832),
	.A2(n25831),
	.B(FE_OCPN7589_n26420),
	.C(n24179));
   O2A1O1Ixp33_ASAP7_75t_SL U24191 (.Y(n24534),
	.A1(n24529),
	.A2(n24528),
	.B(FE_OCPN27514_n25981),
	.C(n24527));
   OAI22xp33_ASAP7_75t_SRAM U24192 (.Y(n26786),
	.A1(w0_3_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_99_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U24193 (.Y(n26209),
	.A1(w2_4_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_36_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   OAI21x1_ASAP7_75t_SL U24194 (.Y(n16050),
	.A1(n15910),
	.A2(n26310),
	.B(n15909));
   OAI21xp5_ASAP7_75t_SL U24195 (.Y(n16222),
	.A1(n16219),
	.A2(n26951),
	.B(n16218));
   NOR2xp33_ASAP7_75t_SRAM U24196 (.Y(n13010),
	.A(dcnt_0_),
	.B(n13007));
   NAND2xp33_ASAP7_75t_SRAM U24197 (.Y(n16489),
	.A(n26538),
	.B(n24506));
   NAND2xp5_ASAP7_75t_L U24198 (.Y(n26678),
	.A(FE_OFN26566_n24208),
	.B(n24206));
   NAND2xp33_ASAP7_75t_SRAM U24199 (.Y(n16530),
	.A(n16527),
	.B(n26615));
   NAND2xp33_ASAP7_75t_SRAM U24200 (.Y(n23527),
	.A(FE_OFN26148_n26245),
	.B(n25128));
   NAND2xp33_ASAP7_75t_SRAM U24201 (.Y(n17674),
	.A(n25076),
	.B(n26243));
   NAND2xp33_ASAP7_75t_SRAM U24202 (.Y(n18788),
	.A(FE_OCPN27394_n26223),
	.B(n24721));
   NAND2xp33_ASAP7_75t_SRAM U24203 (.Y(n21920),
	.A(FE_OCPN27435_n26790),
	.B(n21918));
   NAND2xp33_ASAP7_75t_SRAM U24204 (.Y(n21870),
	.A(n24553),
	.B(n25975));
   NAND3x1_ASAP7_75t_SL U24205 (.Y(n25605),
	.A(FE_OCPN29422_n23397),
	.B(n23368),
	.C(n24559));
   NAND2xp33_ASAP7_75t_SRAM U24206 (.Y(n21813),
	.A(FE_OCPN29390_n26528),
	.B(n26272));
   NAND2xp33_ASAP7_75t_SRAM U24207 (.Y(n23897),
	.A(n26052),
	.B(n27085));
   NAND2xp33_ASAP7_75t_SRAM U24209 (.Y(n18733),
	.A(n18731),
	.B(n26287));
   NAND2xp33_ASAP7_75t_SRAM U24210 (.Y(n23624),
	.A(n25451),
	.B(n26210));
   NAND2xp33_ASAP7_75t_SRAM U24211 (.Y(n17600),
	.A(n24286),
	.B(FE_OFN26058_w3_1));
   NAND2xp5_ASAP7_75t_L U24212 (.Y(n23971),
	.A(n23639),
	.B(n23929));
   NAND2xp33_ASAP7_75t_SRAM U24213 (.Y(n25500),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_78_));
   OAI21xp33_ASAP7_75t_SRAM U24215 (.Y(n24237),
	.A1(text_in_r_70_),
	.A2(n24236),
	.B(n24235));
   NAND2xp33_ASAP7_75t_SRAM U24216 (.Y(n14089),
	.A(n16055),
	.B(FE_OFN28468_ld));
   NAND2xp33_ASAP7_75t_SRAM U24217 (.Y(n15272),
	.A(n16053),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24218 (.Y(n13799),
	.A(FE_OFN27218_n14745),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24219 (.Y(n14009),
	.A(n15902),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24220 (.Y(n16124),
	.A(n16268),
	.B(FE_OFN25_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24221 (.Y(n14743),
	.A(n16048),
	.B(FE_OFN26_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24222 (.Y(n14473),
	.A(n16080),
	.B(FE_OFN25_n16125));
   OAI21xp33_ASAP7_75t_SL U24223 (.Y(n16171),
	.A1(n16168),
	.A2(n16167),
	.B(n16166));
   OAI22xp33_ASAP7_75t_SRAM U24224 (.Y(n13270),
	.A1(n13269),
	.A2(n16285),
	.B1(n16286),
	.B2(n16285));
   NAND2xp33_ASAP7_75t_SRAM U24225 (.Y(n13232),
	.A(FE_OFN28469_ld),
	.B(n13231));
   NAND2xp33_ASAP7_75t_SRAM U24226 (.Y(n13236),
	.A(n13235),
	.B(FE_OFN28457_ld));
   NAND2xp33_ASAP7_75t_SRAM U24227 (.Y(n13200),
	.A(n13199),
	.B(FE_OFN26139_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24228 (.Y(n13040),
	.A(FE_OFN28470_ld),
	.B(n13039));
   NAND2xp33_ASAP7_75t_SRAM U24229 (.Y(n13208),
	.A(n13207),
	.B(FE_OFN22_n16125));
   NAND2xp33_ASAP7_75t_SRAM U24230 (.Y(n13056),
	.A(FE_OFN22_n16125),
	.B(n13055));
   NAND2xp33_ASAP7_75t_SRAM U24231 (.Y(n13062),
	.A(FE_OFN28459_ld),
	.B(n13061));
   NAND2xp33_ASAP7_75t_SRAM U24232 (.Y(n13078),
	.A(FE_OFN28459_ld),
	.B(n13077));
   NAND2xp33_ASAP7_75t_SRAM U24233 (.Y(n13202),
	.A(n13201),
	.B(FE_OFN28463_ld));
   NAND2xp33_ASAP7_75t_SRAM U24234 (.Y(n13098),
	.A(FE_OFN28457_ld),
	.B(n13097));
   NAND2xp33_ASAP7_75t_SRAM U24235 (.Y(n13178),
	.A(n13177),
	.B(FE_OFN28464_ld));
   NAND2xp33_ASAP7_75t_SRAM U24236 (.Y(n13024),
	.A(FE_OFN27_n16125),
	.B(n13023));
   NAND2xp33_ASAP7_75t_SRAM U24237 (.Y(n13180),
	.A(n13179),
	.B(FE_OFN28457_ld));
   NAND2xp33_ASAP7_75t_SRAM U24238 (.Y(n13112),
	.A(FE_OFN28471_ld),
	.B(n13111));
   NAND2xp33_ASAP7_75t_SRAM U24239 (.Y(n13140),
	.A(FE_OFN28460_ld),
	.B(n13139));
   NAND2xp33_ASAP7_75t_SRAM U24240 (.Y(n13118),
	.A(FE_OFN28460_ld),
	.B(n13117));
   NAND2xp33_ASAP7_75t_SRAM U24241 (.Y(n13266),
	.A(n13265),
	.B(FE_OFN28467_ld));
   OAI21xp33_ASAP7_75t_SL U24242 (.Y(n633),
	.A1(n15916),
	.A2(FE_OFN28732_n),
	.B(n15373));
   OAI21xp33_ASAP7_75t_SRAM U24243 (.Y(n533),
	.A1(key_111_),
	.A2(FE_OFN26_n16125),
	.B(n14249));
   OAI21xp33_ASAP7_75t_SRAM U24244 (.Y(n548),
	.A1(key_118_),
	.A2(FE_OFN26_n16125),
	.B(n14184));
   OAI21xp33_ASAP7_75t_SRAM U24245 (.Y(n563),
	.A1(key_124_),
	.A2(FE_OFN28461_ld),
	.B(n13938));
   OAI21xp33_ASAP7_75t_SRAM U24246 (.Y(n578),
	.A1(key_98_),
	.A2(FE_OFN28471_ld),
	.B(n13410));
   OAI21xp33_ASAP7_75t_SRAM U24247 (.Y(n593),
	.A1(key_104_),
	.A2(FE_OFN26_n16125),
	.B(n15657));
   OAI21xp33_ASAP7_75t_SRAM U24248 (.Y(n608),
	.A1(key_113_),
	.A2(FE_OFN26_n16125),
	.B(n14743));
   OAI21xp33_ASAP7_75t_SL U24249 (.Y(n625),
	.A1(n16086),
	.A2(n25596),
	.B(n16085));
   NAND2xp33_ASAP7_75t_SRAM U24250 (.Y(n665),
	.A(n13270),
	.B(FE_OFN28461_ld));
   OAI21xp33_ASAP7_75t_SRAM U24251 (.Y(n693),
	.A1(text_in_13_),
	.A2(FE_OFN28457_ld),
	.B(n13236));
   OAI21xp33_ASAP7_75t_SRAM U24252 (.Y(n723),
	.A1(text_in_28_),
	.A2(FE_OFN28470_ld),
	.B(n13040));
   OAI21xp33_ASAP7_75t_SRAM U24253 (.Y(n753),
	.A1(text_in_43_),
	.A2(FE_OFN22_n16125),
	.B(n13056));
   OAI21xp33_ASAP7_75t_SRAM U24254 (.Y(n783),
	.A1(text_in_58_),
	.A2(FE_OFN28459_ld),
	.B(n13078));
   OAI21xp33_ASAP7_75t_SRAM U24255 (.Y(n813),
	.A1(text_in_73_),
	.A2(FE_OFN28457_ld),
	.B(n13098));
   OAI21xp33_ASAP7_75t_SRAM U24256 (.Y(n843),
	.A1(text_in_88_),
	.A2(FE_OFN27_n16125),
	.B(n13024));
   OAI21xp33_ASAP7_75t_SRAM U24257 (.Y(n873),
	.A1(text_in_103_),
	.A2(FE_OFN28471_ld),
	.B(n13112));
   OAI21xp33_ASAP7_75t_SRAM U24258 (.Y(n903),
	.A1(text_in_118_),
	.A2(FE_OFN28460_ld),
	.B(n13118));
   OAI21xp33_ASAP7_75t_SRAM U24259 (.Y(n27009),
	.A1(n22597),
	.A2(n27006),
	.B(FE_OFN27152_n17315));
   NOR2xp33_ASAP7_75t_SRAM U24260 (.Y(n26974),
	.A(n26973),
	.B(n26972));
   NOR2xp33_ASAP7_75t_SRAM U24261 (.Y(n25085),
	.A(n25083),
	.B(n25082));
   NOR2xp33_ASAP7_75t_SRAM U24262 (.Y(n25055),
	.A(FE_OCPN27423_sa01_0),
	.B(FE_OCPN29475_n25054));
   NOR2xp33_ASAP7_75t_L U24263 (.Y(n23823),
	.A(FE_OCPN28353_n18534),
	.B(n23819));
   OAI21xp33_ASAP7_75t_SL U24264 (.Y(n23248),
	.A1(n23247),
	.A2(n23246),
	.B(n17473));
   NOR2xp33_ASAP7_75t_SRAM U24265 (.Y(n23184),
	.A(n18166),
	.B(n23183));
   OAI21xp33_ASAP7_75t_SL U24266 (.Y(n21825),
	.A1(n21821),
	.A2(FE_OCPN27496_n21820),
	.B(FE_PSN8325_FE_OFN28811_n19170));
   NOR2xp33_ASAP7_75t_SRAM U24267 (.Y(n21609),
	.A(n22156),
	.B(n21608));
   OAI21xp33_ASAP7_75t_SRAM U24268 (.Y(n20579),
	.A1(n22233),
	.A2(n22781),
	.B(FE_OFN25907_sa12_2));
   NOR2xp33_ASAP7_75t_SRAM U24269 (.Y(n19363),
	.A(FE_OCPN28202_n16991),
	.B(FE_OFN27186_sa13_4));
   OAI21xp33_ASAP7_75t_SL U24270 (.Y(n19224),
	.A1(n17445),
	.A2(n22512),
	.B(FE_OCPN27625_sa11_5));
   OAI21xp33_ASAP7_75t_SL U24271 (.Y(n19009),
	.A1(n19000),
	.A2(n20931),
	.B(FE_OCPN27986_n18970));
   NOR2xp33_ASAP7_75t_SRAM U24272 (.Y(n18838),
	.A(FE_OCPN29579_n18837),
	.B(FE_OCPN28423_n18836));
   OAI21xp5_ASAP7_75t_L U24273 (.Y(n20674),
	.A1(n23855),
	.A2(n23831),
	.B(FE_OCPN27580_n));
   OAI21xp33_ASAP7_75t_R U24275 (.Y(n18111),
	.A1(n18108),
	.A2(n18107),
	.B(FE_OCPN27546_sa33_4));
   OAI21xp5_ASAP7_75t_SL U24276 (.Y(n21059),
	.A1(FE_OFN25986_n21012),
	.A2(FE_OCPN27918_n21042),
	.B(n21738));
   OAI21xp5_ASAP7_75t_L U24278 (.Y(n21727),
	.A1(n21715),
	.A2(n21524),
	.B(FE_OFN21730_sa03_3));
   NOR2xp33_ASAP7_75t_SRAM U24279 (.Y(n17844),
	.A(FE_OCPN27556_n17843),
	.B(n16762));
   OAI21xp5_ASAP7_75t_L U24280 (.Y(n17748),
	.A1(FE_OCPN28357_n22882),
	.A2(n20988),
	.B(FE_OCPN8230_n20993));
   OAI21xp5_ASAP7_75t_L U24281 (.Y(n22145),
	.A1(FE_OFN28818_n17602),
	.A2(n20481),
	.B(FE_OFN25917_n21591));
   OAI21xp33_ASAP7_75t_R U24282 (.Y(n17708),
	.A1(n19938),
	.A2(n22368),
	.B(n22392));
   OAI21xp33_ASAP7_75t_SRAM U24283 (.Y(n17490),
	.A1(n23247),
	.A2(n19222),
	.B(n17473));
   OAI22xp33_ASAP7_75t_SRAM U24284 (.Y(n17246),
	.A1(n12998),
	.A2(n24086),
	.B1(FE_OFN28835_n),
	.B2(n24086));
   OAI21xp5_ASAP7_75t_L U24285 (.Y(n16810),
	.A1(FE_OFN16153_n16747),
	.A2(n20301),
	.B(FE_OCPN28298_n));
   OAI21xp33_ASAP7_75t_L U24286 (.Y(n23993),
	.A1(n17221),
	.A2(n24726),
	.B(FE_OFN29204_sa10_2));
   NOR2xp33_ASAP7_75t_L U24287 (.Y(n15798),
	.A(n15876),
	.B(n13726));
   OAI21xp33_ASAP7_75t_L U24288 (.Y(n14847),
	.A1(n14846),
	.A2(n15609),
	.B(FE_OFN26073_n));
   NOR2xp33_ASAP7_75t_SL U24289 (.Y(n14775),
	.A(FE_OFN16352_n14289),
	.B(n14778));
   OAI21xp33_ASAP7_75t_SRAM U24290 (.Y(n14622),
	.A1(FE_OFN26641_w3_14),
	.A2(n13804),
	.B(n15447));
   OAI21xp5_ASAP7_75t_SL U24291 (.Y(n13918),
	.A1(n12994),
	.A2(n13917),
	.B(n14361));
   OAI21xp33_ASAP7_75t_SRAM U24292 (.Y(n13593),
	.A1(FE_OFN25875_n15227),
	.A2(n13581),
	.B(n15185));
   NOR2xp33_ASAP7_75t_L U24293 (.Y(n13381),
	.A(FE_OFN25895_n13662),
	.B(n15187));
   OAI21xp33_ASAP7_75t_SRAM U24294 (.Y(n660),
	.A1(n13274),
	.A2(n16284),
	.B(n13273));
   NAND2xp33_ASAP7_75t_SRAM U24295 (.Y(n22237),
	.A(n23603),
	.B(FE_OCPN29477_sa12_5));
   NAND2xp33_ASAP7_75t_SRAM U24296 (.Y(n19296),
	.A(FE_OCPN27986_n18970),
	.B(FE_OFN29001_n23491));
   OAI22xp33_ASAP7_75t_SRAM U24297 (.Y(n15483),
	.A1(FE_OFN27214_w3_17),
	.A2(n15471),
	.B1(n15729),
	.B2(n15471));
   OAI22xp5_ASAP7_75t_L U24298 (.Y(n15021),
	.A1(n13736),
	.A2(FE_OFN26110_n15848),
	.B1(n15635),
	.B2(FE_OFN26110_n15848));
   OAI22xp33_ASAP7_75t_SL U24299 (.Y(n14962),
	.A1(FE_OFN26564_n),
	.A2(n14926),
	.B1(n15993),
	.B2(n14926));
   NOR3xp33_ASAP7_75t_SRAM U24300 (.Y(n13003),
	.A(dcnt_1_),
	.B(dcnt_0_),
	.C(dcnt_2_));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24301 (.Y(n13000),
	.A1(dcnt_0_),
	.A2(dcnt_1_),
	.B(dcnt_2_),
	.C(n13003));
   NOR2xp33_ASAP7_75t_SRAM U24302 (.Y(n16281),
	.A(dcnt_2_),
	.B(dcnt_3_));
   NOR3xp33_ASAP7_75t_SRAM U24303 (.Y(n13001),
	.A(n13000),
	.B(ld),
	.C(n16281));
   INVxp33_ASAP7_75t_SRAM U24304 (.Y(n13002),
	.A(dcnt_3_));
   NOR2xp33_ASAP7_75t_SRAM U24305 (.Y(n13004),
	.A(n13003),
	.B(n13002));
   NOR3xp33_ASAP7_75t_SRAM U24306 (.Y(n16282),
	.A(n13269),
	.B(ld),
	.C(u0_r0_rcnt_3_));
   NAND3xp33_ASAP7_75t_SRAM U24307 (.Y(n13005),
	.A(u0_r0_rcnt_1_),
	.B(u0_r0_rcnt_0_),
	.C(u0_r0_rcnt_2_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24308 (.Y(n13273),
	.A1(u0_r0_rcnt_1_),
	.A2(u0_r0_rcnt_0_),
	.B(u0_r0_rcnt_2_),
	.C(n13005));
   NOR2xp33_ASAP7_75t_SRAM U24309 (.Y(n13006),
	.A(dcnt_0_),
	.B(dcnt_1_));
   OAI22xp33_ASAP7_75t_SRAM U24310 (.Y(n13008),
	.A1(dcnt_1_),
	.A2(n13006),
	.B1(dcnt_0_),
	.B2(n13006));
   NOR2xp33_ASAP7_75t_SRAM U24311 (.Y(n13009),
	.A(n13008),
	.B(n13007));
   OAI21xp33_ASAP7_75t_SRAM U24312 (.Y(n664),
	.A1(u0_r0_rcnt_2_),
	.A2(n16285),
	.B(n662));
   INVxp33_ASAP7_75t_SRAM U24313 (.Y(n13011),
	.A(text_in_r_105_));
   INVxp33_ASAP7_75t_SRAM U24314 (.Y(n13013),
	.A(text_in_r_123_));
   INVxp33_ASAP7_75t_SRAM U24315 (.Y(n13015),
	.A(text_in_r_119_));
   INVxp33_ASAP7_75t_SRAM U24316 (.Y(n13017),
	.A(text_in_r_89_));
   INVxp33_ASAP7_75t_SRAM U24317 (.Y(n13019),
	.A(text_in_r_126_));
   INVxp33_ASAP7_75t_SRAM U24318 (.Y(n13021),
	.A(text_in_r_90_));
   INVxp33_ASAP7_75t_SRAM U24319 (.Y(n13023),
	.A(text_in_r_88_));
   INVxp33_ASAP7_75t_SRAM U24320 (.Y(n13027),
	.A(text_in_r_106_));
   INVxp33_ASAP7_75t_SRAM U24321 (.Y(n13029),
	.A(text_in_r_91_));
   INVxp33_ASAP7_75t_SRAM U24322 (.Y(n13031),
	.A(text_in_r_107_));
   OAI21xp33_ASAP7_75t_SRAM U24323 (.Y(n921),
	.A1(text_in_127_),
	.A2(FE_OFN28468_ld),
	.B(n13034));
   INVxp33_ASAP7_75t_SRAM U24324 (.Y(n13043),
	.A(text_in_r_21_));
   INVxp33_ASAP7_75t_SRAM U24325 (.Y(n13049),
	.A(text_in_r_38_));
   INVxp33_ASAP7_75t_SRAM U24326 (.Y(n13061),
	.A(text_in_r_50_));
   INVxp33_ASAP7_75t_SRAM U24327 (.Y(n13067),
	.A(text_in_r_34_));
   INVxp33_ASAP7_75t_SRAM U24328 (.Y(n13073),
	.A(text_in_r_55_));
   INVxp33_ASAP7_75t_SRAM U24329 (.Y(n13085),
	.A(text_in_r_66_));
   INVxp33_ASAP7_75t_SRAM U24330 (.Y(n13095),
	.A(text_in_r_72_));
   INVxp33_ASAP7_75t_SRAM U24331 (.Y(n13101),
	.A(text_in_r_74_));
   INVxp33_ASAP7_75t_SRAM U24332 (.Y(n13103),
	.A(text_in_r_75_));
   INVxp33_ASAP7_75t_SRAM U24333 (.Y(n13115),
	.A(text_in_r_104_));
   INVxp33_ASAP7_75t_SRAM U24334 (.Y(n13123),
	.A(text_in_r_84_));
   INVxp33_ASAP7_75t_SRAM U24335 (.Y(n13131),
	.A(text_in_r_124_));
   INVxp33_ASAP7_75t_SRAM U24336 (.Y(n13139),
	.A(text_in_r_110_));
   OAI21xp33_ASAP7_75t_SRAM U24337 (.Y(n691),
	.A1(text_in_12_),
	.A2(FE_OFN28457_ld),
	.B(n13146));
   OAI21xp33_ASAP7_75t_SRAM U24338 (.Y(n697),
	.A1(text_in_15_),
	.A2(FE_OFN28457_ld),
	.B(n13148));
   OAI21xp33_ASAP7_75t_SRAM U24339 (.Y(n685),
	.A1(text_in_9_),
	.A2(FE_OFN28457_ld),
	.B(n13150));
   OAI21xp33_ASAP7_75t_SRAM U24340 (.Y(n689),
	.A1(text_in_11_),
	.A2(FE_OFN28457_ld),
	.B(n13152));
   OAI21xp33_ASAP7_75t_SRAM U24341 (.Y(n695),
	.A1(text_in_14_),
	.A2(FE_OFN28457_ld),
	.B(n13154));
   INVxp33_ASAP7_75t_SRAM U24342 (.Y(n13155),
	.A(text_in_r_10_));
   OAI21xp33_ASAP7_75t_SRAM U24343 (.Y(n687),
	.A1(text_in_10_),
	.A2(FE_OFN28457_ld),
	.B(n13156));
   INVxp33_ASAP7_75t_SRAM U24344 (.Y(n13159),
	.A(text_in_r_4_));
   INVxp33_ASAP7_75t_SRAM U24345 (.Y(n13167),
	.A(text_in_r_111_));
   INVxp33_ASAP7_75t_SRAM U24346 (.Y(n13169),
	.A(text_in_r_101_));
   INVxp33_ASAP7_75t_SRAM U24347 (.Y(n13175),
	.A(text_in_r_78_));
   INVxp33_ASAP7_75t_SRAM U24348 (.Y(n13179),
	.A(text_in_r_95_));
   INVxp33_ASAP7_75t_SRAM U24349 (.Y(n13181),
	.A(text_in_r_61_));
   INVxp33_ASAP7_75t_SRAM U24350 (.Y(n13183),
	.A(text_in_r_24_));
   INVxp33_ASAP7_75t_SRAM U24351 (.Y(n13187),
	.A(text_in_r_47_));
   INVxp33_ASAP7_75t_SRAM U24352 (.Y(n13189),
	.A(text_in_r_53_));
   INVxp33_ASAP7_75t_SRAM U24353 (.Y(n13191),
	.A(text_in_r_26_));
   INVxp33_ASAP7_75t_SRAM U24354 (.Y(n13195),
	.A(text_in_r_32_));
   INVxp33_ASAP7_75t_SRAM U24355 (.Y(n13197),
	.A(text_in_r_116_));
   INVxp33_ASAP7_75t_SRAM U24356 (.Y(n13199),
	.A(text_in_r_20_));
   INVxp33_ASAP7_75t_SRAM U24357 (.Y(n13201),
	.A(text_in_r_65_));
   INVxp33_ASAP7_75t_SRAM U24358 (.Y(n13203),
	.A(text_in_r_93_));
   INVxp33_ASAP7_75t_SRAM U24359 (.Y(n13205),
	.A(text_in_r_48_));
   INVxp33_ASAP7_75t_SRAM U24360 (.Y(n13207),
	.A(text_in_r_35_));
   INVxp33_ASAP7_75t_SRAM U24361 (.Y(n13209),
	.A(text_in_r_52_));
   INVxp33_ASAP7_75t_SRAM U24362 (.Y(n13211),
	.A(text_in_r_56_));
   INVxp33_ASAP7_75t_SRAM U24363 (.Y(n13217),
	.A(text_in_r_33_));
   INVxp33_ASAP7_75t_SRAM U24364 (.Y(n13219),
	.A(text_in_r_115_));
   INVxp33_ASAP7_75t_SRAM U24365 (.Y(n13223),
	.A(text_in_r_19_));
   INVxp33_ASAP7_75t_SRAM U24366 (.Y(n13227),
	.A(text_in_r_7_));
   INVxp33_ASAP7_75t_SRAM U24367 (.Y(n13231),
	.A(text_in_r_6_));
   INVxp33_ASAP7_75t_SRAM U24368 (.Y(n13233),
	.A(text_in_r_16_));
   INVxp33_ASAP7_75t_SRAM U24369 (.Y(n13235),
	.A(text_in_r_13_));
   OAI21xp33_ASAP7_75t_SRAM U24370 (.Y(n671),
	.A1(text_in_2_),
	.A2(FE_OFN28470_ld),
	.B(n13238));
   INVxp33_ASAP7_75t_SRAM U24371 (.Y(n13239),
	.A(text_in_r_36_));
   INVxp33_ASAP7_75t_SRAM U24372 (.Y(n13241),
	.A(text_in_r_17_));
   INVxp33_ASAP7_75t_SRAM U24373 (.Y(n13243),
	.A(text_in_r_113_));
   INVxp33_ASAP7_75t_SRAM U24374 (.Y(n13245),
	.A(text_in_r_109_));
   INVxp33_ASAP7_75t_SRAM U24375 (.Y(n13247),
	.A(text_in_r_96_));
   INVxp33_ASAP7_75t_SRAM U24376 (.Y(n13249),
	.A(text_in_r_97_));
   INVxp33_ASAP7_75t_SRAM U24377 (.Y(n13251),
	.A(text_in_r_100_));
   INVxp33_ASAP7_75t_SRAM U24378 (.Y(n13255),
	.A(text_in_r_1_));
   OAI21xp33_ASAP7_75t_SRAM U24379 (.Y(n669),
	.A1(text_in_1_),
	.A2(FE_OFN28470_ld),
	.B(n13256));
   INVxp33_ASAP7_75t_SRAM U24380 (.Y(n13257),
	.A(text_in_r_0_));
   OAI21xp33_ASAP7_75t_SRAM U24381 (.Y(n667),
	.A1(text_in_0_),
	.A2(FE_OFN28469_ld),
	.B(n13258));
   INVxp33_ASAP7_75t_SRAM U24382 (.Y(n13263),
	.A(text_in_r_42_));
   INVxp33_ASAP7_75t_SRAM U24383 (.Y(n13265),
	.A(text_in_r_125_));
   NAND3xp33_ASAP7_75t_SRAM U24384 (.Y(n13267),
	.A(n16287),
	.B(n16285),
	.C(u0_r0_rcnt_2_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24385 (.Y(n13271),
	.A1(n16285),
	.A2(u0_r0_rcnt_2_),
	.B(n16287),
	.C(n13267));
   NOR3xp33_ASAP7_75t_SRAM U24386 (.Y(n16283),
	.A(u0_r0_rcnt_0_),
	.B(ld),
	.C(u0_r0_rcnt_1_));
   NOR3xp33_ASAP7_75t_SRAM U24387 (.Y(n13268),
	.A(n663),
	.B(n13269),
	.C(n16286));
   OAI21xp33_ASAP7_75t_SRAM U24388 (.Y(n661),
	.A1(n16283),
	.A2(n13268),
	.B(n13273));
   NOR3xp33_ASAP7_75t_SRAM U24389 (.Y(n13274),
	.A(n665),
	.B(n13271),
	.C(n16286));
   INVxp33_ASAP7_75t_SRAM U24390 (.Y(n13272),
	.A(n16283));
   NOR3xp33_ASAP7_75t_SRAM U24391 (.Y(n16284),
	.A(n16287),
	.B(u0_r0_rcnt_2_),
	.C(n13272));
   A2O1A1Ixp33_ASAP7_75t_R U24393 (.Y(n13650),
	.A1(FE_OCPN27656_w3_25),
	.A2(FE_OFN27212_w3_30),
	.B(FE_OFN26049_w3_27),
	.C(n15205));
   NAND3xp33_ASAP7_75t_SL U24397 (.Y(n13673),
	.A(FE_OFN27208_w3_30),
	.B(FE_OCPN27655_w3_25),
	.C(n25675));
   NOR2xp33_ASAP7_75t_SL U24399 (.Y(n15201),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN27207_w3_30));
   NAND2xp33_ASAP7_75t_L U24400 (.Y(n13662),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN26048_w3_27));
   NOR3xp33_ASAP7_75t_L U24401 (.Y(n13646),
	.A(FE_OCPN29428_FE_OFN27131_w3_29),
	.B(FE_OCPN28096_w3_31),
	.C(FE_OFN27130_w3_28));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24402 (.Y(n13275),
	.A1(FE_OCPN29428_FE_OFN27131_w3_29),
	.A2(FE_OFN16201_n15197),
	.B(n13604),
	.C(FE_OCPN28096_w3_31));
   NAND2xp5_ASAP7_75t_SL U24403 (.Y(n13530),
	.A(FE_OFN27211_w3_30),
	.B(FE_OFN26051_w3_27));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24405 (.Y(n13286),
	.A1(n15155),
	.A2(FE_OFN28890_n),
	.B(n15197),
	.C(FE_OFN16451_n));
   A2O1A1Ixp33_ASAP7_75t_R U24406 (.Y(n13294),
	.A1(n15185),
	.A2(n13596),
	.B(n15203),
	.C(n13289));
   A2O1A1Ixp33_ASAP7_75t_R U24407 (.Y(n13292),
	.A1(FE_OFN28817_n),
	.A2(n13613),
	.B(n14504),
	.C(n13291));
   OAI21xp5_ASAP7_75t_L U24408 (.Y(n13301),
	.A1(FE_OCPN27655_w3_25),
	.A2(n14504),
	.B(n15203));
   OAI222xp33_ASAP7_75t_L U24409 (.Y(n13302),
	.A1(n13713),
	.A2(n13301),
	.B1(n15156),
	.B2(n13301),
	.C1(FE_OFN16437_n),
	.C2(n13301));
   OA21x2_ASAP7_75t_SRAM U24410 (.Y(n13304),
	.A1(n15200),
	.A2(n13677),
	.B(n13302));
   A2O1A1Ixp33_ASAP7_75t_R U24411 (.Y(n13318),
	.A1(FE_OFN27212_w3_30),
	.A2(FE_OCPN29547_n15183),
	.B(n13309),
	.C(n13308));
   O2A1O1Ixp33_ASAP7_75t_SL U24412 (.Y(n13316),
	.A1(n14535),
	.A2(n13428),
	.B(n13315),
	.C(n15259));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24413 (.Y(n13319),
	.A1(FE_OFN25893_n15214),
	.A2(FE_OFN28858_FE_OCPN27664_w3_25),
	.B(n14504),
	.C(n15259));
   A2O1A1Ixp33_ASAP7_75t_L U24414 (.Y(n13331),
	.A1(n13595),
	.A2(n13333),
	.B(n13330),
	.C(w0_5_));
   OAI21xp33_ASAP7_75t_SRAM U24415 (.Y(n13335),
	.A1(FE_OCPN8232_FE_OFN27206_w3_30),
	.A2(FE_OFN28891_n),
	.B(FE_OFN25895_n13662));
   NOR2xp33_ASAP7_75t_R U24416 (.Y(n13337),
	.A(FE_OFN25966_n13646),
	.B(n13338));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24417 (.Y(n13336),
	.A1(FE_OFN27209_w3_30),
	.A2(FE_OFN27129_w3_28),
	.B(n15167),
	.C(n15183));
   OA21x2_ASAP7_75t_SRAM U24418 (.Y(n13339),
	.A1(n13336),
	.A2(FE_OCPN29571_n26355),
	.B(n13682));
   A2O1A1Ixp33_ASAP7_75t_L U24419 (.Y(n15223),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OCPN27656_w3_25),
	.B(FE_OFN27207_w3_30),
	.C(n15239));
   NOR2xp33_ASAP7_75t_SRAM U24420 (.Y(n13340),
	.A(n15223),
	.B(n13338));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24422 (.Y(n13346),
	.A1(FE_OFN16206_n15240),
	.A2(FE_OFN25895_n13662),
	.B(n15189),
	.C(n14516));
   NOR3xp33_ASAP7_75t_SRAM U24423 (.Y(n13344),
	.A(n13713),
	.B(FE_OCPN29571_n26355),
	.C(n13343));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24424 (.Y(n13345),
	.A1(n15146),
	.A2(n15209),
	.B(n15224),
	.C(n13344));
   NAND2xp5_ASAP7_75t_L U24425 (.Y(n13350),
	.A(n15155),
	.B(FE_OFN28456_n13348));
   OR2x2_ASAP7_75t_SRAM U24426 (.Y(n13352),
	.A(n15187),
	.B(n15156));
   NAND3xp33_ASAP7_75t_SRAM U24427 (.Y(n13360),
	.A(FE_OFN16206_n15240),
	.B(FE_OFN16159_w3_24),
	.C(FE_OFN16412_w3_26));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24428 (.Y(n13361),
	.A1(FE_OFN28817_n),
	.A2(n13360),
	.B(n15253),
	.C(n13669));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24429 (.Y(n13364),
	.A1(FE_OCPN27665_w3_25),
	.A2(FE_OFN16225_n15195),
	.B(FE_OFN25893_n15214),
	.C(n15259));
   OAI22xp33_ASAP7_75t_L U24430 (.Y(n13481),
	.A1(FE_OFN27210_w3_30),
	.A2(n14559),
	.B1(FE_OFN28929_n15182),
	.B2(n14559));
   OAI21xp33_ASAP7_75t_SL U24431 (.Y(n13540),
	.A1(FE_OFN28859_FE_OCPN27664_w3_25),
	.A2(FE_OFN27212_w3_30),
	.B(FE_OFN28817_n));
   A2O1A1Ixp33_ASAP7_75t_L U24432 (.Y(n13380),
	.A1(n15200),
	.A2(n13502),
	.B(n13379),
	.C(n13378));
   A2O1A1Ixp33_ASAP7_75t_L U24433 (.Y(n13403),
	.A1(FE_OFN26059_n),
	.A2(n13481),
	.B(n13380),
	.C(n15263));
   NOR2xp33_ASAP7_75t_R U24434 (.Y(n13385),
	.A(FE_OFN16437_n),
	.B(n13381));
   NAND2xp33_ASAP7_75t_SL U24435 (.Y(n13384),
	.A(n13665),
	.B(FE_OFN26567_n));
   O2A1O1Ixp33_ASAP7_75t_L U24436 (.Y(n13397),
	.A1(n13390),
	.A2(FE_OFN28453_n13348),
	.B(n13389),
	.C(n15238));
   A2O1A1Ixp33_ASAP7_75t_SL U24437 (.Y(n13393),
	.A1(n15254),
	.A2(n13692),
	.B(n13392),
	.C(n13391));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24438 (.Y(n13395),
	.A1(FE_OFN26049_w3_27),
	.A2(n15156),
	.B(n13394),
	.C(n13393));
   A2O1A1Ixp33_ASAP7_75t_L U24439 (.Y(n13407),
	.A1(n15271),
	.A2(n13409),
	.B(n13406),
	.C(w0_2_));
   NAND2xp33_ASAP7_75t_R U24440 (.Y(n13450),
	.A(n15209),
	.B(FE_OFN28455_n13348));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24441 (.Y(n13424),
	.A1(FE_OFN16437_n),
	.A2(n13420),
	.B(FE_OFN25966_n13646),
	.C(n13670));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24442 (.Y(n13427),
	.A1(FE_OFN27057_n13662),
	.A2(n14504),
	.B(n13636),
	.C(n14515));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24443 (.Y(n13445),
	.A1(FE_OFN16206_n15240),
	.A2(FE_OFN28817_n),
	.B(FE_OFN25875_n15227),
	.C(n13696));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24444 (.Y(n13438),
	.A1(FE_OFN27206_w3_30),
	.A2(FE_OFN28604_n14534),
	.B(n15257),
	.C(n15200));
   O2A1O1Ixp33_ASAP7_75t_SL U24445 (.Y(n13451),
	.A1(FE_OFN27206_w3_30),
	.A2(n14557),
	.B(n13596),
	.C(FE_OFN27085_n));
   OA21x2_ASAP7_75t_L U24446 (.Y(n13455),
	.A1(n15257),
	.A2(n14504),
	.B(n13452));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24447 (.Y(n13460),
	.A1(FE_OCPN28096_w3_31),
	.A2(n14500),
	.B(n13459),
	.C(n14480));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24448 (.Y(n13463),
	.A1(FE_OFN16437_n),
	.A2(n14516),
	.B(n13461),
	.C(n13556));
   A2O1A1Ixp33_ASAP7_75t_L U24449 (.Y(n13477),
	.A1(n13595),
	.A2(n13479),
	.B(n13476),
	.C(w0_1_));
   NOR2xp33_ASAP7_75t_SRAM U24450 (.Y(n13483),
	.A(FE_OFN16437_n),
	.B(FE_OFN25966_n13646));
   NOR2xp33_ASAP7_75t_SRAM U24451 (.Y(n13485),
	.A(n13484),
	.B(FE_OFN25966_n13646));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24452 (.Y(n13497),
	.A1(n15167),
	.A2(n14503),
	.B(n15188),
	.C(n13673));
   AND3x1_ASAP7_75t_SRAM U24453 (.Y(n13505),
	.A(n15205),
	.B(n15197),
	.C(FE_OFN25966_n13646));
   NOR2xp33_ASAP7_75t_R U24454 (.Y(n13504),
	.A(n13499),
	.B(n13505));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24456 (.Y(n13501),
	.A1(FE_OCPN28096_w3_31),
	.A2(n14515),
	.B(n13500),
	.C(FE_OCPN29428_FE_OFN27131_w3_29));
   OAI222xp33_ASAP7_75t_SRAM U24457 (.Y(n13526),
	.A1(n15159),
	.A2(n13514),
	.B1(FE_OFN28717_n15158),
	.B2(n13514),
	.C1(FE_OFN26059_n),
	.C2(n13514));
   OAI21xp5_ASAP7_75t_L U24458 (.Y(n14592),
	.A1(FE_OFN27211_w3_30),
	.A2(FE_OCPN27659_w3_25),
	.B(n15240));
   O2A1O1Ixp33_ASAP7_75t_SL U24459 (.Y(n13528),
	.A1(FE_OCPN27659_w3_25),
	.A2(n14535),
	.B(n13527),
	.C(FE_OFN27206_w3_30));
   A2O1A1Ixp33_ASAP7_75t_L U24460 (.Y(n13532),
	.A1(FE_OFN27222_n14593),
	.A2(n13531),
	.B(n13530),
	.C(n13529));
   A2O1A1Ixp33_ASAP7_75t_SL U24461 (.Y(n13546),
	.A1(n15263),
	.A2(n13548),
	.B(n13545),
	.C(w0_3_));
   NOR2xp33_ASAP7_75t_SRAM U24462 (.Y(n13550),
	.A(FE_OFN26049_w3_27),
	.B(n15155));
   NAND3xp33_ASAP7_75t_SRAM U24463 (.Y(n13557),
	.A(n13556),
	.B(n15156),
	.C(FE_OFN16193_n15200));
   A2O1A1Ixp33_ASAP7_75t_SL U24464 (.Y(n14562),
	.A1(n15145),
	.A2(n14593),
	.B(n13566),
	.C(FE_OFN27210_w3_30));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24465 (.Y(n13569),
	.A1(n14573),
	.A2(FE_OFN27210_w3_30),
	.B(n15179),
	.C(n14562));
   OA21x2_ASAP7_75t_SRAM U24466 (.Y(n13570),
	.A1(n14504),
	.A2(FE_OFN28817_n),
	.B(n13567));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24467 (.Y(n13575),
	.A1(n15159),
	.A2(FE_OFN28717_n15158),
	.B(FE_OFN28453_n13348),
	.C(n13574));
   NOR2xp33_ASAP7_75t_SRAM U24468 (.Y(n13578),
	.A(FE_OFN26552_n14545),
	.B(FE_OCPN29573_n15184));
   NOR2xp33_ASAP7_75t_SRAM U24469 (.Y(n13581),
	.A(FE_OFN25893_n15214),
	.B(n13596));
   A2O1A1Ixp33_ASAP7_75t_L U24470 (.Y(n13647),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OCPN27659_w3_25),
	.B(FE_OFN27207_w3_30),
	.C(FE_OFN16193_n15200));
   NOR2xp33_ASAP7_75t_SRAM U24471 (.Y(n13597),
	.A(FE_OCPN27656_w3_25),
	.B(FE_OFN27044_n15236));
   A2O1A1Ixp33_ASAP7_75t_L U24472 (.Y(n13631),
	.A1(n13634),
	.A2(n13633),
	.B(n13630),
	.C(w0_4_));
   NOR2xp33_ASAP7_75t_R U24473 (.Y(n13641),
	.A(n13437),
	.B(n13642));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24474 (.Y(n13639),
	.A1(n15205),
	.A2(FE_OFN28496_n15201),
	.B(FE_OFN28453_n13348),
	.C(n13638));
   OR2x2_ASAP7_75t_SRAM U24475 (.Y(n13644),
	.A(n13643),
	.B(n13642));
   OA21x2_ASAP7_75t_SRAM U24476 (.Y(n13651),
	.A1(n15201),
	.A2(n13648),
	.B(n13647));
   NOR2xp33_ASAP7_75t_SRAM U24477 (.Y(n13652),
	.A(n13650),
	.B(n13649));
   NOR2xp33_ASAP7_75t_SRAM U24478 (.Y(n13658),
	.A(FE_OCPN29547_n15183),
	.B(n14535));
   A2O1A1Ixp33_ASAP7_75t_R U24479 (.Y(n13674),
	.A1(n15257),
	.A2(n13673),
	.B(n15195),
	.C(n13672));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24480 (.Y(n13718),
	.A1(FE_OCPN29571_n26355),
	.A2(n13715),
	.B(n13714),
	.C(FE_OFN27130_w3_28));
   OAI22xp33_ASAP7_75t_SRAM U24481 (.Y(n13717),
	.A1(n14479),
	.A2(n13716),
	.B1(FE_OFN28455_n13348),
	.B2(n13716));
   OAI22xp33_ASAP7_75t_SRAM U24485 (.Y(n15092),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(n15636),
	.B1(FE_OFN28732_n),
	.B2(n15636));
   NAND3xp33_ASAP7_75t_SRAM U24490 (.Y(n13727),
	.A(n15859),
	.B(n15817),
	.C(FE_OCPN29537_FE_OFN28699_w3_6));
   OAI22xp33_ASAP7_75t_SRAM U24491 (.Y(n13732),
	.A1(FE_OCPN28072_w3_3),
	.A2(n15571),
	.B1(FE_OFN28732_n),
	.B2(n15571));
   NOR2x1p5_ASAP7_75t_SL U24492 (.Y(n15838),
	.A(FE_OFN28661_w3_7),
	.B(n13730));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24493 (.Y(n13731),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(FE_OFN28732_n),
	.B(n15080),
	.C(n15838));
   A2O1A1Ixp33_ASAP7_75t_R U24494 (.Y(n13733),
	.A1(FE_OFN26110_n15848),
	.A2(FE_OCPN28398_n15808),
	.B(n13732),
	.C(n13731));
   OAI21xp5_ASAP7_75t_R U24495 (.Y(n14838),
	.A1(FE_OFN28721_n),
	.A2(n14439),
	.B(n13736));
   OR2x2_ASAP7_75t_SRAM U24496 (.Y(n13737),
	.A(n15876),
	.B(n13775));
   OAI22x1_ASAP7_75t_SL U24498 (.Y(n15028),
	.A1(FE_OFN26591_w3_3),
	.A2(FE_OFN26531_n),
	.B1(FE_OFN26058_w3_1),
	.B2(FE_OFN26531_n));
   OAI21xp33_ASAP7_75t_L U24499 (.Y(n13742),
	.A1(n13729),
	.A2(n13741),
	.B(n15779));
   A2O1A1Ixp33_ASAP7_75t_L U24500 (.Y(n13745),
	.A1(FE_OFN27156_n),
	.A2(n25140),
	.B(n15040),
	.C(n13742));
   OAI21xp5_ASAP7_75t_R U24501 (.Y(n15010),
	.A1(FE_OFN26645_n),
	.A2(n13729),
	.B(n14442));
   NOR2xp33_ASAP7_75t_R U24502 (.Y(n13785),
	.A(n25140),
	.B(FE_OFN28691_n13725));
   NAND2xp33_ASAP7_75t_L U24503 (.Y(n13783),
	.A(FE_OFN28671_FE_OCPN28076),
	.B(n13736));
   O2A1O1Ixp5_ASAP7_75t_L U24504 (.Y(n13792),
	.A1(n13791),
	.A2(n13790),
	.B(n15896),
	.C(n13789));
   NAND3xp33_ASAP7_75t_SRAM U24505 (.Y(n13802),
	.A(n14159),
	.B(n15407),
	.C(n15922));
   NOR2x1p5_ASAP7_75t_SL U24507 (.Y(n15934),
	.A(n24755),
	.B(n14913));
   NOR2x1_ASAP7_75t_L U24509 (.Y(n15924),
	.A(n24755),
	.B(n25782));
   NAND2x2_ASAP7_75t_SL U24510 (.Y(n16012),
	.A(FE_OFN27115_n),
	.B(FE_OCPN29508_FE_OFN16184_w3_9));
   NOR2x1_ASAP7_75t_L U24511 (.Y(n13949),
	.A(FE_OFN26642_w3_14),
	.B(n16012));
   OR2x2_ASAP7_75t_SRAM U24513 (.Y(n13807),
	.A(n25782),
	.B(n14896));
   NOR2xp67_ASAP7_75t_L U24514 (.Y(n14695),
	.A(n14897),
	.B(n13949));
   NOR3x1_ASAP7_75t_L U24515 (.Y(n14924),
	.A(n25782),
	.B(FE_OFN27200_n),
	.C(n24755));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24516 (.Y(n13812),
	.A1(FE_OFN29017_n15921),
	.A2(FE_OFN26635_w3_14),
	.B(n13811),
	.C(n15447));
   NOR2x1p5_ASAP7_75t_SL U24517 (.Y(n14912),
	.A(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(FE_OCPN28408_FE_OFN16433_w3_11));
   NOR2x1_ASAP7_75t_SL U24518 (.Y(n14667),
	.A(n14912),
	.B(FE_OFN26636_w3_14));
   NOR3xp33_ASAP7_75t_SL U24519 (.Y(n16015),
	.A(n14913),
	.B(FE_OCPN29521_n24755),
	.C(n14667));
   NOR2x1_ASAP7_75t_SL U24520 (.Y(n15972),
	.A(FE_OCPN28407_FE_OFN16433_w3_11),
	.B(FE_OFN16459_n));
   OAI22xp5_ASAP7_75t_L U24521 (.Y(n13820),
	.A1(FE_OFN29018_n15921),
	.A2(n13816),
	.B1(FE_OFN109_n15994),
	.B2(n13816));
   OA21x2_ASAP7_75t_R U24522 (.Y(n13821),
	.A1(n14930),
	.A2(n14929),
	.B(n13818));
   NOR2x1p5_ASAP7_75t_SL U24523 (.Y(n15414),
	.A(FE_OFN27115_n),
	.B(FE_OCPN29508_FE_OFN16184_w3_9));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24525 (.Y(n13826),
	.A1(FE_OFN26639_w3_14),
	.A2(FE_OCPN28407_FE_OFN16433_w3_11),
	.B(n16016),
	.C(FE_OFN16459_n));
   A2O1A1Ixp33_ASAP7_75t_R U24526 (.Y(n13827),
	.A1(FE_OFN26624_n15376),
	.A2(FE_OCPN28407_FE_OFN16433_w3_11),
	.B(FE_OFN16459_n),
	.C(n13826));
   NOR2xp33_ASAP7_75t_R U24527 (.Y(n13836),
	.A(n14626),
	.B(n13837));
   NOR2xp33_ASAP7_75t_SRAM U24528 (.Y(n13838),
	.A(n15987),
	.B(n13837));
   NAND2xp5_ASAP7_75t_L U24529 (.Y(n15955),
	.A(FE_OCPN29536_FE_OFN8_w3_14),
	.B(n14912));
   NOR2xp33_ASAP7_75t_R U24530 (.Y(n13843),
	.A(FE_OFN27115_n),
	.B(FE_OCPN29570_n15423));
   NOR3xp33_ASAP7_75t_L U24531 (.Y(n14610),
	.A(FE_OFN109_n15994),
	.B(FE_OFN26642_w3_14),
	.C(FE_OFN28813_n15414));
   A2O1A1Ixp33_ASAP7_75t_L U24532 (.Y(n13845),
	.A1(n15936),
	.A2(n15959),
	.B(FE_OFN26007_n16010),
	.C(n14933));
   NAND2x1p5_ASAP7_75t_SL U24534 (.Y(n15514),
	.A(FE_OFN27096_n),
	.B(FE_OFN27214_w3_17));
   NAND2x1p5_ASAP7_75t_SL U24538 (.Y(n13868),
	.A(n15667),
	.B(FE_OFN28712_n));
   NAND3x2_ASAP7_75t_L U24540 (.Y(n13875),
	.A(w3_21_),
	.B(FE_OFN25909_w3_20),
	.C(w3_23_));
   NAND2x1_ASAP7_75t_SL U24541 (.Y(n15658),
	.A(FE_OFN28683_w3_21),
	.B(FE_OFN28712_n));
   NOR2xp33_ASAP7_75t_SRAM U24542 (.Y(n13872),
	.A(n14371),
	.B(n15739));
   OAI22xp33_ASAP7_75t_L U24545 (.Y(n15665),
	.A1(FE_OFN26091_n24663),
	.A2(n15347),
	.B1(FE_OFN26539_w3_19),
	.B2(n15347));
   NOR3x2_ASAP7_75t_SL U24546 (.Y(n13916),
	.A(FE_OFN29087_n),
	.B(FE_OFN28976_n),
	.C(FE_OCPN27987_FE_OFN4_w3_22));
   OAI21xp33_ASAP7_75t_SRAM U24547 (.Y(n13894),
	.A1(FE_OFN26053_n25415),
	.A2(n15296),
	.B(n13889));
   NOR2x1_ASAP7_75t_L U24549 (.Y(n15485),
	.A(FE_OFN28_w3_23),
	.B(FE_OFN28683_w3_21));
   O2A1O1Ixp5_ASAP7_75t_SL U24550 (.Y(n13891),
	.A1(FE_OFN27214_w3_17),
	.A2(FE_OFN26053_n25415),
	.B(FE_OFN6_w3_22),
	.C(n15739));
   OAI21xp33_ASAP7_75t_SRAM U24551 (.Y(n13893),
	.A1(FE_OFN26538_w3_19),
	.A2(FE_OCPN8264_n13890),
	.B(n13892));
   O2A1O1Ixp5_ASAP7_75t_SL U24552 (.Y(n15512),
	.A1(FE_OFN26535_w3_19),
	.A2(FE_OFN28977_n),
	.B(n15514),
	.C(FE_OFN27151_n));
   NOR2x1p5_ASAP7_75t_SL U24553 (.Y(n15713),
	.A(FE_OFN28551_FE_OFN26114_n),
	.B(n15512));
   NAND2xp5_ASAP7_75t_L U24554 (.Y(n13902),
	.A(n12994),
	.B(n14361));
   O2A1O1Ixp5_ASAP7_75t_SL U24556 (.Y(n15517),
	.A1(FE_OFN26539_w3_19),
	.A2(FE_OFN28706_n),
	.B(FE_OFN5_w3_22),
	.C(n15341));
   O2A1O1Ixp5_ASAP7_75t_SL U24558 (.Y(n15349),
	.A1(FE_OFN5_w3_22),
	.A2(FE_OFN26053_n25415),
	.B(FE_PSN8292_FE_OFN26041_w3_17),
	.C(n14369));
   A2O1A1Ixp33_ASAP7_75t_SL U24559 (.Y(n13934),
	.A1(n13936),
	.A2(n13867),
	.B(n13933),
	.C(n26375));
   NOR2xp33_ASAP7_75t_SRAM U24561 (.Y(n13940),
	.A(n16000),
	.B(n13941));
   O2A1O1Ixp5_ASAP7_75t_SL U24562 (.Y(n15963),
	.A1(FE_OFN27115_n),
	.A2(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(n16012),
	.C(FE_OCPN29535_FE_OFN8_w3_14));
   OAI22xp5_ASAP7_75t_R U24563 (.Y(n13952),
	.A1(n15936),
	.A2(FE_OFN29018_n15921),
	.B1(n15956),
	.B2(FE_OFN29018_n15921));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24564 (.Y(n15984),
	.A1(FE_OFN27115_n),
	.A2(FE_OCPN29508_FE_OFN16184_w3_9),
	.B(FE_OCPN29534_FE_OFN8_w3_14),
	.C(n15963));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24565 (.Y(n13950),
	.A1(FE_PSN8271_n15924),
	.A2(n13949),
	.B(n13985),
	.C(FE_OFN28715_w3_15));
   AND2x2_ASAP7_75t_R U24567 (.Y(n13962),
	.A(n13959),
	.B(n13958));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24568 (.Y(n13994),
	.A1(FE_OFN26635_w3_14),
	.A2(n15447),
	.B(FE_OFN26007_n16010),
	.C(FE_OFN29018_n15921));
   NOR2xp33_ASAP7_75t_R U24569 (.Y(n13969),
	.A(FE_OFN16459_n),
	.B(FE_OFN109_n15994));
   NOR2xp33_ASAP7_75t_SRAM U24570 (.Y(n13968),
	.A(FE_PSN8271_n15924),
	.B(n13969));
   NOR2xp33_ASAP7_75t_SRAM U24571 (.Y(n13970),
	.A(FE_OFN28856_n15450),
	.B(n13969));
   A2O1A1Ixp33_ASAP7_75t_R U24573 (.Y(n13978),
	.A1(n16000),
	.A2(n15999),
	.B(n16016),
	.C(n15998));
   OAI22xp33_ASAP7_75t_SRAM U24574 (.Y(n13984),
	.A1(FE_OCPN28296_n15386),
	.A2(FE_OFN109_n15994),
	.B1(FE_OFN26635_w3_14),
	.B2(FE_OFN109_n15994));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24575 (.Y(n13990),
	.A1(FE_OFN29017_n15921),
	.A2(FE_OFN27135_n15992),
	.B(n13984),
	.C(n15936));
   A2O1A1Ixp33_ASAP7_75t_L U24576 (.Y(n14000),
	.A1(n14971),
	.A2(n14002),
	.B(n13999),
	.C(w0_21_));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24577 (.Y(n14014),
	.A1(FE_OFN16426_w3_20),
	.A2(n15744),
	.B(n14013),
	.C(n25961));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24578 (.Y(n14028),
	.A1(FE_OFN5_w3_22),
	.A2(FE_OFN28623_n13874),
	.B(n14015),
	.C(n14014));
   NOR2xp33_ASAP7_75t_R U24579 (.Y(n14020),
	.A(n15485),
	.B(n14017));
   NOR2xp33_ASAP7_75t_SRAM U24581 (.Y(n14022),
	.A(n14021),
	.B(n14017));
   NOR2xp33_ASAP7_75t_R U24582 (.Y(n14035),
	.A(FE_OCPN28404_n13874),
	.B(n14036));
   OAI22xp33_ASAP7_75t_L U24583 (.Y(n15319),
	.A1(FE_OFN26091_n24663),
	.A2(n13916),
	.B1(FE_OFN28624_n13874),
	.B2(n13916));
   OAI21xp33_ASAP7_75t_L U24584 (.Y(n14303),
	.A1(FE_OFN26091_n24663),
	.A2(n15536),
	.B(n15674));
   A2O1A1Ixp33_ASAP7_75t_SL U24586 (.Y(n14085),
	.A1(n14087),
	.A2(n13867),
	.B(n14084),
	.C(n26811));
   OA21x2_ASAP7_75t_SRAM U24587 (.Y(n14094),
	.A1(n16016),
	.A2(n14159),
	.B(n14694));
   OA21x2_ASAP7_75t_SRAM U24588 (.Y(n14103),
	.A1(n15382),
	.A2(n15385),
	.B(n14623));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24589 (.Y(n14109),
	.A1(n15924),
	.A2(n14915),
	.B(n14108),
	.C(FE_OCPN29427_w3_15));
   NAND2xp5_ASAP7_75t_L U24590 (.Y(n14113),
	.A(n15455),
	.B(n14112));
   NOR2x1_ASAP7_75t_L U24591 (.Y(n15927),
	.A(FE_OCPN29536_FE_OFN8_w3_14),
	.B(n15972));
   OR3x1_ASAP7_75t_SRAM U24592 (.Y(n14119),
	.A(n16016),
	.B(n13804),
	.C(n14667));
   A2O1A1Ixp33_ASAP7_75t_SL U24593 (.Y(n14173),
	.A1(n15946),
	.A2(n14136),
	.B(n16026),
	.C(n14135));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24594 (.Y(n14170),
	.A1(FE_OCPN29536_FE_OFN8_w3_14),
	.A2(FE_OFN28856_n15450),
	.B(n14924),
	.C(n14137));
   OAI21xp33_ASAP7_75t_SRAM U24595 (.Y(n14150),
	.A1(FE_OCPN29534_FE_OFN8_w3_14),
	.A2(FE_OFN27115_n),
	.B(n15948));
   NOR2xp33_ASAP7_75t_SL U24596 (.Y(n14144),
	.A(FE_OFN28659_n15934),
	.B(n14927));
   OAI21xp5_ASAP7_75t_L U24597 (.Y(n15453),
	.A1(FE_OFN26642_w3_14),
	.A2(n14912),
	.B(n14159));
   A2O1A1Ixp33_ASAP7_75t_SL U24598 (.Y(n14167),
	.A1(FE_OFN26624_n15376),
	.A2(n14914),
	.B(n14166),
	.C(n14165));
   A2O1A1Ixp33_ASAP7_75t_SL U24599 (.Y(n14180),
	.A1(n14183),
	.A2(n14182),
	.B(n14179),
	.C(w0_22_));
   NOR3xp33_ASAP7_75t_SRAM U24600 (.Y(n14185),
	.A(FE_OFN25900_w3_4),
	.B(FE_OFN28695_n),
	.C(FE_OFN28661_w3_7));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24601 (.Y(n14831),
	.A1(n24831),
	.A2(FE_OCPN27978_w3_3),
	.B(FE_OFN28721_n),
	.C(n15842));
   NAND3xp33_ASAP7_75t_SRAM U24602 (.Y(n14188),
	.A(n14439),
	.B(n15569),
	.C(FE_OFN28695_n));
   A2O1A1Ixp33_ASAP7_75t_R U24603 (.Y(n14248),
	.A1(n15834),
	.A2(n14193),
	.B(n13730),
	.C(n14192));
   OAI21xp5_ASAP7_75t_L U24604 (.Y(n15020),
	.A1(FE_OFN28747_n),
	.A2(FE_OFN16195_n13771),
	.B(n14214));
   OAI21xp33_ASAP7_75t_SRAM U24605 (.Y(n15797),
	.A1(FE_OFN28747_n),
	.A2(n15817),
	.B(FE_OFN25912_n15848));
   A2O1A1Ixp33_ASAP7_75t_L U24606 (.Y(n14195),
	.A1(n15034),
	.A2(FE_OFN25897_w3_4),
	.B(n14194),
	.C(n15857));
   AND2x2_ASAP7_75t_SRAM U24607 (.Y(n14204),
	.A(n15823),
	.B(n15635));
   OAI22xp33_ASAP7_75t_SRAM U24608 (.Y(n14202),
	.A1(n15578),
	.A2(FE_OFN26084_n15106),
	.B1(n15876),
	.B2(FE_OFN26084_n15106));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24609 (.Y(n14240),
	.A1(n14439),
	.A2(FE_OFN28721_n),
	.B(n14845),
	.C(n14209));
   NAND2xp5_ASAP7_75t_SL U24610 (.Y(n14218),
	.A(n14212),
	.B(n14215));
   A2O1A1Ixp33_ASAP7_75t_SL U24611 (.Y(n15851),
	.A1(FE_OCPN8254_w3_3),
	.A2(n24831),
	.B(n15862),
	.C(FE_OFN28699_w3_6));
   A2O1A1Ixp33_ASAP7_75t_SL U24612 (.Y(n15847),
	.A1(FE_OFN29209_FE_OCPN27978_w3_3),
	.A2(FE_OFN28732_n),
	.B(FE_OFN28829_n),
	.C(n14985));
   NAND2xp33_ASAP7_75t_L U24613 (.Y(n14220),
	.A(FE_OFN28699_w3_6),
	.B(n15859));
   O2A1O1Ixp33_ASAP7_75t_SL U24614 (.Y(n14241),
	.A1(n14240),
	.A2(n14239),
	.B(n15896),
	.C(n14238));
   A2O1A1Ixp33_ASAP7_75t_SL U24615 (.Y(n14246),
	.A1(FE_OFN16411_n15884),
	.A2(n14248),
	.B(n14245),
	.C(w0_15_));
   A2O1A1Ixp33_ASAP7_75t_SL U24616 (.Y(n15899),
	.A1(FE_OFN16411_n15884),
	.A2(n14248),
	.B(n14247),
	.C(n14246));
   O2A1O1Ixp33_ASAP7_75t_SL U24617 (.Y(n15496),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(n15714),
	.B(n14766),
	.C(FE_OFN16352_n14289));
   O2A1O1Ixp33_ASAP7_75t_SL U24618 (.Y(n14327),
	.A1(FE_OFN28481_n15298),
	.A2(n14263),
	.B(n14361),
	.C(n14262));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24619 (.Y(n14265),
	.A1(FE_OFN4_w3_22),
	.A2(FE_OFN25915_n15514),
	.B(n13916),
	.C(n14264));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24620 (.Y(n14267),
	.A1(FE_OFN28976_n),
	.A2(n14806),
	.B(n14266),
	.C(FE_OFN28623_n13874));
   OAI22xp5_ASAP7_75t_L U24621 (.Y(n14398),
	.A1(FE_OFN26535_w3_19),
	.A2(n13868),
	.B1(FE_OFN28977_n),
	.B2(n13868));
   A2O1A1Ixp33_ASAP7_75t_L U24622 (.Y(n14278),
	.A1(n15694),
	.A2(n15719),
	.B(FE_OFN16352_n14289),
	.C(n14277));
   A2O1A1Ixp33_ASAP7_75t_SL U24623 (.Y(n14290),
	.A1(FE_OFN26091_n24663),
	.A2(FE_OFN28706_n),
	.B(FE_OFN26539_w3_19),
	.C(n15290));
   OA21x2_ASAP7_75t_L U24624 (.Y(n14293),
	.A1(n14795),
	.A2(n13875),
	.B(n14290));
   A2O1A1Ixp33_ASAP7_75t_SL U24625 (.Y(n14297),
	.A1(FE_OFN28977_n),
	.A2(FE_OFN27151_n),
	.B(n13916),
	.C(FE_OFN26535_w3_19));
   NOR2xp33_ASAP7_75t_SRAM U24626 (.Y(n14309),
	.A(FE_OFN27066_n13869),
	.B(n14310));
   NOR2xp33_ASAP7_75t_SRAM U24627 (.Y(n14311),
	.A(FE_OFN27214_w3_17),
	.B(n14310));
   OA21x2_ASAP7_75t_SRAM U24629 (.Y(n14353),
	.A1(n15674),
	.A2(FE_OFN16210_n13876),
	.B(n14351));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24630 (.Y(n14357),
	.A1(FE_OFN6_w3_22),
	.A2(n14778),
	.B(FE_OFN25915_n15514),
	.C(n15528));
   OAI21xp33_ASAP7_75t_L U24631 (.Y(n14773),
	.A1(FE_OFN6_w3_22),
	.A2(FE_OFN28623_n13874),
	.B(n14361));
   NOR2x1_ASAP7_75t_L U24632 (.Y(n15479),
	.A(FE_OFN26053_n25415),
	.B(n13868));
   OAI22xp33_ASAP7_75t_R U24633 (.Y(n14748),
	.A1(FE_OFN6_w3_22),
	.A2(n15534),
	.B1(FE_OFN27082_n25377),
	.B2(n15534));
   A2O1A1Ixp33_ASAP7_75t_L U24634 (.Y(n14370),
	.A1(FE_OCPN27928_FE_OFN4_w3_22),
	.A2(FE_OFN28706_n),
	.B(n14369),
	.C(n12994));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24635 (.Y(n14395),
	.A1(FE_OFN27151_n),
	.A2(FE_OFN25915_n15514),
	.B(n13916),
	.C(n15528));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24636 (.Y(n14399),
	.A1(n14398),
	.A2(n14397),
	.B(n15744),
	.C(n14396));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24637 (.Y(n14420),
	.A1(FE_OFN28662_w3_7),
	.A2(n13726),
	.B(FE_OFN28691_n13725),
	.C(n15589));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24638 (.Y(n14418),
	.A1(FE_OFN16195_n13771),
	.A2(FE_OFN28889_n15845),
	.B(n14417),
	.C(n14996));
   A2O1A1Ixp33_ASAP7_75t_SL U24639 (.Y(n15002),
	.A1(FE_OCPN27985_n24831),
	.A2(FE_OFN28699_w3_6),
	.B(FE_OFN25887_w3_3),
	.C(n15838));
   OAI22xp33_ASAP7_75t_R U24640 (.Y(n15568),
	.A1(FE_OFN28829_n),
	.A2(n14996),
	.B1(FE_OFN26057_w3_1),
	.B2(n14996));
   A2O1A1Ixp33_ASAP7_75t_L U24641 (.Y(n14427),
	.A1(FE_OFN26645_n),
	.A2(n15817),
	.B(n15813),
	.C(n15607));
   A2O1A1Ixp33_ASAP7_75t_L U24642 (.Y(n14436),
	.A1(FE_OFN25928_n15779),
	.A2(n15002),
	.B(n13741),
	.C(n14435));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24643 (.Y(n14464),
	.A1(FE_OFN28699_w3_6),
	.A2(n15862),
	.B(n15033),
	.C(n15619));
   OAI21xp5_ASAP7_75t_R U24644 (.Y(n14976),
	.A1(FE_OFN28721_n),
	.A2(n13736),
	.B(n14440));
   OAI22xp33_ASAP7_75t_L U24645 (.Y(n15843),
	.A1(n24831),
	.A2(FE_OFN26531_n),
	.B1(FE_OFN26591_w3_3),
	.B2(FE_OFN26531_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24646 (.Y(n14445),
	.A1(FE_OCPN27978_w3_3),
	.A2(FE_OFN28721_n),
	.B(n15843),
	.C(n15859));
   A2O1A1Ixp33_ASAP7_75t_L U24647 (.Y(n14443),
	.A1(FE_OCPN27978_w3_3),
	.A2(FE_OFN28732_n),
	.B(n15808),
	.C(n14441));
   OAI222xp33_ASAP7_75t_SL U24648 (.Y(n14448),
	.A1(FE_OFN26531_n),
	.A2(n15028),
	.B1(FE_OFN26058_w3_1),
	.B2(n15028),
	.C1(FE_OFN26591_w3_3),
	.C2(n15028));
   NOR2xp33_ASAP7_75t_L U24649 (.Y(n14451),
	.A(n14985),
	.B(n14452));
   OAI22xp33_ASAP7_75t_L U24650 (.Y(n15567),
	.A1(FE_OFN28721_n),
	.A2(n14986),
	.B1(FE_OCPN27978_w3_3),
	.B2(n14986));
   NOR2xp33_ASAP7_75t_SL U24651 (.Y(n14463),
	.A(n14462),
	.B(n14461));
   NOR2xp33_ASAP7_75t_SRAM U24652 (.Y(n14476),
	.A(FE_OFN27129_w3_28),
	.B(n15146));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24653 (.Y(n14482),
	.A1(FE_OFN27061_n15239),
	.A2(FE_OCPN29571_n26355),
	.B(n14481),
	.C(n14480));
   O2A1O1Ixp33_ASAP7_75t_L U24654 (.Y(n14551),
	.A1(n25675),
	.A2(FE_OCPN27655_w3_25),
	.B(FE_OFN27209_w3_30),
	.C(n15146));
   A2O1A1Ixp33_ASAP7_75t_L U24655 (.Y(n14505),
	.A1(n15203),
	.A2(n14504),
	.B(n14551),
	.C(n14503));
   NAND2xp33_ASAP7_75t_L U24656 (.Y(n14518),
	.A(n14515),
	.B(FE_OFN25875_n15227));
   NAND2xp33_ASAP7_75t_L U24657 (.Y(n14517),
	.A(n14544),
	.B(FE_OFN25875_n15227));
   OR2x2_ASAP7_75t_SRAM U24658 (.Y(n14522),
	.A(FE_OFN28602_n14534),
	.B(n15200));
   NAND2xp33_ASAP7_75t_SRAM U24659 (.Y(n14536),
	.A(FE_OFN27057_n13662),
	.B(FE_OFN28456_n13348));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24660 (.Y(n14550),
	.A1(n15155),
	.A2(FE_OFN26051_w3_27),
	.B(n15197),
	.C(FE_OFN16225_n15195));
   NOR2xp33_ASAP7_75t_R U24661 (.Y(n14549),
	.A(FE_OFN25966_n13646),
	.B(n14550));
   AND2x2_ASAP7_75t_R U24662 (.Y(n14552),
	.A(n14548),
	.B(n14547));
   NOR2xp33_ASAP7_75t_R U24663 (.Y(n14553),
	.A(n14551),
	.B(n14550));
   NOR2xp33_ASAP7_75t_L U24664 (.Y(n14558),
	.A(n14557),
	.B(n14556));
   A2O1A1Ixp33_ASAP7_75t_SL U24665 (.Y(n14563),
	.A1(FE_OFN28817_n),
	.A2(n15257),
	.B(n15203),
	.C(n14562));
   NOR2xp33_ASAP7_75t_R U24666 (.Y(n14577),
	.A(FE_OFN16193_n15200),
	.B(n14578));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24667 (.Y(n14576),
	.A1(FE_OFN27211_w3_30),
	.A2(FE_OCPN27659_w3_25),
	.B(n13596),
	.C(n14535));
   A2O1A1Ixp33_ASAP7_75t_SL U24668 (.Y(n14590),
	.A1(n14589),
	.A2(n14588),
	.B(n15238),
	.C(n14587));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24669 (.Y(n14596),
	.A1(FE_OFN27057_n13662),
	.A2(FE_OFN27222_n14593),
	.B(n14592),
	.C(n15238));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24670 (.Y(n14609),
	.A1(n16000),
	.A2(n15959),
	.B(FE_OFN26007_n16010),
	.C(n14608));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24671 (.Y(n14621),
	.A1(n14611),
	.A2(n14610),
	.B(FE_OCPN29564_n16012),
	.C(n14609));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24672 (.Y(n14656),
	.A1(FE_OFN26641_w3_14),
	.A2(n15447),
	.B(n13844),
	.C(n16015));
   AND2x2_ASAP7_75t_SRAM U24673 (.Y(n14631),
	.A(n14630),
	.B(n14919));
   NAND3xp33_ASAP7_75t_L U24674 (.Y(n14653),
	.A(n14637),
	.B(n14931),
	.C(n14636));
   A2O1A1Ixp33_ASAP7_75t_SL U24675 (.Y(n14652),
	.A1(n14695),
	.A2(n15956),
	.B(n14651),
	.C(n14650));
   NOR2xp33_ASAP7_75t_SRAM U24676 (.Y(n14668),
	.A(FE_OFN16459_n),
	.B(n16016));
   AND2x2_ASAP7_75t_SRAM U24677 (.Y(n14673),
	.A(n14670),
	.B(n14669));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24678 (.Y(n14677),
	.A1(FE_OFN26642_w3_14),
	.A2(FE_OCPN29509_FE_OFN16184_w3_9),
	.B(FE_OFN28758_n15422),
	.C(n15383));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24679 (.Y(n14737),
	.A1(FE_OFN26642_w3_14),
	.A2(FE_OFN28856_n15450),
	.B(FE_OFN25920_n15995),
	.C(FE_OFN26007_n16010));
   NOR2xp33_ASAP7_75t_SRAM U24680 (.Y(n14680),
	.A(FE_OFN27115_n),
	.B(FE_OFN26003_n15992));
   NOR2xp33_ASAP7_75t_SRAM U24681 (.Y(n14681),
	.A(FE_OFN26635_w3_14),
	.B(FE_OFN26003_n15992));
   NOR2xp33_ASAP7_75t_R U24682 (.Y(n14684),
	.A(n14695),
	.B(n14685));
   A2O1A1Ixp33_ASAP7_75t_L U24683 (.Y(n15970),
	.A1(FE_OCPN28296_n15386),
	.A2(FE_OFN26636_w3_14),
	.B(n15374),
	.C(n13844));
   OA21x2_ASAP7_75t_R U24684 (.Y(n14687),
	.A1(n14941),
	.A2(n15398),
	.B(n15970));
   NOR2xp33_ASAP7_75t_R U24685 (.Y(n14688),
	.A(n14686),
	.B(n14685));
   NOR2xp33_ASAP7_75t_SRAM U24686 (.Y(n14701),
	.A(n14695),
	.B(n14702));
   NOR2xp33_ASAP7_75t_R U24687 (.Y(n14704),
	.A(n13844),
	.B(n14702));
   O2A1O1Ixp33_ASAP7_75t_L U24688 (.Y(n15315),
	.A1(FE_OCPN27929_FE_OFN4_w3_22),
	.A2(FE_OFN27082_n25377),
	.B(n14747),
	.C(n13875));
   OR2x2_ASAP7_75t_R U24689 (.Y(n14753),
	.A(n14748),
	.B(n15315));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24690 (.Y(n14772),
	.A1(FE_OFN25915_n15514),
	.A2(n15501),
	.B(FE_OFN28551_FE_OFN26114_n),
	.C(n15534));
   OR2x2_ASAP7_75t_R U24691 (.Y(n14780),
	.A(n15477),
	.B(n14779));
   OAI21xp33_ASAP7_75t_R U24692 (.Y(n14814),
	.A1(n15714),
	.A2(FE_OFN16210_n13876),
	.B(n14789));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24693 (.Y(n14791),
	.A1(FE_OFN27066_n13869),
	.A2(n15471),
	.B(FE_PSN8334_n15539),
	.C(n14790));
   OAI21xp33_ASAP7_75t_L U24694 (.Y(n15709),
	.A1(FE_OFN27214_w3_17),
	.A2(FE_OFN26114_n),
	.B(n14795));
   A2O1A1Ixp33_ASAP7_75t_SL U24695 (.Y(n15046),
	.A1(FE_OCPN28072_w3_3),
	.A2(FE_OFN28732_n),
	.B(n15571),
	.C(n15838));
   OAI21xp33_ASAP7_75t_SRAM U24696 (.Y(n14849),
	.A1(n14986),
	.A2(n15813),
	.B(n14845));
   OAI22xp33_ASAP7_75t_SRAM U24697 (.Y(n14856),
	.A1(FE_OFN28671_FE_OCPN28076),
	.A2(n15033),
	.B1(FE_OCPN8254_w3_3),
	.B2(n15033));
   A2O1A1Ixp33_ASAP7_75t_L U24698 (.Y(n14865),
	.A1(FE_OFN27124_w3_1),
	.A2(n15834),
	.B(FE_OFN26084_n15106),
	.C(n14864));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24699 (.Y(n14898),
	.A1(FE_OCPN29506_FE_OFN16184_w3_9),
	.A2(FE_OFN29017_n15921),
	.B(FE_OFN28758_n15422),
	.C(n14897));
   OAI22xp33_ASAP7_75t_SRAM U24700 (.Y(n14910),
	.A1(FE_OFN112_n15994),
	.A2(n14905),
	.B1(n14904),
	.B2(n14905));
   INVxp33_ASAP7_75t_L U24701 (.Y(n14921),
	.A(n15438));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24702 (.Y(n14937),
	.A1(n14930),
	.A2(n14929),
	.B(n14928),
	.C(n14927));
   OAI21xp33_ASAP7_75t_SRAM U24703 (.Y(n14935),
	.A1(n14932),
	.A2(FE_OFN109_n15994),
	.B(n14931));
   NOR2xp33_ASAP7_75t_R U24704 (.Y(n14934),
	.A(FE_PSN8324_n15987),
	.B(n14933));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24705 (.Y(n14949),
	.A1(n24755),
	.A2(FE_OCPN29534_FE_OFN8_w3_14),
	.B(n15414),
	.C(n15922));
   INVxp67_ASAP7_75t_L U24706 (.Y(n14943),
	.A(n14942));
   NAND2xp33_ASAP7_75t_L U24707 (.Y(n14946),
	.A(n14945),
	.B(n14944));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24708 (.Y(n14978),
	.A1(n15857),
	.A2(FE_OFN26073_n),
	.B(n15872),
	.C(n15626));
   OA21x2_ASAP7_75t_SRAM U24709 (.Y(n14981),
	.A1(n14977),
	.A2(FE_OFN28889_n15845),
	.B(n14978));
   NOR2xp33_ASAP7_75t_SRAM U24710 (.Y(n14987),
	.A(n15871),
	.B(n14988));
   OAI22xp33_ASAP7_75t_SRAM U24711 (.Y(n15788),
	.A1(FE_OFN28695_n),
	.A2(n14986),
	.B1(n13766),
	.B2(n14986));
   NOR2xp33_ASAP7_75t_SRAM U24712 (.Y(n14991),
	.A(n14989),
	.B(n14988));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24713 (.Y(n15018),
	.A1(n24831),
	.A2(n15596),
	.B(n15000),
	.C(n15884));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24714 (.Y(n15016),
	.A1(n15884),
	.A2(FE_OFN26532_n13766),
	.B(n15015),
	.C(FE_OFN25912_n15848));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24715 (.Y(n15029),
	.A1(n13729),
	.A2(FE_OFN28889_n15845),
	.B(n15870),
	.C(n15028));
   NOR2xp33_ASAP7_75t_L U24716 (.Y(n15038),
	.A(n15124),
	.B(n15032));
   NOR2xp33_ASAP7_75t_R U24717 (.Y(n15035),
	.A(FE_OFN26532_n13766),
	.B(n13741));
   NOR2xp33_ASAP7_75t_SRAM U24718 (.Y(n15043),
	.A(n15041),
	.B(n15064));
   A2O1A1Ixp33_ASAP7_75t_L U24720 (.Y(n15047),
	.A1(FE_OFN29052_w3_5),
	.A2(n13741),
	.B(n15045),
	.C(FE_OFN25897_w3_4));
   OAI222xp33_ASAP7_75t_SRAM U24721 (.Y(n15073),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(n15809),
	.B1(n15859),
	.B2(n15809),
	.C1(n15627),
	.C2(n15809));
   A2O1A1Ixp33_ASAP7_75t_L U24722 (.Y(n15057),
	.A1(n15896),
	.A2(n15059),
	.B(FE_OFN16235_n15055),
	.C(FE_OFN43_w0_10));
   NOR2xp33_ASAP7_75t_SRAM U24723 (.Y(n15063),
	.A(n15787),
	.B(n15064));
   O2A1O1Ixp33_ASAP7_75t_SL U24724 (.Y(n15062),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(n15627),
	.B(n15626),
	.C(FE_OFN26084_n15106));
   NOR2xp33_ASAP7_75t_R U24725 (.Y(n15066),
	.A(FE_OCPN28072_w3_3),
	.B(n15064));
   OAI22xp33_ASAP7_75t_R U24726 (.Y(n15598),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(n15080),
	.B1(FE_OFN28732_n),
	.B2(n15080));
   NOR2xp33_ASAP7_75t_L U24727 (.Y(n15095),
	.A(n15838),
	.B(n15595));
   OR2x2_ASAP7_75t_R U24728 (.Y(n15096),
	.A(n15635),
	.B(n15595));
   NOR3xp33_ASAP7_75t_SRAM U24729 (.Y(n15101),
	.A(n15876),
	.B(FE_OFN29052_w3_5),
	.C(FE_OCPN29500_FE_OFN28662_w3_7));
   OR2x2_ASAP7_75t_SRAM U24730 (.Y(n15111),
	.A(n15617),
	.B(n15639));
   NAND2xp5_ASAP7_75t_L U24731 (.Y(n15123),
	.A(n15117),
	.B(n15120));
   NOR2xp33_ASAP7_75t_SRAM U24732 (.Y(n15121),
	.A(n15119),
	.B(n15118));
   A2O1A1Ixp33_ASAP7_75t_L U24733 (.Y(n15129),
	.A1(n15128),
	.A2(n24831),
	.B(n15619),
	.C(n15884));
   O2A1O1Ixp33_ASAP7_75t_SL U24734 (.Y(n15133),
	.A1(n15132),
	.A2(n15131),
	.B(n15896),
	.C(n15130));
   A2O1A1Ixp33_ASAP7_75t_SL U24735 (.Y(n16097),
	.A1(FE_OFN16411_n15884),
	.A2(n15142),
	.B(n15141),
	.C(n15140));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24736 (.Y(n15149),
	.A1(FE_OFN27208_w3_30),
	.A2(n15145),
	.B(FE_OFN28817_n),
	.C(n15203));
   NOR2xp33_ASAP7_75t_SRAM U24737 (.Y(n15148),
	.A(n15146),
	.B(n15149));
   OR3x1_ASAP7_75t_SRAM U24738 (.Y(n15150),
	.A(FE_OFN28890_n),
	.B(n15155),
	.C(n14535));
   NOR2xp33_ASAP7_75t_R U24739 (.Y(n15151),
	.A(FE_OFN16437_n),
	.B(n15149));
   NOR2xp33_ASAP7_75t_SRAM U24740 (.Y(n15161),
	.A(n15154),
	.B(n15162));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24741 (.Y(n15157),
	.A1(FE_OFN26049_w3_27),
	.A2(n15156),
	.B(n15155),
	.C(FE_OFN26059_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24742 (.Y(n15160),
	.A1(n15159),
	.A2(FE_OFN28717_n15158),
	.B(FE_OFN16225_n15195),
	.C(n15157));
   NOR2xp33_ASAP7_75t_SRAM U24743 (.Y(n15164),
	.A(FE_OFN28890_n),
	.B(n15162));
   NOR2xp33_ASAP7_75t_SRAM U24744 (.Y(n15173),
	.A(n15171),
	.B(n15170));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24745 (.Y(n15186),
	.A1(FE_OFN16206_n15240),
	.A2(n15185),
	.B(FE_OCPN29573_n15184),
	.C(FE_OCPN29547_n15183));
   OA21x2_ASAP7_75t_R U24746 (.Y(n15190),
	.A1(n15187),
	.A2(n14516),
	.B(n15186));
   NAND3xp33_ASAP7_75t_SRAM U24747 (.Y(n15198),
	.A(n15205),
	.B(n15197),
	.C(FE_OFN28456_n13348));
   A2O1A1Ixp33_ASAP7_75t_R U24748 (.Y(n15208),
	.A1(FE_OFN26049_w3_27),
	.A2(FE_OCPN27659_w3_25),
	.B(n15199),
	.C(n15198));
   NOR2xp33_ASAP7_75t_SRAM U24749 (.Y(n15207),
	.A(FE_OFN16193_n15200),
	.B(n15208));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24750 (.Y(n15202),
	.A1(FE_OFN27207_w3_30),
	.A2(FE_OFN26051_w3_27),
	.B(n15201),
	.C(n15240));
   A2O1A1Ixp33_ASAP7_75t_SL U24751 (.Y(n15206),
	.A1(n15205),
	.A2(FE_OFN28496_n15201),
	.B(n15203),
	.C(n15202));
   NOR2xp33_ASAP7_75t_SRAM U24752 (.Y(n15211),
	.A(n15209),
	.B(n15208));
   O2A1O1Ixp5_ASAP7_75t_SL U24753 (.Y(n15245),
	.A1(n15234),
	.A2(FE_OFN25893_n15214),
	.B(n15232),
	.C(n15238));
   NOR2xp33_ASAP7_75t_SL U24754 (.Y(n15244),
	.A(n15235),
	.B(n15245));
   NOR2xp33_ASAP7_75t_SL U24755 (.Y(n15248),
	.A(n15246),
	.B(n15245));
   NOR2xp33_ASAP7_75t_SRAM U24756 (.Y(n15285),
	.A(FE_OCPN29329_n15517),
	.B(n15286));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24757 (.Y(n15307),
	.A1(FE_OCPN29578_FE_OFN27214_w3_17),
	.A2(FE_OFN27096_n),
	.B(FE_OCPN27928_FE_OFN4_w3_22),
	.C(FE_PSN8334_n15539));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24758 (.Y(n15312),
	.A1(FE_OFN27214_w3_17),
	.A2(FE_OFN29087_n),
	.B(FE_OCPN27987_FE_OFN4_w3_22),
	.C(n15719));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24759 (.Y(n15323),
	.A1(n15680),
	.A2(FE_OCPN8264_n13890),
	.B(n15738),
	.C(n15501));
   NAND2xp33_ASAP7_75t_SRAM U24760 (.Y(n15331),
	.A(n15713),
	.B(FE_OFN28600_n14289));
   NOR2xp33_ASAP7_75t_R U24761 (.Y(n15329),
	.A(FE_OCPN28404_n13874),
	.B(FE_OCPN28278_n15512));
   A2O1A1Ixp33_ASAP7_75t_SL U24762 (.Y(n15342),
	.A1(n15667),
	.A2(n15341),
	.B(n15340),
	.C(FE_OFN16426_w3_20));
   A2O1A1Ixp33_ASAP7_75t_SL U24764 (.Y(n15352),
	.A1(n15683),
	.A2(n15351),
	.B(n15350),
	.C(n13867));
   A2O1A1Ixp33_ASAP7_75t_SL U24765 (.Y(n15355),
	.A1(n15354),
	.A2(n15353),
	.B(n15704),
	.C(n15352));
   NOR2xp33_ASAP7_75t_R U24766 (.Y(n15368),
	.A(key_5_),
	.B(FE_OFN26_n16125));
   NOR2xp33_ASAP7_75t_SRAM U24767 (.Y(n15377),
	.A(n16016),
	.B(n15375));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24768 (.Y(n15395),
	.A1(FE_OCPN29583_n15422),
	.A2(n15414),
	.B(n15934),
	.C(n15379));
   NOR2xp33_ASAP7_75t_SRAM U24769 (.Y(n15388),
	.A(n15381),
	.B(n15389));
   A2O1A1Ixp33_ASAP7_75t_L U24770 (.Y(n15387),
	.A1(FE_OCPN28296_n15386),
	.A2(FE_OCPN29536_FE_OFN8_w3_14),
	.B(n15385),
	.C(n15384));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24771 (.Y(n15401),
	.A1(FE_OFN28883_n),
	.A2(n15447),
	.B(n15446),
	.C(FE_OFN26007_n16010));
   NOR2xp33_ASAP7_75t_SRAM U24772 (.Y(n15400),
	.A(n13844),
	.B(n15401));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24773 (.Y(n15399),
	.A1(FE_OFN26635_w3_14),
	.A2(n15447),
	.B(n15398),
	.C(n15397));
   NOR2xp33_ASAP7_75t_SRAM U24774 (.Y(n15404),
	.A(n15402),
	.B(n15401));
   O2A1O1Ixp33_ASAP7_75t_L U24776 (.Y(n15415),
	.A1(FE_OFN28813_n15414),
	.A2(FE_OFN28544_n13805),
	.B(n15413),
	.C(n15993));
   OR3x1_ASAP7_75t_L U24777 (.Y(n15426),
	.A(FE_OCPN29570_n15423),
	.B(FE_OFN26642_w3_14),
	.C(FE_OCPN29509_FE_OFN16184_w3_9));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24778 (.Y(n15448),
	.A1(n15447),
	.A2(n15446),
	.B(FE_OFN26007_n16010),
	.C(n15445));
   OAI21xp33_ASAP7_75t_R U24779 (.Y(n15452),
	.A1(FE_OFN26624_n15376),
	.A2(n15451),
	.B(FE_OFN28856_n15450));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24780 (.Y(n15456),
	.A1(n15455),
	.A2(FE_OCPN28408_FE_OFN16433_w3_11),
	.B(n15953),
	.C(n15454));
   A2O1A1Ixp33_ASAP7_75t_SL U24781 (.Y(n15482),
	.A1(FE_OFN28628_n15667),
	.A2(n15477),
	.B(n15476),
	.C(FE_OFN26614_n));
   OAI22xp33_ASAP7_75t_SRAM U24782 (.Y(n15481),
	.A1(FE_OFN27066_n13869),
	.A2(n15479),
	.B1(n15478),
	.B2(n15479));
   O2A1O1Ixp5_ASAP7_75t_SRAM U24783 (.Y(n15489),
	.A1(FE_OCPN27929_FE_OFN4_w3_22),
	.A2(n15694),
	.B(n15719),
	.C(n13875));
   NAND2xp33_ASAP7_75t_L U24784 (.Y(n15493),
	.A(n15528),
	.B(n14061));
   A2O1A1Ixp33_ASAP7_75t_SL U24785 (.Y(n15504),
	.A1(FE_OFN28551_FE_OFN26114_n),
	.A2(FE_OFN27082_n25377),
	.B(n15503),
	.C(n15502));
   NAND2xp33_ASAP7_75t_SRAM U24786 (.Y(n15537),
	.A(n15536),
	.B(FE_OFN25981_n13868));
   NAND2xp33_ASAP7_75t_SRAM U24787 (.Y(n15543),
	.A(n15694),
	.B(n15719));
   OA21x2_ASAP7_75t_L U24788 (.Y(n15546),
	.A1(n15480),
	.A2(n15543),
	.B(n15542));
   A2O1A1Ixp33_ASAP7_75t_L U24789 (.Y(n15750),
	.A1(FE_OFN27096_n),
	.A2(FE_OFN27082_n25377),
	.B(FE_OFN27151_n),
	.C(n15760));
   NOR2xp33_ASAP7_75t_R U24790 (.Y(n15547),
	.A(n15750),
	.B(n15545));
   OA21x2_ASAP7_75t_SRAM U24791 (.Y(n15579),
	.A1(FE_OCPN28398_n15808),
	.A2(n25140),
	.B(n15575));
   NOR2xp33_ASAP7_75t_SRAM U24792 (.Y(n15580),
	.A(n15578),
	.B(n15577));
   OAI21xp33_ASAP7_75t_R U24793 (.Y(n15588),
	.A1(n25140),
	.A2(FE_OFN28691_n13725),
	.B(n15585));
   A2O1A1Ixp33_ASAP7_75t_R U24794 (.Y(n15593),
	.A1(n15857),
	.A2(n15592),
	.B(n15591),
	.C(FE_OFN26073_n));
   NOR2xp33_ASAP7_75t_L U24795 (.Y(n15624),
	.A(FE_OFN16411_n15884),
	.B(n15646));
   OAI21xp5_ASAP7_75t_L U24796 (.Y(n15597),
	.A1(FE_OCPN28072_w3_3),
	.A2(FE_OFN27156_n),
	.B(n15596));
   OA21x2_ASAP7_75t_SL U24797 (.Y(n15602),
	.A1(n15598),
	.A2(n13725),
	.B(n15597));
   A2O1A1Ixp33_ASAP7_75t_R U24798 (.Y(n15616),
	.A1(FE_OFN28721_n),
	.A2(n15817),
	.B(n15814),
	.C(n15615));
   O2A1O1Ixp33_ASAP7_75t_R U24799 (.Y(n15628),
	.A1(FE_OCPN29537_FE_OFN28699_w3_6),
	.A2(n15627),
	.B(n15626),
	.C(FE_OFN25928_n15779));
   NOR2xp33_ASAP7_75t_SL U24800 (.Y(n15649),
	.A(n15647),
	.B(n15646));
   A2O1A1Ixp33_ASAP7_75t_L U24801 (.Y(n15654),
	.A1(n15896),
	.A2(n15656),
	.B(n15653),
	.C(w0_8_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24802 (.Y(n15670),
	.A1(FE_OFN26091_n24663),
	.A2(FE_OFN28624_n13874),
	.B(n13916),
	.C(FE_OFN28827_n15683));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24803 (.Y(n15669),
	.A1(n15694),
	.A2(FE_OFN28712_n),
	.B(n15668),
	.C(n15667));
   A2O1A1Ixp33_ASAP7_75t_L U24804 (.Y(n15695),
	.A1(FE_OFN6_w3_22),
	.A2(n15694),
	.B(n13875),
	.C(n15693));
   OAI22xp33_ASAP7_75t_R U24806 (.Y(n15712),
	.A1(FE_OFN28977_n),
	.A2(n13916),
	.B1(FE_OFN26053_n25415),
	.B2(n13916));
   NOR2xp33_ASAP7_75t_SRAM U24807 (.Y(n15790),
	.A(n15788),
	.B(n15791));
   NOR2xp33_ASAP7_75t_SRAM U24808 (.Y(n15794),
	.A(n15792),
	.B(n15791));
   NOR2xp33_ASAP7_75t_SRAM U24809 (.Y(n15800),
	.A(n15799),
	.B(n15798));
   OR2x2_ASAP7_75t_SRAM U24810 (.Y(n15801),
	.A(n14996),
	.B(FE_OCPN28398_n15808));
   OA21x2_ASAP7_75t_SRAM U24811 (.Y(n15830),
	.A1(n15034),
	.A2(n15825),
	.B(n15824));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24812 (.Y(n15839),
	.A1(FE_OFN16195_n13771),
	.A2(FE_OFN28831_n15838),
	.B(n15837),
	.C(FE_OFN28671_FE_OCPN28076));
   NOR3xp33_ASAP7_75t_SRAM U24813 (.Y(n15840),
	.A(n13725),
	.B(FE_OFN28699_w3_6),
	.C(FE_OFN28732_n));
   OAI21xp5_ASAP7_75t_R U24814 (.Y(n15885),
	.A1(n15808),
	.A2(n15856),
	.B(n15855));
   OR2x2_ASAP7_75t_R U24815 (.Y(n15877),
	.A(n15876),
	.B(n15875));
   A2O1A1Ixp33_ASAP7_75t_SL U24816 (.Y(n15893),
	.A1(n15896),
	.A2(n15895),
	.B(n15892),
	.C(w0_11_));
   A2O1A1Ixp33_ASAP7_75t_SL U24817 (.Y(n15912),
	.A1(n25140),
	.A2(FE_OFN26_n16125),
	.B(n15911),
	.C(n16050));
   A2O1A1Ixp33_ASAP7_75t_SL U24818 (.Y(n15914),
	.A1(FE_OFN26139_n16125),
	.A2(n23937),
	.B(n15913),
	.C(n15915));
   OA21x2_ASAP7_75t_SRAM U24819 (.Y(n15930),
	.A1(n15927),
	.A2(n15926),
	.B(n15925));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24820 (.Y(n15935),
	.A1(FE_OFN26633_w3_14),
	.A2(FE_OCPN29506_FE_OFN16184_w3_9),
	.B(FE_OCPN28408_FE_OFN16433_w3_11),
	.C(n13844));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24821 (.Y(n15937),
	.A1(n15936),
	.A2(n15956),
	.B(FE_OFN26007_n16010),
	.C(n15935));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24822 (.Y(n15960),
	.A1(n16000),
	.A2(n15959),
	.B(n15958),
	.C(n15957));
   OA21x2_ASAP7_75t_R U24823 (.Y(n15979),
	.A1(n15976),
	.A2(n15975),
	.B(n15974));
   OR2x2_ASAP7_75t_R U24824 (.Y(n15991),
	.A(FE_OFN16305_n15984),
	.B(n15985));
   NOR2xp33_ASAP7_75t_SRAM U24825 (.Y(n15989),
	.A(n15986),
	.B(n15985));
   OAI22xp33_ASAP7_75t_SRAM U24826 (.Y(n16001),
	.A1(n16000),
	.A2(FE_OFN28898_n13805),
	.B1(n15999),
	.B2(FE_OFN28898_n13805));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24827 (.Y(n16013),
	.A1(FE_OFN16417_n),
	.A2(FE_OCPN29564_n16012),
	.B(FE_OFN27136_n15992),
	.C(FE_OFN26007_n16010));
   A2O1A1Ixp33_ASAP7_75t_L U24828 (.Y(n16061),
	.A1(FE_OFN26073_n),
	.A2(FE_OFN26_n16125),
	.B(n16060),
	.C(n16078));
   A2O1A1Ixp33_ASAP7_75t_L U24829 (.Y(n16071),
	.A1(FE_OFN26_n16125),
	.A2(FE_OCPN29502_w3_23),
	.B(n16070),
	.C(FE_OCPN29550_n16114));
   A2O1A1Ixp33_ASAP7_75t_SL U24830 (.Y(n16093),
	.A1(FE_OFN25_n16125),
	.A2(FE_PSN8297_FE_OFN8_w3_14),
	.B(n16092),
	.C(n16094));
   A2O1A1Ixp33_ASAP7_75t_SL U24831 (.Y(n16109),
	.A1(FE_OFN26_n16125),
	.A2(n25961),
	.B(n16108),
	.C(n16110));
   A2O1A1Ixp33_ASAP7_75t_L U24832 (.Y(n16112),
	.A1(FE_OFN28470_ld),
	.A2(FE_OFN27129_w3_28),
	.B(n16111),
	.C(FE_OFN16246_n16113));
   A2O1A1Ixp33_ASAP7_75t_SL U24833 (.Y(n16129),
	.A1(FE_OFN25_n16125),
	.A2(FE_OFN26129_w3_15),
	.B(n16128),
	.C(n16148));
   A2O1A1Ixp33_ASAP7_75t_SL U24834 (.Y(n16147),
	.A1(FE_OFN28674_n),
	.A2(FE_OFN26_n16125),
	.B(n16146),
	.C(n16172));
   A2O1A1Ixp33_ASAP7_75t_L U24835 (.Y(n16161),
	.A1(n24470),
	.A2(FE_OFN28470_ld),
	.B(n16160),
	.C(FE_OFN16251_n16162));
   OAI21xp33_ASAP7_75t_SL U24836 (.Y(n634),
	.A1(FE_OFN16251_n16162),
	.A2(n24470),
	.B(n16161));
   A2O1A1Ixp33_ASAP7_75t_SL U24837 (.Y(n16181),
	.A1(FE_OFN27_n16125),
	.A2(FE_OCPN29520_n24755),
	.B(n16180),
	.C(n16201));
   A2O1A1Ixp33_ASAP7_75t_SL U24838 (.Y(n16188),
	.A1(FE_OCPN29428_FE_OFN27131_w3_29),
	.A2(FE_OFN28470_ld),
	.B(n16187),
	.C(FE_OFN16253_n16189));
   A2O1A1Ixp33_ASAP7_75t_SL U24839 (.Y(n16196),
	.A1(FE_OFN26163_w3_13),
	.A2(FE_OFN28457_ld),
	.B(n16195),
	.C(n16240));
   A2O1A1Ixp33_ASAP7_75t_SL U24840 (.Y(n16230),
	.A1(w2_27_),
	.A2(FE_OFN22_n16125),
	.B(n16216),
	.C(n16215));
   A2O1A1Ixp33_ASAP7_75t_SL U24841 (.Y(n16221),
	.A1(n25051),
	.A2(FE_OFN25_n16125),
	.B(n16220),
	.C(n16222));
   A2O1A1Ixp33_ASAP7_75t_SL U24842 (.Y(n16227),
	.A1(FE_OFN27_n16125),
	.A2(FE_OCPN28408_FE_OFN16433_w3_11),
	.B(n16226),
	.C(n16265));
   NOR2xp33_ASAP7_75t_SRAM U24843 (.Y(n16228),
	.A(key_27_),
	.B(FE_OFN28472_ld));
   A2O1A1Ixp33_ASAP7_75t_SL U24844 (.Y(n16229),
	.A1(FE_OFN28472_ld),
	.A2(FE_OFN28890_n),
	.B(n16228),
	.C(FE_OFN16287_n16230));
   A2O1A1Ixp33_ASAP7_75t_SL U24845 (.Y(n16246),
	.A1(FE_OFN28461_ld),
	.A2(FE_OFN16421_n23974),
	.B(n16245),
	.C(n16247));
   NOR2xp33_ASAP7_75t_SRAM U24846 (.Y(n16252),
	.A(key_16_),
	.B(FE_OFN28463_ld));
   NOR2xp33_ASAP7_75t_SRAM U24847 (.Y(n16251),
	.A(w3_16_),
	.B(ld));
   A2O1A1Ixp33_ASAP7_75t_L U24848 (.Y(n16260),
	.A1(FE_OFN16159_w3_24),
	.A2(FE_OFN28470_ld),
	.B(n16259),
	.C(FE_OFN16370_n16261));
   A2O1A1Ixp33_ASAP7_75t_SL U24849 (.Y(n16270),
	.A1(FE_OFN25961_w3_8),
	.A2(FE_OFN26_n16125),
	.B(n16269),
	.C(n16271));
   NOR2xp33_ASAP7_75t_SRAM U24850 (.Y(n16280),
	.A(ld),
	.B(dcnt_1_));
   NAND3xp33_ASAP7_75t_SRAM U24851 (.Y(n923),
	.A(n16281),
	.B(n16280),
	.C(dcnt_0_));
   NAND3xp33_ASAP7_75t_SRAM U24852 (.Y(n655),
	.A(n16282),
	.B(n16286),
	.C(u0_r0_rcnt_2_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24853 (.Y(n657),
	.A1(n16287),
	.A2(u0_r0_rcnt_2_),
	.B(n16284),
	.C(n16283));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24854 (.Y(n658),
	.A1(n16285),
	.A2(n16287),
	.B(n16284),
	.C(FE_OFN28468_ld));
   NOR2xp33_ASAP7_75t_SRAM U24855 (.Y(n16288),
	.A(n16286),
	.B(n665));
   NAND3xp33_ASAP7_75t_SRAM U24856 (.Y(n656),
	.A(n16288),
	.B(n16287),
	.C(u0_r0_rcnt_2_));
   INVx4_ASAP7_75t_SL U24857 (.Y(n20868),
	.A(FE_OCPN27697_n16309));
   NOR2x1_ASAP7_75t_L U24858 (.Y(n20064),
	.A(FE_OFN26629_sa31_4),
	.B(FE_OFN28669_sa31_5));
   NAND3x2_ASAP7_75t_SL U24859 (.Y(n21948),
	.A(n20868),
	.B(FE_OCPN27444_n20064),
	.C(n16493));
   NOR2x1_ASAP7_75t_L U24860 (.Y(n16303),
	.A(FE_OFN29136_n),
	.B(n16329));
   NOR3x2_ASAP7_75t_SL U24861 (.Y(n20050),
	.A(FE_OFN28669_sa31_5),
	.B(n16493),
	.C(FE_OCPN29526_sa31_4));
   NAND3x2_ASAP7_75t_SL U24862 (.Y(n21981),
	.A(FE_OFN29145_sa31_1),
	.B(FE_OFN26095_n16293),
	.C(FE_OFN28516_FE_OFN27192_sa31_2));
   NAND2x1p5_ASAP7_75t_L U24863 (.Y(n20853),
	.A(n16493),
	.B(n20064));
   NAND2x1p5_ASAP7_75t_SL U24864 (.Y(n21939),
	.A(FE_OFN100_sa31_1),
	.B(FE_OFN26095_n16293));
   NOR3x1_ASAP7_75t_SL U24865 (.Y(n20078),
	.A(n20853),
	.B(FE_OFN28719_n20025),
	.C(n21939));
   NOR2xp33_ASAP7_75t_L U24866 (.Y(n16291),
	.A(n20876),
	.B(n20078));
   NAND3x2_ASAP7_75t_SL U24867 (.Y(n21980),
	.A(FE_OCPN29526_sa31_4),
	.B(FE_OFN28669_sa31_5),
	.C(FE_OFN28840_n));
   NOR2x1_ASAP7_75t_SL U24868 (.Y(n26293),
	.A(FE_OFN26096_n16294),
	.B(n20076));
   NAND2x1_ASAP7_75t_SL U24870 (.Y(n16497),
	.A(FE_OFN28516_FE_OFN27192_sa31_2),
	.B(n16295));
   NAND2x1p5_ASAP7_75t_L U24871 (.Y(n16340),
	.A(n16298),
	.B(FE_OFN28669_sa31_5));
   NOR3x1_ASAP7_75t_SL U24872 (.Y(n16512),
	.A(FE_OFN26095_n16293),
	.B(FE_OFN28753_sa31_2),
	.C(FE_OFN29147_sa31_1));
   NOR2x1_ASAP7_75t_SL U24873 (.Y(n21977),
	.A(FE_OFN28719_n20025),
	.B(n16349));
   NOR2x1p5_ASAP7_75t_SL U24874 (.Y(n16348),
	.A(FE_OFN28516_FE_OFN27192_sa31_2),
	.B(n16329));
   A2O1A1Ixp33_ASAP7_75t_L U24875 (.Y(n16302),
	.A1(n21940),
	.A2(FE_OFN29117_n),
	.B(FE_OCPN28394_FE_OFN27043_n),
	.C(n26007));
   NOR2x1p5_ASAP7_75t_SL U24876 (.Y(n26291),
	.A(FE_OFN26015_sa31_3),
	.B(n16394));
   NAND2xp5_ASAP7_75t_SL U24877 (.Y(n25316),
	.A(n20868),
	.B(n26291));
   NOR2x1p5_ASAP7_75t_SL U24878 (.Y(n20841),
	.A(n16493),
	.B(n16394));
   NOR2x1p5_ASAP7_75t_SL U24879 (.Y(n26292),
	.A(FE_OFN28719_n20025),
	.B(n21939));
   NAND2x1p5_ASAP7_75t_SL U24880 (.Y(n16321),
	.A(FE_OCPN29482_FE_OFN26014_sa31_3),
	.B(FE_OCPN29526_sa31_4));
   NAND2xp33_ASAP7_75t_SL U24881 (.Y(n16326),
	.A(n26292),
	.B(n16299));
   NOR2xp33_ASAP7_75t_L U24882 (.Y(n16304),
	.A(FE_OCPN28334_n16497),
	.B(n20853));
   NAND2x1p5_ASAP7_75t_L U24883 (.Y(n20842),
	.A(n16493),
	.B(n24181));
   NOR2x1_ASAP7_75t_L U24884 (.Y(n20027),
	.A(n20854),
	.B(n20842));
   NOR2xp33_ASAP7_75t_L U24885 (.Y(n16396),
	.A(n20027),
	.B(n20837));
   NAND3xp33_ASAP7_75t_SL U24886 (.Y(n16310),
	.A(n16338),
	.B(n16396),
	.C(n16341));
   NAND3xp33_ASAP7_75t_SL U24887 (.Y(n26400),
	.A(n16300),
	.B(n26292),
	.C(FE_OFN26060_sa31_4));
   NOR2xp33_ASAP7_75t_L U24888 (.Y(n16314),
	.A(FE_OFN28808_n26291),
	.B(n20049));
   NAND2xp5_ASAP7_75t_R U24889 (.Y(n21933),
	.A(FE_OCPN27516_n26292),
	.B(n21989));
   NOR2x1_ASAP7_75t_L U24890 (.Y(n27070),
	.A(FE_OCPN28314_n20842),
	.B(FE_OCPN28008_n16290));
   NOR2xp33_ASAP7_75t_SL U24891 (.Y(n16313),
	.A(n20078),
	.B(n27070));
   AND3x1_ASAP7_75t_SL U24892 (.Y(n16315),
	.A(n21933),
	.B(n21932),
	.C(n16313));
   NAND2x1p5_ASAP7_75t_SL U24893 (.Y(n20074),
	.A(FE_OFN26060_sa31_4),
	.B(n16300));
   OAI21x1_ASAP7_75t_L U24894 (.Y(n24184),
	.A1(FE_OCPN7597_n21981),
	.A2(n20074),
	.B(n16407));
   NOR2x1_ASAP7_75t_L U24896 (.Y(n18062),
	.A(FE_OCPN28394_FE_OFN27043_n),
	.B(n20074));
   NOR2x1_ASAP7_75t_L U24897 (.Y(n21938),
	.A(n20059),
	.B(n18062));
   NOR2x1_ASAP7_75t_L U24898 (.Y(n18098),
	.A(n24184),
	.B(n16322));
   NAND3xp33_ASAP7_75t_R U24899 (.Y(n16323),
	.A(FE_OFN28618_n25322),
	.B(n16398),
	.C(n20075));
   NAND2x1_ASAP7_75t_SL U24900 (.Y(n27072),
	.A(n18098),
	.B(n16324));
   NOR2x1_ASAP7_75t_L U24901 (.Y(n16327),
	.A(n18071),
	.B(n16391));
   NOR2x1_ASAP7_75t_L U24902 (.Y(n25319),
	.A(FE_OFN28516_FE_OFN27192_sa31_2),
	.B(n16330));
   NAND3xp33_ASAP7_75t_R U24903 (.Y(n16337),
	.A(n16335),
	.B(n20874),
	.C(n20034));
   NOR2x1_ASAP7_75t_R U24904 (.Y(n26401),
	.A(FE_OCPN29483_FE_OFN26014_sa31_3),
	.B(n20081));
   NAND2x1p5_ASAP7_75t_L U24905 (.Y(n25317),
	.A(n20841),
	.B(n16295));
   NAND3xp33_ASAP7_75t_L U24906 (.Y(n16336),
	.A(FE_PSN8293_n25317),
	.B(n25316),
	.C(n18094));
   NOR3xp33_ASAP7_75t_SL U24907 (.Y(n16339),
	.A(n16337),
	.B(n26401),
	.C(n16336));
   NAND2x1p5_ASAP7_75t_SL U24909 (.Y(n20083),
	.A(n26291),
	.B(n26292));
   A2O1A1Ixp33_ASAP7_75t_R U24910 (.Y(n16347),
	.A1(FE_OCPN28394_FE_OFN27043_n),
	.A2(n16408),
	.B(FE_OCPN28314_n20842),
	.C(FE_OCPN27780_n20083));
   NAND2xp5_ASAP7_75t_L U24911 (.Y(n16385),
	.A(n20868),
	.B(n16299));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24912 (.Y(n16354),
	.A1(n26942),
	.A2(n26907),
	.B(n26904),
	.C(w2_2_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24913 (.Y(n439),
	.A1(n26942),
	.A2(n26907),
	.B(n16355),
	.C(n16354));
   NOR2xp33_ASAP7_75t_L U24914 (.Y(n16357),
	.A(FE_OCPN27316_n25849),
	.B(n20043));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24915 (.Y(n16356),
	.A1(n16295),
	.A2(n20050),
	.B(n20876),
	.C(FE_OFN16415_sa31_2));
   NOR2xp33_ASAP7_75t_SRAM U24916 (.Y(n16360),
	.A(FE_OCPN28314_n20842),
	.B(n21939));
   NOR2xp33_ASAP7_75t_SRAM U24917 (.Y(n16366),
	.A(n24181),
	.B(n24194));
   INVxp33_ASAP7_75t_SRAM U24918 (.Y(n16365),
	.A(n24184));
   NOR2xp33_ASAP7_75t_SRAM U24919 (.Y(n16368),
	.A(FE_OFN27043_n),
	.B(n24194));
   NAND2x1p5_ASAP7_75t_SL U24920 (.Y(n20882),
	.A(FE_OFN28710_n20841),
	.B(n20868));
   OAI21xp5_ASAP7_75t_SL U24921 (.Y(n21945),
	.A1(FE_OCPN7597_n21981),
	.A2(FE_OFN29117_n),
	.B(n20882));
   NOR2x1p5_ASAP7_75t_L U24922 (.Y(n20023),
	.A(n21980),
	.B(FE_OCPN28394_FE_OFN27043_n));
   NAND2xp5_ASAP7_75t_SL U24923 (.Y(n20048),
	.A(n21936),
	.B(n25322));
   NOR3x1_ASAP7_75t_SL U24924 (.Y(n24189),
	.A(n21945),
	.B(n20023),
	.C(n20048));
   NAND3xp33_ASAP7_75t_SRAM U24925 (.Y(n16415),
	.A(n24191),
	.B(n16371),
	.C(n24189));
   NAND2x1_ASAP7_75t_SL U24926 (.Y(n21964),
	.A(n18069),
	.B(n20832));
   NOR2xp33_ASAP7_75t_SL U24927 (.Y(n16379),
	.A(FE_OFN28808_n26291),
	.B(n26009));
   AND2x2_ASAP7_75t_R U24928 (.Y(n16380),
	.A(n21938),
	.B(n20066));
   NOR2xp33_ASAP7_75t_SL U24929 (.Y(n16381),
	.A(FE_OFN29032_FE_OCPN27728_n21981),
	.B(n26009));
   NOR2xp33_ASAP7_75t_SRAM U24931 (.Y(n16393),
	.A(FE_OCPN27316_n25849),
	.B(n25848));
   NAND2xp5_ASAP7_75t_SL U24932 (.Y(n20068),
	.A(n21948),
	.B(n16385));
   NOR3xp33_ASAP7_75t_SL U24933 (.Y(n16386),
	.A(n20068),
	.B(n18072),
	.C(n18071));
   NAND2xp5_ASAP7_75t_SL U24934 (.Y(n16388),
	.A(n24189),
	.B(n16386));
   NOR3xp33_ASAP7_75t_SL U24935 (.Y(n20836),
	.A(n16388),
	.B(n26401),
	.C(n16387));
   O2A1O1Ixp33_ASAP7_75t_SRAM U24936 (.Y(n16389),
	.A1(FE_OFN28753_sa31_2),
	.A2(sa31_1_),
	.B(FE_OFN26095_n16293),
	.C(n20074));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24937 (.Y(n16390),
	.A1(FE_OFN28753_sa31_2),
	.A2(sa31_1_),
	.B(FE_OFN26095_n16293),
	.C(n16389));
   NOR2xp33_ASAP7_75t_SRAM U24938 (.Y(n16409),
	.A(FE_OCPN7617_n26009),
	.B(n26008));
   OAI21xp5_ASAP7_75t_L U24939 (.Y(n18076),
	.A1(FE_OCPN28334_n16497),
	.A2(FE_OFN29047_n21980),
	.B(n21948));
   NOR2x1_ASAP7_75t_L U24940 (.Y(n16494),
	.A(n20023),
	.B(n18062));
   NOR2x1_ASAP7_75t_SL U24942 (.Y(n16523),
	.A(n16499),
	.B(FE_OFN26570_n20866));
   AND3x1_ASAP7_75t_SL U24943 (.Y(n16401),
	.A(n16494),
	.B(n20865),
	.C(n16523));
   NOR2xp33_ASAP7_75t_L U24944 (.Y(n16402),
	.A(n16299),
	.B(n18076));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24945 (.Y(n16413),
	.A1(n26407),
	.A2(n16415),
	.B(n16412),
	.C(w2_4_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24946 (.Y(n438),
	.A1(n26407),
	.A2(n16415),
	.B(n16414),
	.C(n16413));
   NOR2xp33_ASAP7_75t_SRAM U24947 (.Y(n23571),
	.A(sa33_6_),
	.B(n16468));
   NOR2x1p5_ASAP7_75t_L U24948 (.Y(n17416),
	.A(FE_OCPN29391_FE_OFN29162_sa33_2),
	.B(n16416));
   NAND2x1p5_ASAP7_75t_L U24950 (.Y(n16947),
	.A(n16928),
	.B(FE_OCPN29438_sa33_2));
   NAND3xp33_ASAP7_75t_SRAM U24951 (.Y(n16419),
	.A(FE_OFN25938_sa33_3),
	.B(n16418),
	.C(FE_OFN28679_sa33_5));
   NAND3xp33_ASAP7_75t_L U24952 (.Y(n16426),
	.A(n16855),
	.B(n18129),
	.C(n16419));
   NOR2x1_ASAP7_75t_SL U24953 (.Y(n16873),
	.A(FE_OFN28727_sa33_1),
	.B(FE_OFN28643_sa33_0));
   NAND2x1p5_ASAP7_75t_L U24955 (.Y(n16872),
	.A(FE_OFN26078_sa33_2),
	.B(n16422));
   NAND2x1p5_ASAP7_75t_SL U24956 (.Y(n23556),
	.A(FE_OFN28679_sa33_5),
	.B(FE_OCPN27544_sa33_4));
   NAND2x1p5_ASAP7_75t_SL U24957 (.Y(n16925),
	.A(FE_OFN16430_sa33_3),
	.B(n16417));
   A2O1A1Ixp33_ASAP7_75t_SL U24959 (.Y(n16476),
	.A1(n16925),
	.A2(n16673),
	.B(FE_OFN26545_n16447),
	.C(n16448));
   NAND3xp33_ASAP7_75t_L U24960 (.Y(n16913),
	.A(FE_OFN29134_sa33_0),
	.B(FE_OFN28727_sa33_1),
	.C(FE_OFN29162_sa33_2));
   NAND2x1_ASAP7_75t_L U24961 (.Y(n16677),
	.A(FE_OFN28694_sa33_4),
	.B(FE_OFN28679_sa33_5));
   NOR3xp33_ASAP7_75t_SRAM U24962 (.Y(n16443),
	.A(FE_OFN28541_n16476),
	.B(n24485),
	.C(n16433));
   NOR2x1_ASAP7_75t_L U24963 (.Y(n16937),
	.A(FE_OFN29164_sa33_2),
	.B(n18134));
   NOR2x1_ASAP7_75t_SL U24964 (.Y(n16909),
	.A(FE_OFN28679_sa33_5),
	.B(FE_OCPN27568_sa33_3));
   NOR2x1_ASAP7_75t_SL U24965 (.Y(n16831),
	.A(FE_OFN29134_sa33_0),
	.B(FE_OFN26062_n16435));
   NAND3xp33_ASAP7_75t_L U24966 (.Y(n16442),
	.A(n16437),
	.B(n16471),
	.C(n23531));
   NOR3xp33_ASAP7_75t_SRAM U24967 (.Y(n16439),
	.A(FE_OCPN28127_n16872),
	.B(FE_OFN26055_n),
	.C(FE_OFN27062_n16438));
   NOR2x1_ASAP7_75t_SL U24968 (.Y(n16929),
	.A(n16429),
	.B(n16436));
   NAND3xp33_ASAP7_75t_L U24969 (.Y(n16441),
	.A(n16440),
	.B(n24619),
	.C(n23542));
   NOR2xp33_ASAP7_75t_SL U24970 (.Y(n18442),
	.A(FE_OCPN28141_n),
	.B(n18426));
   A2O1A1Ixp33_ASAP7_75t_L U24971 (.Y(n16451),
	.A1(FE_OCPN29299_FE_OFN29232_n16875),
	.A2(FE_OCPN28127_n16872),
	.B(n16429),
	.C(n18442));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24972 (.Y(n16454),
	.A1(FE_OFN28998_n16923),
	.A2(FE_OCPN27555_n16422),
	.B(n18415),
	.C(FE_OFN29164_sa33_2));
   NOR2x1p5_ASAP7_75t_SL U24973 (.Y(n24613),
	.A(n16947),
	.B(n16429));
   NOR2xp33_ASAP7_75t_SL U24974 (.Y(n16460),
	.A(n16430),
	.B(n24613));
   NOR2x1p5_ASAP7_75t_SL U24975 (.Y(n16853),
	.A(n16421),
	.B(n16872));
   INVxp67_ASAP7_75t_L U24976 (.Y(n16456),
	.A(n16455));
   NOR2xp67_ASAP7_75t_L U24977 (.Y(n16458),
	.A(n18430),
	.B(n24296));
   NAND3x1_ASAP7_75t_SL U24978 (.Y(n16465),
	.A(n16895),
	.B(n18129),
	.C(n16894));
   NOR3x1_ASAP7_75t_SL U24979 (.Y(n16730),
	.A(n16465),
	.B(n24297),
	.C(n24300));
   NOR3xp33_ASAP7_75t_R U24980 (.Y(n16467),
	.A(n18434),
	.B(n24327),
	.C(n17425));
   NOR2x1_ASAP7_75t_L U24981 (.Y(n23537),
	.A(n16874),
	.B(FE_OCPN27460_n16913));
   NOR2x1_ASAP7_75t_SL U24982 (.Y(n26122),
	.A(FE_OCPN28127_n16872),
	.B(n16429));
   NOR2x1_ASAP7_75t_L U24983 (.Y(n16859),
	.A(n16874),
	.B(FE_OFN29208_n16436));
   NAND3xp33_ASAP7_75t_L U24984 (.Y(n16466),
	.A(n23551),
	.B(n16910),
	.C(n23529));
   NAND3xp33_ASAP7_75t_SL U24985 (.Y(n16478),
	.A(n16471),
	.B(n16470),
	.C(n16729));
   NOR3x1_ASAP7_75t_SL U24986 (.Y(n23546),
	.A(n16474),
	.B(n23552),
	.C(n23530));
   NAND3xp33_ASAP7_75t_SL U24987 (.Y(n16938),
	.A(n16475),
	.B(n23528),
	.C(n23546));
   NOR2x1p5_ASAP7_75t_SL U24988 (.Y(n16936),
	.A(FE_OCPN27604_n16421),
	.B(FE_OFN29208_n16436));
   NOR2x1_ASAP7_75t_SL U24989 (.Y(n16846),
	.A(FE_OCPN27593_n16908),
	.B(n16936));
   NAND3xp33_ASAP7_75t_L U24990 (.Y(n16477),
	.A(n24487),
	.B(n16724),
	.C(n16846));
   A2O1A1Ixp33_ASAP7_75t_SL U24991 (.Y(n26537),
	.A1(n16890),
	.A2(n16487),
	.B(n24331),
	.C(n16486));
   A2O1A1Ixp33_ASAP7_75t_SRAM U24992 (.Y(n16488),
	.A1(n23571),
	.A2(FE_OFN16275_n26536),
	.B(FE_OCPN29481_n26537),
	.C(w0_6_));
   NOR2xp33_ASAP7_75t_SRAM U24994 (.Y(n16492),
	.A(n27072),
	.B(n27071));
   NAND3xp33_ASAP7_75t_R U24995 (.Y(n16506),
	.A(n16494),
	.B(n21979),
	.C(n26007));
   OAI21xp5_ASAP7_75t_L U24996 (.Y(n21928),
	.A1(FE_OCPN28334_n16497),
	.A2(FE_OFN29047_n21980),
	.B(n20856));
   NAND3xp33_ASAP7_75t_R U24997 (.Y(n16505),
	.A(n16504),
	.B(n20054),
	.C(n16503));
   NOR3xp33_ASAP7_75t_SL U24998 (.Y(n26044),
	.A(n16506),
	.B(n21951),
	.C(n16505));
   AOI21xp5_ASAP7_75t_SL U24999 (.Y(n27080),
	.A1(n25847),
	.A2(n16511),
	.B(n26315));
   OAI22xp5_ASAP7_75t_L U25000 (.Y(n21925),
	.A1(FE_OFN29016_n16512),
	.A2(n20023),
	.B1(n16299),
	.B2(n20023));
   OAI21xp33_ASAP7_75t_R U25001 (.Y(n16522),
	.A1(n20074),
	.A2(FE_OCPN7597_n21981),
	.B(n21925));
   A2O1A1Ixp33_ASAP7_75t_R U25002 (.Y(n25816),
	.A1(n20868),
	.A2(n16300),
	.B(n25319),
	.C(FE_OFN26060_sa31_4));
   NAND3xp33_ASAP7_75t_SRAM U25003 (.Y(n16514),
	.A(FE_PSN8295_FE_OFN28669_sa31_5),
	.B(n26292),
	.C(FE_OCPN29483_FE_OFN26014_sa31_3));
   NAND3xp33_ASAP7_75t_SL U25004 (.Y(n16517),
	.A(n25316),
	.B(n16514),
	.C(n16513));
   NOR3xp33_ASAP7_75t_SL U25005 (.Y(n16518),
	.A(n16517),
	.B(n16516),
	.C(n16515));
   NAND3xp33_ASAP7_75t_SL U25006 (.Y(n26046),
	.A(n16525),
	.B(n16524),
	.C(n16523));
   OAI22xp33_ASAP7_75t_SRAM U25007 (.Y(n16526),
	.A1(n26407),
	.A2(FE_OCPN28438_n27080),
	.B1(n26046),
	.B2(FE_OCPN28438_n27080));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25008 (.Y(n16528),
	.A1(n26045),
	.A2(n26044),
	.B(n27168),
	.C(n16526));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25009 (.Y(n16529),
	.A1(n26942),
	.A2(n16531),
	.B(n16528),
	.C(w2_7_));
   NOR3x1_ASAP7_75t_L U25010 (.Y(n16575),
	.A(FE_OCPN28145_n16535),
	.B(FE_OFN28749_n),
	.C(FE_OCPN28053_sa10_1));
   NOR2xp33_ASAP7_75t_SRAM U25011 (.Y(n16537),
	.A(n16575),
	.B(FE_PSN8338_n19791));
   NOR2x1_ASAP7_75t_SL U25012 (.Y(n17216),
	.A(FE_OCPN28053_sa10_1),
	.B(FE_OCPN28145_n16535));
   NOR2x2_ASAP7_75t_SL U25013 (.Y(n19766),
	.A(FE_OFN26160_sa10_4),
	.B(FE_OFN130_sa10_5));
   NAND2x2_ASAP7_75t_SL U25014 (.Y(n23982),
	.A(FE_OFN27196_n),
	.B(n19766));
   NOR2xp33_ASAP7_75t_SRAM U25015 (.Y(n16536),
	.A(n23044),
	.B(n19672));
   NOR2x1p5_ASAP7_75t_SL U25016 (.Y(n16597),
	.A(FE_OCPN28053_sa10_1),
	.B(FE_OFN29161_n));
   NAND2x1p5_ASAP7_75t_SL U25017 (.Y(n23036),
	.A(FE_OFN29255_n),
	.B(n16597));
   NAND2x1p5_ASAP7_75t_SL U25018 (.Y(n19669),
	.A(FE_OCPN28157_n16534),
	.B(n24959));
   NOR2x1p5_ASAP7_75t_SL U25020 (.Y(n19756),
	.A(FE_OFN26587_n23011),
	.B(FE_OFN28916_sa10_4));
   NOR2xp33_ASAP7_75t_SRAM U25021 (.Y(n16539),
	.A(n19756),
	.B(FE_PSN8338_n19791));
   NOR2x1_ASAP7_75t_L U25022 (.Y(n19630),
	.A(FE_OCPN28323_FE_OFN16427_sa10_3),
	.B(n16647));
   NOR2x1p5_ASAP7_75t_SL U25023 (.Y(n24955),
	.A(FE_OFN27196_n),
	.B(n16647));
   NAND2x1p5_ASAP7_75t_SL U25024 (.Y(n23120),
	.A(n24955),
	.B(n24959));
   NAND3x2_ASAP7_75t_SL U25025 (.Y(n16616),
	.A(FE_OCPN29407_FE_OFN142_sa10_0),
	.B(n24955),
	.C(FE_OFN29043_n));
   A2O1A1Ixp33_ASAP7_75t_SL U25027 (.Y(n16543),
	.A1(n23982),
	.A2(n23012),
	.B(n16533),
	.C(n17201));
   NOR3xp33_ASAP7_75t_SRAM U25028 (.Y(n16546),
	.A(FE_OFN27094_n24956),
	.B(n23027),
	.C(n24976));
   NOR2x1_ASAP7_75t_SL U25029 (.Y(n23035),
	.A(FE_OFN28749_n),
	.B(FE_OCPN28145_n16535));
   NAND3xp33_ASAP7_75t_L U25030 (.Y(n16545),
	.A(n17219),
	.B(n21885),
	.C(n19653));
   NAND3xp33_ASAP7_75t_SRAM U25031 (.Y(n16607),
	.A(n24965),
	.B(n16546),
	.C(n24964));
   NOR2x1_ASAP7_75t_L U25032 (.Y(n16640),
	.A(n23981),
	.B(FE_OFN28832_n19789));
   NAND2x1p5_ASAP7_75t_SL U25033 (.Y(n17191),
	.A(FE_OCPN28052_sa10_1),
	.B(n23035));
   NOR2x1_ASAP7_75t_L U25034 (.Y(n21892),
	.A(n17191),
	.B(n19677));
   OAI222xp33_ASAP7_75t_R U25035 (.Y(n17200),
	.A1(FE_OCPN28052_sa10_1),
	.A2(n21888),
	.B1(FE_OCPN28157_n16534),
	.B2(n21888),
	.C1(n23035),
	.C2(n21888));
   NAND3xp33_ASAP7_75t_R U25036 (.Y(n16562),
	.A(n17210),
	.B(n16550),
	.C(n17226));
   A2O1A1Ixp33_ASAP7_75t_SL U25037 (.Y(n19767),
	.A1(n23980),
	.A2(FE_OFN27196_n),
	.B(n23948),
	.C(FE_OFN26161_sa10_4));
   NAND3xp33_ASAP7_75t_L U25038 (.Y(n16554),
	.A(n19767),
	.B(n23129),
	.C(n19683));
   NOR2x1_ASAP7_75t_L U25039 (.Y(n17221),
	.A(n23981),
	.B(n16552));
   OAI21xp33_ASAP7_75t_L U25040 (.Y(n23143),
	.A1(FE_OCPN29424_FE_OFN26039_sa10_2),
	.A2(n16616),
	.B(n19637));
   NOR2xp33_ASAP7_75t_SRAM U25041 (.Y(n16574),
	.A(n24943),
	.B(n24941));
   NOR3xp33_ASAP7_75t_SRAM U25042 (.Y(n16565),
	.A(n16610),
	.B(FE_OCPN28053_sa10_1),
	.C(FE_OCPN28145_n16535));
   NOR3xp33_ASAP7_75t_SL U25043 (.Y(n16570),
	.A(n17186),
	.B(FE_OCPN28358_n21899),
	.C(n19672));
   NAND3xp33_ASAP7_75t_SRAM U25044 (.Y(n16582),
	.A(n17216),
	.B(FE_OFN28912_n16534),
	.C(FE_OFN28751_n));
   OAI21xp5_ASAP7_75t_L U25045 (.Y(n21873),
	.A1(n19677),
	.A2(n16533),
	.B(n19644));
   NAND3xp33_ASAP7_75t_SL U25047 (.Y(n16568),
	.A(n16637),
	.B(n16582),
	.C(n16566));
   OAI21xp33_ASAP7_75t_R U25048 (.Y(n16567),
	.A1(n23982),
	.A2(n16533),
	.B(n17201));
   A2O1A1Ixp33_ASAP7_75t_SL U25049 (.Y(n24736),
	.A1(n21902),
	.A2(n19677),
	.B(n16648),
	.C(n23128));
   NOR2x1_ASAP7_75t_L U25050 (.Y(n16661),
	.A(n19772),
	.B(n24736));
   NOR3xp33_ASAP7_75t_SRAM U25051 (.Y(n16573),
	.A(n24952),
	.B(n24953),
	.C(n21874));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25052 (.Y(n16601),
	.A1(n16574),
	.A2(n16573),
	.B(n25139),
	.C(n16618));
   NOR2xp33_ASAP7_75t_SL U25054 (.Y(n16577),
	.A(n16576),
	.B(FE_OFN25956_n16575));
   NOR2xp33_ASAP7_75t_SL U25055 (.Y(n16585),
	.A(n16542),
	.B(n19663));
   NAND2xp5_ASAP7_75t_SL U25056 (.Y(n16591),
	.A(n16587),
	.B(n16586));
   NOR2x1_ASAP7_75t_L U25057 (.Y(n23043),
	.A(FE_OFN28751_n),
	.B(n16588));
   NOR2x1p5_ASAP7_75t_SL U25058 (.Y(n21893),
	.A(n23982),
	.B(n17191));
   NAND3xp33_ASAP7_75t_SL U25059 (.Y(n16633),
	.A(n16591),
	.B(n16590),
	.C(n23994));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25060 (.Y(n16605),
	.A1(n24974),
	.A2(n16607),
	.B(n16604),
	.C(FE_OFN16179_w3_19));
   OR2x2_ASAP7_75t_R U25061 (.Y(n16631),
	.A(FE_OFN25956_n16575),
	.B(n19677));
   NOR2xp33_ASAP7_75t_L U25062 (.Y(n23024),
	.A(n23996),
	.B(n23995));
   NOR2x1_ASAP7_75t_L U25063 (.Y(n19758),
	.A(n16610),
	.B(FE_OFN25956_n16575));
   OAI222xp33_ASAP7_75t_SL U25064 (.Y(n21886),
	.A1(FE_OFN27196_n),
	.A2(n19758),
	.B1(n19787),
	.B2(n19758),
	.C1(FE_OCPN28040_n19766),
	.C2(n19758));
   NOR2x1p5_ASAP7_75t_SL U25065 (.Y(n23133),
	.A(n16648),
	.B(n23012));
   NOR2xp33_ASAP7_75t_SRAM U25066 (.Y(n16622),
	.A(FE_OCPN27900_n23949),
	.B(n19670));
   NAND3xp33_ASAP7_75t_R U25067 (.Y(n16625),
	.A(n16637),
	.B(n19647),
	.C(n17217));
   NAND3xp33_ASAP7_75t_SRAM U25068 (.Y(n16636),
	.A(n16631),
	.B(n16630),
	.C(n16629));
   NAND3xp33_ASAP7_75t_R U25069 (.Y(n16634),
	.A(n23121),
	.B(n19647),
	.C(n16632));
   NOR2xp33_ASAP7_75t_SRAM U25070 (.Y(n16638),
	.A(n23138),
	.B(n23139));
   NOR2x1_ASAP7_75t_L U25071 (.Y(n21884),
	.A(n19663),
	.B(n16640));
   NAND3xp33_ASAP7_75t_SL U25072 (.Y(n16645),
	.A(n21884),
	.B(n16642),
	.C(n16641));
   NOR2xp33_ASAP7_75t_R U25073 (.Y(n16643),
	.A(FE_OFN27196_n),
	.B(FE_OCPN27636_sa10_4));
   OAI21xp5_ASAP7_75t_SL U25074 (.Y(n24892),
	.A1(n21902),
	.A2(n16533),
	.B(n16646));
   NOR3xp33_ASAP7_75t_L U25075 (.Y(n16649),
	.A(n24892),
	.B(n16653),
	.C(n23043));
   NOR2xp33_ASAP7_75t_SL U25076 (.Y(n16658),
	.A(n19787),
	.B(n23133));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25078 (.Y(n16671),
	.A1(FE_OCPN29587_n26857),
	.A2(FE_OFN29242_n26856),
	.B(FE_OCPN27377_n26853),
	.C(n26831));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25079 (.Y(n300),
	.A1(FE_OCPN29587_n26857),
	.A2(FE_OFN29242_n26856),
	.B(n16672),
	.C(n16671));
   NOR3xp33_ASAP7_75t_SRAM U25080 (.Y(n16683),
	.A(n24299),
	.B(n24297),
	.C(FE_OCPN28078_n24296));
   OAI21xp33_ASAP7_75t_SRAM U25081 (.Y(n16682),
	.A1(n16946),
	.A2(n24300),
	.B(FE_OCPN27544_sa33_4));
   NOR3xp33_ASAP7_75t_SL U25082 (.Y(n18142),
	.A(n16676),
	.B(FE_OFN28679_sa33_5),
	.C(n16947));
   NOR2x1_ASAP7_75t_L U25083 (.Y(n16832),
	.A(n18142),
	.B(n18109));
   NAND3xp33_ASAP7_75t_SRAM U25084 (.Y(n16678),
	.A(n16726),
	.B(n23550),
	.C(n16832));
   NAND3xp33_ASAP7_75t_R U25085 (.Y(n16834),
	.A(n16418),
	.B(n16417),
	.C(FE_OFN16430_sa33_3));
   NAND3xp33_ASAP7_75t_SL U25086 (.Y(n16688),
	.A(n18406),
	.B(n16686),
	.C(n16685));
   NAND2xp5_ASAP7_75t_SL U25087 (.Y(n18121),
	.A(n16427),
	.B(n17416));
   OAI21xp5_ASAP7_75t_SL U25088 (.Y(n16931),
	.A1(FE_OCPN27604_n16421),
	.A2(FE_OCPN27460_n16913),
	.B(n18121));
   NOR3x1_ASAP7_75t_L U25089 (.Y(n23560),
	.A(n16931),
	.B(n16936),
	.C(n24324));
   NAND2xp5_ASAP7_75t_SL U25090 (.Y(n16687),
	.A(n16893),
	.B(n23560));
   NOR2xp33_ASAP7_75t_SRAM U25091 (.Y(n16700),
	.A(n16430),
	.B(n18431));
   NOR2xp33_ASAP7_75t_L U25092 (.Y(n16693),
	.A(FE_OFN29101_n16418),
	.B(n17405));
   NOR2xp33_ASAP7_75t_SL U25093 (.Y(n16695),
	.A(n16430),
	.B(n17405));
   NAND3x1_ASAP7_75t_SL U25094 (.Y(n18443),
	.A(n16699),
	.B(n18128),
	.C(n16698));
   NOR2xp33_ASAP7_75t_SRAM U25095 (.Y(n16702),
	.A(n16873),
	.B(n18431));
   NOR2xp33_ASAP7_75t_SRAM U25096 (.Y(n16712),
	.A(n16946),
	.B(n16867));
   NOR2xp33_ASAP7_75t_R U25097 (.Y(n16713),
	.A(FE_OFN28999_n16923),
	.B(n16867));
   NAND3x1_ASAP7_75t_SL U25098 (.Y(n16930),
	.A(n18129),
	.B(FE_OFN16369_n16717),
	.C(n16716));
   NAND3xp33_ASAP7_75t_L U25099 (.Y(n16718),
	.A(n16918),
	.B(n23550),
	.C(n18121));
   NOR3xp33_ASAP7_75t_SL U25100 (.Y(n16741),
	.A(n16930),
	.B(n16728),
	.C(n23544));
   NAND3xp33_ASAP7_75t_SL U25101 (.Y(n16857),
	.A(n16725),
	.B(n16724),
	.C(n16846));
   NAND3xp33_ASAP7_75t_SL U25102 (.Y(n16739),
	.A(n16730),
	.B(n16729),
	.C(n26360));
   OAI21xp33_ASAP7_75t_SRAM U25103 (.Y(n16734),
	.A1(n16947),
	.A2(FE_OCPN27604_n16421),
	.B(n16953));
   NOR3xp33_ASAP7_75t_SRAM U25104 (.Y(n16735),
	.A(n16734),
	.B(n23535),
	.C(n18443));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25105 (.Y(n16743),
	.A1(n16742),
	.A2(n16741),
	.B(n24331),
	.C(n16740));
   NAND3xp33_ASAP7_75t_SL U25106 (.Y(n16767),
	.A(FE_OFN28698_sa21_1),
	.B(FE_OCPN27367_sa21_0),
	.C(sa21_2_));
   NAND2x1_ASAP7_75t_SL U25107 (.Y(n16806),
	.A(n16783),
	.B(FE_OFN25989_sa21_4));
   NOR2xp33_ASAP7_75t_R U25108 (.Y(n16752),
	.A(FE_OFN16153_n16747),
	.B(n16768));
   NAND2x1_ASAP7_75t_SL U25109 (.Y(n17881),
	.A(sa21_2_),
	.B(FE_OFN28698_sa21_1));
   NAND2x1p5_ASAP7_75t_L U25110 (.Y(n19867),
	.A(n16748),
	.B(FE_OFN16447_n16749));
   NOR2x1_ASAP7_75t_SL U25111 (.Y(n20007),
	.A(FE_OFN28698_sa21_1),
	.B(n16751));
   NAND2xp5_ASAP7_75t_SL U25112 (.Y(n23928),
	.A(FE_OCPN27328_sa21_2),
	.B(FE_OCPN29519_n));
   NOR2xp33_ASAP7_75t_SRAM U25114 (.Y(n16754),
	.A(n16763),
	.B(n16768));
   NOR2x1_ASAP7_75t_SL U25115 (.Y(n24257),
	.A(FE_OFN28678_sa21_3),
	.B(n22329));
   NAND2x1p5_ASAP7_75t_SL U25116 (.Y(n25351),
	.A(FE_OFN27157_n23928),
	.B(FE_OFN28779_n24257));
   NAND2x1_ASAP7_75t_SL U25117 (.Y(n17843),
	.A(FE_OFN28698_sa21_1),
	.B(FE_OCPN29450_sa21_0));
   NAND3xp33_ASAP7_75t_SL U25119 (.Y(n16759),
	.A(FE_OCPN27774_n25351),
	.B(n25350),
	.C(n20303));
   NAND2xp5_ASAP7_75t_SL U25120 (.Y(n23640),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(FE_OCPN28299_n));
   NOR2x1p5_ASAP7_75t_SL U25121 (.Y(n19979),
	.A(FE_OFN28678_sa21_3),
	.B(FE_OFN25989_sa21_4));
   NAND2x1p5_ASAP7_75t_L U25123 (.Y(n16762),
	.A(FE_OCPN27289_sa21_5),
	.B(n19979));
   NAND2x1p5_ASAP7_75t_SL U25124 (.Y(n17860),
	.A(FE_OFN28678_sa21_3),
	.B(n16763));
   NOR3x1_ASAP7_75t_SL U25125 (.Y(n23925),
	.A(n17860),
	.B(FE_OCPN29580_n),
	.C(FE_OCPN27556_n17843));
   NOR2x1_ASAP7_75t_R U25126 (.Y(n24881),
	.A(FE_OCPN27246_n22663),
	.B(n22662));
   A2O1A1Ixp33_ASAP7_75t_L U25127 (.Y(n16764),
	.A1(n23633),
	.A2(FE_OFN28820_n),
	.B(n16762),
	.C(n20298));
   NAND3xp33_ASAP7_75t_SRAM U25129 (.Y(n16770),
	.A(FE_OFN25993_n16767),
	.B(FE_OFN28985_sa21_5),
	.C(FE_OCPN29293_FE_OFN28678_sa21_3));
   NAND2x1p5_ASAP7_75t_SL U25130 (.Y(n19982),
	.A(FE_OCPN29265_FE_OFN28698_sa21_1),
	.B(n16760));
   NOR3xp33_ASAP7_75t_L U25131 (.Y(n16769),
	.A(n23661),
	.B(n23643),
	.C(FE_OCPN29279_n25353));
   OAI22xp33_ASAP7_75t_L U25132 (.Y(n22703),
	.A1(FE_OCPN27642_n16758),
	.A2(n16768),
	.B1(FE_OFN28779_n24257),
	.B2(n16768));
   AND3x1_ASAP7_75t_L U25133 (.Y(n19888),
	.A(n16770),
	.B(n16769),
	.C(n22703));
   NAND2x1p5_ASAP7_75t_L U25134 (.Y(n23650),
	.A(n16790),
	.B(FE_OCPN27642_n16758));
   NAND2xp5_ASAP7_75t_L U25135 (.Y(n22666),
	.A(FE_OCPN27616_n16760),
	.B(FE_OFN16447_n16749));
   NOR2x1_ASAP7_75t_L U25136 (.Y(n22679),
	.A(FE_OCPN29265_FE_OFN28698_sa21_1),
	.B(n22666));
   NAND2x1_ASAP7_75t_L U25137 (.Y(n22669),
	.A(n16771),
	.B(FE_OFN29023_n16750));
   NOR2x1_ASAP7_75t_SL U25138 (.Y(n16774),
	.A(FE_OCPN29414_n),
	.B(n16801));
   NOR2x1_ASAP7_75t_SL U25139 (.Y(n19886),
	.A(n19968),
	.B(n22349));
   NOR2xp33_ASAP7_75t_L U25140 (.Y(n16779),
	.A(n19967),
	.B(FE_OCPN27553_n19975));
   NAND3xp33_ASAP7_75t_L U25142 (.Y(n16781),
	.A(n19886),
	.B(n19881),
	.C(n19879));
   NAND2x1p5_ASAP7_75t_L U25143 (.Y(n19877),
	.A(n25350),
	.B(n17852));
   NOR3xp33_ASAP7_75t_SL U25144 (.Y(n16782),
	.A(n16781),
	.B(n19877),
	.C(n19876));
   NAND2x1p5_ASAP7_75t_R U25145 (.Y(n23656),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(FE_OCPN27631_n16774));
   NAND3xp33_ASAP7_75t_L U25146 (.Y(n19974),
	.A(FE_OCPN27289_sa21_5),
	.B(n19979),
	.C(n16748));
   NOR2xp33_ASAP7_75t_L U25147 (.Y(n16784),
	.A(FE_OFN25989_sa21_4),
	.B(FE_OFN62_sa21_3));
   NOR2x1_ASAP7_75t_L U25148 (.Y(n22331),
	.A(n16762),
	.B(n19982));
   O2A1O1Ixp33_ASAP7_75t_SRAM U25149 (.Y(n19864),
	.A1(FE_OFN29023_n16750),
	.A2(FE_OCPN28298_n),
	.B(FE_OCPN27690_n16757),
	.C(n22331));
   NAND3xp33_ASAP7_75t_SRAM U25150 (.Y(n16786),
	.A(n22353),
	.B(n23625),
	.C(n19864));
   NAND2x1p5_ASAP7_75t_L U25151 (.Y(n19973),
	.A(n16757),
	.B(FE_OCPN29512_n16750));
   NAND2x1p5_ASAP7_75t_SL U25152 (.Y(n25355),
	.A(n16790),
	.B(n16771));
   NAND3x2_ASAP7_75t_L U25153 (.Y(n16809),
	.A(n19973),
	.B(n19884),
	.C(n25355));
   NAND3xp33_ASAP7_75t_SL U25154 (.Y(n20315),
	.A(FE_OCPN27616_n16760),
	.B(FE_OFN28779_n24257),
	.C(FE_OCPN29265_FE_OFN28698_sa21_1));
   NOR2xp33_ASAP7_75t_SRAM U25155 (.Y(n16794),
	.A(FE_OCPN27553_n19975),
	.B(n17833));
   NAND2x1_ASAP7_75t_L U25156 (.Y(n20002),
	.A(n16808),
	.B(FE_OCPN27642_n16758));
   NOR3xp33_ASAP7_75t_SL U25157 (.Y(n23649),
	.A(n20318),
	.B(n22331),
	.C(n20325));
   NOR2x1_ASAP7_75t_L U25158 (.Y(n22696),
	.A(n17860),
	.B(n22662));
   NOR3xp33_ASAP7_75t_SL U25159 (.Y(n16807),
	.A(n22696),
	.B(n19892),
	.C(n22676));
   NAND3xp33_ASAP7_75t_SL U25160 (.Y(n20314),
	.A(n20009),
	.B(n23656),
	.C(n20327));
   OAI21xp5_ASAP7_75t_SL U25161 (.Y(n19896),
	.A1(n19982),
	.A2(n17860),
	.B(n19867));
   OAI21xp5_ASAP7_75t_L U25162 (.Y(n20334),
	.A1(n19982),
	.A2(n16762),
	.B(n22690));
   NOR2xp33_ASAP7_75t_SRAM U25163 (.Y(n16819),
	.A(FE_OFN16447_n16749),
	.B(n19890));
   O2A1O1Ixp5_ASAP7_75t_SL U25164 (.Y(n16826),
	.A1(n20011),
	.A2(n16825),
	.B(n26829),
	.C(n16824));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25165 (.Y(n16829),
	.A1(n25575),
	.A2(n24749),
	.B(FE_OCPN7631_n24750),
	.C(FE_OCPN28407_FE_OFN16433_w3_11));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25166 (.Y(n419),
	.A1(n25575),
	.A2(n24749),
	.B(n16830),
	.C(n16829));
   NAND2xp33_ASAP7_75t_SRAM U25167 (.Y(n16836),
	.A(n17408),
	.B(n18406));
   OAI21xp33_ASAP7_75t_SRAM U25168 (.Y(n16835),
	.A1(n16874),
	.A2(FE_OCPN28127_n16872),
	.B(n16834));
   NOR3xp33_ASAP7_75t_SRAM U25169 (.Y(n16849),
	.A(n16836),
	.B(n18144),
	.C(n16835));
   NOR2xp33_ASAP7_75t_SRAM U25170 (.Y(n16845),
	.A(n24300),
	.B(FE_OFN16241_n23552));
   NOR2xp33_ASAP7_75t_SRAM U25171 (.Y(n16839),
	.A(n18430),
	.B(n18107));
   NAND3xp33_ASAP7_75t_L U25172 (.Y(n16844),
	.A(n16868),
	.B(n16839),
	.C(n18149));
   A2O1A1Ixp33_ASAP7_75t_L U25173 (.Y(n18140),
	.A1(n16946),
	.A2(FE_OCPN29487_FE_OFN28694_sa33_4),
	.B(n16852),
	.C(FE_PSN8337_n16909));
   OAI22xp33_ASAP7_75t_SRAM U25174 (.Y(n18130),
	.A1(n16854),
	.A2(n16853),
	.B1(n16418),
	.B2(n16853));
   NOR3xp33_ASAP7_75t_SRAM U25175 (.Y(n16902),
	.A(n24326),
	.B(FE_OFN29040_n17404),
	.C(n24324));
   A2O1A1Ixp33_ASAP7_75t_L U25176 (.Y(n18120),
	.A1(n16417),
	.A2(n16946),
	.B(n18431),
	.C(FE_OFN25938_sa33_3));
   NOR3xp33_ASAP7_75t_SRAM U25177 (.Y(n16901),
	.A(n24325),
	.B(n24328),
	.C(n24327));
   NOR2xp33_ASAP7_75t_L U25179 (.Y(n16877),
	.A(FE_OFN28999_n16923),
	.B(n23539));
   OR2x2_ASAP7_75t_L U25180 (.Y(n16878),
	.A(n16946),
	.B(n23539));
   NAND3xp33_ASAP7_75t_SRAM U25181 (.Y(n16889),
	.A(n18406),
	.B(n16888),
	.C(n16887));
   NAND3xp33_ASAP7_75t_L U25182 (.Y(n24334),
	.A(n18123),
	.B(n16891),
	.C(n16890));
   NAND3xp33_ASAP7_75t_SRAM U25183 (.Y(n16897),
	.A(n18121),
	.B(n23528),
	.C(n16893));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25184 (.Y(n16905),
	.A1(n24610),
	.A2(n16907),
	.B(n16904),
	.C(w0_5_));
   A2O1A1Ixp33_ASAP7_75t_L U25185 (.Y(n16951),
	.A1(n16424),
	.A2(n16909),
	.B(FE_OCPN27593_n16908),
	.C(FE_OCPN29487_FE_OFN28694_sa33_4));
   NAND3xp33_ASAP7_75t_SRAM U25186 (.Y(n16911),
	.A(n16951),
	.B(n23528),
	.C(n16910));
   NOR3xp33_ASAP7_75t_SRAM U25187 (.Y(n16921),
	.A(n16912),
	.B(FE_OCPN28141_n),
	.C(FE_OFN28918_n16949));
   NAND3xp33_ASAP7_75t_SRAM U25188 (.Y(n16920),
	.A(n18405),
	.B(n16919),
	.C(n16918));
   NAND3xp33_ASAP7_75t_SL U25189 (.Y(n16926),
	.A(n18124),
	.B(n16921),
	.C(n18437));
   NOR2xp33_ASAP7_75t_SRAM U25190 (.Y(n16939),
	.A(FE_OCPN27555_n16422),
	.B(n24297));
   INVxp33_ASAP7_75t_SRAM U25191 (.Y(n16940),
	.A(n24613));
   NOR2xp33_ASAP7_75t_SRAM U25192 (.Y(n16941),
	.A(FE_OFN28592_n16427),
	.B(n24297));
   NAND3xp33_ASAP7_75t_SL U25193 (.Y(n16950),
	.A(n17423),
	.B(n16944),
	.C(n17408));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25194 (.Y(n16948),
	.A1(n16947),
	.A2(FE_OFN26545_n16447),
	.B(FE_OCPN27604_n16421),
	.C(n16945));
   AND3x1_ASAP7_75t_R U25195 (.Y(n16955),
	.A(n16953),
	.B(n16952),
	.C(n16951));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25196 (.Y(n16972),
	.A1(n23571),
	.A2(n16974),
	.B(FE_OCPN28024_n26427),
	.C(w0_0_));
   NAND2xp5_ASAP7_75t_SL U25197 (.Y(n20526),
	.A(FE_OFN28478_sa13_2),
	.B(n16977));
   NOR2x1p5_ASAP7_75t_SL U25198 (.Y(n19409),
	.A(FE_OCPN27836_n16976),
	.B(FE_OCPN28204_n20526));
   NOR2x1p5_ASAP7_75t_SL U25199 (.Y(n17159),
	.A(FE_OFN16268_sa13_3),
	.B(n16981));
   NAND2x2_ASAP7_75t_SL U25200 (.Y(n19360),
	.A(n16982),
	.B(FE_OFN26061_n));
   NAND2x1_ASAP7_75t_SL U25201 (.Y(n19372),
	.A(FE_OFN28801_n16978),
	.B(FE_OCPN28212_n16980));
   NOR2x1p5_ASAP7_75t_SL U25202 (.Y(n17170),
	.A(FE_OFN16268_sa13_3),
	.B(FE_OFN27065_n17059));
   NOR2x1p5_ASAP7_75t_L U25203 (.Y(n20514),
	.A(FE_OFN28478_sa13_2),
	.B(n16982));
   NAND2x1p5_ASAP7_75t_SL U25204 (.Y(n17121),
	.A(FE_OFN16181_sa13_5),
	.B(FE_OFN16268_sa13_3));
   NOR2x1p5_ASAP7_75t_SL U25205 (.Y(n25868),
	.A(FE_OFN28862_n),
	.B(n17121));
   NOR3x1_ASAP7_75t_SL U25206 (.Y(n17001),
	.A(FE_OFN28725_n16982),
	.B(FE_OCPN29426_FE_OFN16444_sa13_1),
	.C(FE_OFN28478_sa13_2));
   NAND2xp5_ASAP7_75t_SL U25207 (.Y(n19361),
	.A(FE_OFN27186_sa13_4),
	.B(n17159));
   NAND2x1_ASAP7_75t_SL U25208 (.Y(n17079),
	.A(FE_OFN16444_sa13_1),
	.B(n16982));
   NAND3xp33_ASAP7_75t_SL U25209 (.Y(n16985),
	.A(FE_OFN28913_n18247),
	.B(n19424),
	.C(n19423));
   NAND2x2_ASAP7_75t_SL U25210 (.Y(n17115),
	.A(FE_OFN16268_sa13_3),
	.B(n25545));
   NAND3xp33_ASAP7_75t_L U25211 (.Y(n16984),
	.A(FE_OFN28979_n),
	.B(n16983),
	.C(FE_OFN16181_sa13_5));
   NOR3x2_ASAP7_75t_SL U25212 (.Y(n16996),
	.A(FE_OFN16268_sa13_3),
	.B(FE_OFN16181_sa13_5),
	.C(FE_OFN27186_sa13_4));
   NAND3xp33_ASAP7_75t_SL U25213 (.Y(n18257),
	.A(FE_OCPN27761_n16977),
	.B(FE_OFN29234_n16996),
	.C(FE_OFN29173_n));
   NAND3x1_ASAP7_75t_SL U25214 (.Y(n16991),
	.A(FE_OFN28478_sa13_2),
	.B(FE_OFN28725_n16982),
	.C(FE_OCPN29426_FE_OFN16444_sa13_1));
   OAI21xp5_ASAP7_75t_SL U25215 (.Y(n17116),
	.A1(FE_OCPN27836_n16976),
	.A2(FE_OCPN28202_n16991),
	.B(n18263));
   NOR2xp33_ASAP7_75t_L U25216 (.Y(n16990),
	.A(n17171),
	.B(n17116));
   NAND2xp5_ASAP7_75t_SL U25219 (.Y(n24165),
	.A(n16983),
	.B(n16996));
   NOR2x1_ASAP7_75t_L U25221 (.Y(n18283),
	.A(n16989),
	.B(n16997));
   NOR2x1_ASAP7_75t_SL U25222 (.Y(n17017),
	.A(n18283),
	.B(n16998));
   NOR3xp33_ASAP7_75t_SRAM U25223 (.Y(n17000),
	.A(n16999),
	.B(n19430),
	.C(n18267));
   NAND2x2_ASAP7_75t_L U25224 (.Y(n25285),
	.A(FE_OFN28801_n16978),
	.B(n19399));
   NOR2xp33_ASAP7_75t_SL U25225 (.Y(n17003),
	.A(n16983),
	.B(n24155));
   NAND2x1p5_ASAP7_75t_SL U25226 (.Y(n17161),
	.A(n25868),
	.B(n16983));
   A2O1A1Ixp33_ASAP7_75t_SL U25227 (.Y(n17008),
	.A1(FE_OCPN29490_n17001),
	.A2(n19360),
	.B(FE_OCPN29446_n17115),
	.C(n17089));
   NAND3xp33_ASAP7_75t_R U25228 (.Y(n17015),
	.A(n20532),
	.B(n20510),
	.C(n18926));
   NAND2x1_ASAP7_75t_SL U25229 (.Y(n18940),
	.A(n17170),
	.B(n16980));
   NOR2xp33_ASAP7_75t_SRAM U25230 (.Y(n17018),
	.A(n17082),
	.B(n19381));
   NOR2xp67_ASAP7_75t_SL U25231 (.Y(n17026),
	.A(n20506),
	.B(n17019));
   NOR2xp33_ASAP7_75t_SRAM U25232 (.Y(n17022),
	.A(FE_OCPN29510_n16996),
	.B(n19410));
   NAND2x1_ASAP7_75t_SL U25234 (.Y(n19374),
	.A(n25285),
	.B(n17161));
   NOR3xp33_ASAP7_75t_L U25235 (.Y(n18930),
	.A(FE_OCPN28204_n20526),
	.B(FE_OFN28862_n),
	.C(n17121));
   NAND2x1p5_ASAP7_75t_R U25236 (.Y(n27102),
	.A(FE_OFN128_sa13_7),
	.B(n19359));
   NOR2xp33_ASAP7_75t_R U25237 (.Y(n17035),
	.A(FE_OFN29173_n),
	.B(n25875));
   NOR2xp33_ASAP7_75t_R U25238 (.Y(n17037),
	.A(n24156),
	.B(n25875));
   NOR3x1_ASAP7_75t_SL U25239 (.Y(n25197),
	.A(n18286),
	.B(n18269),
	.C(n20490));
   NAND2x1_ASAP7_75t_R U25240 (.Y(n26959),
	.A(FE_OFN128_sa13_7),
	.B(FE_OFN16389_n19359));
   INVxp33_ASAP7_75t_SRAM U25241 (.Y(n17041),
	.A(n25225));
   NAND3xp33_ASAP7_75t_SRAM U25242 (.Y(n17044),
	.A(n25222),
	.B(n25221),
	.C(n17041));
   NOR2xp33_ASAP7_75t_SL U25243 (.Y(n25219),
	.A(n20527),
	.B(n17042));
   OAI21xp5_ASAP7_75t_L U25244 (.Y(n25218),
	.A1(FE_OCPN28202_n16991),
	.A2(FE_OCPN27836_n16976),
	.B(n17102));
   NOR3xp33_ASAP7_75t_SRAM U25245 (.Y(n17051),
	.A(n17044),
	.B(FE_OFN16220_n25219),
	.C(FE_OFN29228_n25218));
   NOR2xp33_ASAP7_75t_SL U25246 (.Y(n18242),
	.A(n24156),
	.B(n19409));
   NOR2xp33_ASAP7_75t_SL U25247 (.Y(n17046),
	.A(n20491),
	.B(n18954));
   OAI21xp5_ASAP7_75t_L U25249 (.Y(n17165),
	.A1(FE_OFN28583_n17001),
	.A2(FE_OCPN29446_n17115),
	.B(n17146));
   O2A1O1Ixp33_ASAP7_75t_R U25250 (.Y(n17048),
	.A1(FE_OFN16162_n25869),
	.A2(FE_OCPN27761_n16977),
	.B(n16996),
	.C(n19434));
   OAI21xp33_ASAP7_75t_SRAM U25251 (.Y(n17062),
	.A1(FE_OCPN29490_n17001),
	.A2(FE_OFN27065_n17059),
	.B(n17058));
   O2A1O1Ixp5_ASAP7_75t_SL U25252 (.Y(n17061),
	.A1(n19399),
	.A2(n17060),
	.B(FE_OFN28801_n16978),
	.C(n19379));
   NOR3x2_ASAP7_75t_SL U25253 (.Y(n20513),
	.A(FE_OCPN29446_n17115),
	.B(FE_OFN28809_n),
	.C(FE_OCPN29340_n17079));
   NOR3xp33_ASAP7_75t_SRAM U25254 (.Y(n17063),
	.A(n17062),
	.B(FE_OFN28622_n25870),
	.C(FE_OCPN8206_n25544));
   NAND3xp33_ASAP7_75t_SRAM U25255 (.Y(n17113),
	.A(n25551),
	.B(n17063),
	.C(n25549));
   NAND3xp33_ASAP7_75t_SL U25256 (.Y(n17081),
	.A(n20525),
	.B(FE_OCPN8228_n24165),
	.C(n18261));
   NOR3xp33_ASAP7_75t_R U25257 (.Y(n17067),
	.A(FE_OCPN28204_n20526),
	.B(FE_OFN28862_n),
	.C(n17103));
   NOR2x1_ASAP7_75t_L U25258 (.Y(n17075),
	.A(n20522),
	.B(n20523));
   NAND3x1_ASAP7_75t_SL U25259 (.Y(n18947),
	.A(n16983),
	.B(FE_OCPN28121_n16975),
	.C(FE_OFN28491_sa13_3));
   NAND3x1_ASAP7_75t_SL U25262 (.Y(n17114),
	.A(n17080),
	.B(n19385),
	.C(n17132));
   NOR2x1_ASAP7_75t_L U25263 (.Y(n18921),
	.A(FE_OFN28862_n),
	.B(n17142));
   NOR3xp33_ASAP7_75t_SRAM U25264 (.Y(n17084),
	.A(n17083),
	.B(n17082),
	.C(n19381));
   A2O1A1Ixp33_ASAP7_75t_SL U25265 (.Y(n17131),
	.A1(FE_OFN16162_n25869),
	.A2(FE_OCPN28121_n16975),
	.B(n18269),
	.C(FE_OFN28979_n));
   NOR2xp33_ASAP7_75t_SRAM U25266 (.Y(n17086),
	.A(n19430),
	.B(n19379));
   NOR2xp33_ASAP7_75t_SRAM U25267 (.Y(n17088),
	.A(n18286),
	.B(n20513));
   NAND2x1_ASAP7_75t_SL U25268 (.Y(n18960),
	.A(n17089),
	.B(n19385));
   NOR2xp33_ASAP7_75t_R U25269 (.Y(n17090),
	.A(n19399),
	.B(n18960));
   NOR2xp33_ASAP7_75t_SL U25271 (.Y(n17092),
	.A(n17091),
	.B(n18960));
   OAI22xp33_ASAP7_75t_SRAM U25272 (.Y(n17108),
	.A1(n25555),
	.A2(n27095),
	.B1(n25554),
	.B2(n27095));
   NAND3xp33_ASAP7_75t_SL U25273 (.Y(n17097),
	.A(n25197),
	.B(n17095),
	.C(n18926));
   NOR2xp33_ASAP7_75t_L U25274 (.Y(n17096),
	.A(n19410),
	.B(n18921));
   NOR2xp33_ASAP7_75t_SRAM U25275 (.Y(n17106),
	.A(FE_OFN28548_n27092),
	.B(n25539));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25276 (.Y(n325),
	.A1(n26915),
	.A2(n17113),
	.B(n17112),
	.C(n17111));
   O2A1O1Ixp5_ASAP7_75t_SL U25277 (.Y(n24166),
	.A1(FE_OFN28801_n16978),
	.A2(FE_OFN29074_n17170),
	.B(n16983),
	.C(n17114));
   NOR2xp33_ASAP7_75t_SRAM U25278 (.Y(n19382),
	.A(FE_OCPN29490_n17001),
	.B(n17115));
   NOR2xp33_ASAP7_75t_SRAM U25279 (.Y(n24163),
	.A(n19410),
	.B(n19382));
   NAND3xp33_ASAP7_75t_SRAM U25280 (.Y(n17119),
	.A(FE_OCPN7613_n24166),
	.B(n24163),
	.C(n25197));
   NAND2xp33_ASAP7_75t_SRAM U25281 (.Y(n17118),
	.A(n18924),
	.B(n25872));
   NAND3xp33_ASAP7_75t_L U25282 (.Y(n24157),
	.A(n17162),
	.B(n17117),
	.C(FE_OFN29035_n17116));
   NOR3xp33_ASAP7_75t_SRAM U25283 (.Y(n17127),
	.A(n17119),
	.B(n17118),
	.C(n24157));
   NAND3xp33_ASAP7_75t_SRAM U25284 (.Y(n17184),
	.A(n17127),
	.B(n24165),
	.C(n24164));
   A2O1A1Ixp33_ASAP7_75t_L U25285 (.Y(n18262),
	.A1(n16980),
	.A2(n16975),
	.B(n19379),
	.C(FE_OFN28979_n));
   OAI21xp33_ASAP7_75t_L U25286 (.Y(n18277),
	.A1(FE_OCPN27836_n16976),
	.A2(FE_OFN28738_n16989),
	.B(n18256));
   NOR2xp33_ASAP7_75t_SRAM U25287 (.Y(n17133),
	.A(n16983),
	.B(n18283));
   NOR2xp33_ASAP7_75t_SRAM U25288 (.Y(n17135),
	.A(FE_OFN28801_n16978),
	.B(n18283));
   NOR2x1_ASAP7_75t_SL U25289 (.Y(n17141),
	.A(n20495),
	.B(n25287));
   NOR3xp33_ASAP7_75t_SL U25291 (.Y(n17143),
	.A(n19408),
	.B(n18954),
	.C(FE_OCPN27589_n25987));
   NOR2xp33_ASAP7_75t_L U25292 (.Y(n17153),
	.A(n16983),
	.B(n17154));
   A2O1A1Ixp33_ASAP7_75t_SL U25293 (.Y(n20521),
	.A1(FE_OFN28738_n16989),
	.A2(FE_OCPN28202_n16991),
	.B(FE_OCPN5143_n19361),
	.C(n18940));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25295 (.Y(n17160),
	.A1(FE_OFN28801_n16978),
	.A2(FE_OCPN27761_n16977),
	.B(n18283),
	.C(FE_OFN28809_n));
   OAI22xp33_ASAP7_75t_SRAM U25296 (.Y(n17179),
	.A1(FE_OCPN29425_n24172),
	.A2(n27102),
	.B1(n24171),
	.B2(n27102));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25297 (.Y(n17182),
	.A1(n26915),
	.A2(n17184),
	.B(n17181),
	.C(w2_21_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25298 (.Y(n311),
	.A1(n26915),
	.A2(n17184),
	.B(n17183),
	.C(n17182));
   NOR2xp33_ASAP7_75t_SRAM U25299 (.Y(n17187),
	.A(n23995),
	.B(n17186));
   A2O1A1Ixp33_ASAP7_75t_L U25300 (.Y(n19665),
	.A1(n17216),
	.A2(FE_OCPN28157_n16534),
	.B(n24726),
	.C(FE_OFN29255_n));
   NOR3xp33_ASAP7_75t_SRAM U25301 (.Y(n17192),
	.A(n17191),
	.B(FE_OFN130_sa10_5),
	.C(FE_OFN27196_n));
   NOR3xp33_ASAP7_75t_L U25302 (.Y(n17193),
	.A(n17192),
	.B(n24958),
	.C(n23997));
   NAND3xp33_ASAP7_75t_L U25303 (.Y(n17199),
	.A(n19665),
	.B(n19660),
	.C(n21877));
   NOR2xp33_ASAP7_75t_L U25304 (.Y(n17195),
	.A(n19791),
	.B(n21893));
   NOR2x1_ASAP7_75t_L U25305 (.Y(n24896),
	.A(n19754),
	.B(FE_OFN29154_n19753));
   NAND2x1_ASAP7_75t_SL U25306 (.Y(n19679),
	.A(n19669),
	.B(n17201));
   NOR2xp33_ASAP7_75t_R U25307 (.Y(n17204),
	.A(n23980),
	.B(n23137));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25308 (.Y(n17233),
	.A1(FE_OCPN29586_n26857),
	.A2(n25044),
	.B(FE_OCPN29433_n25040),
	.C(FE_OFN51_w3_18));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25309 (.Y(n339),
	.A1(FE_OCPN29586_n26857),
	.A2(n25044),
	.B(n17234),
	.C(n17233));
   NOR2x1p5_ASAP7_75t_SL U25310 (.Y(n17271),
	.A(FE_OCPN29302_sa00_4),
	.B(FE_OCPN27224_sa00_5));
   NAND2x1p5_ASAP7_75t_SL U25311 (.Y(n17282),
	.A(n19149),
	.B(FE_OCPN29302_sa00_4));
   NOR2x1_ASAP7_75t_SL U25312 (.Y(n18631),
	.A(FE_OFN28744_FE_OCPN27908),
	.B(FE_OFN28514_sa00_1));
   NAND2x1p5_ASAP7_75t_SL U25313 (.Y(n18651),
	.A(FE_PSN8275_FE_OCPN27818_n17267),
	.B(n18631));
   NOR2xp33_ASAP7_75t_R U25315 (.Y(n17240),
	.A(FE_OFN28835_n),
	.B(n19840));
   NOR2x1_ASAP7_75t_SL U25316 (.Y(n21151),
	.A(FE_OCPN29302_sa00_4),
	.B(sa00_5_));
   NAND2xp5_ASAP7_75t_SL U25317 (.Y(n19098),
	.A(FE_OCPN29463_n),
	.B(n21151));
   NAND2x1p5_ASAP7_75t_SL U25318 (.Y(n17237),
	.A(FE_OFN29249_n),
	.B(n17271));
   A2O1A1Ixp33_ASAP7_75t_L U25321 (.Y(n17239),
	.A1(FE_OCPN28250_n19573),
	.A2(FE_OCPN27649_n17236),
	.B(FE_OCPN27951_n19098),
	.C(n19113));
   NOR2xp33_ASAP7_75t_SRAM U25322 (.Y(n17242),
	.A(n19122),
	.B(n19840));
   NAND3xp33_ASAP7_75t_SRAM U25324 (.Y(n17250),
	.A(FE_OCPN29376_n24099),
	.B(n19574),
	.C(n17246));
   A2O1A1Ixp33_ASAP7_75t_L U25325 (.Y(n24102),
	.A1(n19116),
	.A2(FE_OCPN29346_n12998),
	.B(FE_OCPN27703_n19847),
	.C(FE_OCPN27908_FE_OFN16156_sa00_2));
   NOR2x1_ASAP7_75t_SL U25327 (.Y(n21445),
	.A(FE_OCPN29385_n),
	.B(n18640));
   NOR3xp33_ASAP7_75t_SRAM U25329 (.Y(n17257),
	.A(n17250),
	.B(n24517),
	.C(FE_OFN28556_n24516));
   NOR2x1p5_ASAP7_75t_SL U25330 (.Y(n19834),
	.A(FE_OCPN29463_n),
	.B(FE_OCPN29260_sa00_5));
   NAND3xp33_ASAP7_75t_SL U25331 (.Y(n17261),
	.A(n18739),
	.B(n19834),
	.C(FE_OCPN29302_sa00_4));
   NAND3xp33_ASAP7_75t_L U25332 (.Y(n17256),
	.A(n18629),
	.B(FE_OCPN29553_n19602),
	.C(n21181));
   NOR2xp33_ASAP7_75t_SRAM U25333 (.Y(n17253),
	.A(n21150),
	.B(n19818));
   NAND2xp5_ASAP7_75t_L U25334 (.Y(n18773),
	.A(n17254),
	.B(FE_OCPN28021_n21445));
   NAND3xp33_ASAP7_75t_SRAM U25336 (.Y(n17314),
	.A(n24100),
	.B(n17257),
	.C(n25258));
   NAND3xp33_ASAP7_75t_SRAM U25337 (.Y(n17259),
	.A(n24085),
	.B(FE_OFN28767_n26103),
	.C(n18632));
   AND3x1_ASAP7_75t_SRAM U25338 (.Y(n17258),
	.A(FE_OCPN29542_n21151),
	.B(FE_OCPN27679_n18631),
	.C(FE_OCPN29396_n19149));
   NAND3xp33_ASAP7_75t_SRAM U25339 (.Y(n24093),
	.A(n21468),
	.B(FE_OCPN29553_n19602),
	.C(n19114));
   OAI21xp5_ASAP7_75t_SL U25340 (.Y(n18623),
	.A1(FE_OCPN27951_n19098),
	.A2(FE_OCPN27649_n17236),
	.B(n17260));
   NAND3xp33_ASAP7_75t_SL U25341 (.Y(n18770),
	.A(n19116),
	.B(FE_OCPN29346_n12998),
	.C(FE_OCPN27908_FE_OFN16156_sa00_2));
   NOR3xp33_ASAP7_75t_SL U25343 (.Y(n17269),
	.A(n21165),
	.B(FE_OFN29027_n19135),
	.C(n19588));
   NAND3xp33_ASAP7_75t_R U25344 (.Y(n19614),
	.A(FE_OFN42_sa00_0),
	.B(n17266),
	.C(n17245));
   OAI22xp33_ASAP7_75t_L U25345 (.Y(n17268),
	.A1(FE_OCPN29346_n12998),
	.A2(n19605),
	.B1(FE_OFN28835_n),
	.B2(n19605));
   NAND3xp33_ASAP7_75t_L U25346 (.Y(n17270),
	.A(n17269),
	.B(n19614),
	.C(n17268));
   A2O1A1Ixp33_ASAP7_75t_SL U25347 (.Y(n24089),
	.A1(n19097),
	.A2(FE_OCPN27518_n17251),
	.B(FE_OCPN27951_n19098),
	.C(FE_OCPN29376_n24099));
   NAND2xp5_ASAP7_75t_L U25348 (.Y(n19615),
	.A(FE_OCPN28021_n21445),
	.B(n12998));
   OAI22xp33_ASAP7_75t_SRAM U25349 (.Y(n19104),
	.A1(FE_OCPN28021_n21445),
	.A2(n21150),
	.B1(FE_OCPN28389_n21479),
	.B2(n21150));
   AND3x1_ASAP7_75t_L U25350 (.Y(n17309),
	.A(n17272),
	.B(n19615),
	.C(n19104));
   NAND3xp33_ASAP7_75t_L U25351 (.Y(n17295),
	.A(FE_PSN8312_n21442),
	.B(n18764),
	.C(n24101));
   NOR2xp33_ASAP7_75t_L U25352 (.Y(n17277),
	.A(FE_OFN28744_FE_OCPN27908),
	.B(n19090));
   A2O1A1Ixp33_ASAP7_75t_SL U25353 (.Y(n17276),
	.A1(n17275),
	.A2(FE_OCPN29415_n17237),
	.B(FE_OFN29062_n18651),
	.C(n21441));
   NOR2xp33_ASAP7_75t_L U25354 (.Y(n17279),
	.A(n19847),
	.B(n19090));
   NOR2x1p5_ASAP7_75t_SL U25355 (.Y(n21455),
	.A(FE_OFN26651_n19573),
	.B(n17275));
   NAND3x1_ASAP7_75t_SL U25357 (.Y(n19142),
	.A(n19825),
	.B(n17293),
	.C(n21472));
   NOR3xp33_ASAP7_75t_L U25358 (.Y(n17299),
	.A(n17297),
	.B(n21439),
	.C(FE_OFN28958_n17261));
   NOR2x1_ASAP7_75t_L U25359 (.Y(n19129),
	.A(FE_OCPN27951_n19098),
	.B(FE_OCPN28250_n19573));
   A2O1A1Ixp33_ASAP7_75t_L U25360 (.Y(n17302),
	.A1(FE_OFN28796_n17301),
	.A2(FE_OCPN27338_n19149),
	.B(n21154),
	.C(FE_OCPN29542_n21151));
   NOR2xp33_ASAP7_75t_L U25361 (.Y(n17303),
	.A(n19129),
	.B(n19596));
   NAND3xp33_ASAP7_75t_SL U25362 (.Y(n17306),
	.A(n21463),
	.B(n17304),
	.C(n17303));
   A2O1A1Ixp33_ASAP7_75t_R U25363 (.Y(n24529),
	.A1(n24626),
	.A2(n24625),
	.B(n26777),
	.C(n17310));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25365 (.Y(n17312),
	.A1(n27127),
	.A2(n17314),
	.B(n24529),
	.C(w0_26_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25366 (.Y(n324),
	.A1(n27127),
	.A2(n17314),
	.B(n17313),
	.C(n17312));
   NAND2x2_ASAP7_75t_L U25367 (.Y(n21561),
	.A(FE_OCPN27423_sa01_0),
	.B(FE_OFN125_sa01_1));
   NOR2x1p5_ASAP7_75t_SL U25368 (.Y(n18671),
	.A(FE_OFN25950_sa01_2),
	.B(n21561));
   NAND2x2_ASAP7_75t_SL U25369 (.Y(n22450),
	.A(n17326),
	.B(n21553));
   NAND2x1p5_ASAP7_75t_SL U25370 (.Y(n18710),
	.A(FE_OCPN27423_sa01_0),
	.B(n18707));
   NOR2x1_ASAP7_75t_SL U25371 (.Y(n18726),
	.A(n22450),
	.B(n18710));
   NOR2xp33_ASAP7_75t_SRAM U25372 (.Y(n17320),
	.A(FE_OCPN29455_n18671),
	.B(n18726));
   NAND2x1p5_ASAP7_75t_L U25374 (.Y(n18684),
	.A(FE_OFN26054_sa01_3),
	.B(n17326));
   NOR2xp33_ASAP7_75t_SRAM U25375 (.Y(n17323),
	.A(n17321),
	.B(n18726));
   NAND3xp33_ASAP7_75t_SL U25376 (.Y(n22598),
	.A(FE_OCPN28217_sa01_5),
	.B(n17326),
	.C(FE_OFN16141_sa01_3));
   NOR2x1p5_ASAP7_75t_SL U25377 (.Y(n26454),
	.A(FE_OCPN27423_sa01_0),
	.B(n17345));
   NAND3xp33_ASAP7_75t_SL U25378 (.Y(n17328),
	.A(n17327),
	.B(n23104),
	.C(n20415));
   NOR2x1p5_ASAP7_75t_SL U25379 (.Y(n20409),
	.A(FE_OCPN27399_n22598),
	.B(FE_OCPN8237_n21561));
   NAND2x1_ASAP7_75t_L U25380 (.Y(n26452),
	.A(FE_OFN27152_n17315),
	.B(n20409));
   NAND3x1_ASAP7_75t_SL U25381 (.Y(n21534),
	.A(FE_OCPN29408_n22461),
	.B(FE_OCPN27871_n17317),
	.C(FE_OFN26054_sa01_3));
   NAND3x1_ASAP7_75t_SL U25382 (.Y(n21549),
	.A(n26452),
	.B(n18721),
	.C(n21534));
   NOR2x1p5_ASAP7_75t_SL U25383 (.Y(n17359),
	.A(FE_OFN28672_sa01_2),
	.B(FE_OFN28718_sa01_1));
   NOR2x1p5_ASAP7_75t_SL U25385 (.Y(n18714),
	.A(FE_OFN27072_n18671),
	.B(FE_OFN27052_n21551));
   OAI22xp33_ASAP7_75t_R U25386 (.Y(n17332),
	.A1(n17329),
	.A2(n18714),
	.B1(FE_OCPN8219_n22197),
	.B2(n18714));
   NOR2x1p5_ASAP7_75t_SL U25387 (.Y(n23059),
	.A(FE_OCPN29429_FE_OFN16141_sa01_3),
	.B(n17389));
   NOR2x1p5_ASAP7_75t_L U25388 (.Y(n20387),
	.A(n17330),
	.B(n18667));
   OAI22xp5_ASAP7_75t_L U25389 (.Y(n21559),
	.A1(n26454),
	.A2(n20387),
	.B1(FE_OFN29135_n21551),
	.B2(n20387));
   NAND3xp33_ASAP7_75t_SL U25390 (.Y(n17333),
	.A(n17332),
	.B(n24396),
	.C(n21559));
   NOR2x1p5_ASAP7_75t_SL U25391 (.Y(n27006),
	.A(FE_OCPN27399_n22598),
	.B(n18667));
   NOR2x1p5_ASAP7_75t_L U25392 (.Y(n18717),
	.A(FE_OCPN29320_n22461),
	.B(n17330));
   NAND3xp33_ASAP7_75t_SRAM U25393 (.Y(n17334),
	.A(n17331),
	.B(n17329),
	.C(FE_OFN28672_sa01_2));
   OAI21x1_ASAP7_75t_L U25394 (.Y(n24390),
	.A1(n17335),
	.A2(n17329),
	.B(FE_OCPN27988_n26454));
   A2O1A1Ixp33_ASAP7_75t_SL U25395 (.Y(n22193),
	.A1(FE_OCPN29333_n17330),
	.A2(FE_OFN27052_n21551),
	.B(FE_OFN26648_n22197),
	.C(n24390));
   NOR2x1_ASAP7_75t_L U25396 (.Y(n22602),
	.A(n17318),
	.B(n18667));
   NOR2x1_ASAP7_75t_L U25397 (.Y(n22196),
	.A(FE_OCPN28000_n22450),
	.B(n23107));
   NOR2xp33_ASAP7_75t_R U25398 (.Y(n17336),
	.A(n17386),
	.B(n22196));
   NOR2xp33_ASAP7_75t_L U25399 (.Y(n17338),
	.A(FE_OFN26054_sa01_3),
	.B(n22196));
   NAND3xp33_ASAP7_75t_SL U25400 (.Y(n17342),
	.A(n23102),
	.B(n17341),
	.C(n18675));
   NOR2x1_ASAP7_75t_SL U25401 (.Y(n26998),
	.A(n17355),
	.B(n17342));
   NAND3x1_ASAP7_75t_SL U25402 (.Y(n24225),
	.A(n18685),
	.B(n23079),
	.C(n26998));
   NOR2xp33_ASAP7_75t_SRAM U25403 (.Y(n17344),
	.A(n17343),
	.B(n24225));
   NAND3xp33_ASAP7_75t_SL U25404 (.Y(n27003),
	.A(n21553),
	.B(n26454),
	.C(n17326));
   NOR3xp33_ASAP7_75t_L U25405 (.Y(n17346),
	.A(FE_OCPN28380_n22433),
	.B(n21563),
	.C(n22584));
   OA21x2_ASAP7_75t_SL U25406 (.Y(n22198),
	.A1(FE_OFN26648_n22197),
	.A2(FE_OFN25878_n17329),
	.B(n17346));
   NOR2xp33_ASAP7_75t_SL U25407 (.Y(n17348),
	.A(n17386),
	.B(FE_OFN16252_n27003));
   NOR3x1_ASAP7_75t_SL U25408 (.Y(n26459),
	.A(n17354),
	.B(FE_OCPN8222_n27006),
	.C(n17353));
   NOR2xp33_ASAP7_75t_SRAM U25409 (.Y(n17358),
	.A(FE_OFN29135_n21551),
	.B(n18726));
   NOR2xp33_ASAP7_75t_SRAM U25410 (.Y(n17360),
	.A(n17359),
	.B(n18726));
   NOR2x1p5_ASAP7_75t_SL U25411 (.Y(n22436),
	.A(n17318),
	.B(FE_OFN27072_n18671));
   NOR2xp33_ASAP7_75t_SRAM U25412 (.Y(n17363),
	.A(n21553),
	.B(n22436));
   AND2x4_ASAP7_75t_SL U25413 (.Y(n20361),
	.A(FE_OCPN28310_n22585),
	.B(n22414));
   NOR2xp33_ASAP7_75t_R U25414 (.Y(n17364),
	.A(FE_OCPN29388_n22461),
	.B(n22436));
   OR2x2_ASAP7_75t_R U25416 (.Y(n23078),
	.A(n22598),
	.B(FE_OCPN29406_n18710));
   A2O1A1Ixp33_ASAP7_75t_SL U25417 (.Y(n22415),
	.A1(FE_OFN28594_n26454),
	.A2(FE_OFN26054_sa01_3),
	.B(n18714),
	.C(FE_OCPN27871_n17317));
   NOR3xp33_ASAP7_75t_SL U25418 (.Y(n17370),
	.A(n22451),
	.B(n22582),
	.C(n22602));
   NAND3xp33_ASAP7_75t_SL U25419 (.Y(n17371),
	.A(n23079),
	.B(n23078),
	.C(n17370));
   NOR2x1p5_ASAP7_75t_SL U25420 (.Y(n23087),
	.A(FE_OFN27152_n17315),
	.B(n22191));
   NOR2x1p5_ASAP7_75t_L U25421 (.Y(n23099),
	.A(n22450),
	.B(FE_OFN27072_n18671));
   OAI21xp33_ASAP7_75t_SRAM U25422 (.Y(n17379),
	.A1(FE_OFN27072_n18671),
	.A2(FE_OCPN29333_n17330),
	.B(n25063));
   NOR2xp33_ASAP7_75t_SRAM U25423 (.Y(n17372),
	.A(n21563),
	.B(FE_OCPN28380_n22433));
   NAND2xp5_ASAP7_75t_R U25424 (.Y(n18677),
	.A(n17329),
	.B(FE_OCPN27988_n26454));
   NOR2x1_ASAP7_75t_SL U25425 (.Y(n23062),
	.A(FE_OCPN27399_n22598),
	.B(FE_OFN26648_n22197));
   NOR2x1p5_ASAP7_75t_SL U25426 (.Y(n22438),
	.A(n23107),
	.B(FE_OCPN29334_n17330));
   NOR3xp33_ASAP7_75t_SL U25427 (.Y(n17374),
	.A(n22601),
	.B(n20404),
	.C(n22438));
   NAND2xp5_ASAP7_75t_L U25428 (.Y(n27004),
	.A(sa01_6_),
	.B(n17392));
   NOR3xp33_ASAP7_75t_SRAM U25429 (.Y(n17380),
	.A(FE_OCPN28365_n21549),
	.B(n23062),
	.C(FE_OCPN8236_n22438));
   NOR2xp33_ASAP7_75t_L U25430 (.Y(n22416),
	.A(n17386),
	.B(n23099));
   NOR2xp33_ASAP7_75t_R U25431 (.Y(n22418),
	.A(FE_OCPN27871_n17317),
	.B(n23099));
   NOR2x1_ASAP7_75t_L U25432 (.Y(n18672),
	.A(n18698),
	.B(n18717));
   NAND3xp33_ASAP7_75t_L U25433 (.Y(n21541),
	.A(FE_OFN28736_FE_OCPN28216_sa01_5),
	.B(n17386),
	.C(FE_OFN26054_sa01_3));
   NAND3xp33_ASAP7_75t_SL U25434 (.Y(n17391),
	.A(n18672),
	.B(n21541),
	.C(n17388));
   NOR2x1_ASAP7_75t_L U25435 (.Y(n18704),
	.A(n23093),
	.B(n22602));
   NAND3xp33_ASAP7_75t_SL U25436 (.Y(n17390),
	.A(n22183),
	.B(n18677),
	.C(n18704));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25437 (.Y(n17395),
	.A1(n26282),
	.A2(n24126),
	.B(n24123),
	.C(w1_29_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25438 (.Y(n396),
	.A1(n26282),
	.A2(n24126),
	.B(n17396),
	.C(n17395));
   NOR2xp33_ASAP7_75t_SRAM U25439 (.Y(n17397),
	.A(n16430),
	.B(n17398));
   NOR2xp33_ASAP7_75t_SRAM U25440 (.Y(n17399),
	.A(FE_OFN29164_sa33_2),
	.B(FE_OCPN27555_n16422));
   NOR2xp33_ASAP7_75t_SRAM U25441 (.Y(n17401),
	.A(n17399),
	.B(n17398));
   NOR3xp33_ASAP7_75t_SRAM U25442 (.Y(n17406),
	.A(n18430),
	.B(n17405),
	.C(n18433));
   NOR3xp33_ASAP7_75t_R U25443 (.Y(n17409),
	.A(n18144),
	.B(n17407),
	.C(n23539));
   NAND3xp33_ASAP7_75t_SRAM U25444 (.Y(n17413),
	.A(n23533),
	.B(n18405),
	.C(n17412));
   OAI21xp5_ASAP7_75t_L U25445 (.Y(n17419),
	.A1(FE_OCPN27666_n17418),
	.A2(FE_OCPN27604_n16421),
	.B(n17417));
   NOR2x1_ASAP7_75t_L U25446 (.Y(n26120),
	.A(n24617),
	.B(n17419));
   OAI222xp33_ASAP7_75t_SL U25447 (.Y(n17428),
	.A1(FE_OFN29164_sa33_2),
	.A2(n24613),
	.B1(FE_OCPN27555_n16422),
	.B2(n24613),
	.C1(FE_OFN28998_n16923),
	.C2(n24613));
   NAND3xp33_ASAP7_75t_L U25448 (.Y(n17431),
	.A(n17428),
	.B(n23550),
	.C(n23551));
   NAND3xp33_ASAP7_75t_SRAM U25449 (.Y(n17433),
	.A(n23533),
	.B(n17432),
	.C(n18140));
   NOR2xp33_ASAP7_75t_SL U25450 (.Y(n17435),
	.A(n24325),
	.B(n17433));
   NOR2xp33_ASAP7_75t_SRAM U25451 (.Y(n17434),
	.A(n23553),
	.B(n18430));
   OA222x2_ASAP7_75t_SL U25452 (.Y(n17436),
	.A1(n18105),
	.A2(n23548),
	.B1(n17435),
	.B2(n23548),
	.C1(n17434),
	.C2(n23548));
   NOR2x1_ASAP7_75t_SL U25453 (.Y(n17441),
	.A(n17440),
	.B(n17439));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25454 (.Y(n17442),
	.A1(n26770),
	.A2(n24309),
	.B(n24310),
	.C(w0_1_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25455 (.Y(n378),
	.A1(n26770),
	.A2(n24309),
	.B(n17443),
	.C(n17442));
   NOR2x1_ASAP7_75t_SL U25456 (.Y(n21341),
	.A(n19170),
	.B(FE_OCPN29504_sa11_4));
   NOR2x1_ASAP7_75t_L U25457 (.Y(n19223),
	.A(FE_OCPN27242_sa11_1),
	.B(FE_OFN28507_sa11_0));
   NAND2xp5_ASAP7_75t_SL U25459 (.Y(n17501),
	.A(FE_OCPN27242_sa11_1),
	.B(FE_OFN28507_sa11_0));
   NAND3xp33_ASAP7_75t_SRAM U25460 (.Y(n17450),
	.A(FE_OCPN27848_n23255),
	.B(n23254),
	.C(n22486));
   NAND2x2_ASAP7_75t_SL U25461 (.Y(n17494),
	.A(n19170),
	.B(FE_OCPN27625_sa11_5));
   NAND3xp33_ASAP7_75t_L U25462 (.Y(n17454),
	.A(FE_OFN28507_sa11_0),
	.B(sa11_2_),
	.C(FE_OCPN27242_sa11_1));
   NOR2x1_ASAP7_75t_SL U25464 (.Y(n19172),
	.A(FE_OCPN27625_sa11_5),
	.B(FE_OCPN27365_sa11_4));
   NAND2x1p5_ASAP7_75t_SL U25465 (.Y(n21819),
	.A(FE_OFN28811_n19170),
	.B(n21815));
   NOR3xp33_ASAP7_75t_SRAM U25466 (.Y(n17461),
	.A(n17450),
	.B(n17449),
	.C(n17469));
   NAND2x1_ASAP7_75t_SL U25467 (.Y(n21814),
	.A(FE_OCPN27512_sa11_2),
	.B(n19223));
   NOR2x1p5_ASAP7_75t_L U25468 (.Y(n19206),
	.A(FE_OCPN27242_sa11_1),
	.B(FE_OFN28508_sa11_0));
   NOR2xp67_ASAP7_75t_SL U25469 (.Y(n23252),
	.A(FE_OFN28507_sa11_0),
	.B(FE_OCPN27512_sa11_2));
   NOR3x1_ASAP7_75t_SL U25470 (.Y(n17464),
	.A(FE_OCPN29504_sa11_4),
	.B(n19170),
	.C(FE_OCPN27625_sa11_5));
   NAND2xp5_ASAP7_75t_SL U25471 (.Y(n23266),
	.A(FE_OCPN27625_sa11_5),
	.B(n21341));
   NOR2x1_ASAP7_75t_L U25472 (.Y(n21822),
	.A(FE_OCPN29378_n23266),
	.B(n21374));
   NOR2x1_ASAP7_75t_SL U25473 (.Y(n25786),
	.A(FE_OCPN28006_n17454),
	.B(FE_OCPN27601_n17475));
   OAI22xp33_ASAP7_75t_SRAM U25474 (.Y(n23260),
	.A1(FE_OCPN27730_n17464),
	.A2(n25786),
	.B1(FE_OFN29061_n22505),
	.B2(n25786));
   NOR3xp33_ASAP7_75t_SRAM U25475 (.Y(n17460),
	.A(n17455),
	.B(n21822),
	.C(n17493));
   NAND2x1p5_ASAP7_75t_SL U25476 (.Y(n17510),
	.A(n19172),
	.B(FE_OFN26554_n19170));
   NAND2x1p5_ASAP7_75t_SL U25478 (.Y(n22487),
	.A(n21366),
	.B(n17445));
   NAND2x1_ASAP7_75t_L U25479 (.Y(n21393),
	.A(n17473),
	.B(n23247));
   NOR3x1_ASAP7_75t_SL U25480 (.Y(n21860),
	.A(n17494),
	.B(FE_OFN28874_FE_OCPN27551_sa11_4),
	.C(FE_OCPN28006_n17454));
   NOR2x1p5_ASAP7_75t_SL U25481 (.Y(n26071),
	.A(FE_OCPN27584_n22497),
	.B(n17457));
   NAND3xp33_ASAP7_75t_SRAM U25483 (.Y(n17458),
	.A(FE_OFN28874_FE_OCPN27551_sa11_4),
	.B(FE_OCPN27414_n23359),
	.C(FE_PSN8325_FE_OFN28811_n19170));
   NOR2x1_ASAP7_75t_L U25485 (.Y(n21817),
	.A(FE_OFN28996_n17464),
	.B(FE_OCPN28006_n17454));
   NOR2xp33_ASAP7_75t_SL U25486 (.Y(n21859),
	.A(n21817),
	.B(n21372));
   NOR2x1p5_ASAP7_75t_SL U25487 (.Y(n21365),
	.A(FE_OCPN27228_sa11_2),
	.B(n21818));
   NOR2xp33_ASAP7_75t_SRAM U25488 (.Y(n17465),
	.A(FE_OCPN27228_sa11_2),
	.B(FE_OFN138_sa11_0));
   NAND2xp5_ASAP7_75t_SL U25489 (.Y(n23392),
	.A(FE_OCPN27242_sa11_1),
	.B(n23252));
   NOR2x1p5_ASAP7_75t_L U25490 (.Y(n21358),
	.A(FE_OCPN27601_n17475),
	.B(FE_OCPN28447_n23392));
   NAND2xp5_ASAP7_75t_SL U25491 (.Y(n17468),
	.A(FE_PSN8325_FE_OFN28811_n19170),
	.B(n21821));
   NAND2xp33_ASAP7_75t_SL U25492 (.Y(n21841),
	.A(n19162),
	.B(FE_OCPN29513_n17447));
   NAND3xp33_ASAP7_75t_L U25493 (.Y(n17474),
	.A(n21841),
	.B(n23254),
	.C(n26064));
   NOR2x1_ASAP7_75t_SL U25494 (.Y(n23375),
	.A(FE_OCPN27313_n21845),
	.B(n21814));
   NAND3x2_ASAP7_75t_SL U25495 (.Y(n23380),
	.A(FE_OCPN27866_n),
	.B(FE_OCPN28038_n23252),
	.C(n21366));
   NAND3xp33_ASAP7_75t_L U25496 (.Y(n17476),
	.A(n23372),
	.B(n23380),
	.C(n19176));
   NOR2x1_ASAP7_75t_SL U25497 (.Y(n22512),
	.A(FE_OCPN27601_n17475),
	.B(n21814));
   NOR2xp33_ASAP7_75t_SRAM U25499 (.Y(n17484),
	.A(n17444),
	.B(n21817));
   A2O1A1Ixp33_ASAP7_75t_SL U25500 (.Y(n17483),
	.A1(FE_OCPN27730_n17464),
	.A2(FE_OCPN28038_n23252),
	.B(n22500),
	.C(FE_OCPN27866_n));
   NAND2x1_ASAP7_75t_SL U25501 (.Y(n19229),
	.A(n23372),
	.B(n23380));
   NOR2xp33_ASAP7_75t_R U25502 (.Y(n17486),
	.A(FE_OFN29034_FE_OCPN27414_n23359),
	.B(n21817));
   A2O1A1Ixp33_ASAP7_75t_R U25503 (.Y(n21413),
	.A1(FE_OCPN27730_n17464),
	.A2(FE_OCPN27903_n19223),
	.B(n21406),
	.C(n17473));
   NOR2x1_ASAP7_75t_SL U25504 (.Y(n23374),
	.A(n21819),
	.B(n19166));
   NOR2xp33_ASAP7_75t_SRAM U25505 (.Y(n17491),
	.A(n21358),
	.B(n23374));
   NAND3xp33_ASAP7_75t_R U25506 (.Y(n17492),
	.A(n21413),
	.B(n17491),
	.C(n17490));
   NOR3x1_ASAP7_75t_L U25507 (.Y(n19192),
	.A(n21814),
	.B(FE_OFN28874_FE_OCPN27551_sa11_4),
	.C(n17494));
   NOR2x1p5_ASAP7_75t_SL U25508 (.Y(n21349),
	.A(FE_OFN29169_n17510),
	.B(FE_OCPN27592_n17501));
   NAND3xp33_ASAP7_75t_SL U25509 (.Y(n17504),
	.A(n17502),
	.B(n23284),
	.C(n21850));
   A2O1A1Ixp33_ASAP7_75t_SL U25510 (.Y(n17507),
	.A1(FE_OCPN28006_n17454),
	.A2(FE_OCPN28447_n23392),
	.B(FE_OCPN27757_n21819),
	.C(n23372));
   A2O1A1Ixp33_ASAP7_75t_L U25511 (.Y(n17513),
	.A1(FE_OCPN27313_n21845),
	.A2(FE_OCPN27757_n21819),
	.B(n21374),
	.C(n26065));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25512 (.Y(n17511),
	.A1(FE_OFN94_sa11_5),
	.A2(n19171),
	.B(n21854),
	.C(FE_OFN26554_n19170));
   NOR3xp33_ASAP7_75t_SL U25513 (.Y(n24627),
	.A(n17518),
	.B(n17517),
	.C(n17516));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25514 (.Y(n17519),
	.A1(n26082),
	.A2(n24633),
	.B(n24630),
	.C(w0_18_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25515 (.Y(n349),
	.A1(n26082),
	.A2(n24633),
	.B(n17520),
	.C(n17519));
   NAND2x1p5_ASAP7_75t_SL U25517 (.Y(n17592),
	.A(FE_OFN27148_sa32_3),
	.B(FE_OFN69_sa32_4));
   NOR2x1p5_ASAP7_75t_L U25518 (.Y(n22392),
	.A(FE_OCPN29459_n),
	.B(n17592));
   NOR2x1_ASAP7_75t_L U25520 (.Y(n24868),
	.A(n18836),
	.B(FE_OCPN27420_n18794));
   NOR2x1p5_ASAP7_75t_SL U25521 (.Y(n19911),
	.A(FE_OFN28696_sa32_4),
	.B(FE_OCPN27499_FE_OFN16151_sa32_5));
   NOR2x1p5_ASAP7_75t_SL U25522 (.Y(n19940),
	.A(FE_OFN28892_n),
	.B(n18793));
   NOR2xp33_ASAP7_75t_L U25523 (.Y(n17522),
	.A(n17564),
	.B(n18793));
   NOR3xp33_ASAP7_75t_SL U25524 (.Y(n24644),
	.A(FE_OCPN27499_FE_OFN16151_sa32_5),
	.B(FE_OFN27148_sa32_3),
	.C(FE_OFN28696_sa32_4));
   NAND2x1p5_ASAP7_75t_SL U25525 (.Y(n18837),
	.A(FE_OFN28696_sa32_4),
	.B(FE_OCPN27499_FE_OFN16151_sa32_5));
   NOR2xp33_ASAP7_75t_SRAM U25526 (.Y(n17528),
	.A(n17560),
	.B(n18846));
   NOR2x1_ASAP7_75t_L U25527 (.Y(n17563),
	.A(FE_OFN16463_sa32_0),
	.B(FE_OCPN29304_n17526));
   NAND2x1_ASAP7_75t_SL U25528 (.Y(n18829),
	.A(FE_OFN28892_n),
	.B(n17563));
   NOR2xp33_ASAP7_75t_R U25529 (.Y(n17531),
	.A(FE_OCPN28229_n17529),
	.B(n18846));
   NOR3x2_ASAP7_75t_SL U25530 (.Y(n19938),
	.A(FE_OFN26035_n),
	.B(FE_OFN28892_n),
	.C(FE_OFN16463_sa32_0));
   NAND2x2_ASAP7_75t_SL U25531 (.Y(n18828),
	.A(FE_OFN28696_sa32_4),
	.B(n19725));
   AND3x1_ASAP7_75t_SL U25532 (.Y(n17537),
	.A(n17723),
	.B(n17535),
	.C(n17703));
   NOR2xp33_ASAP7_75t_SRAM U25533 (.Y(n17538),
	.A(FE_OCPN28229_n17529),
	.B(n24868));
   NOR2x1p5_ASAP7_75t_SL U25534 (.Y(n20096),
	.A(FE_OCPN27882_n18829),
	.B(n17542));
   NAND2xp5_ASAP7_75t_SL U25535 (.Y(n25028),
	.A(FE_OFN27148_sa32_3),
	.B(n19911));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25536 (.Y(n17543),
	.A1(n17521),
	.A2(n17560),
	.B(n19926),
	.C(FE_OFN28893_n));
   NOR2x1p5_ASAP7_75t_SL U25537 (.Y(n19921),
	.A(FE_OCPN29298_n25028),
	.B(FE_OCPN27882_n18829));
   NOR2x1_ASAP7_75t_L U25538 (.Y(n17551),
	.A(n17693),
	.B(n19921));
   NAND3xp33_ASAP7_75t_SRAM U25539 (.Y(n17547),
	.A(n17521),
	.B(n17525),
	.C(FE_OFN28893_n));
   NOR2xp33_ASAP7_75t_SRAM U25540 (.Y(n17548),
	.A(FE_OFN28893_n),
	.B(n17521));
   NAND3x1_ASAP7_75t_SL U25541 (.Y(n17552),
	.A(n18338),
	.B(n18321),
	.C(n17551));
   NOR2x1_ASAP7_75t_SL U25542 (.Y(n23900),
	.A(n19954),
	.B(n17552));
   NAND3x1_ASAP7_75t_SL U25543 (.Y(n20094),
	.A(FE_OCPN29449_n17521),
	.B(n22392),
	.C(FE_OFN28893_n));
   NOR2x1p5_ASAP7_75t_SL U25544 (.Y(n20107),
	.A(FE_OFN26577_n),
	.B(n18828));
   NAND3xp33_ASAP7_75t_SL U25545 (.Y(n17554),
	.A(n20111),
	.B(n18839),
	.C(n20098));
   NOR2xp33_ASAP7_75t_L U25546 (.Y(n20104),
	.A(n18836),
	.B(n18818));
   NOR2xp33_ASAP7_75t_SRAM U25547 (.Y(n17570),
	.A(n22399),
	.B(n19908));
   A2O1A1Ixp33_ASAP7_75t_SL U25548 (.Y(n18819),
	.A1(n17521),
	.A2(FE_OFN28893_n),
	.B(n17675),
	.C(n17525));
   NAND3xp33_ASAP7_75t_SRAM U25549 (.Y(n17568),
	.A(n18839),
	.B(n19951),
	.C(n18819));
   NOR3xp33_ASAP7_75t_L U25550 (.Y(n17569),
	.A(n17568),
	.B(FE_OCPN27490_n18798),
	.C(n17567));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25551 (.Y(n17577),
	.A1(FE_OCPN29449_n17521),
	.A2(n17560),
	.B(n19921),
	.C(FE_OCPN29421_FE_OFN16128_sa32_2));
   NOR2xp33_ASAP7_75t_L U25552 (.Y(n17576),
	.A(n17572),
	.B(n17571));
   NAND2xp5_ASAP7_75t_SL U25553 (.Y(n24864),
	.A(n17578),
	.B(n22390));
   NAND3xp33_ASAP7_75t_L U25554 (.Y(n17583),
	.A(n17581),
	.B(n24872),
	.C(n17708));
   NAND3xp33_ASAP7_75t_SL U25555 (.Y(n17590),
	.A(n18336),
	.B(n22397),
	.C(n20094));
   NOR2x1_ASAP7_75t_SL U25556 (.Y(n19922),
	.A(FE_OCPN27937_n18841),
	.B(n17590));
   NOR3xp33_ASAP7_75t_SRAM U25557 (.Y(n17594),
	.A(n22366),
	.B(n19732),
	.C(n19698));
   NAND3xp33_ASAP7_75t_L U25558 (.Y(n17595),
	.A(n19922),
	.B(n17594),
	.C(n18820));
   O2A1O1Ixp5_ASAP7_75t_SL U25559 (.Y(n23902),
	.A1(n19723),
	.A2(n17598),
	.B(n17580),
	.C(n17597));
   A2O1A1Ixp33_ASAP7_75t_SL U25560 (.Y(n24996),
	.A1(n23900),
	.A2(n23898),
	.B(n23899),
	.C(n23902));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25561 (.Y(n17599),
	.A1(n22405),
	.A2(n24289),
	.B(n24996),
	.C(FE_OFN16423_n24831));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25562 (.Y(n413),
	.A1(n22405),
	.A2(n24289),
	.B(n17600),
	.C(n17599));
   NOR2x1p5_ASAP7_75t_SL U25563 (.Y(n25108),
	.A(n17618),
	.B(n18364));
   NOR2x1p5_ASAP7_75t_SL U25565 (.Y(n17630),
	.A(FE_OFN28901_sa30_4),
	.B(FE_OCPN29412_sa30_5));
   NAND2x1p5_ASAP7_75t_SL U25566 (.Y(n18473),
	.A(FE_OCPN29399_sa30_3),
	.B(n17630));
   NAND2x1p5_ASAP7_75t_SL U25567 (.Y(n19051),
	.A(n17601),
	.B(FE_OFN16247_sa30_1));
   NAND2x1p5_ASAP7_75t_SL U25568 (.Y(n20429),
	.A(FE_OFN28895_sa30_2),
	.B(n17603));
   NOR2x1_ASAP7_75t_SL U25569 (.Y(n17646),
	.A(FE_OFN26597_n),
	.B(FE_OCPN28049_sa30_0));
   NAND2x1p5_ASAP7_75t_SL U25570 (.Y(n21625),
	.A(FE_OCPN29368_FE_OFN16247_sa30_1),
	.B(n17646));
   NOR2x1_ASAP7_75t_SL U25572 (.Y(n19037),
	.A(n20471),
	.B(n18473));
   NOR3x1_ASAP7_75t_SL U25573 (.Y(n21591),
	.A(n17618),
	.B(FE_OCPN29431_sa30_3),
	.C(FE_OFN28901_sa30_4));
   OAI21xp33_ASAP7_75t_SL U25574 (.Y(n18393),
	.A1(n18381),
	.A2(n21625),
	.B(n20449));
   NAND2x1p5_ASAP7_75t_SL U25575 (.Y(n20428),
	.A(FE_OFN28901_sa30_4),
	.B(n22632));
   NAND3xp33_ASAP7_75t_SL U25576 (.Y(n22133),
	.A(FE_OCPN28049_sa30_0),
	.B(FE_OFN16247_sa30_1),
	.C(FE_OFN26597_n));
   NOR2xp33_ASAP7_75t_L U25579 (.Y(n18453),
	.A(n21608),
	.B(n22159));
   NAND3x1_ASAP7_75t_SL U25580 (.Y(n26027),
	.A(FE_OFN28901_sa30_4),
	.B(n17618),
	.C(FE_OCPN29431_sa30_3));
   NAND2x1p5_ASAP7_75t_L U25581 (.Y(n21627),
	.A(FE_OFN28901_sa30_4),
	.B(n17618));
   NAND2x1_ASAP7_75t_L U25582 (.Y(n18503),
	.A(n17618),
	.B(FE_OFN16333_sa30_4));
   NOR2x1p5_ASAP7_75t_SL U25583 (.Y(n22613),
	.A(n20428),
	.B(FE_OFN29121_n26026));
   NOR3x1_ASAP7_75t_SL U25584 (.Y(n21603),
	.A(n17605),
	.B(n26023),
	.C(n22613));
   NAND3xp33_ASAP7_75t_SRAM U25585 (.Y(n17614),
	.A(n18453),
	.B(n20478),
	.C(n21603));
   NOR3x1_ASAP7_75t_SL U25586 (.Y(n22125),
	.A(FE_OFN16247_sa30_1),
	.B(FE_OFN26597_n),
	.C(FE_OCPN28049_sa30_0));
   NOR2x1p5_ASAP7_75t_SL U25587 (.Y(n24780),
	.A(FE_OFN28895_sa30_2),
	.B(n18352));
   NAND2x1_ASAP7_75t_L U25588 (.Y(n22621),
	.A(n24780),
	.B(n25108));
   NOR2x1_ASAP7_75t_L U25589 (.Y(n22168),
	.A(FE_OCPN27829_n25102),
	.B(n21626));
   NOR2xp33_ASAP7_75t_SRAM U25590 (.Y(n17613),
	.A(n22168),
	.B(n22169));
   NOR2x1_ASAP7_75t_SL U25591 (.Y(n24791),
	.A(n20429),
	.B(FE_PSN8270_n26027));
   A2O1A1Ixp33_ASAP7_75t_R U25592 (.Y(n17608),
	.A1(FE_OCPN28378_n22632),
	.A2(FE_OFN28610_n22125),
	.B(n24791),
	.C(n18463));
   NOR2x1_ASAP7_75t_L U25593 (.Y(n21607),
	.A(FE_OCPN29413_sa30_5),
	.B(n18381));
   NOR2x1_ASAP7_75t_SL U25594 (.Y(n18365),
	.A(n20428),
	.B(FE_OCPN27829_n25102));
   OAI22xp33_ASAP7_75t_L U25595 (.Y(n18488),
	.A1(FE_OFN29094_n21607),
	.A2(n18365),
	.B1(n17602),
	.B2(n18365));
   NAND3xp33_ASAP7_75t_L U25596 (.Y(n17612),
	.A(n17608),
	.B(n18488),
	.C(n22145));
   A2O1A1Ixp33_ASAP7_75t_SL U25597 (.Y(n24787),
	.A1(n24780),
	.A2(n22632),
	.B(n18368),
	.C(FE_OFN28901_sa30_4));
   NOR2xp33_ASAP7_75t_SL U25598 (.Y(n17610),
	.A(FE_OCPN27764_n22152),
	.B(n17609));
   NOR2x1p5_ASAP7_75t_SL U25599 (.Y(n18497),
	.A(FE_OCPN29400_sa30_3),
	.B(n18503));
   NOR2xp33_ASAP7_75t_SRAM U25600 (.Y(n17615),
	.A(n25082),
	.B(n18506));
   NOR2x1_ASAP7_75t_SL U25601 (.Y(n24785),
	.A(n22629),
	.B(n18365));
   NAND3xp33_ASAP7_75t_SRAM U25602 (.Y(n17628),
	.A(n24137),
	.B(n17615),
	.C(n24785));
   NAND2xp5_ASAP7_75t_SL U25603 (.Y(n18501),
	.A(FE_OFN28818_n17602),
	.B(FE_OFN29094_n21607));
   NOR2x1_ASAP7_75t_SL U25604 (.Y(n21619),
	.A(n21604),
	.B(FE_OFN29121_n26026));
   NAND2xp5_ASAP7_75t_SL U25605 (.Y(n19049),
	.A(n24780),
	.B(n17630));
   NOR2x1p5_ASAP7_75t_L U25606 (.Y(n18458),
	.A(FE_OCPN29399_sa30_3),
	.B(n19049));
   NAND2xp5_ASAP7_75t_L U25607 (.Y(n17627),
	.A(n17626),
	.B(n17625));
   NAND3xp33_ASAP7_75t_SL U25608 (.Y(n20437),
	.A(n18489),
	.B(n22151),
	.C(n17627));
   NOR3xp33_ASAP7_75t_SRAM U25609 (.Y(n17672),
	.A(n17628),
	.B(n24128),
	.C(FE_OFN28619_n20437));
   NOR2x1_ASAP7_75t_SL U25610 (.Y(n18455),
	.A(n22161),
	.B(n22152));
   NOR2xp33_ASAP7_75t_SRAM U25611 (.Y(n17631),
	.A(n17630),
	.B(n22613));
   NOR2xp33_ASAP7_75t_SRAM U25612 (.Y(n17633),
	.A(FE_OFN28637_n25102),
	.B(n22613));
   NOR2xp33_ASAP7_75t_R U25613 (.Y(n17640),
	.A(n22629),
	.B(n18368));
   OAI21xp33_ASAP7_75t_L U25614 (.Y(n17638),
	.A1(n20429),
	.A2(FE_PSN8272_n20428),
	.B(n19047));
   NOR3xp33_ASAP7_75t_SL U25615 (.Y(n17642),
	.A(n17641),
	.B(n25082),
	.C(n25118));
   A2O1A1Ixp33_ASAP7_75t_L U25616 (.Y(n18496),
	.A1(FE_OCPN8207_n18497),
	.A2(FE_OCPN7643_n17646),
	.B(n17645),
	.C(FE_OCPN29368_FE_OFN16247_sa30_1));
   A2O1A1Ixp33_ASAP7_75t_R U25617 (.Y(n17658),
	.A1(n20471),
	.A2(FE_OCPN27829_n25102),
	.B(FE_PSN8272_n20428),
	.C(n17653));
   NOR2x1_ASAP7_75t_L U25618 (.Y(n21613),
	.A(n22169),
	.B(FE_OCPN29289_n22162));
   NAND2xp5_ASAP7_75t_L U25619 (.Y(n17654),
	.A(n22130),
	.B(n20427));
   NOR2x1_ASAP7_75t_L U25620 (.Y(n22155),
	.A(n21619),
	.B(n17654));
   NAND3xp33_ASAP7_75t_SL U25621 (.Y(n20460),
	.A(n17655),
	.B(n22132),
	.C(n22155));
   NOR2xp33_ASAP7_75t_R U25622 (.Y(n17656),
	.A(n20471),
	.B(n18503));
   NOR3x1_ASAP7_75t_L U25623 (.Y(n22624),
	.A(n21625),
	.B(FE_OCPN29400_sa30_3),
	.C(FE_OCPN8240_n17618));
   NOR2xp33_ASAP7_75t_SL U25624 (.Y(n17660),
	.A(n22624),
	.B(n24791));
   NOR2xp33_ASAP7_75t_R U25625 (.Y(n17664),
	.A(FE_OFN25917_n21591),
	.B(n26023));
   NOR2xp33_ASAP7_75t_SRAM U25626 (.Y(n17666),
	.A(FE_OCPN28057_n17603),
	.B(n26023));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25627 (.Y(n17673),
	.A1(FE_OFN16164_n25081),
	.A2(n25080),
	.B(n25077),
	.C(FE_OFN58_w1_4));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25628 (.Y(n309),
	.A1(FE_OFN16164_n25081),
	.A2(n25080),
	.B(n17674),
	.C(n17673));
   NAND2x1_ASAP7_75t_SL U25629 (.Y(n24648),
	.A(n17684),
	.B(n17683));
   NOR2xp33_ASAP7_75t_SL U25630 (.Y(n17685),
	.A(n20106),
	.B(n17716));
   AND2x2_ASAP7_75t_SRAM U25631 (.Y(n17686),
	.A(n24645),
	.B(n24646));
   OAI21xp5_ASAP7_75t_L U25632 (.Y(n17689),
	.A1(FE_OCPN29298_n25028),
	.A2(FE_OCPN29323_n19721),
	.B(n22377));
   NAND2xp33_ASAP7_75t_SRAM U25633 (.Y(n17699),
	.A(n19934),
	.B(n24853));
   NOR2x1_ASAP7_75t_L U25634 (.Y(n20108),
	.A(FE_OFN16232_n17691),
	.B(n19908));
   NAND3xp33_ASAP7_75t_SL U25635 (.Y(n17694),
	.A(n18302),
	.B(n20108),
	.C(n25022));
   OAI21xp33_ASAP7_75t_SRAM U25637 (.Y(n17701),
	.A1(n18827),
	.A2(n18837),
	.B(n18330));
   NOR2xp33_ASAP7_75t_SRAM U25638 (.Y(n24863),
	.A(FE_OCPN28245_n),
	.B(n17700));
   NOR3xp33_ASAP7_75t_SRAM U25639 (.Y(n17730),
	.A(n17701),
	.B(n24863),
	.C(n17722));
   OAI222xp33_ASAP7_75t_SRAM U25640 (.Y(n17720),
	.A1(n17731),
	.A2(n17584),
	.B1(n17702),
	.B2(n17584),
	.C1(n17730),
	.C2(n17584));
   NAND3xp33_ASAP7_75t_SRAM U25641 (.Y(n17709),
	.A(FE_OFN16231_n17691),
	.B(n18336),
	.C(n17703));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25642 (.Y(n17706),
	.A1(FE_OFN26035_n),
	.A2(n18847),
	.B(FE_OCPN27792_n18333),
	.C(FE_OFN16463_sa32_0));
   NOR3xp33_ASAP7_75t_L U25643 (.Y(n17705),
	.A(n17722),
	.B(n20104),
	.C(n18846));
   NOR2xp33_ASAP7_75t_SRAM U25644 (.Y(n17707),
	.A(n19703),
	.B(n19704));
   NAND3xp33_ASAP7_75t_R U25645 (.Y(n17726),
	.A(n18839),
	.B(n17712),
	.C(n17711));
   NOR2xp33_ASAP7_75t_SRAM U25646 (.Y(n17718),
	.A(n17726),
	.B(n17727));
   OAI22xp33_ASAP7_75t_SRAM U25647 (.Y(n17715),
	.A1(FE_OCPN27267_n18794),
	.A2(FE_OFN26577_n),
	.B1(n18828),
	.B2(FE_OFN26577_n));
   NOR3xp33_ASAP7_75t_SRAM U25648 (.Y(n17717),
	.A(n17722),
	.B(FE_OFN28633_n17716),
	.C(n17715));
   NOR3xp33_ASAP7_75t_SRAM U25649 (.Y(n17721),
	.A(n17720),
	.B(n17733),
	.C(n17719));
   NAND2xp33_ASAP7_75t_R U25650 (.Y(n17738),
	.A(n17721),
	.B(n24913));
   NOR3xp33_ASAP7_75t_SRAM U25651 (.Y(n17724),
	.A(n17722),
	.B(n20107),
	.C(n20106));
   NAND3xp33_ASAP7_75t_SRAM U25652 (.Y(n17725),
	.A(n17724),
	.B(n20094),
	.C(n17723));
   AND3x1_ASAP7_75t_SRAM U25653 (.Y(n17729),
	.A(n19934),
	.B(n24853),
	.C(n17728));
   NAND3xp33_ASAP7_75t_L U25654 (.Y(n17734),
	.A(n17731),
	.B(n17730),
	.C(n17729));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25655 (.Y(n17737),
	.A1(n22405),
	.A2(FE_OFN26030_n25368),
	.B(FE_OCPN28100_n25470),
	.C(FE_OFN26531_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25656 (.Y(n282),
	.A1(n22405),
	.A2(FE_OFN26030_n25368),
	.B(n17738),
	.C(n17737));
   NOR2x1_ASAP7_75t_L U25657 (.Y(n20169),
	.A(FE_OCPN27261_sa02_0),
	.B(FE_OCPN27585_sa02_1));
   NOR2x1_ASAP7_75t_L U25658 (.Y(n22089),
	.A(n17763),
	.B(n17740));
   NAND2x1p5_ASAP7_75t_L U25659 (.Y(n22076),
	.A(FE_OCPN27634_n20169),
	.B(n22089));
   NOR2x1p5_ASAP7_75t_SL U25660 (.Y(n17799),
	.A(FE_OFN16234_sa02_2),
	.B(FE_OCPN27572_sa02_1));
   NAND2xp5_ASAP7_75t_SL U25662 (.Y(n20155),
	.A(FE_OFN16234_sa02_2),
	.B(n20169));
   NAND2x1p5_ASAP7_75t_SL U25663 (.Y(n20196),
	.A(n17763),
	.B(n22543));
   NOR2x1_ASAP7_75t_SL U25665 (.Y(n25531),
	.A(FE_OCPN27573_n20196),
	.B(FE_OCPN29545_n22529));
   NOR2xp67_ASAP7_75t_L U25666 (.Y(n17742),
	.A(n17763),
	.B(FE_OCPN8269_FE_OFN16136_sa02_5));
   NOR3xp33_ASAP7_75t_SRAM U25667 (.Y(n17743),
	.A(n25525),
	.B(n25531),
	.C(n25530));
   NAND3xp33_ASAP7_75t_SRAM U25668 (.Y(n17745),
	.A(n22076),
	.B(n22075),
	.C(n17743));
   NOR2x1_ASAP7_75t_L U25669 (.Y(n22882),
	.A(FE_OFN16234_sa02_2),
	.B(sa02_1_));
   NOR3xp33_ASAP7_75t_SRAM U25670 (.Y(n17767),
	.A(n17745),
	.B(FE_OCPN29318_n25524),
	.C(n25523));
   NAND2x1_ASAP7_75t_SL U25671 (.Y(n22527),
	.A(FE_OCPN27261_sa02_0),
	.B(FE_OCPN27572_sa02_1));
   NOR2x1p5_ASAP7_75t_SL U25672 (.Y(n22094),
	.A(FE_OCPN29436_n22080),
	.B(n22527));
   NOR2x1_ASAP7_75t_SL U25674 (.Y(n20161),
	.A(FE_OFN27058_n22094),
	.B(n22526));
   NAND3xp33_ASAP7_75t_R U25675 (.Y(n25529),
	.A(n19257),
	.B(n20127),
	.C(FE_OCPN27689_n20172));
   NOR2xp33_ASAP7_75t_SL U25676 (.Y(n17751),
	.A(FE_OFN25998_n17781),
	.B(n17798));
   NOR2x1_ASAP7_75t_SL U25677 (.Y(n20988),
	.A(n20195),
	.B(n22529));
   INVxp67_ASAP7_75t_SL U25678 (.Y(n17749),
	.A(n17748));
   NOR2xp33_ASAP7_75t_SL U25680 (.Y(n17753),
	.A(FE_OFN108_n26971),
	.B(n17798));
   NAND2x1p5_ASAP7_75t_SL U25681 (.Y(n20962),
	.A(n17760),
	.B(n17761));
   NOR2x1_ASAP7_75t_L U25682 (.Y(n22086),
	.A(n20176),
	.B(n22881));
   OAI21xp33_ASAP7_75t_R U25683 (.Y(n17762),
	.A1(FE_OCPN27574_n20196),
	.A2(FE_OFN27058_n22094),
	.B(n22086));
   NAND3x1_ASAP7_75t_SL U25684 (.Y(n25536),
	.A(n20997),
	.B(n17764),
	.C(n22557));
   NOR3xp33_ASAP7_75t_SRAM U25685 (.Y(n17766),
	.A(n25529),
	.B(n25528),
	.C(n25536));
   NAND3xp33_ASAP7_75t_SL U25686 (.Y(n22070),
	.A(FE_OCPN27570_n17791),
	.B(FE_PSN8323_n22543),
	.C(FE_OFN28730_FE_OCPN28416_sa02_3));
   NOR2xp33_ASAP7_75t_SL U25687 (.Y(n25526),
	.A(n22095),
	.B(n25212));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25688 (.Y(n17769),
	.A1(n17763),
	.A2(FE_OFN28665_FE_OCPN27566),
	.B(n17760),
	.C(n17768));
   NAND3xp33_ASAP7_75t_SL U25689 (.Y(n17773),
	.A(n17770),
	.B(n17769),
	.C(n22074));
   NOR3x1_ASAP7_75t_L U25690 (.Y(n20982),
	.A(FE_OFN29148_n),
	.B(FE_OFN28665_FE_OCPN27566),
	.C(n17771));
   OAI21xp5_ASAP7_75t_L U25691 (.Y(n20206),
	.A1(n22529),
	.A2(n20962),
	.B(n22902));
   NOR2x1p5_ASAP7_75t_L U25692 (.Y(n20995),
	.A(FE_OFN27058_n22094),
	.B(FE_OFN29144_n17747));
   NOR2x1_ASAP7_75t_SL U25693 (.Y(n19274),
	.A(n20981),
	.B(n20995));
   NOR2x1p5_ASAP7_75t_R U25694 (.Y(n22540),
	.A(FE_OFN28961_n17744),
	.B(FE_OCPN27573_n20196));
   NOR2x1p5_ASAP7_75t_SL U25695 (.Y(n22085),
	.A(n25297),
	.B(n22540));
   NOR2x1p5_ASAP7_75t_SL U25696 (.Y(n20978),
	.A(FE_OCPN27573_n20196),
	.B(FE_OFN27058_n22094));
   NAND3x1_ASAP7_75t_SL U25697 (.Y(n26968),
	.A(n22085),
	.B(n17776),
	.C(n22877));
   NAND3xp33_ASAP7_75t_L U25698 (.Y(n17777),
	.A(n17807),
	.B(n17775),
	.C(n22105));
   NOR2x1_ASAP7_75t_L U25699 (.Y(n20186),
	.A(FE_OFN29184_n17744),
	.B(FE_OCPN27624_n26971));
   OAI22xp33_ASAP7_75t_SL U25700 (.Y(n22890),
	.A1(FE_OCPN29469_n17747),
	.A2(n25531),
	.B1(FE_OFN28844_FE_OCPN27570_n17791),
	.B2(n25531));
   NOR2xp33_ASAP7_75t_SRAM U25701 (.Y(n17787),
	.A(n20161),
	.B(n25523));
   OAI21xp5_ASAP7_75t_SL U25702 (.Y(n20994),
	.A1(FE_OFN28665_FE_OCPN27566),
	.A2(n20153),
	.B(n22062));
   NAND3xp33_ASAP7_75t_R U25703 (.Y(n17783),
	.A(n20137),
	.B(FE_OCPN28303_n20961),
	.C(FE_OFN97_n20994));
   NAND3xp33_ASAP7_75t_SL U25704 (.Y(n22532),
	.A(n20190),
	.B(n17782),
	.C(n25213));
   O2A1O1Ixp33_ASAP7_75t_SRAM U25705 (.Y(n17784),
	.A1(FE_OFN28812_FE_OCPN27261_sa02_0),
	.A2(FE_OCPN29341_FE_OFN29148_n),
	.B(n22083),
	.C(n20195));
   NAND3xp33_ASAP7_75t_R U25706 (.Y(n17819),
	.A(n17787),
	.B(n17786),
	.C(n17785));
   NAND3xp33_ASAP7_75t_L U25707 (.Y(n19255),
	.A(FE_PSN8323_n22543),
	.B(FE_OCPN27384_n22888),
	.C(FE_OFN28730_FE_OCPN28416_sa02_3));
   NOR2xp67_ASAP7_75t_SL U25708 (.Y(n20214),
	.A(n25530),
	.B(n22540));
   NOR2xp33_ASAP7_75t_R U25709 (.Y(n17789),
	.A(n20978),
	.B(n20194));
   NOR2x1_ASAP7_75t_SL U25710 (.Y(n20189),
	.A(n17791),
	.B(n17790));
   NOR2xp33_ASAP7_75t_L U25711 (.Y(n17793),
	.A(n20189),
	.B(n20168));
   OR2x2_ASAP7_75t_L U25712 (.Y(n17794),
	.A(FE_OFN28704_FE_OCPN27740_sa02_4),
	.B(n20168));
   NAND3xp33_ASAP7_75t_L U25713 (.Y(n17814),
	.A(n22075),
	.B(n20198),
	.C(n17796));
   NOR2xp33_ASAP7_75t_SRAM U25714 (.Y(n17797),
	.A(n26971),
	.B(n20155));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25715 (.Y(n19280),
	.A1(n17761),
	.A2(FE_OCPN27570_n17791),
	.B(n17797),
	.C(FE_OFN28703_FE_OCPN27740_sa02_4));
   NOR2xp33_ASAP7_75t_SL U25716 (.Y(n20197),
	.A(n20196),
	.B(n20155));
   NOR2xp33_ASAP7_75t_L U25717 (.Y(n17810),
	.A(n17808),
	.B(n20144));
   NAND2xp5_ASAP7_75t_SL U25718 (.Y(n17813),
	.A(n17812),
	.B(n17811));
   NAND3x1_ASAP7_75t_SL U25719 (.Y(n21001),
	.A(n17813),
	.B(n20953),
	.C(n20190));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25720 (.Y(n17822),
	.A1(n27216),
	.A2(n27215),
	.B(n27212),
	.C(w2_26_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25721 (.Y(n314),
	.A1(n27216),
	.A2(n27215),
	.B(n17823),
	.C(n17822));
   NOR2xp33_ASAP7_75t_SRAM U25722 (.Y(n17825),
	.A(FE_OFN27157_n23928),
	.B(FE_OCPN29279_n25353));
   INVxp33_ASAP7_75t_SRAM U25723 (.Y(n17824),
	.A(n17872));
   OR2x2_ASAP7_75t_SRAM U25724 (.Y(n17826),
	.A(FE_OCPN28298_n),
	.B(FE_OCPN29279_n25353));
   NOR2xp33_ASAP7_75t_SRAM U25725 (.Y(n17834),
	.A(n16771),
	.B(n22676));
   NOR2xp33_ASAP7_75t_R U25726 (.Y(n17835),
	.A(FE_OFN28529_n16774),
	.B(n22676));
   NAND3xp33_ASAP7_75t_SRAM U25727 (.Y(n17842),
	.A(n17838),
	.B(n23656),
	.C(n19863));
   NOR2xp33_ASAP7_75t_SRAM U25728 (.Y(n17840),
	.A(FE_OCPN27246_n22663),
	.B(FE_OFN27140_n20007));
   NOR3xp33_ASAP7_75t_SRAM U25729 (.Y(n17841),
	.A(n20329),
	.B(n17840),
	.C(n20305));
   NOR3xp33_ASAP7_75t_L U25730 (.Y(n17853),
	.A(FE_OCPN5079_n20287),
	.B(n17844),
	.C(FE_OFN28970_n19890));
   NOR2xp33_ASAP7_75t_R U25731 (.Y(n17846),
	.A(FE_OFN29023_n16750),
	.B(n22675));
   NOR2xp33_ASAP7_75t_SRAM U25732 (.Y(n17848),
	.A(n16771),
	.B(n22675));
   NAND2x1p5_ASAP7_75t_SL U25733 (.Y(n24919),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(FE_OFN28779_n24257));
   NAND3xp33_ASAP7_75t_SL U25734 (.Y(n17858),
	.A(n20312),
	.B(n19884),
	.C(n22715));
   NOR3x1_ASAP7_75t_L U25735 (.Y(n24281),
	.A(n17858),
	.B(n17857),
	.C(n17856));
   NOR2xp33_ASAP7_75t_R U25736 (.Y(n17861),
	.A(FE_OFN28823_n17860),
	.B(n19982));
   AND2x2_ASAP7_75t_L U25737 (.Y(n22697),
	.A(n17863),
	.B(n23626));
   NAND3xp33_ASAP7_75t_L U25738 (.Y(n17870),
	.A(n19972),
	.B(n19889),
	.C(n22333));
   NOR2xp33_ASAP7_75t_R U25739 (.Y(n17875),
	.A(FE_OFN16447_n16749),
	.B(FE_OCPN29321_n17876));
   NOR2xp33_ASAP7_75t_SL U25740 (.Y(n17877),
	.A(FE_OFN28914_n20007),
	.B(FE_OCPN29321_n17876));
   NAND3x1_ASAP7_75t_SL U25741 (.Y(n25589),
	.A(n17880),
	.B(n22669),
	.C(n19901));
   NOR3xp33_ASAP7_75t_R U25742 (.Y(n17882),
	.A(n16762),
	.B(FE_OFN28903_sa21_0),
	.C(n17881));
   NAND3xp33_ASAP7_75t_L U25743 (.Y(n17883),
	.A(n22354),
	.B(n20002),
	.C(n22351));
   NOR2xp33_ASAP7_75t_R U25744 (.Y(n17885),
	.A(n22694),
	.B(n23643));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25745 (.Y(n17895),
	.A1(n26829),
	.A2(n23971),
	.B(FE_OFN29031_n23968),
	.C(w3_10_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25746 (.Y(n420),
	.A1(n26829),
	.A2(n23971),
	.B(n17896),
	.C(n17895));
   NAND2x1p5_ASAP7_75t_L U25747 (.Y(n20554),
	.A(FE_OFN25908_sa12_2),
	.B(n17953));
   NOR2x1p5_ASAP7_75t_SL U25749 (.Y(n20593),
	.A(n19538),
	.B(FE_OFN28676_sa12_5));
   NAND2x1p5_ASAP7_75t_SL U25750 (.Y(n17952),
	.A(n22721),
	.B(FE_OFN28764_n17928));
   NOR2x2_ASAP7_75t_SL U25751 (.Y(n24364),
	.A(FE_OFN28476_sa12_0),
	.B(n17952));
   NAND2x1p5_ASAP7_75t_L U25752 (.Y(n25398),
	.A(FE_OFN28739_n17898),
	.B(n24364));
   NAND2x1_ASAP7_75t_SL U25753 (.Y(n17971),
	.A(FE_OCPN29499_FE_OFN16131_sa12_1),
	.B(FE_OFN29225_sa12_0));
   AND3x1_ASAP7_75t_R U25754 (.Y(n20817),
	.A(n19552),
	.B(n25398),
	.C(n20561));
   NAND3xp33_ASAP7_75t_L U25755 (.Y(n22224),
	.A(n17928),
	.B(FE_OFN29225_sa12_0),
	.C(FE_OCPN27888_sa12_2));
   NOR3xp33_ASAP7_75t_SL U25756 (.Y(n23208),
	.A(FE_OFN26158_n22224),
	.B(FE_OCPN29492_sa12_4),
	.C(FE_OCPN29477_sa12_5));
   NOR2xp33_ASAP7_75t_SRAM U25757 (.Y(n17902),
	.A(n19546),
	.B(n17954));
   NAND2xp5_ASAP7_75t_SL U25758 (.Y(n17923),
	.A(sa12_0_),
	.B(FE_OFN16131_sa12_1));
   NOR3x2_ASAP7_75t_SL U25760 (.Y(n24362),
	.A(FE_OFN73_sa12_5),
	.B(FE_OCPN29493_sa12_4),
	.C(FE_OCPN29486_sa12_3));
   NAND2xp5_ASAP7_75t_SL U25761 (.Y(n20542),
	.A(n19539),
	.B(n24362));
   OR2x2_ASAP7_75t_SRAM U25762 (.Y(n17903),
	.A(n17953),
	.B(n17954));
   NAND2xp5_ASAP7_75t_SL U25763 (.Y(n23216),
	.A(FE_OCPN29492_sa12_4),
	.B(n20593));
   A2O1A1Ixp33_ASAP7_75t_R U25764 (.Y(n20550),
	.A1(n17906),
	.A2(n24364),
	.B(n20583),
	.C(FE_OCPN29485_sa12_3));
   NOR2x1_ASAP7_75t_SL U25765 (.Y(n22742),
	.A(FE_OCPN27368_sa12_3),
	.B(n19509));
   NOR2x1_ASAP7_75t_L U25767 (.Y(n22233),
	.A(FE_OCPN27253_n17923),
	.B(n23217));
   OAI21xp5_ASAP7_75t_SL U25768 (.Y(n22749),
	.A1(n22233),
	.A2(n23206),
	.B(FE_OFN25907_sa12_2));
   NOR2x1_ASAP7_75t_L U25769 (.Y(n20806),
	.A(n19527),
	.B(FE_OCPN29324_n23216));
   NOR2x1_ASAP7_75t_SL U25770 (.Y(n22776),
	.A(FE_OFN28764_n17928),
	.B(FE_OFN28476_sa12_0));
   OAI21xp5_ASAP7_75t_SL U25771 (.Y(n17939),
	.A1(n23217),
	.A2(n19502),
	.B(n22236));
   NAND2xp5_ASAP7_75t_SL U25772 (.Y(n20595),
	.A(FE_OFN29075_n22745),
	.B(n24362));
   OAI222xp33_ASAP7_75t_L U25773 (.Y(n17920),
	.A1(FE_OCPN5137_n23600),
	.A2(n23214),
	.B1(FE_OCPN28386_n17899),
	.B2(n23214),
	.C1(FE_OFN28764_n17928),
	.C2(n23214));
   NAND3xp33_ASAP7_75t_L U25774 (.Y(n17922),
	.A(n20790),
	.B(n20795),
	.C(n17920));
   NAND3x1_ASAP7_75t_SL U25775 (.Y(n22778),
	.A(n17906),
	.B(FE_OCPN29559_n17900),
	.C(FE_OCPN27429_sa12_3));
   A2O1A1Ixp33_ASAP7_75t_SL U25776 (.Y(n17925),
	.A1(n19502),
	.A2(n19510),
	.B(FE_OCPN29324_n23216),
	.C(n22778));
   NAND2x1p5_ASAP7_75t_R U25777 (.Y(n22251),
	.A(FE_OCPN29559_n17900),
	.B(n24362));
   NAND2xp33_ASAP7_75t_SL U25778 (.Y(n17932),
	.A(FE_OCPN27368_sa12_3),
	.B(n17931));
   NOR2x1_ASAP7_75t_SL U25779 (.Y(n22750),
	.A(n20554),
	.B(n20555));
   NAND2xp5_ASAP7_75t_L U25781 (.Y(n23612),
	.A(n17898),
	.B(FE_OCPN29559_n17900));
   NAND2xp5_ASAP7_75t_L U25782 (.Y(n19562),
	.A(n23600),
	.B(FE_OCPN29559_n17900));
   NOR2xp33_ASAP7_75t_SRAM U25783 (.Y(n17940),
	.A(n19546),
	.B(n20583));
   NAND2xp5_ASAP7_75t_L U25784 (.Y(n17945),
	.A(n19512),
	.B(n20542));
   NOR2x1_ASAP7_75t_L U25785 (.Y(n24585),
	.A(n22726),
	.B(n17945));
   OAI22xp33_ASAP7_75t_R U25786 (.Y(n22728),
	.A1(n24364),
	.A2(n20784),
	.B1(FE_OFN29211_n23587),
	.B2(n20784));
   A2O1A1Ixp33_ASAP7_75t_SL U25787 (.Y(n22725),
	.A1(n17906),
	.A2(FE_OFN29075_n22745),
	.B(n23214),
	.C(FE_OCPN27429_sa12_3));
   NOR3x1_ASAP7_75t_L U25788 (.Y(n23581),
	.A(FE_OFN26158_n22224),
	.B(FE_OCPN29494_sa12_4),
	.C(n17949));
   A2O1A1Ixp33_ASAP7_75t_SL U25789 (.Y(n17950),
	.A1(FE_OCPN5137_n23600),
	.A2(FE_OCPN28386_n17899),
	.B(n23581),
	.C(FE_OFN28764_n17928));
   NAND3x1_ASAP7_75t_SL U25790 (.Y(n26596),
	.A(n22252),
	.B(n22228),
	.C(n20824));
   A2O1A1Ixp33_ASAP7_75t_SL U25791 (.Y(n22253),
	.A1(FE_OCPN28198_n22776),
	.A2(FE_OCPN27729_n24362),
	.B(n22781),
	.C(FE_OFN25908_sa12_2));
   NOR2xp33_ASAP7_75t_R U25792 (.Y(n17965),
	.A(FE_OFN28834_FE_OCPN28371_n17900),
	.B(n22734));
   NAND3xp33_ASAP7_75t_SL U25793 (.Y(n24051),
	.A(n19543),
	.B(n17969),
	.C(n22266));
   A2O1A1Ixp33_ASAP7_75t_SL U25794 (.Y(n17981),
	.A1(FE_OFN28651_FE_OFN26140_n23585),
	.A2(n17980),
	.B(n24377),
	.C(n17979));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25796 (.Y(n17983),
	.A1(n26139),
	.A2(n25178),
	.B(n25748),
	.C(w1_18_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25797 (.Y(n402),
	.A1(n26139),
	.A2(n25178),
	.B(n17984),
	.C(n17983));
   NOR2x1p5_ASAP7_75t_SL U25798 (.Y(n21317),
	.A(FE_OFN29199_FE_OCPN27726_n),
	.B(n18034));
   NOR2x1p5_ASAP7_75t_SL U25799 (.Y(n18860),
	.A(FE_OCPN27405_sa03_4),
	.B(n17992));
   NAND2x1p5_ASAP7_75t_SL U25800 (.Y(n21012),
	.A(FE_OFN29158_n18860),
	.B(FE_OFN27125_n21057));
   NAND2x2_ASAP7_75t_SL U25801 (.Y(n18875),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2),
	.B(n18045));
   NOR2xp67_ASAP7_75t_L U25802 (.Y(n21310),
	.A(FE_OFN28689_sa03_5),
	.B(sa03_3_));
   NOR2x1_ASAP7_75t_L U25803 (.Y(n23455),
	.A(n18875),
	.B(FE_OCPN27998_n18019));
   NOR2x1_ASAP7_75t_SL U25804 (.Y(n21500),
	.A(FE_OCPN27726_n),
	.B(FE_OFN141_sa03_1));
   NAND2xp5_ASAP7_75t_SL U25805 (.Y(n21048),
	.A(n21500),
	.B(FE_OCPN29517_n));
   NAND2x1p5_ASAP7_75t_SL U25806 (.Y(n18029),
	.A(FE_OCPN27405_sa03_4),
	.B(FE_OFN21730_sa03_3));
   O2A1O1Ixp5_ASAP7_75t_SL U25808 (.Y(n23449),
	.A1(FE_OCPN27990_FE_OFN16132_sa03_5),
	.A2(n18029),
	.B(FE_OFN28953_n18011),
	.C(n18875));
   NOR2xp33_ASAP7_75t_SRAM U25809 (.Y(n17994),
	.A(n23450),
	.B(n23449));
   NAND2x1p5_ASAP7_75t_SL U25810 (.Y(n21511),
	.A(n17995),
	.B(FE_OFN29199_FE_OCPN27726_n));
   NOR2xp33_ASAP7_75t_SL U25812 (.Y(n18858),
	.A(FE_OFN28689_sa03_5),
	.B(n21726));
   NOR2x1p5_ASAP7_75t_SL U25813 (.Y(n21304),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2),
	.B(FE_OFN141_sa03_1));
   NAND2x1p5_ASAP7_75t_L U25814 (.Y(n23457),
	.A(n21327),
	.B(FE_OFN27125_n21057));
   A2O1A1Ixp33_ASAP7_75t_SL U25816 (.Y(n23417),
	.A1(n21327),
	.A2(n21708),
	.B(n21734),
	.C(FE_OFN21730_sa03_3));
   NOR3xp33_ASAP7_75t_SL U25817 (.Y(n18001),
	.A(n18000),
	.B(n18858),
	.C(FE_OFN29175_n21755));
   NAND2x1p5_ASAP7_75t_SL U25818 (.Y(n23439),
	.A(FE_OFN29123_n),
	.B(FE_OFN29158_n18860));
   NOR2x1_ASAP7_75t_SL U25819 (.Y(n21738),
	.A(FE_OCPN27393_sa03_0),
	.B(n18040));
   NOR2xp33_ASAP7_75t_SRAM U25820 (.Y(n18003),
	.A(n21738),
	.B(n21023));
   NOR2xp33_ASAP7_75t_SRAM U25821 (.Y(n18005),
	.A(n21295),
	.B(n21023));
   NOR2x1_ASAP7_75t_SL U25823 (.Y(n21747),
	.A(FE_OFN28677_n17998),
	.B(FE_OCPN27733_n17996));
   NAND3xp33_ASAP7_75t_L U25824 (.Y(n18010),
	.A(n18009),
	.B(n19487),
	.C(n21727));
   NOR2x1_ASAP7_75t_SL U25825 (.Y(n21015),
	.A(n23457),
	.B(FE_OCPN27675_n17986));
   NOR2xp33_ASAP7_75t_L U25826 (.Y(n18012),
	.A(n21015),
	.B(n21513));
   NAND3xp33_ASAP7_75t_L U25827 (.Y(n18027),
	.A(n23462),
	.B(n21045),
	.C(n18013));
   A2O1A1Ixp33_ASAP7_75t_R U25828 (.Y(n18018),
	.A1(FE_OCPN27483_FE_OFN16132_sa03_5),
	.A2(FE_OFN21730_sa03_3),
	.B(FE_OCPN27405_sa03_4),
	.C(n18014));
   NAND3xp33_ASAP7_75t_SL U25829 (.Y(n18017),
	.A(FE_OCPN27405_sa03_4),
	.B(n23431),
	.C(FE_OFN28689_sa03_5));
   NOR2x2_ASAP7_75t_SL U25830 (.Y(n21027),
	.A(FE_OCPN29283_n23439),
	.B(n21511));
   NOR3x1_ASAP7_75t_L U25831 (.Y(n23447),
	.A(FE_OCPN27998_n18019),
	.B(FE_OCPN27393_sa03_0),
	.C(n18040));
   NOR2x1p5_ASAP7_75t_SL U25832 (.Y(n19485),
	.A(n23447),
	.B(n17989));
   NAND2xp5_ASAP7_75t_L U25833 (.Y(n18020),
	.A(FE_OCPN5195_FE_OFN25874_sa03_2),
	.B(n21500));
   NOR2x1p5_ASAP7_75t_SL U25834 (.Y(n21729),
	.A(FE_OCPN29283_n23439),
	.B(FE_OCPN28184_n18020));
   OAI21xp5_ASAP7_75t_SL U25835 (.Y(n18023),
	.A1(FE_OFN29179_n),
	.A2(n21726),
	.B(n19483));
   NAND2x1p5_ASAP7_75t_SL U25836 (.Y(n21049),
	.A(n21531),
	.B(FE_OFN28635_n21034));
   NOR2xp33_ASAP7_75t_L U25837 (.Y(n18026),
	.A(FE_OCPN28431_n21734),
	.B(n18025));
   NAND2xp5_ASAP7_75t_R U25838 (.Y(n21035),
	.A(n21738),
	.B(FE_OFN28655_FE_OFN25986_n21012));
   NOR2x1_ASAP7_75t_L U25839 (.Y(n21301),
	.A(FE_OCPN28184_n18020),
	.B(n21725));
   OAI21xp33_ASAP7_75t_L U25840 (.Y(n18032),
	.A1(FE_OCPN28184_n18020),
	.A2(n17996),
	.B(n21034));
   NOR3xp33_ASAP7_75t_SL U25841 (.Y(n18033),
	.A(n18032),
	.B(n21296),
	.C(n18904));
   NAND3x1_ASAP7_75t_SL U25842 (.Y(n18036),
	.A(n21291),
	.B(n18033),
	.C(n23414));
   NOR2x1_ASAP7_75t_L U25843 (.Y(n21724),
	.A(n21502),
	.B(n21525));
   NOR2x1_ASAP7_75t_R U25844 (.Y(n19456),
	.A(n18859),
	.B(n21751));
   NAND3xp33_ASAP7_75t_SRAM U25845 (.Y(n18042),
	.A(n21059),
	.B(n18041),
	.C(n19456));
   OAI22xp33_ASAP7_75t_SRAM U25846 (.Y(n18050),
	.A1(FE_OFN25986_n21012),
	.A2(n18008),
	.B1(n21738),
	.B2(n18008));
   NOR3xp33_ASAP7_75t_L U25847 (.Y(n18047),
	.A(n21297),
	.B(FE_OCPN28431_n21734),
	.C(n21505));
   NAND2xp5_ASAP7_75t_L U25848 (.Y(n23418),
	.A(FE_OCPN28214_n21500),
	.B(FE_OFN25986_n21012));
   NOR3xp33_ASAP7_75t_L U25849 (.Y(n18052),
	.A(n19462),
	.B(n21513),
	.C(FE_OCPN27975_n18871));
   NOR2xp33_ASAP7_75t_SRAM U25850 (.Y(n18053),
	.A(n19492),
	.B(n21278));
   NOR3xp33_ASAP7_75t_L U25851 (.Y(n18056),
	.A(n18055),
	.B(n21504),
	.C(n18054));
   NAND3xp33_ASAP7_75t_SL U25852 (.Y(n18057),
	.A(n19470),
	.B(n18056),
	.C(n23462));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25854 (.Y(n18059),
	.A1(FE_OFN16148_n25466),
	.A2(n23916),
	.B(FE_OFN26578_n23913),
	.C(FE_OFN25934_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25855 (.Y(n318),
	.A1(FE_OFN16148_n25466),
	.A2(n23916),
	.B(n18060),
	.C(n18059));
   NOR2xp33_ASAP7_75t_SRAM U25856 (.Y(n18064),
	.A(n18062),
	.B(n18061));
   NAND3xp33_ASAP7_75t_R U25857 (.Y(n18067),
	.A(n18064),
	.B(n18063),
	.C(n21986));
   NAND3xp33_ASAP7_75t_SRAM U25858 (.Y(n18077),
	.A(n25815),
	.B(n25817),
	.C(n25816));
   NAND3xp33_ASAP7_75t_L U25859 (.Y(n18090),
	.A(n18083),
	.B(n18082),
	.C(n21925));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25860 (.Y(n18102),
	.A1(n21961),
	.A2(FE_OFN16334_n25823),
	.B(FE_OFN28528_n25241),
	.C(w2_6_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25861 (.Y(n273),
	.A1(n21961),
	.A2(FE_OFN16334_n25823),
	.B(n18103),
	.C(n18102));
   NOR3xp33_ASAP7_75t_SRAM U25862 (.Y(n18106),
	.A(FE_OFN28936_n18104),
	.B(n18114),
	.C(n24297));
   NOR2xp33_ASAP7_75t_SRAM U25863 (.Y(n18110),
	.A(n18109),
	.B(n23530));
   NOR3xp33_ASAP7_75t_L U25864 (.Y(n26091),
	.A(n18113),
	.B(n18443),
	.C(n18112));
   NOR2xp33_ASAP7_75t_SRAM U25865 (.Y(n18115),
	.A(FE_OFN29101_n16418),
	.B(n18415));
   NOR2xp33_ASAP7_75t_SRAM U25866 (.Y(n18117),
	.A(n16430),
	.B(n18415));
   NAND3xp33_ASAP7_75t_SRAM U25867 (.Y(n18127),
	.A(n18122),
	.B(n18121),
	.C(n18120));
   NOR3xp33_ASAP7_75t_L U25868 (.Y(n18139),
	.A(n18137),
	.B(n18136),
	.C(n18135));
   NAND3xp33_ASAP7_75t_R U25869 (.Y(n18153),
	.A(n18140),
	.B(n18139),
	.C(n18138));
   NOR2xp33_ASAP7_75t_SRAM U25870 (.Y(n18148),
	.A(n18433),
	.B(n18144));
   NOR3xp33_ASAP7_75t_SRAM U25871 (.Y(n18147),
	.A(n18146),
	.B(n18145),
	.C(n18426));
   OAI21x1_ASAP7_75t_L U25872 (.Y(n26087),
	.A1(n18155),
	.A2(n24331),
	.B(n18154));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25874 (.Y(n18156),
	.A1(n23571),
	.A2(FE_OFN28546_n26091),
	.B(FE_OFN25973_n26087),
	.C(w0_3_));
   NOR2x1p5_ASAP7_75t_SL U25875 (.Y(n21793),
	.A(FE_OCPN29269_sa22_1),
	.B(n23183));
   NAND2x1_ASAP7_75t_SL U25876 (.Y(n18206),
	.A(FE_OFN28688_sa22_2),
	.B(n21793));
   NAND2x1p5_ASAP7_75t_SL U25878 (.Y(n18169),
	.A(FE_OFN16135_sa22_4),
	.B(n18164));
   NAND2x1p5_ASAP7_75t_SL U25879 (.Y(n22310),
	.A(FE_OCPN29269_sa22_1),
	.B(FE_OCPN29281_sa22_0));
   NOR2x1_ASAP7_75t_L U25880 (.Y(n22293),
	.A(FE_OCPN29269_sa22_1),
	.B(FE_OFN29152_sa22_0));
   NAND2x1p5_ASAP7_75t_SL U25881 (.Y(n23303),
	.A(FE_OFN28688_sa22_2),
	.B(n22293));
   NOR3xp33_ASAP7_75t_SL U25882 (.Y(n23307),
	.A(FE_OFN29152_sa22_0),
	.B(FE_OFN28688_sa22_2),
	.C(FE_OCPN29269_sa22_1));
   NAND2x1p5_ASAP7_75t_SL U25885 (.Y(n22855),
	.A(n21793),
	.B(FE_OFN54_sa22_2));
   NOR2xp33_ASAP7_75t_SRAM U25888 (.Y(n18170),
	.A(n18199),
	.B(n18217));
   OAI21xp33_ASAP7_75t_SRAM U25889 (.Y(n18175),
	.A1(FE_OFN25987_n23322),
	.A2(FE_OCPN29478_n23306),
	.B(n22285));
   NOR3xp33_ASAP7_75t_SRAM U25890 (.Y(n18180),
	.A(n26880),
	.B(n24694),
	.C(n18175));
   NAND3xp33_ASAP7_75t_SRAM U25891 (.Y(n18240),
	.A(n24701),
	.B(n18180),
	.C(n24699));
   NOR2xp33_ASAP7_75t_R U25892 (.Y(n18182),
	.A(n18162),
	.B(FE_OFN16304_n22808));
   NOR2xp33_ASAP7_75t_R U25893 (.Y(n18183),
	.A(n23315),
	.B(FE_OFN16304_n22808));
   NAND2x2_ASAP7_75t_SL U25894 (.Y(n18186),
	.A(FE_OCPN29308_n),
	.B(n18176));
   INVxp33_ASAP7_75t_SRAM U25895 (.Y(n18189),
	.A(n26870));
   NOR2x1_ASAP7_75t_R U25896 (.Y(n22857),
	.A(FE_OCPN29305_n23302),
	.B(FE_OFN26548_n18206));
   NAND2xp5_ASAP7_75t_SL U25897 (.Y(n18216),
	.A(n23315),
	.B(n18177));
   NAND3xp33_ASAP7_75t_SRAM U25898 (.Y(n18196),
	.A(n18189),
	.B(n24702),
	.C(n26872));
   NOR2x1_ASAP7_75t_L U25899 (.Y(n22278),
	.A(n18166),
	.B(FE_OFN26548_n18206));
   NOR2x1p5_ASAP7_75t_SL U25900 (.Y(n21764),
	.A(FE_OCPN28037_n22855),
	.B(n18178));
   NAND3xp33_ASAP7_75t_R U25901 (.Y(n21788),
	.A(n23308),
	.B(n18199),
	.C(FE_RN_0_0));
   NOR3x1_ASAP7_75t_SL U25902 (.Y(n22850),
	.A(n21769),
	.B(FE_PSN8315_FE_OFN16135_sa22_4),
	.C(n21123));
   NAND3xp33_ASAP7_75t_R U25903 (.Y(n18193),
	.A(n21126),
	.B(n21788),
	.C(n18191));
   NOR2x2_ASAP7_75t_SL U25904 (.Y(n23161),
	.A(n18166),
	.B(FE_OFN25987_n23322));
   NOR3xp33_ASAP7_75t_SRAM U25905 (.Y(n18235),
	.A(n18196),
	.B(n26876),
	.C(n26875));
   NOR3xp33_ASAP7_75t_SRAM U25906 (.Y(n18212),
	.A(n23298),
	.B(FE_OFN26009_n18213),
	.C(n23185));
   NOR2xp33_ASAP7_75t_R U25907 (.Y(n18202),
	.A(n22795),
	.B(n23161));
   INVxp33_ASAP7_75t_SRAM U25908 (.Y(n18201),
	.A(n22321));
   A2O1A1Ixp33_ASAP7_75t_R U25909 (.Y(n22798),
	.A1(FE_OCPN27750_n22293),
	.A2(n23336),
	.B(n21771),
	.C(FE_OCPN27673_n18163));
   NAND3xp33_ASAP7_75t_L U25910 (.Y(n18210),
	.A(n24702),
	.B(FE_OFN28939_n21129),
	.C(n22798));
   NOR2x1_ASAP7_75t_L U25911 (.Y(n22796),
	.A(n18166),
	.B(n23303));
   NOR2xp67_ASAP7_75t_L U25912 (.Y(n18205),
	.A(n22796),
	.B(n21764));
   NOR2x1_ASAP7_75t_L U25913 (.Y(n18204),
	.A(n23323),
	.B(n23169));
   NOR2x1_ASAP7_75t_SL U25914 (.Y(n20720),
	.A(FE_OFN26548_n18206),
	.B(FE_OCPN27719_n23306));
   NOR2x1_ASAP7_75t_L U25915 (.Y(n26871),
	.A(n21770),
	.B(n23160));
   NAND3xp33_ASAP7_75t_SL U25916 (.Y(n18218),
	.A(FE_OFN28966_n23329),
	.B(n23192),
	.C(n22296));
   NOR2xp33_ASAP7_75t_SL U25917 (.Y(n18221),
	.A(FE_OCPN27947_n18177),
	.B(n21122));
   NAND2x1p5_ASAP7_75t_SL U25918 (.Y(n23197),
	.A(n18223),
	.B(n18222));
   NAND3x1_ASAP7_75t_SL U25919 (.Y(n18225),
	.A(n18215),
	.B(n18224),
	.C(n23197));
   NOR3x1_ASAP7_75t_SL U25920 (.Y(n20745),
	.A(n18225),
	.B(n22827),
	.C(FE_OCPN29585_n22281));
   NAND3xp33_ASAP7_75t_R U25921 (.Y(n18230),
	.A(n23328),
	.B(n22854),
	.C(n20773));
   NAND3xp33_ASAP7_75t_R U25922 (.Y(n18229),
	.A(n21120),
	.B(n21118),
	.C(n18228));
   OAI22xp5_ASAP7_75t_L U25923 (.Y(n23327),
	.A1(FE_OCPN29557_n18161),
	.A2(n24694),
	.B1(FE_OFN27173_n),
	.B2(n24694));
   NAND3xp33_ASAP7_75t_L U25924 (.Y(n18231),
	.A(n22295),
	.B(n23327),
	.C(n22270));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25925 (.Y(n18237),
	.A1(n26874),
	.A2(n18235),
	.B(n26889),
	.C(n26882));
   NAND3xp33_ASAP7_75t_SRAM U25926 (.Y(n18246),
	.A(n18242),
	.B(n18241),
	.C(n18268));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25927 (.Y(n18244),
	.A1(FE_OFN26170_n19361),
	.A2(FE_OFN28479_sa13_2),
	.B(FE_OFN28801_n16978),
	.C(FE_OCPN27761_n16977));
   NAND3xp33_ASAP7_75t_SRAM U25928 (.Y(n18245),
	.A(n25285),
	.B(n25221),
	.C(n18244));
   NOR2xp33_ASAP7_75t_R U25929 (.Y(n18248),
	.A(n16983),
	.B(FE_OFN132_n18247));
   NOR2xp33_ASAP7_75t_SRAM U25930 (.Y(n18250),
	.A(FE_OFN28801_n16978),
	.B(FE_OFN132_n18247));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25931 (.Y(n18259),
	.A1(FE_OFN28775_n16992),
	.A2(FE_OFN28738_n16989),
	.B(FE_OCPN8242_n20527),
	.C(n18256));
   NOR3xp33_ASAP7_75t_R U25932 (.Y(n18295),
	.A(n18259),
	.B(n20502),
	.C(n18258));
   NAND2xp33_ASAP7_75t_SL U25933 (.Y(n18274),
	.A(n20531),
	.B(n20532));
   NAND3xp33_ASAP7_75t_SRAM U25935 (.Y(n18289),
	.A(n18924),
	.B(n25221),
	.C(n18925));
   NOR2xp33_ASAP7_75t_SL U25936 (.Y(n18293),
	.A(n18292),
	.B(n18291));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25938 (.Y(n18296),
	.A1(n26915),
	.A2(n26914),
	.B(FE_OFN28473_n26911),
	.C(w2_18_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25939 (.Y(n330),
	.A1(n26915),
	.A2(n26914),
	.B(n18297),
	.C(n18296));
   NOR2xp33_ASAP7_75t_R U25940 (.Y(n20118),
	.A(FE_OFN28991_n19938),
	.B(n18818));
   NOR2xp33_ASAP7_75t_L U25941 (.Y(n20092),
	.A(n20118),
	.B(n19908));
   NOR2xp33_ASAP7_75t_L U25942 (.Y(n18300),
	.A(n19921),
	.B(FE_OCPN27792_n18333));
   NOR3xp33_ASAP7_75t_SRAM U25943 (.Y(n18301),
	.A(n22385),
	.B(FE_OCPN27937_n18841),
	.C(FE_OCPN27490_n18798));
   NAND3xp33_ASAP7_75t_SRAM U25944 (.Y(n18305),
	.A(n20092),
	.B(n18301),
	.C(n19924));
   NOR3xp33_ASAP7_75t_R U25945 (.Y(n25026),
	.A(n18805),
	.B(n19728),
	.C(n18307));
   NAND3x1_ASAP7_75t_L U25946 (.Y(n18312),
	.A(n18309),
	.B(n22372),
	.C(n20111));
   NOR3xp33_ASAP7_75t_SL U25947 (.Y(n18313),
	.A(n18312),
	.B(n19926),
	.C(n18311));
   NAND3xp33_ASAP7_75t_SL U25948 (.Y(n18314),
	.A(n18811),
	.B(n18313),
	.C(n18325));
   NOR2xp33_ASAP7_75t_SRAM U25949 (.Y(n18315),
	.A(FE_OCPN28434_n17546),
	.B(n18842));
   NOR2xp33_ASAP7_75t_SRAM U25950 (.Y(n18316),
	.A(n18298),
	.B(n18842));
   NAND3xp33_ASAP7_75t_L U25951 (.Y(n18345),
	.A(n25024),
	.B(n18319),
	.C(n25022));
   NAND3xp33_ASAP7_75t_SL U25952 (.Y(n18323),
	.A(n18336),
	.B(n19943),
	.C(n18814));
   NAND3xp33_ASAP7_75t_SL U25953 (.Y(n18337),
	.A(n20093),
	.B(n19951),
	.C(n19720));
   A2O1A1Ixp33_ASAP7_75t_SL U25954 (.Y(n25020),
	.A1(n19956),
	.A2(n18344),
	.B(n23899),
	.C(n18343));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25955 (.Y(n18347),
	.A1(n17580),
	.A2(n18349),
	.B(n25143),
	.C(FE_OFN140_w3_2));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25956 (.Y(n412),
	.A1(n17580),
	.A2(n18349),
	.B(n18348),
	.C(n18347));
   NOR2xp33_ASAP7_75t_SRAM U25957 (.Y(n18353),
	.A(FE_OFN27176_n),
	.B(n24779));
   NOR2x1_ASAP7_75t_L U25958 (.Y(n26029),
	.A(FE_PSN8270_n26027),
	.B(n21625));
   NOR2xp33_ASAP7_75t_SRAM U25959 (.Y(n18355),
	.A(n18495),
	.B(n24779));
   NAND3xp33_ASAP7_75t_SRAM U25960 (.Y(n18403),
	.A(n24579),
	.B(n24580),
	.C(n24581));
   NOR2x1p5_ASAP7_75t_L U25961 (.Y(n22139),
	.A(n18473),
	.B(n21625));
   NOR2xp33_ASAP7_75t_L U25962 (.Y(n18359),
	.A(FE_OFN29121_n26026),
	.B(FE_OFN28790_n));
   NAND3xp33_ASAP7_75t_SL U25963 (.Y(n18361),
	.A(n18388),
	.B(n18360),
	.C(n25113));
   NOR3xp33_ASAP7_75t_SL U25964 (.Y(n22639),
	.A(n18361),
	.B(n18373),
	.C(n18506));
   NOR3xp33_ASAP7_75t_SRAM U25965 (.Y(n18366),
	.A(n22640),
	.B(n18458),
	.C(n18365));
   NOR2xp33_ASAP7_75t_SL U25966 (.Y(n18487),
	.A(n22168),
	.B(n21586));
   NAND3xp33_ASAP7_75t_L U25967 (.Y(n18367),
	.A(n18455),
	.B(n18366),
	.C(n18487));
   AND3x1_ASAP7_75t_SL U25968 (.Y(n18375),
	.A(n24785),
	.B(n22151),
	.C(n19056));
   A2O1A1Ixp33_ASAP7_75t_L U25969 (.Y(n18480),
	.A1(FE_OFN26597_n),
	.A2(n17606),
	.B(n19037),
	.C(n18379));
   NAND3xp33_ASAP7_75t_R U25970 (.Y(n18380),
	.A(n24780),
	.B(FE_OCPN28378_n22632),
	.C(FE_OFN28901_sa30_4));
   NAND3xp33_ASAP7_75t_SL U25971 (.Y(n18383),
	.A(n18480),
	.B(n18380),
	.C(n18499));
   NAND2x1p5_ASAP7_75t_SL U25972 (.Y(n26028),
	.A(n19078),
	.B(n18384));
   NOR2x1_ASAP7_75t_SL U25973 (.Y(n18386),
	.A(n18385),
	.B(n26028));
   NOR2x1_ASAP7_75t_L U25974 (.Y(n18397),
	.A(n26687),
	.B(n18386));
   NAND2x1p5_ASAP7_75t_SL U25975 (.Y(n25105),
	.A(FE_OFN29094_n21607),
	.B(FE_OCPN28057_n17603));
   NOR2x1_ASAP7_75t_SL U25976 (.Y(n18508),
	.A(FE_OFN28896_sa30_2),
	.B(n25105));
   NAND3xp33_ASAP7_75t_SRAM U25977 (.Y(n19033),
	.A(FE_OCPN29431_sa30_3),
	.B(n17618),
	.C(n17602));
   NAND3xp33_ASAP7_75t_L U25978 (.Y(n18391),
	.A(n20469),
	.B(n19033),
	.C(n18388));
   NOR2xp33_ASAP7_75t_L U25979 (.Y(n18389),
	.A(n18458),
	.B(n21590));
   NAND3xp33_ASAP7_75t_SL U25980 (.Y(n19075),
	.A(n18392),
	.B(n19036),
	.C(n22646));
   A2O1A1Ixp33_ASAP7_75t_SL U25981 (.Y(n26442),
	.A1(n18485),
	.A2(n18399),
	.B(n26926),
	.C(n18398));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25982 (.Y(n18401),
	.A1(FE_OFN16164_n25081),
	.A2(n18403),
	.B(FE_OCPN29458_n26442),
	.C(w1_7_));
   NAND3xp33_ASAP7_75t_SRAM U25983 (.Y(n24618),
	.A(n18406),
	.B(n18405),
	.C(n18404));
   NOR2xp33_ASAP7_75t_SRAM U25984 (.Y(n18407),
	.A(FE_OCPN27555_n16422),
	.B(n24613));
   NOR2xp33_ASAP7_75t_SRAM U25985 (.Y(n18409),
	.A(FE_OFN28592_n16427),
	.B(n24613));
   NOR2xp33_ASAP7_75t_SRAM U25986 (.Y(n18417),
	.A(FE_OCPN7607_n23539),
	.B(n18415));
   NAND3xp33_ASAP7_75t_SRAM U25987 (.Y(n18419),
	.A(n18417),
	.B(n24614),
	.C(n18416));
   NOR3xp33_ASAP7_75t_SRAM U25989 (.Y(n18427),
	.A(n18426),
	.B(FE_OFN27090_n23558),
	.C(FE_OCPN28141_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25992 (.Y(n18450),
	.A1(n26770),
	.A2(n26769),
	.B(n26766),
	.C(FE_OFN48_w0_2));
   A2O1A1Ixp33_ASAP7_75t_SRAM U25993 (.Y(n377),
	.A1(n26770),
	.A2(n26769),
	.B(n18451),
	.C(n18450));
   NAND2xp5_ASAP7_75t_L U25994 (.Y(n26025),
	.A(FE_OFN28637_n25102),
	.B(FE_OCPN8207_n18497));
   NOR2xp33_ASAP7_75t_SRAM U25995 (.Y(n18454),
	.A(n17601),
	.B(FE_OFN16200_sa30_2));
   NAND2xp5_ASAP7_75t_R U25996 (.Y(n18498),
	.A(n18454),
	.B(n25108));
   A2O1A1Ixp33_ASAP7_75t_R U25997 (.Y(n20453),
	.A1(n17603),
	.A2(FE_OFN28895_sa30_2),
	.B(n18458),
	.C(FE_OCPN8207_n18497));
   NOR2x1_ASAP7_75t_SL U25998 (.Y(n18461),
	.A(n18460),
	.B(n18459));
   NAND3x1_ASAP7_75t_SL U25999 (.Y(n24789),
	.A(n22130),
	.B(n18462),
	.C(n18461));
   NOR2xp33_ASAP7_75t_SRAM U26000 (.Y(n18465),
	.A(FE_OCPN29399_sa30_3),
	.B(FE_OFN16333_sa30_4));
   NOR2xp33_ASAP7_75t_SRAM U26001 (.Y(n18468),
	.A(n24779),
	.B(n24781));
   NAND3xp33_ASAP7_75t_SRAM U26002 (.Y(n18469),
	.A(n18468),
	.B(n22621),
	.C(n24802));
   NOR2xp33_ASAP7_75t_SRAM U26003 (.Y(n18470),
	.A(FE_OCPN29496_n24789),
	.B(n18469));
   NAND3xp33_ASAP7_75t_SRAM U26004 (.Y(n18520),
	.A(n24787),
	.B(n18470),
	.C(n24785));
   NAND3xp33_ASAP7_75t_SRAM U26005 (.Y(n18477),
	.A(n24127),
	.B(n18471),
	.C(n22151));
   OAI21xp5_ASAP7_75t_L U26006 (.Y(n21597),
	.A1(FE_OFN25901_n22133),
	.A2(FE_OCPN27966_n18473),
	.B(n22626));
   NOR3xp33_ASAP7_75t_SRAM U26007 (.Y(n18514),
	.A(n18477),
	.B(n24791),
	.C(n26022));
   NAND2xp5_ASAP7_75t_L U26008 (.Y(n19054),
	.A(n17603),
	.B(FE_OCPN8207_n18497));
   NOR3xp33_ASAP7_75t_SL U26009 (.Y(n19042),
	.A(n20439),
	.B(n22629),
	.C(n18508));
   NAND3xp33_ASAP7_75t_SL U26010 (.Y(n18494),
	.A(n18488),
	.B(n18487),
	.C(n19042));
   NOR2xp33_ASAP7_75t_SRAM U26011 (.Y(n18491),
	.A(n20450),
	.B(n22641));
   OAI22xp5_ASAP7_75t_L U26012 (.Y(n25115),
	.A1(n17602),
	.A2(n22613),
	.B1(n18495),
	.B2(n22613));
   OAI22xp5_ASAP7_75t_L U26013 (.Y(n22138),
	.A1(FE_OCPN8207_n18497),
	.A2(n22139),
	.B1(FE_OCPN28057_n17603),
	.B2(n22139));
   OAI222xp33_ASAP7_75t_SRAM U26014 (.Y(n18512),
	.A1(n18511),
	.A2(n26926),
	.B1(n25104),
	.B2(n26926),
	.C1(n24760),
	.C2(n26926));
   A2O1A1Ixp33_ASAP7_75t_R U26015 (.Y(n18517),
	.A1(n18514),
	.A2(n24794),
	.B(n26687),
	.C(n18513));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26016 (.Y(n18518),
	.A1(n25081),
	.A2(n18520),
	.B(n18517),
	.C(w1_0_));
   OAI21xp33_ASAP7_75t_L U26017 (.Y(n21674),
	.A1(FE_OFN28815_n18523),
	.A2(n18544),
	.B(n21637));
   NOR3x2_ASAP7_75t_SL U26018 (.Y(n23869),
	.A(FE_OFN29223_sa20_0),
	.B(FE_OCPN27371_sa20_2),
	.C(FE_OCPN29380_sa20_1));
   NOR3xp33_ASAP7_75t_SL U26019 (.Y(n23875),
	.A(FE_OCPN27633_sa20_5),
	.B(n18536),
	.C(FE_OFN29178_sa20_4));
   NAND2xp5_ASAP7_75t_SL U26020 (.Y(n18588),
	.A(FE_OFN29081_n18526),
	.B(FE_OCPN27715_n23875));
   NOR3xp33_ASAP7_75t_SRAM U26021 (.Y(n18543),
	.A(n18528),
	.B(FE_OFN28607_n23884),
	.C(n21658));
   NOR2x2_ASAP7_75t_SL U26022 (.Y(n21195),
	.A(n18536),
	.B(FE_OCPN27558_sa20_4));
   NOR2x1_ASAP7_75t_SL U26023 (.Y(n21691),
	.A(n20654),
	.B(n18531));
   NAND2x1p5_ASAP7_75t_L U26025 (.Y(n18571),
	.A(n18536),
	.B(FE_OCPN27633_sa20_5));
   NAND3xp33_ASAP7_75t_SL U26026 (.Y(n23837),
	.A(FE_OCPN27558_sa20_4),
	.B(FE_OCPN27633_sa20_5),
	.C(n18536));
   NAND2x1p5_ASAP7_75t_SL U26027 (.Y(n18534),
	.A(FE_OCPN28163_FE_OFN99_sa20_5),
	.B(n21195));
   NOR2x1p5_ASAP7_75t_SL U26028 (.Y(n23814),
	.A(FE_OFN28815_n18523),
	.B(FE_OCPN28353_n18534));
   OAI22xp33_ASAP7_75t_L U26029 (.Y(n18537),
	.A1(n20685),
	.A2(n23814),
	.B1(FE_OFN28986_n18597),
	.B2(n23814));
   NAND2x1_ASAP7_75t_L U26030 (.Y(n21664),
	.A(FE_OFN28988_n18597),
	.B(FE_OCPN27715_n23875));
   NOR2x1p5_ASAP7_75t_L U26031 (.Y(n23740),
	.A(FE_OCPN27891_n18561),
	.B(n18530));
   NAND3xp33_ASAP7_75t_SL U26032 (.Y(n26322),
	.A(n18543),
	.B(n18542),
	.C(n18541));
   NAND3x1_ASAP7_75t_SL U26033 (.Y(n18566),
	.A(n21239),
	.B(n21684),
	.C(n25328));
   INVxp33_ASAP7_75t_SRAM U26034 (.Y(n18550),
	.A(n23694));
   NOR3xp33_ASAP7_75t_R U26035 (.Y(n18560),
	.A(n23764),
	.B(n23791),
	.C(n18550));
   NAND2x2_ASAP7_75t_SL U26036 (.Y(n23838),
	.A(FE_OCPN29584_n),
	.B(n18532));
   NAND3xp33_ASAP7_75t_L U26037 (.Y(n23833),
	.A(n18529),
	.B(FE_OCPN27715_n23875),
	.C(FE_OFN29131_FE_OCPN27371_sa20_2));
   OAI21xp33_ASAP7_75t_L U26039 (.Y(n20660),
	.A1(n18530),
	.A2(FE_OCPN27891_n18561),
	.B(n21664));
   NAND2xp33_ASAP7_75t_SL U26040 (.Y(n18555),
	.A(n18554),
	.B(n21637));
   NOR2x1_ASAP7_75t_SL U26041 (.Y(n23719),
	.A(n18561),
	.B(n20670));
   NOR2x1_ASAP7_75t_L U26042 (.Y(n21648),
	.A(FE_OFN28815_n18523),
	.B(n23711));
   NOR2xp67_ASAP7_75t_L U26043 (.Y(n20653),
	.A(n18530),
	.B(n23711));
   NAND3x2_ASAP7_75t_L U26045 (.Y(n25188),
	.A(FE_OFN29081_n18526),
	.B(FE_OFN29200_n18521),
	.C(FE_OCPN27542_sa20_3));
   NOR2xp33_ASAP7_75t_SRAM U26046 (.Y(n18576),
	.A(n21669),
	.B(n21682));
   NAND3xp33_ASAP7_75t_L U26047 (.Y(n21665),
	.A(n18532),
	.B(FE_OCPN27715_n23875),
	.C(FE_OFN29091_n));
   AND3x1_ASAP7_75t_SL U26048 (.Y(n21200),
	.A(n18579),
	.B(n21235),
	.C(n20644));
   AND2x2_ASAP7_75t_R U26049 (.Y(n18590),
	.A(n18588),
	.B(n21637));
   NAND2xp5_ASAP7_75t_L U26050 (.Y(n23755),
	.A(n18583),
	.B(FE_OFN29081_n18526));
   NAND3xp33_ASAP7_75t_L U26051 (.Y(n21256),
	.A(n23833),
	.B(n23755),
	.C(n23716));
   O2A1O1Ixp33_ASAP7_75t_SL U26052 (.Y(n18610),
	.A1(n23798),
	.A2(n18609),
	.B(n27207),
	.C(n18608));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26054 (.Y(n18612),
	.A1(n26323),
	.A2(n26322),
	.B(FE_OCPN7642_n26319),
	.C(w2_11_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26055 (.Y(n363),
	.A1(n26323),
	.A2(n26322),
	.B(n18613),
	.C(n18612));
   NOR2xp33_ASAP7_75t_SRAM U26056 (.Y(n18615),
	.A(n19609),
	.B(FE_PSN8318_n21455));
   NOR2xp33_ASAP7_75t_SRAM U26057 (.Y(n18617),
	.A(FE_OCPN29346_n12998),
	.B(FE_PSN8318_n21455));
   NAND3xp33_ASAP7_75t_SRAM U26059 (.Y(n18622),
	.A(FE_OCPN27500_n19834),
	.B(FE_OFN28835_n),
	.C(FE_OFN29172_sa00_4));
   NAND3xp33_ASAP7_75t_SRAM U26060 (.Y(n21474),
	.A(FE_PSN8286_FE_OCPN29260_sa00_5),
	.B(FE_OCPN29295_n18739),
	.C(FE_PSN8285_FE_OCPN29463_n));
   NAND3xp33_ASAP7_75t_L U26061 (.Y(n18624),
	.A(n18622),
	.B(n21474),
	.C(n18632));
   NOR3xp33_ASAP7_75t_SRAM U26062 (.Y(n18625),
	.A(n19118),
	.B(FE_OCPN27588_n19824),
	.C(n21148));
   NAND3xp33_ASAP7_75t_SRAM U26063 (.Y(n18634),
	.A(n18652),
	.B(n18756),
	.C(n24085));
   OAI21xp5_ASAP7_75t_L U26065 (.Y(n18638),
	.A1(n19097),
	.A2(n19817),
	.B(n26103));
   NOR2xp33_ASAP7_75t_SRAM U26066 (.Y(n18644),
	.A(FE_OFN16216_n19573),
	.B(FE_OCPN27703_n19847));
   NOR2xp33_ASAP7_75t_SRAM U26067 (.Y(n18646),
	.A(FE_OCPN29542_n21151),
	.B(FE_OCPN27703_n19847));
   O2A1O1Ixp5_ASAP7_75t_SL U26068 (.Y(n18662),
	.A1(n19611),
	.A2(n18661),
	.B(n26637),
	.C(n18660));
   OAI21x1_ASAP7_75t_SL U26069 (.Y(n27056),
	.A1(n18663),
	.A2(n21493),
	.B(n18662));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26070 (.Y(n18664),
	.A1(n27127),
	.A2(n25255),
	.B(FE_OCPN7658_n27056),
	.C(FE_OFN64_w0_31));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26071 (.Y(n296),
	.A1(n27127),
	.A2(n25255),
	.B(n18665),
	.C(n18664));
   NOR3xp33_ASAP7_75t_SRAM U26072 (.Y(n18670),
	.A(n18668),
	.B(n22582),
	.C(n20391));
   NAND3xp33_ASAP7_75t_R U26073 (.Y(n18674),
	.A(n18670),
	.B(n22605),
	.C(n21557));
   NAND3xp33_ASAP7_75t_SRAM U26074 (.Y(n18673),
	.A(n20367),
	.B(n22470),
	.C(n18672));
   NOR3xp33_ASAP7_75t_L U26075 (.Y(n18676),
	.A(n18674),
	.B(n23076),
	.C(n18673));
   NAND2xp5_ASAP7_75t_SL U26076 (.Y(n22469),
	.A(n17321),
	.B(FE_OFN28594_n26454));
   NOR3xp33_ASAP7_75t_L U26077 (.Y(n18692),
	.A(n23069),
	.B(n18678),
	.C(n20366));
   NOR2xp33_ASAP7_75t_L U26078 (.Y(n18679),
	.A(n17321),
	.B(n18717));
   NOR2xp33_ASAP7_75t_L U26079 (.Y(n18682),
	.A(n20404),
	.B(n21571));
   AND3x1_ASAP7_75t_SL U26080 (.Y(n18689),
	.A(n22596),
	.B(n18687),
	.C(n21552));
   NAND3x1_ASAP7_75t_SL U26081 (.Y(n18697),
	.A(n18692),
	.B(FE_OFN29000_n18698),
	.C(n23113));
   OAI21xp5_ASAP7_75t_L U26082 (.Y(n20388),
	.A1(FE_OCPN29334_n17330),
	.A2(FE_OFN27072_n18671),
	.B(n22457));
   NOR2x1_ASAP7_75t_L U26083 (.Y(n23092),
	.A(n18693),
	.B(n17318));
   NAND3xp33_ASAP7_75t_SL U26084 (.Y(n22599),
	.A(n18695),
	.B(n18694),
	.C(n22590));
   NOR3x1_ASAP7_75t_SL U26085 (.Y(n24404),
	.A(n18697),
	.B(n18696),
	.C(n22579));
   AND2x2_ASAP7_75t_SL U26086 (.Y(n18700),
	.A(n26451),
	.B(FE_OCPN28310_n22585));
   NOR2xp33_ASAP7_75t_SL U26087 (.Y(n18701),
	.A(n17321),
	.B(n21544));
   NAND3xp33_ASAP7_75t_SL U26088 (.Y(n18712),
	.A(n18706),
	.B(n18705),
	.C(n18704));
   A2O1A1Ixp33_ASAP7_75t_L U26089 (.Y(n21539),
	.A1(FE_OCPN29409_n22461),
	.A2(n21553),
	.B(n27006),
	.C(n17326));
   A2O1A1Ixp33_ASAP7_75t_SL U26090 (.Y(n24391),
	.A1(FE_OCPN29388_n22461),
	.A2(FE_OFN16141_sa01_3),
	.B(n18714),
	.C(FE_OCPN27871_n17317));
   NOR3xp33_ASAP7_75t_SRAM U26091 (.Y(n24395),
	.A(n22435),
	.B(n18717),
	.C(n23075));
   NOR2xp33_ASAP7_75t_L U26092 (.Y(n18720),
	.A(FE_OCPN28301_n22448),
	.B(n22447));
   NAND3xp33_ASAP7_75t_R U26093 (.Y(n18725),
	.A(n22588),
	.B(n18721),
	.C(n18720));
   NOR3xp33_ASAP7_75t_SL U26094 (.Y(n23073),
	.A(n18723),
	.B(n20365),
	.C(n18722));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26095 (.Y(n18732),
	.A1(n26282),
	.A2(FE_OCPN29352_n25173),
	.B(FE_OCPN7598_n25174),
	.C(w1_26_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26096 (.Y(n394),
	.A1(n26282),
	.A2(FE_OCPN29352_n25173),
	.B(n18733),
	.C(n18732));
   NAND3x1_ASAP7_75t_SL U26097 (.Y(n26226),
	.A(n18738),
	.B(n18737),
	.C(n19598));
   NOR2x1p5_ASAP7_75t_SL U26098 (.Y(n19601),
	.A(n26101),
	.B(n21455));
   OAI21x1_ASAP7_75t_SL U26099 (.Y(n19091),
	.A1(FE_OCPN27649_n17236),
	.A2(FE_OCPN27951_n19098),
	.B(n18765));
   NOR2x1p5_ASAP7_75t_SL U26100 (.Y(n19154),
	.A(n18746),
	.B(n18745));
   NAND3x1_ASAP7_75t_SL U26101 (.Y(n19841),
	.A(n18748),
	.B(n18747),
	.C(n19154));
   NOR2x1_ASAP7_75t_SL U26102 (.Y(n18749),
	.A(n19117),
	.B(n19841));
   NAND2x1_ASAP7_75t_SL U26103 (.Y(n21164),
	.A(n18749),
	.B(n18766));
   NAND3xp33_ASAP7_75t_R U26104 (.Y(n18754),
	.A(n18752),
	.B(n21442),
	.C(n19854));
   OAI21xp5_ASAP7_75t_SL U26105 (.Y(n19610),
	.A1(n19817),
	.A2(FE_OCPN27649_n17236),
	.B(n24092));
   A2O1A1Ixp33_ASAP7_75t_SL U26106 (.Y(n19575),
	.A1(FE_OCPN27951_n19098),
	.A2(n17275),
	.B(FE_OCPN27649_n17236),
	.C(n18758));
   NOR3xp33_ASAP7_75t_SL U26107 (.Y(n18762),
	.A(n19138),
	.B(n19575),
	.C(n19848));
   NOR3xp33_ASAP7_75t_SRAM U26108 (.Y(n18760),
	.A(FE_OFN29079_FE_OCPN27518_n17251),
	.B(FE_OFN29172_sa00_4),
	.C(FE_PSN8286_FE_OCPN29260_sa00_5));
   A2O1A1Ixp33_ASAP7_75t_L U26110 (.Y(n21482),
	.A1(FE_OCPN27500_n19834),
	.A2(FE_PSN8282_n21154),
	.B(FE_OCPN27588_n19824),
	.C(FE_OFN29172_sa00_4));
   NAND3xp33_ASAP7_75t_SRAM U26111 (.Y(n18772),
	.A(n19132),
	.B(n18770),
	.C(n21482));
   OA21x2_ASAP7_75t_R U26112 (.Y(n19123),
	.A1(FE_OFN29079_FE_OCPN27518_n17251),
	.A2(n19817),
	.B(n18773));
   NOR2xp33_ASAP7_75t_SRAM U26113 (.Y(n18777),
	.A(FE_OCPN29346_n12998),
	.B(n18776));
   O2A1O1Ixp5_ASAP7_75t_SL U26114 (.Y(n18784),
	.A1(n19610),
	.A2(n18783),
	.B(n27127),
	.C(n18782));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26115 (.Y(n18787),
	.A1(FE_OFN16170_n26637),
	.A2(n26226),
	.B(FE_OFN29180_n26222),
	.C(w0_27_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26116 (.Y(n323),
	.A1(FE_OFN16170_n26637),
	.A2(n26226),
	.B(n18788),
	.C(n18787));
   NOR2xp33_ASAP7_75t_R U26117 (.Y(n24856),
	.A(FE_OCPN28229_n17529),
	.B(n20095));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26118 (.Y(n18802),
	.A1(n18793),
	.A2(n18827),
	.B(FE_OCPN29298_n25028),
	.C(n24866));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26119 (.Y(n18796),
	.A1(n18818),
	.A2(FE_OCPN27420_n18794),
	.B(FE_OCPN28423_n18836),
	.C(n22386));
   NOR3xp33_ASAP7_75t_SL U26120 (.Y(n19738),
	.A(n18796),
	.B(n19907),
	.C(n18795));
   NOR3xp33_ASAP7_75t_SL U26121 (.Y(n18803),
	.A(n18802),
	.B(n19908),
	.C(n19935));
   NOR2xp33_ASAP7_75t_SRAM U26122 (.Y(n18806),
	.A(FE_OCPN28434_n17546),
	.B(n22399));
   NOR2xp33_ASAP7_75t_SRAM U26123 (.Y(n18808),
	.A(n17527),
	.B(n22399));
   NAND3xp33_ASAP7_75t_R U26124 (.Y(n18817),
	.A(n18812),
	.B(n19720),
	.C(n18811));
   NAND3xp33_ASAP7_75t_L U26125 (.Y(n18816),
	.A(n18815),
	.B(n18814),
	.C(n18813));
   NAND3xp33_ASAP7_75t_SL U26126 (.Y(n18821),
	.A(n18820),
	.B(n18819),
	.C(n23900));
   NAND3xp33_ASAP7_75t_SL U26128 (.Y(n19730),
	.A(n18824),
	.B(n18823),
	.C(n22379));
   NAND3xp33_ASAP7_75t_L U26129 (.Y(n18831),
	.A(FE_OFN28965_n24869),
	.B(n18826),
	.C(n18825));
   NOR3xp33_ASAP7_75t_R U26130 (.Y(n19910),
	.A(n18832),
	.B(FE_OFN27148_sa32_3),
	.C(n18837));
   NOR2xp33_ASAP7_75t_SRAM U26131 (.Y(n18840),
	.A(n19921),
	.B(n18838));
   O2A1O1Ixp33_ASAP7_75t_SL U26132 (.Y(n18854),
	.A1(FE_OFN28609_n19730),
	.A2(n18853),
	.B(n17580),
	.C(n18852));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26133 (.Y(n18856),
	.A1(n22405),
	.A2(FE_OCPN27940_n26842),
	.B(n26839),
	.C(FE_OFN16313_w3_0));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26134 (.Y(n414),
	.A1(n22405),
	.A2(FE_OCPN27940_n26842),
	.B(n18857),
	.C(n18856));
   OAI21xp5_ASAP7_75t_L U26135 (.Y(n19448),
	.A1(n21706),
	.A2(FE_OCPN27948_FE_OFN26173_n21511),
	.B(FE_OFN16294_n19461));
   NOR3xp33_ASAP7_75t_SRAM U26136 (.Y(n18863),
	.A(n21731),
	.B(FE_OCPN27611_n23426),
	.C(n21747));
   NAND3xp33_ASAP7_75t_L U26137 (.Y(n18865),
	.A(n21282),
	.B(n18863),
	.C(n18862));
   NOR2x1_ASAP7_75t_SL U26138 (.Y(n21275),
	.A(n21278),
	.B(n23451));
   OAI22xp5_ASAP7_75t_L U26139 (.Y(n18866),
	.A1(n21708),
	.A2(n21017),
	.B1(FE_OFN28656_FE_OFN25986_n21012),
	.B2(n21017));
   NOR3x1_ASAP7_75t_SL U26140 (.Y(n21071),
	.A(n18870),
	.B(n18869),
	.C(n18868));
   INVxp33_ASAP7_75t_SRAM U26141 (.Y(n21269),
	.A(FE_OCPN27599_n18875));
   NAND3xp33_ASAP7_75t_R U26142 (.Y(n18877),
	.A(n21510),
	.B(n18876),
	.C(n21077));
   NOR2xp33_ASAP7_75t_SL U26143 (.Y(n18881),
	.A(FE_OCPN27617_n18016),
	.B(n21518));
   NOR2xp33_ASAP7_75t_R U26144 (.Y(n18883),
	.A(FE_OCPN28214_n21500),
	.B(n21518));
   OAI21xp33_ASAP7_75t_L U26145 (.Y(n18909),
	.A1(FE_OCPN28184_n18020),
	.A2(FE_OFN28954_n18011),
	.B(n18886));
   OAI21xp5_ASAP7_75t_SL U26146 (.Y(n18891),
	.A1(n23457),
	.A2(FE_OFN28588_n21048),
	.B(n21059));
   OAI21xp5_ASAP7_75t_SL U26147 (.Y(n21728),
	.A1(FE_OCPN29283_n23439),
	.A2(FE_OFN28677_n17998),
	.B(n21719));
   NAND3xp33_ASAP7_75t_SL U26148 (.Y(n18893),
	.A(n21064),
	.B(n18892),
	.C(n21014));
   NOR2xp33_ASAP7_75t_SL U26149 (.Y(n18894),
	.A(n21733),
	.B(n23450));
   NOR2xp33_ASAP7_75t_SRAM U26150 (.Y(n18899),
	.A(FE_OCPN27998_n18019),
	.B(FE_OCPN28184_n18020));
   NAND3xp33_ASAP7_75t_SL U26151 (.Y(n18901),
	.A(n23429),
	.B(n21718),
	.C(n18900));
   O2A1O1Ixp5_ASAP7_75t_SL U26152 (.Y(n18910),
	.A1(n18909),
	.A2(n18908),
	.B(n26819),
	.C(n18907));
   NAND2xp33_ASAP7_75t_SRAM U26154 (.Y(n18913),
	.A(FE_OCPN27682_n25414),
	.B(FE_OFN26120_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26155 (.Y(n18912),
	.A1(FE_OFN16148_n25466),
	.A2(n18914),
	.B(FE_OFN28902_n25414),
	.C(FE_OFN27100_n25675));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26156 (.Y(n317),
	.A1(FE_OFN16148_n25466),
	.A2(n18914),
	.B(n18913),
	.C(n18912));
   NOR2xp33_ASAP7_75t_SRAM U26157 (.Y(n18920),
	.A(n25885),
	.B(n18917));
   NAND3x1_ASAP7_75t_SL U26158 (.Y(n18929),
	.A(n18923),
	.B(n25222),
	.C(n19438));
   NAND2xp5_ASAP7_75t_L U26159 (.Y(n18927),
	.A(n18926),
	.B(n19414));
   NOR3x1_ASAP7_75t_SL U26160 (.Y(n25864),
	.A(n18929),
	.B(n18928),
	.C(n18927));
   NAND3xp33_ASAP7_75t_SRAM U26161 (.Y(n25866),
	.A(n25995),
	.B(n25994),
	.C(n18931));
   NOR3xp33_ASAP7_75t_SRAM U26162 (.Y(n18933),
	.A(n25866),
	.B(FE_OCPN29525_n18947),
	.C(n25996));
   OAI222xp33_ASAP7_75t_SRAM U26163 (.Y(n18963),
	.A1(n25997),
	.A2(n26959),
	.B1(n18933),
	.B2(n26959),
	.C1(n26001),
	.C2(n26959));
   O2A1O1Ixp5_ASAP7_75t_SRAM U26164 (.Y(n18945),
	.A1(FE_OFN16396_n25869),
	.A2(FE_OCPN27761_n16977),
	.B(FE_OCPN8213_FE_OFN29234_n16996),
	.C(FE_OFN28919_n24155));
   NOR2x1_ASAP7_75t_L U26165 (.Y(n25887),
	.A(n18943),
	.B(n18942));
   NOR2xp33_ASAP7_75t_SL U26166 (.Y(n18948),
	.A(FE_OCPN27859_n25868),
	.B(n19410));
   NAND3xp33_ASAP7_75t_SL U26167 (.Y(n18961),
	.A(n25988),
	.B(n18952),
	.C(n18951));
   NOR2xp33_ASAP7_75t_SRAM U26168 (.Y(n18953),
	.A(FE_OFN28801_n16978),
	.B(n18954));
   NAND2x1p5_ASAP7_75t_SL U26169 (.Y(n25293),
	.A(n24172),
	.B(n18959));
   NOR2x1p5_ASAP7_75t_SL U26170 (.Y(n22009),
	.A(FE_OCPN27627_sa23_1),
	.B(n22950));
   NAND2x1p5_ASAP7_75t_SL U26171 (.Y(n20235),
	.A(FE_OFN29191_sa23_2),
	.B(n22009));
   NOR2x1p5_ASAP7_75t_L U26172 (.Y(n23472),
	.A(n20241),
	.B(n20235));
   NOR2x1_ASAP7_75t_SL U26174 (.Y(n22964),
	.A(FE_OCPN27803_sa23_4),
	.B(FE_OFN27078_sa23_5));
   NAND2x1p5_ASAP7_75t_L U26175 (.Y(n20920),
	.A(FE_OFN27126_sa23_3),
	.B(n22964));
   NOR2x1_ASAP7_75t_SL U26176 (.Y(n20224),
	.A(FE_OCPN29488_FE_OFN25883_n22945),
	.B(FE_OCPN28266_n20920));
   NOR3xp33_ASAP7_75t_SL U26177 (.Y(n23487),
	.A(FE_OCPN27627_sa23_1),
	.B(FE_OFN29191_sa23_2),
	.C(FE_OFN29189_sa23_0));
   NOR3xp33_ASAP7_75t_L U26178 (.Y(n26557),
	.A(n23472),
	.B(n20224),
	.C(n20255));
   NAND3x1_ASAP7_75t_SL U26179 (.Y(n20913),
	.A(FE_OFN29189_sa23_0),
	.B(FE_OCPN27627_sa23_1),
	.C(FE_OFN29191_sa23_2));
   NOR2x1p5_ASAP7_75t_L U26180 (.Y(n20933),
	.A(FE_OCPN29489_sa23_3),
	.B(FE_OCPN27803_sa23_4));
   A2O1A1Ixp33_ASAP7_75t_L U26181 (.Y(n18972),
	.A1(FE_OFN29187_FE_OCPN27571_n20235),
	.A2(FE_OFN25889_n20913),
	.B(n22980),
	.C(FE_OCPN5191_n20272));
   NOR2x1_ASAP7_75t_SL U26182 (.Y(n26664),
	.A(FE_OCPN29373_FE_OFN29191_sa23_2),
	.B(n22970));
   NOR3xp33_ASAP7_75t_SL U26183 (.Y(n22995),
	.A(FE_OFN27078_sa23_5),
	.B(FE_OCPN29489_sa23_3),
	.C(FE_OCPN29440_sa23_4));
   NAND2x1_ASAP7_75t_L U26184 (.Y(n20922),
	.A(FE_OCPN28112_n26664),
	.B(FE_OFN27056_n22995));
   NAND2x1p5_ASAP7_75t_SL U26185 (.Y(n26559),
	.A(n20922),
	.B(n20242));
   NOR2xp67_ASAP7_75t_L U26187 (.Y(n25095),
	.A(FE_OCPN27288_n25091),
	.B(FE_OCPN28266_n20920));
   NAND3xp33_ASAP7_75t_SL U26188 (.Y(n20907),
	.A(n20933),
	.B(n26664),
	.C(FE_OFN27078_sa23_5));
   NAND3xp33_ASAP7_75t_SL U26189 (.Y(n19329),
	.A(FE_OCPN29373_FE_OFN29191_sa23_2),
	.B(FE_OCPN27986_n18970),
	.C(n19313));
   NAND2xp33_ASAP7_75t_SL U26190 (.Y(n26558),
	.A(n25097),
	.B(n20934));
   NOR3xp33_ASAP7_75t_SRAM U26191 (.Y(n18979),
	.A(n25100),
	.B(n26559),
	.C(n26558));
   NOR2xp33_ASAP7_75t_SRAM U26193 (.Y(n18973),
	.A(FE_OFN27056_n22995),
	.B(n25093));
   NAND2xp33_ASAP7_75t_SRAM U26194 (.Y(n18977),
	.A(n18973),
	.B(n18974));
   NOR2xp33_ASAP7_75t_SRAM U26195 (.Y(n18975),
	.A(n19019),
	.B(n25093));
   NAND2xp33_ASAP7_75t_SRAM U26196 (.Y(n18976),
	.A(n18975),
	.B(n18974));
   NAND2x1_ASAP7_75t_SL U26198 (.Y(n22979),
	.A(FE_OCPN27627_sa23_1),
	.B(n18971));
   NOR2x1_ASAP7_75t_L U26199 (.Y(n19013),
	.A(n22980),
	.B(FE_OCPN28363_n22979));
   NOR2xp33_ASAP7_75t_SRAM U26200 (.Y(n18980),
	.A(FE_OFN16248_n20235),
	.B(n19013));
   OAI22xp33_ASAP7_75t_SL U26201 (.Y(n18985),
	.A1(FE_OCPN28363_n22979),
	.A2(FE_OCPN28071_n25092),
	.B1(FE_OFN25889_n20913),
	.B2(FE_OCPN28071_n25092));
   NOR2xp33_ASAP7_75t_SL U26202 (.Y(n20903),
	.A(n20241),
	.B(FE_OCPN28107_n23504));
   NOR2x1_ASAP7_75t_SL U26203 (.Y(n23490),
	.A(FE_OFN25883_n22945),
	.B(n25092));
   NAND3xp33_ASAP7_75t_SRAM U26204 (.Y(n18999),
	.A(n22943),
	.B(n23501),
	.C(n20257));
   NAND2xp5_ASAP7_75t_L U26205 (.Y(n26148),
	.A(n20907),
	.B(n22019));
   OAI22xp5_ASAP7_75t_SL U26206 (.Y(n26147),
	.A1(FE_OFN29001_n23491),
	.A2(FE_OCPN28086_n22034),
	.B1(FE_OCPN28112_n26664),
	.B2(FE_OCPN28086_n22034));
   NOR2xp33_ASAP7_75t_SL U26208 (.Y(n18992),
	.A(n19019),
	.B(n22033));
   NOR3x1_ASAP7_75t_L U26209 (.Y(n23473),
	.A(n22971),
	.B(FE_OCPN29441_sa23_4),
	.C(FE_OCPN27954_n22945));
   NOR2xp67_ASAP7_75t_L U26210 (.Y(n20909),
	.A(n22010),
	.B(FE_OCPN28363_n22979));
   NOR2x1_ASAP7_75t_L U26211 (.Y(n20916),
	.A(FE_OFN28562_n19342),
	.B(n26154));
   NAND2xp5_ASAP7_75t_R U26212 (.Y(n19001),
	.A(FE_OFN29026_n20911),
	.B(FE_OFN28752_n));
   NOR2x1_ASAP7_75t_SL U26213 (.Y(n19020),
	.A(n22004),
	.B(n22041));
   NAND2x1_ASAP7_75t_SL U26214 (.Y(n19321),
	.A(n25717),
	.B(n26556));
   NOR3x1_ASAP7_75t_SL U26215 (.Y(n23482),
	.A(n19321),
	.B(n23496),
	.C(n19013));
   NOR2x1_ASAP7_75t_SL U26216 (.Y(n22954),
	.A(n20260),
	.B(n26559));
   NOR2xp33_ASAP7_75t_L U26217 (.Y(n19002),
	.A(FE_OFN27078_sa23_5),
	.B(n22990));
   NAND3xp33_ASAP7_75t_SL U26218 (.Y(n19003),
	.A(n23482),
	.B(n22954),
	.C(n20943));
   OAI21xp33_ASAP7_75t_SL U26219 (.Y(n20901),
	.A1(FE_OFN29187_FE_OCPN27571_n20235),
	.A2(FE_OCPN28266_n20920),
	.B(n22006));
   NOR3xp33_ASAP7_75t_SL U26220 (.Y(n22975),
	.A(n19003),
	.B(FE_OFN26127_n22925),
	.C(n20901));
   NAND3xp33_ASAP7_75t_SL U26221 (.Y(n19004),
	.A(n22941),
	.B(n26163),
	.C(n22975));
   NAND3xp33_ASAP7_75t_SL U26222 (.Y(n20904),
	.A(FE_OCPN27986_n18970),
	.B(FE_OCPN28381_n26660),
	.C(FE_OCPN29374_FE_OFN29191_sa23_2));
   NOR3x1_ASAP7_75t_SL U26223 (.Y(n22051),
	.A(n19004),
	.B(n20224),
	.C(n23474));
   NOR3xp33_ASAP7_75t_SL U26224 (.Y(n19007),
	.A(n23499),
	.B(n23490),
	.C(n20942));
   NAND3xp33_ASAP7_75t_SL U26225 (.Y(n20899),
	.A(n18971),
	.B(FE_OCPN27727_n22964),
	.C(FE_OCPN29551_n));
   OAI22xp5_ASAP7_75t_L U26227 (.Y(n22987),
	.A1(FE_OCPN28112_n26664),
	.A2(n25093),
	.B1(n19313),
	.B2(n25093));
   NOR2xp33_ASAP7_75t_SRAM U26229 (.Y(n19294),
	.A(n20241),
	.B(FE_OCPN27288_n25091));
   NOR3xp33_ASAP7_75t_SL U26230 (.Y(n19014),
	.A(n20227),
	.B(n19294),
	.C(n20909));
   NOR2x1p5_ASAP7_75t_SL U26231 (.Y(n22935),
	.A(n22980),
	.B(FE_OCPN29488_FE_OFN25883_n22945));
   NOR2xp33_ASAP7_75t_SL U26232 (.Y(n22934),
	.A(FE_OFN29026_n20911),
	.B(n22935));
   NOR2xp33_ASAP7_75t_SRAM U26233 (.Y(n19024),
	.A(n25095),
	.B(n23473));
   AOI21x1_ASAP7_75t_R U26234 (.Y(n23002),
	.A1(FE_OFN28580_n23491),
	.A2(n19019),
	.B(n22926));
   NAND2xp5_ASAP7_75t_SL U26235 (.Y(n19022),
	.A(n23002),
	.B(n19020));
   NAND2xp5_ASAP7_75t_L U26236 (.Y(n20223),
	.A(FE_OCPN28112_n26664),
	.B(FE_OFN29001_n23491));
   NAND3xp33_ASAP7_75t_L U26237 (.Y(n19021),
	.A(n22941),
	.B(n23501),
	.C(n20223));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26238 (.Y(n19030),
	.A1(n26249),
	.A2(n19032),
	.B(FE_OCPN5105_n25099),
	.C(w1_11_));
   NOR2xp33_ASAP7_75t_SRAM U26239 (.Y(n19086),
	.A(sa30_6_),
	.B(n19060));
   NAND3xp33_ASAP7_75t_SRAM U26240 (.Y(n19034),
	.A(n19072),
	.B(FE_OCPN28241_n22142),
	.C(n19033));
   NAND3xp33_ASAP7_75t_R U26241 (.Y(n19041),
	.A(n19036),
	.B(n19035),
	.C(FE_OFN16326_n19058));
   NAND3xp33_ASAP7_75t_SL U26242 (.Y(n22143),
	.A(n20456),
	.B(n19043),
	.C(n19042));
   NOR2xp33_ASAP7_75t_SL U26243 (.Y(n19045),
	.A(n19044),
	.B(n25083));
   NAND3xp33_ASAP7_75t_SL U26244 (.Y(n19048),
	.A(n22145),
	.B(n22146),
	.C(n22136));
   NOR2x1_ASAP7_75t_L U26245 (.Y(n24030),
	.A(n22143),
	.B(n19048));
   NAND3xp33_ASAP7_75t_SL U26246 (.Y(n19050),
	.A(n19049),
	.B(FE_PSN8311_n25105),
	.C(n25113));
   OAI21xp33_ASAP7_75t_SRAM U26247 (.Y(n19073),
	.A1(FE_OFN25901_n22133),
	.A2(FE_PSN8270_n26027),
	.B(FE_OCPN28241_n22142));
   NOR3xp33_ASAP7_75t_L U26248 (.Y(n19055),
	.A(n19050),
	.B(FE_OCPN27764_n22152),
	.C(n19073));
   OAI21xp33_ASAP7_75t_SRAM U26249 (.Y(n19052),
	.A1(n20428),
	.A2(n19051),
	.B(n22633));
   NOR2xp33_ASAP7_75t_SRAM U26250 (.Y(n19053),
	.A(n26029),
	.B(n19052));
   NAND3xp33_ASAP7_75t_L U26251 (.Y(n19059),
	.A(n19055),
	.B(n19054),
	.C(n19053));
   NOR2xp33_ASAP7_75t_R U26252 (.Y(n19068),
	.A(FE_OCPN27829_n25102),
	.B(n19066));
   NOR2xp33_ASAP7_75t_SRAM U26253 (.Y(n19074),
	.A(n20450),
	.B(n22613));
   A2O1A1Ixp33_ASAP7_75t_L U26254 (.Y(n26685),
	.A1(n19083),
	.A2(n19082),
	.B(n24800),
	.C(n19081));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26255 (.Y(n19084),
	.A1(n19086),
	.A2(n26690),
	.B(FE_OCPN27753_n26685),
	.C(w1_6_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26256 (.Y(n275),
	.A1(n19086),
	.A2(n26690),
	.B(n19085),
	.C(n19084));
   NOR3xp33_ASAP7_75t_L U26257 (.Y(n19092),
	.A(n19089),
	.B(n19117),
	.C(n19088));
   NAND2xp5_ASAP7_75t_SL U26258 (.Y(n21163),
	.A(n19095),
	.B(n19094));
   OAI22xp5_ASAP7_75t_L U26259 (.Y(n19100),
	.A1(FE_OCPN27500_n19834),
	.A2(n24087),
	.B1(FE_OCPN28021_n21445),
	.B2(n24087));
   A2O1A1Ixp33_ASAP7_75t_SL U26260 (.Y(n19099),
	.A1(FE_OCPN27500_n19834),
	.A2(n19609),
	.B(n19818),
	.C(FE_OFN29172_sa00_4));
   NAND3xp33_ASAP7_75t_SL U26261 (.Y(n19102),
	.A(n19100),
	.B(FE_OFN28767_n26103),
	.C(n19099));
   NOR2xp33_ASAP7_75t_SRAM U26262 (.Y(n19108),
	.A(FE_OFN26146_n18774),
	.B(n19845));
   NAND3xp33_ASAP7_75t_R U26263 (.Y(n24526),
	.A(n19112),
	.B(n19132),
	.C(n19111));
   NOR2xp33_ASAP7_75t_L U26264 (.Y(n19120),
	.A(FE_OFN28835_n),
	.B(n19121));
   NOR2xp33_ASAP7_75t_L U26265 (.Y(n19124),
	.A(n19122),
	.B(n19121));
   NAND3xp33_ASAP7_75t_SRAM U26266 (.Y(n19130),
	.A(n19128),
	.B(n19127),
	.C(n19591));
   NOR2x1_ASAP7_75t_SL U26267 (.Y(n19133),
	.A(n21147),
	.B(FE_OFN28942_n21456));
   NOR2xp33_ASAP7_75t_SRAM U26270 (.Y(n19146),
	.A(n17254),
	.B(n19144));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26271 (.Y(n19159),
	.A1(n27127),
	.A2(FE_OCPN7622_n24526),
	.B(FE_OCPN27402_n24523),
	.C(w0_25_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26272 (.Y(n345),
	.A1(n27127),
	.A2(FE_OCPN7622_n24526),
	.B(n19160),
	.C(n19159));
   NOR2xp33_ASAP7_75t_R U26273 (.Y(n19163),
	.A(FE_OCPN28006_n17454),
	.B(FE_OCPN27313_n21845));
   NOR2xp33_ASAP7_75t_L U26274 (.Y(n19165),
	.A(FE_OFN28630_n23385),
	.B(n24544));
   NOR2xp33_ASAP7_75t_L U26275 (.Y(n19177),
	.A(FE_OFN29061_n22505),
	.B(n21817));
   NOR2xp33_ASAP7_75t_R U26276 (.Y(n23355),
	.A(FE_OCPN27625_sa11_5),
	.B(FE_OFN26554_n19170));
   NAND3xp33_ASAP7_75t_L U26277 (.Y(n19173),
	.A(n21815),
	.B(n19171),
	.C(FE_OFN28811_n19170));
   AND3x4_ASAP7_75t_SL U26278 (.Y(n19178),
	.A(n19176),
	.B(n19175),
	.C(n19174));
   NOR2xp33_ASAP7_75t_L U26279 (.Y(n19179),
	.A(FE_OCPN27562_n17447),
	.B(n21817));
   NAND2x1_ASAP7_75t_SL U26280 (.Y(n24560),
	.A(n19181),
	.B(n19180));
   NOR2xp33_ASAP7_75t_SRAM U26281 (.Y(n19182),
	.A(FE_OFN29061_n22505),
	.B(FE_PSN8304_n24565));
   NOR2xp33_ASAP7_75t_SRAM U26282 (.Y(n19184),
	.A(FE_OFN29171_n17510),
	.B(FE_PSN8304_n24565));
   NOR2xp33_ASAP7_75t_SL U26283 (.Y(n19187),
	.A(FE_OCPN27730_n17464),
	.B(n19217));
   NOR2xp33_ASAP7_75t_L U26284 (.Y(n19189),
	.A(FE_OFN29061_n22505),
	.B(n19217));
   NAND3xp33_ASAP7_75t_SRAM U26285 (.Y(n19196),
	.A(n25787),
	.B(n19195),
	.C(n24559));
   NOR3xp33_ASAP7_75t_SRAM U26286 (.Y(n19238),
	.A(n19196),
	.B(FE_PSN8302_n24562),
	.C(n24561));
   NOR3x1_ASAP7_75t_SL U26287 (.Y(n19197),
	.A(n25786),
	.B(n23375),
	.C(n23374));
   OAI21xp5_ASAP7_75t_SL U26288 (.Y(n23246),
	.A1(FE_OCPN27757_n21819),
	.A2(FE_OCPN28006_n17454),
	.B(n23378));
   O2A1O1Ixp33_ASAP7_75t_SRAM U26289 (.Y(n19205),
	.A1(n22505),
	.A2(n17453),
	.B(n21366),
	.C(n23267));
   NOR2xp33_ASAP7_75t_R U26290 (.Y(n19216),
	.A(FE_OFN29137_FE_OCPN27228_sa11_2),
	.B(n19217));
   NAND2x1_ASAP7_75t_SL U26291 (.Y(n21426),
	.A(n25795),
	.B(n24560));
   NOR2xp33_ASAP7_75t_R U26292 (.Y(n19219),
	.A(n21349),
	.B(n19217));
   INVxp67_ASAP7_75t_L U26293 (.Y(n19225),
	.A(n19224));
   NAND3xp33_ASAP7_75t_SL U26294 (.Y(n19236),
	.A(n19213),
	.B(n19235),
	.C(n23283));
   A2O1A1Ixp33_ASAP7_75t_R U26295 (.Y(n26802),
	.A1(n24560),
	.A2(n19238),
	.B(n26078),
	.C(n24569));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26296 (.Y(n19239),
	.A1(n23400),
	.A2(FE_OFN16395_n26801),
	.B(n26802),
	.C(FE_OFN49_w0_23));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26297 (.Y(n271),
	.A1(n23400),
	.A2(FE_OFN16395_n26801),
	.B(n19240),
	.C(n19239));
   NOR2xp33_ASAP7_75t_SRAM U26298 (.Y(n19241),
	.A(FE_OFN28844_FE_OCPN27570_n17791),
	.B(n20978));
   NOR2xp33_ASAP7_75t_R U26300 (.Y(n19243),
	.A(FE_PSN8313_FE_OCPN29469_n17747),
	.B(n20978));
   NOR2xp33_ASAP7_75t_SRAM U26301 (.Y(n19246),
	.A(FE_PSN8313_FE_OCPN29469_n17747),
	.B(n25210));
   OAI21xp5_ASAP7_75t_SL U26302 (.Y(n22063),
	.A1(FE_OCPN27919_n20155),
	.A2(FE_OCPN29533_n26971),
	.B(n22075));
   NAND3xp33_ASAP7_75t_SRAM U26303 (.Y(n19248),
	.A(FE_OCPN27566_FE_OFN16138_sa02_5),
	.B(FE_OCPN29546_n),
	.C(FE_OFN28730_FE_OCPN28416_sa02_3));
   A2O1A1Ixp33_ASAP7_75t_L U26304 (.Y(n19251),
	.A1(FE_OFN28704_FE_OCPN27740_sa02_4),
	.A2(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(FE_OCPN27566_FE_OFN16138_sa02_5),
	.C(n19250));
   NAND3xp33_ASAP7_75t_SL U26305 (.Y(n19252),
	.A(n20198),
	.B(n20954),
	.C(n19251));
   NOR3xp33_ASAP7_75t_SRAM U26306 (.Y(n19254),
	.A(n25212),
	.B(n25217),
	.C(n25211));
   NOR3xp33_ASAP7_75t_L U26307 (.Y(n25200),
	.A(n20135),
	.B(n20161),
	.C(n22894));
   NAND3xp33_ASAP7_75t_SRAM U26308 (.Y(n19260),
	.A(n25200),
	.B(n25206),
	.C(n25204));
   NOR3xp33_ASAP7_75t_SRAM U26309 (.Y(n19259),
	.A(n19272),
	.B(FE_OCPN27972_n20988),
	.C(n20981));
   NAND3xp33_ASAP7_75t_L U26310 (.Y(n19258),
	.A(n19257),
	.B(n22554),
	.C(n19256));
   NOR2xp33_ASAP7_75t_L U26311 (.Y(n19266),
	.A(n19264),
	.B(n22564));
   NAND3xp33_ASAP7_75t_SL U26312 (.Y(n25273),
	.A(n21004),
	.B(n19270),
	.C(n19269));
   NOR3xp33_ASAP7_75t_SL U26313 (.Y(n19273),
	.A(n22088),
	.B(n22899),
	.C(n19272));
   NAND2x1_ASAP7_75t_SL U26314 (.Y(n22064),
	.A(n19274),
	.B(n20955));
   OAI21xp33_ASAP7_75t_SL U26315 (.Y(n22563),
	.A1(FE_OCPN7645_n20962),
	.A2(FE_OCPN29545_n22529),
	.B(n22084));
   NOR3xp33_ASAP7_75t_L U26316 (.Y(n19278),
	.A(n19281),
	.B(n22064),
	.C(n22563));
   NOR2xp33_ASAP7_75t_R U26317 (.Y(n19277),
	.A(n22893),
	.B(n19276));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26318 (.Y(n19279),
	.A1(FE_OCPN29546_n),
	.A2(FE_OFN28730_FE_OCPN28416_sa02_3),
	.B(n22095),
	.C(FE_OCPN27566_FE_OFN16138_sa02_5));
   NOR3xp33_ASAP7_75t_SL U26319 (.Y(n19283),
	.A(n19282),
	.B(n21001),
	.C(n19281));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26321 (.Y(n19286),
	.A1(n27216),
	.A2(n25837),
	.B(n25834),
	.C(w2_30_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26322 (.Y(n284),
	.A1(n27216),
	.A2(n25837),
	.B(n19287),
	.C(n19286));
   INVx1_ASAP7_75t_R U26323 (.Y(n19289),
	.A(n23496));
   NAND2xp33_ASAP7_75t_SL U26324 (.Y(n19292),
	.A(n19288),
	.B(n19289));
   NOR2xp33_ASAP7_75t_R U26325 (.Y(n19290),
	.A(n19019),
	.B(n20931));
   NAND2xp33_ASAP7_75t_R U26326 (.Y(n19291),
	.A(n19290),
	.B(n19289));
   NAND3xp33_ASAP7_75t_SL U26327 (.Y(n20230),
	.A(FE_OFN27165_n),
	.B(n19325),
	.C(n26549));
   NAND2xp33_ASAP7_75t_SRAM U26328 (.Y(n19297),
	.A(n19296),
	.B(n22953));
   NAND3xp33_ASAP7_75t_SRAM U26329 (.Y(n19299),
	.A(n19298),
	.B(n20250),
	.C(n25097));
   NOR3xp33_ASAP7_75t_SRAM U26330 (.Y(n19300),
	.A(n24044),
	.B(n20230),
	.C(n19299));
   NOR2xp33_ASAP7_75t_SRAM U26331 (.Y(n19301),
	.A(n22980),
	.B(FE_OCPN27288_n25091));
   NAND2xp5_ASAP7_75t_SL U26332 (.Y(n22008),
	.A(FE_OCPN28098_n20907),
	.B(FE_OFN26557_n19302));
   A2O1A1Ixp33_ASAP7_75t_L U26333 (.Y(n22985),
	.A1(n20933),
	.A2(FE_OFN29026_n20911),
	.B(n20260),
	.C(FE_OCPN27482_sa23_5));
   NOR2x1_ASAP7_75t_SL U26334 (.Y(n19308),
	.A(n26149),
	.B(n20251));
   NAND2xp5_ASAP7_75t_L U26335 (.Y(n22030),
	.A(n19313),
	.B(n26664));
   NOR2xp33_ASAP7_75t_L U26336 (.Y(n19316),
	.A(n18971),
	.B(n22035));
   NAND2xp5_ASAP7_75t_SL U26337 (.Y(n20932),
	.A(n23511),
	.B(n20922));
   NOR2xp33_ASAP7_75t_SRAM U26338 (.Y(n19322),
	.A(n20928),
	.B(n19321));
   NAND3xp33_ASAP7_75t_SRAM U26339 (.Y(n19330),
	.A(n20242),
	.B(FE_OFN26557_n19302),
	.C(n19325));
   NOR2xp33_ASAP7_75t_SRAM U26340 (.Y(n19326),
	.A(FE_OFN29189_sa23_0),
	.B(n22951));
   NAND3xp33_ASAP7_75t_SRAM U26341 (.Y(n19328),
	.A(n19326),
	.B(FE_OCPN27727_n22964),
	.C(FE_OFN27126_sa23_3));
   NOR2xp33_ASAP7_75t_L U26342 (.Y(n19327),
	.A(FE_OCPN28071_n25092),
	.B(FE_OCPN28363_n22979));
   NAND3xp33_ASAP7_75t_R U26343 (.Y(n19340),
	.A(n26163),
	.B(FE_OCPN29548_n25717),
	.C(n20934));
   OAI22xp33_ASAP7_75t_L U26344 (.Y(n19338),
	.A1(n19019),
	.A2(n22935),
	.B1(n19000),
	.B2(n22935));
   NAND2xp33_ASAP7_75t_R U26345 (.Y(n19347),
	.A(n20237),
	.B(n19343));
   NOR2x1_ASAP7_75t_L U26346 (.Y(n19345),
	.A(n22976),
	.B(n22002));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26347 (.Y(n19356),
	.A1(n26249),
	.A2(n19358),
	.B(n19355),
	.C(w1_13_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26348 (.Y(n287),
	.A1(n26249),
	.A2(n19358),
	.B(n19357),
	.C(n19356));
   NOR2xp33_ASAP7_75t_SRAM U26349 (.Y(n19398),
	.A(FE_OFN128_sa13_7),
	.B(FE_OFN16389_n19359));
   NAND3xp33_ASAP7_75t_SRAM U26350 (.Y(n19397),
	.A(n25887),
	.B(n25561),
	.C(n25562));
   NOR3xp33_ASAP7_75t_SL U26351 (.Y(n25566),
	.A(n19375),
	.B(n19374),
	.C(n19373));
   NOR2xp33_ASAP7_75t_SRAM U26352 (.Y(n19377),
	.A(FE_OFN27186_sa13_4),
	.B(FE_OCPN29490_n17001));
   NOR3xp33_ASAP7_75t_SL U26353 (.Y(n19390),
	.A(n25282),
	.B(n19379),
	.C(n19405));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26354 (.Y(n19395),
	.A1(n19398),
	.A2(n19397),
	.B(n19394),
	.C(w2_23_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26355 (.Y(n310),
	.A1(n19398),
	.A2(n19397),
	.B(n19396),
	.C(n19395));
   NOR2xp33_ASAP7_75t_SRAM U26356 (.Y(n19400),
	.A(n19399),
	.B(n25990));
   NOR2xp33_ASAP7_75t_SRAM U26357 (.Y(n19401),
	.A(FE_OFN28801_n16978),
	.B(n25990));
   NOR3xp33_ASAP7_75t_SRAM U26358 (.Y(n19406),
	.A(FE_OCPN8210_n25287),
	.B(FE_OCPN28115_n25293),
	.C(n19404));
   NOR3xp33_ASAP7_75t_R U26359 (.Y(n25279),
	.A(n19409),
	.B(FE_OCPN27589_n25987),
	.C(n19408));
   NOR3xp33_ASAP7_75t_SL U26360 (.Y(n19412),
	.A(FE_OCPN29525_n18947),
	.B(n19411),
	.C(n19410));
   OAI22xp33_ASAP7_75t_SRAM U26361 (.Y(n25280),
	.A1(FE_OFN26170_n19361),
	.A2(n20529),
	.B1(FE_OFN16162_n25869),
	.B2(n20529));
   OAI222xp33_ASAP7_75t_SRAM U26362 (.Y(n19439),
	.A1(n25880),
	.A2(n27102),
	.B1(n19417),
	.B2(n27102),
	.C1(n25280),
	.C2(n27102));
   NOR2xp33_ASAP7_75t_SRAM U26363 (.Y(n19418),
	.A(FE_OCPN29510_n16996),
	.B(FE_OFN16220_n25219));
   NOR2xp33_ASAP7_75t_R U26364 (.Y(n19420),
	.A(FE_OFN16396_n25869),
	.B(FE_OFN16220_n25219));
   NAND2xp5_ASAP7_75t_SRAM U26365 (.Y(n19432),
	.A(n19431),
	.B(n20500));
   NOR3xp33_ASAP7_75t_SL U26366 (.Y(n19437),
	.A(n19433),
	.B(n20506),
	.C(n19432));
   NOR2xp33_ASAP7_75t_SRAM U26367 (.Y(n19436),
	.A(n19435),
	.B(n19434));
   OAI22xp5_ASAP7_75t_L U26368 (.Y(n23416),
	.A1(n21738),
	.A2(n21729),
	.B1(n21295),
	.B2(n21729));
   NOR2xp33_ASAP7_75t_R U26369 (.Y(n19451),
	.A(FE_OFN25986_n21012),
	.B(n21027));
   NOR2xp33_ASAP7_75t_R U26370 (.Y(n19453),
	.A(FE_OFN28589_n21048),
	.B(n21027));
   NOR2xp33_ASAP7_75t_SRAM U26371 (.Y(n19460),
	.A(n24440),
	.B(n24839));
   NAND3xp33_ASAP7_75t_SRAM U26372 (.Y(n19501),
	.A(n24835),
	.B(n19460),
	.C(n24834));
   NAND3xp33_ASAP7_75t_R U26373 (.Y(n19474),
	.A(n19463),
	.B(FE_OCPN8262_n21726),
	.C(n21280));
   NOR2xp33_ASAP7_75t_L U26374 (.Y(n19465),
	.A(n18045),
	.B(n21751));
   NOR2xp33_ASAP7_75t_R U26375 (.Y(n19467),
	.A(FE_OCPN27617_n18016),
	.B(n21751));
   NAND3x1_ASAP7_75t_SL U26376 (.Y(n23423),
	.A(n19472),
	.B(n19471),
	.C(n19470));
   NOR3xp33_ASAP7_75t_SRAM U26377 (.Y(n19476),
	.A(n21058),
	.B(n19475),
	.C(n21502));
   NOR3xp33_ASAP7_75t_SRAM U26378 (.Y(n19486),
	.A(n21043),
	.B(n21068),
	.C(FE_OCPN28431_n21734));
   NAND3xp33_ASAP7_75t_SL U26379 (.Y(n19491),
	.A(n19487),
	.B(n19486),
	.C(n19485));
   NOR2x1_ASAP7_75t_L U26380 (.Y(n23443),
	.A(FE_OCPN27998_n18019),
	.B(FE_OFN28588_n21048));
   NOR3x1_ASAP7_75t_SL U26381 (.Y(n19498),
	.A(n19497),
	.B(n19496),
	.C(n19495));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26382 (.Y(n19499),
	.A1(n26819),
	.A2(n19501),
	.B(n24837),
	.C(n26798));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26383 (.Y(n335),
	.A1(n26819),
	.A2(n19501),
	.B(n19500),
	.C(n19499));
   OAI21xp33_ASAP7_75t_L U26384 (.Y(n24052),
	.A1(FE_OFN25907_sa12_2),
	.A2(n19512),
	.B(n22251));
   NOR2xp33_ASAP7_75t_L U26385 (.Y(n19513),
	.A(n20591),
	.B(n24052));
   OAI22xp33_ASAP7_75t_L U26386 (.Y(n23608),
	.A1(n19546),
	.A2(n24370),
	.B1(n22745),
	.B2(n24370));
   NOR2xp33_ASAP7_75t_SRAM U26387 (.Y(n19519),
	.A(n22233),
	.B(n22781));
   NOR2x1_ASAP7_75t_SL U26388 (.Y(n23588),
	.A(FE_OFN25907_sa12_2),
	.B(n22722));
   OAI22xp33_ASAP7_75t_R U26389 (.Y(n19518),
	.A1(n23587),
	.A2(n23588),
	.B1(n23603),
	.B2(n23588));
   NOR2xp33_ASAP7_75t_R U26390 (.Y(n19521),
	.A(FE_OFN29075_n22745),
	.B(n22718));
   NOR2xp33_ASAP7_75t_L U26391 (.Y(n19530),
	.A(n20796),
	.B(n24055));
   NAND3xp33_ASAP7_75t_SL U26392 (.Y(n19535),
	.A(n19534),
	.B(n19540),
	.C(n20602));
   NOR3xp33_ASAP7_75t_L U26393 (.Y(n19544),
	.A(n19542),
	.B(n22719),
	.C(n25737));
   NAND2xp5_ASAP7_75t_SL U26394 (.Y(n22759),
	.A(n23587),
	.B(n24364));
   NOR2xp33_ASAP7_75t_SL U26395 (.Y(n19561),
	.A(n22726),
	.B(n20806));
   OAI21x1_ASAP7_75t_L U26396 (.Y(n23238),
	.A1(FE_OFN26158_n22224),
	.A2(FE_OCPN29324_n23216),
	.B(n19562));
   OAI22xp5_ASAP7_75t_L U26397 (.Y(n24586),
	.A1(FE_OCPN29477_sa12_5),
	.A2(n23238),
	.B1(n22724),
	.B2(n23238));
   O2A1O1Ixp5_ASAP7_75t_SL U26398 (.Y(n19568),
	.A1(n22247),
	.A2(n19567),
	.B(n26139),
	.C(n19566));
   OAI21x1_ASAP7_75t_SL U26399 (.Y(n25681),
	.A1(n19569),
	.A2(n26607),
	.B(n19568));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26400 (.Y(n19570),
	.A1(n25682),
	.A2(n25680),
	.B(n25681),
	.C(w1_19_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26401 (.Y(n400),
	.A1(n25682),
	.A2(n25680),
	.B(n19571),
	.C(n19570));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26402 (.Y(n19576),
	.A1(FE_OCPN28250_n19573),
	.A2(FE_OCPN27649_n17236),
	.B(FE_OCPN28270_n17237),
	.C(n19572));
   NOR2xp33_ASAP7_75t_SRAM U26403 (.Y(n19580),
	.A(FE_PSN8282_n21154),
	.B(n19578));
   NAND3xp33_ASAP7_75t_SL U26404 (.Y(n19587),
	.A(n21495),
	.B(n19583),
	.C(n19601));
   NAND3x1_ASAP7_75t_SL U26405 (.Y(n27126),
	.A(n19590),
	.B(n21441),
	.C(n19589));
   NAND3xp33_ASAP7_75t_SRAM U26406 (.Y(n19597),
	.A(n19595),
	.B(n19831),
	.C(n21155));
   NOR3xp33_ASAP7_75t_L U26407 (.Y(n19607),
	.A(n19606),
	.B(n19605),
	.C(n19604));
   OAI222xp33_ASAP7_75t_R U26408 (.Y(n21461),
	.A1(FE_OCPN27500_n19834),
	.A2(n26100),
	.B1(n19609),
	.B2(n26100),
	.C1(FE_OFN29172_sa00_4),
	.C2(n26100));
   A2O1A1Ixp33_ASAP7_75t_SL U26409 (.Y(n27123),
	.A1(n19621),
	.A2(n19620),
	.B(n26777),
	.C(n19619));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26410 (.Y(n19622),
	.A1(n27127),
	.A2(n27126),
	.B(n27122),
	.C(w0_28_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26411 (.Y(n295),
	.A1(n27127),
	.A2(n27126),
	.B(n19623),
	.C(n19622));
   A2O1A1Ixp33_ASAP7_75t_L U26412 (.Y(n19624),
	.A1(n16533),
	.A2(FE_OFN28832_n19789),
	.B(n23981),
	.C(n21886));
   NOR3xp33_ASAP7_75t_SL U26413 (.Y(n23956),
	.A(n19624),
	.B(n23139),
	.C(n24943));
   NOR2xp33_ASAP7_75t_SRAM U26414 (.Y(n19627),
	.A(FE_OCPN27900_n23949),
	.B(n19625));
   NAND3xp33_ASAP7_75t_SRAM U26416 (.Y(n19639),
	.A(n23956),
	.B(n23950),
	.C(n19628));
   NOR2xp33_ASAP7_75t_R U26417 (.Y(n19629),
	.A(n23980),
	.B(n23995));
   NOR2xp33_ASAP7_75t_SRAM U26418 (.Y(n19632),
	.A(n19630),
	.B(n23995));
   NOR3xp33_ASAP7_75t_L U26419 (.Y(n19643),
	.A(n19672),
	.B(n24958),
	.C(n23141));
   NAND3xp33_ASAP7_75t_L U26420 (.Y(n21891),
	.A(n23120),
	.B(n19644),
	.C(n19643));
   NOR3xp33_ASAP7_75t_SRAM U26421 (.Y(n19693),
	.A(n19645),
	.B(FE_OFN28586_n24736),
	.C(n21891));
   NOR2xp33_ASAP7_75t_SRAM U26422 (.Y(n19655),
	.A(FE_OFN28807_n24944),
	.B(n23995));
   NOR2xp33_ASAP7_75t_L U26423 (.Y(n19648),
	.A(n23980),
	.B(n21893));
   NOR2xp33_ASAP7_75t_L U26424 (.Y(n19650),
	.A(n16542),
	.B(n21893));
   AND3x1_ASAP7_75t_SL U26425 (.Y(n19656),
	.A(n21882),
	.B(n19654),
	.C(n19653));
   NOR2xp33_ASAP7_75t_SRAM U26426 (.Y(n19657),
	.A(FE_OCPN28157_n16534),
	.B(n23995));
   NOR2xp33_ASAP7_75t_SRAM U26427 (.Y(n19666),
	.A(n19661),
	.B(n23131));
   NAND3xp33_ASAP7_75t_SRAM U26428 (.Y(n19662),
	.A(n23035),
	.B(FE_OFN28912_n16534),
	.C(FE_OCPN28053_sa10_1));
   NAND3xp33_ASAP7_75t_R U26429 (.Y(n19675),
	.A(n19669),
	.B(n19668),
	.C(n23135));
   OAI222xp33_ASAP7_75t_SL U26430 (.Y(n19685),
	.A1(n23980),
	.A2(n21906),
	.B1(FE_OFN25959_n23011),
	.B2(n21906),
	.C1(FE_OFN27196_n),
	.C2(n21906));
   NOR2xp33_ASAP7_75t_L U26431 (.Y(n19678),
	.A(n16533),
	.B(n19677));
   NOR2xp33_ASAP7_75t_R U26432 (.Y(n19681),
	.A(FE_OFN28605_n23949),
	.B(n19678));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26433 (.Y(n19695),
	.A1(n26857),
	.A2(n19640),
	.B(FE_OCPN27478_n25011),
	.C(n25377));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26434 (.Y(n338),
	.A1(n26857),
	.A2(n19640),
	.B(n19696),
	.C(n19695));
   NAND3xp33_ASAP7_75t_L U26435 (.Y(n19702),
	.A(n24872),
	.B(n19697),
	.C(n22393));
   NOR3xp33_ASAP7_75t_SRAM U26436 (.Y(n19709),
	.A(n19702),
	.B(n19701),
	.C(n19950));
   OR2x2_ASAP7_75t_SRAM U26437 (.Y(n19708),
	.A(n19940),
	.B(n19703));
   NOR2xp33_ASAP7_75t_SRAM U26438 (.Y(n19706),
	.A(n17525),
	.B(n19703));
   NOR2xp33_ASAP7_75t_SRAM U26439 (.Y(n19711),
	.A(n17560),
	.B(n19712));
   NOR2xp33_ASAP7_75t_SRAM U26440 (.Y(n19715),
	.A(n19713),
	.B(n19712));
   NOR3xp33_ASAP7_75t_L U26441 (.Y(n19737),
	.A(n19729),
	.B(n20106),
	.C(n19728));
   O2A1O1Ixp5_ASAP7_75t_SL U26442 (.Y(n19749),
	.A1(n19748),
	.A2(n19747),
	.B(n22405),
	.C(n19746));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26443 (.Y(n19751),
	.A1(n25367),
	.A2(n25366),
	.B(FE_OFN29160_n25363),
	.C(FE_OFN16278_w3_5));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26444 (.Y(n285),
	.A1(n25367),
	.A2(n25366),
	.B(n19752),
	.C(n19751));
   NOR3xp33_ASAP7_75t_R U26445 (.Y(n19764),
	.A(n24892),
	.B(FE_OFN57_n19754),
	.C(FE_OFN29154_n19753));
   NOR3xp33_ASAP7_75t_SRAM U26446 (.Y(n19763),
	.A(n24895),
	.B(n24901),
	.C(n24894));
   NOR2xp33_ASAP7_75t_R U26447 (.Y(n19796),
	.A(n19787),
	.B(n19758));
   NOR2xp67_ASAP7_75t_SL U26448 (.Y(n19755),
	.A(n21893),
	.B(n21888));
   AND3x1_ASAP7_75t_SL U26449 (.Y(n19797),
	.A(n19769),
	.B(n19770),
	.C(n19755));
   AND3x1_ASAP7_75t_SRAM U26450 (.Y(n19759),
	.A(n19797),
	.B(n23126),
	.C(n21884));
   NOR2xp33_ASAP7_75t_R U26451 (.Y(n19798),
	.A(n23148),
	.B(n19758));
   NAND3xp33_ASAP7_75t_SRAM U26452 (.Y(n19773),
	.A(n19771),
	.B(n19770),
	.C(n19769));
   NOR2xp33_ASAP7_75t_R U26454 (.Y(n19790),
	.A(n19787),
	.B(n19791));
   OA21x2_ASAP7_75t_SRAM U26455 (.Y(n19792),
	.A1(n21902),
	.A2(FE_OFN28832_n19789),
	.B(n19788));
   NOR2xp33_ASAP7_75t_SRAM U26456 (.Y(n19793),
	.A(n16542),
	.B(n19791));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26457 (.Y(n19809),
	.A1(n26857),
	.A2(n24678),
	.B(FE_OCPN8243_n24899),
	.C(FE_OFN34_w3_22));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26458 (.Y(n291),
	.A1(n26857),
	.A2(n24678),
	.B(n19810),
	.C(n19809));
   NOR2xp33_ASAP7_75t_SRAM U26459 (.Y(n19814),
	.A(n26100),
	.B(FE_OFN28783_n26099));
   NAND3xp33_ASAP7_75t_SRAM U26460 (.Y(n19815),
	.A(FE_OFN30_n25256),
	.B(FE_OFN28767_n26103),
	.C(n19814));
   NOR2xp33_ASAP7_75t_R U26461 (.Y(n19820),
	.A(FE_OFN26146_n18774),
	.B(n24097));
   INVxp67_ASAP7_75t_L U26462 (.Y(n19819),
	.A(n19818));
   OR2x2_ASAP7_75t_SRAM U26463 (.Y(n19822),
	.A(FE_OCPN29284_n19821),
	.B(n24097));
   NAND3xp33_ASAP7_75t_L U26464 (.Y(n19830),
	.A(n19827),
	.B(n19826),
	.C(n19825));
   NOR3xp33_ASAP7_75t_SRAM U26465 (.Y(n19832),
	.A(n21438),
	.B(n21439),
	.C(FE_OCPN27703_n19847));
   NAND3xp33_ASAP7_75t_L U26466 (.Y(n19857),
	.A(n19833),
	.B(n19832),
	.C(n19831));
   NAND3xp33_ASAP7_75t_SRAM U26467 (.Y(n19837),
	.A(FE_OCPN27500_n19834),
	.B(n21166),
	.C(FE_OCPN29302_sa00_4));
   NAND3xp33_ASAP7_75t_L U26468 (.Y(n19838),
	.A(n19837),
	.B(FE_OCPN27843_n18750),
	.C(n19835));
   NOR3xp33_ASAP7_75t_SL U26469 (.Y(n19853),
	.A(n19846),
	.B(n19845),
	.C(n19844));
   A2O1A1Ixp33_ASAP7_75t_SL U26471 (.Y(n26113),
	.A1(n19860),
	.A2(n19859),
	.B(n21493),
	.C(n19858));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26472 (.Y(n19861),
	.A1(n27127),
	.A2(n24543),
	.B(FE_OCPN27314_n26113),
	.C(w0_24_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26473 (.Y(n351),
	.A1(n27127),
	.A2(n24543),
	.B(n19862),
	.C(n19861));
   NAND3xp33_ASAP7_75t_L U26474 (.Y(n24277),
	.A(n19864),
	.B(n23656),
	.C(n19863));
   NAND3xp33_ASAP7_75t_SL U26475 (.Y(n19866),
	.A(n20008),
	.B(n23626),
	.C(n19865));
   OAI21xp33_ASAP7_75t_L U26476 (.Y(n23657),
	.A1(FE_OFN28820_n),
	.A2(FE_OCPN27246_n22663),
	.B(n25350));
   NOR2xp33_ASAP7_75t_SRAM U26477 (.Y(n19904),
	.A(n25579),
	.B(n25581));
   NAND2x1_ASAP7_75t_SL U26478 (.Y(n20005),
	.A(n19872),
	.B(n24919));
   NAND2x1p5_ASAP7_75t_SL U26479 (.Y(n25580),
	.A(n19873),
	.B(n22667));
   NOR3xp33_ASAP7_75t_R U26482 (.Y(n19887),
	.A(n19885),
	.B(n22676),
	.C(n24881));
   NAND3xp33_ASAP7_75t_SRAM U26483 (.Y(n19898),
	.A(n19972),
	.B(n19889),
	.C(FE_OFN25968_n22668));
   O2A1O1Ixp5_ASAP7_75t_SL U26485 (.Y(n19902),
	.A1(FE_OCPN27629_n25589),
	.A2(n25588),
	.B(n26829),
	.C(n25574));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26487 (.Y(n19905),
	.A1(n25575),
	.A2(n25382),
	.B(FE_OFN28960_n25379),
	.C(w3_8_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26488 (.Y(n421),
	.A1(n25575),
	.A2(n25382),
	.B(n19906),
	.C(n19905));
   NOR2xp33_ASAP7_75t_SRAM U26489 (.Y(n19909),
	.A(FE_OCPN29524_n25029),
	.B(n19910));
   OAI22xp33_ASAP7_75t_SRAM U26490 (.Y(n19923),
	.A1(FE_OCPN28229_n17529),
	.A2(n19921),
	.B1(n22392),
	.B2(n19921));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26491 (.Y(n19933),
	.A1(FE_OCPN27499_FE_OFN16151_sa32_5),
	.A2(n17527),
	.B(n19932),
	.C(FE_OCPN28245_n));
   NAND3xp33_ASAP7_75t_SRAM U26492 (.Y(n19937),
	.A(n19934),
	.B(n24853),
	.C(n19933));
   NAND3xp33_ASAP7_75t_SRAM U26493 (.Y(n19942),
	.A(FE_OFN69_sa32_4),
	.B(n19940),
	.C(FE_OFN27148_sa32_3));
   O2A1O1Ixp33_ASAP7_75t_SL U26494 (.Y(n19961),
	.A1(FE_OFN16349_n19960),
	.A2(n19959),
	.B(n22405),
	.C(n19958));
   A2O1A1Ixp33_ASAP7_75t_SL U26495 (.Y(n26351),
	.A1(n20114),
	.A2(n19962),
	.B(n23899),
	.C(n19961));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26497 (.Y(n19963),
	.A1(n17580),
	.A2(n24830),
	.B(FE_OCPN27491_n26351),
	.C(FE_OFN25979_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26498 (.Y(n315),
	.A1(n17580),
	.A2(n24830),
	.B(n19964),
	.C(n19963));
   NOR2xp33_ASAP7_75t_L U26499 (.Y(n19966),
	.A(FE_OFN16267_sa21_4),
	.B(n23628));
   NOR2xp33_ASAP7_75t_R U26500 (.Y(n19965),
	.A(FE_OCPN8266_sa21_2),
	.B(n19966));
   NOR2xp33_ASAP7_75t_SRAM U26501 (.Y(n19969),
	.A(FE_OFN29044_n19967),
	.B(n19966));
   NOR3xp33_ASAP7_75t_L U26502 (.Y(n19976),
	.A(n22678),
	.B(FE_OCPN27553_n19975),
	.C(n22341));
   A2O1A1Ixp33_ASAP7_75t_SL U26503 (.Y(n20300),
	.A1(n19979),
	.A2(n16771),
	.B(FE_OCPN27508_n20339),
	.C(FE_OCPN27289_sa21_5));
   NOR2xp33_ASAP7_75t_SRAM U26504 (.Y(n19991),
	.A(FE_OFN168_n24268),
	.B(n24272));
   NOR3x1_ASAP7_75t_SL U26505 (.Y(n24921),
	.A(n19990),
	.B(n22676),
	.C(n22696));
   NOR2xp33_ASAP7_75t_SRAM U26506 (.Y(n19994),
	.A(n24256),
	.B(FE_OFN28920_n24254));
   NAND3xp33_ASAP7_75t_SRAM U26507 (.Y(n19995),
	.A(FE_OFN29215_n24262),
	.B(n24919),
	.C(n19994));
   AND3x1_ASAP7_75t_SRAM U26508 (.Y(n19997),
	.A(n20009),
	.B(n23656),
	.C(n20300));
   NOR2xp33_ASAP7_75t_R U26509 (.Y(n19998),
	.A(FE_OFN28981_n16767),
	.B(n25581));
   O2A1O1Ixp5_ASAP7_75t_SRAM U26510 (.Y(n20018),
	.A1(n24267),
	.A2(n24266),
	.B(n26829),
	.C(FE_OCPN7653_n24270));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26511 (.Y(n20020),
	.A1(n25575),
	.A2(n25475),
	.B(n25472),
	.C(FE_OCPN29427_w3_15));
   NOR2xp33_ASAP7_75t_SRAM U26512 (.Y(n20038),
	.A(n20050),
	.B(n21968));
   NOR3xp33_ASAP7_75t_SL U26513 (.Y(n20022),
	.A(n20840),
	.B(n20078),
	.C(n26290));
   OAI21xp5_ASAP7_75t_SL U26514 (.Y(n20024),
	.A1(FE_OCPN28061_n20076),
	.A2(n20853),
	.B(n20022));
   OAI21x1_ASAP7_75t_SL U26515 (.Y(n20056),
	.A1(n25317),
	.A2(FE_OFN29136_n),
	.B(n20083));
   NOR2xp33_ASAP7_75t_SL U26516 (.Y(n20030),
	.A(n20028),
	.B(n20027));
   NAND3xp33_ASAP7_75t_SL U26518 (.Y(n20036),
	.A(n20035),
	.B(n20034),
	.C(n20847));
   NOR3xp33_ASAP7_75t_SL U26519 (.Y(n20037),
	.A(n20036),
	.B(n21963),
	.C(n21964));
   NAND2x1_ASAP7_75t_SL U26520 (.Y(n21942),
	.A(n21984),
	.B(n20037));
   NOR3xp33_ASAP7_75t_SRAM U26521 (.Y(n20044),
	.A(n26401),
	.B(n20059),
	.C(n26402));
   NAND3xp33_ASAP7_75t_L U26522 (.Y(n20045),
	.A(n20044),
	.B(n26399),
	.C(n26406));
   NOR2xp33_ASAP7_75t_SRAM U26523 (.Y(n20058),
	.A(n20050),
	.B(n20059));
   NAND3xp33_ASAP7_75t_SRAM U26524 (.Y(n20057),
	.A(n20053),
	.B(n20052),
	.C(n20051));
   NOR2xp33_ASAP7_75t_SRAM U26525 (.Y(n20061),
	.A(n20060),
	.B(n20059));
   NAND3xp33_ASAP7_75t_SRAM U26526 (.Y(n20069),
	.A(n20066),
	.B(n21979),
	.C(n20882));
   NOR3xp33_ASAP7_75t_L U26527 (.Y(n20072),
	.A(n20069),
	.B(n20068),
	.C(n20067));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26528 (.Y(n20082),
	.A1(FE_OCPN28314_n20842),
	.A2(n20074),
	.B(FE_OCPN28008_n16290),
	.C(n20073));
   A2O1A1Ixp33_ASAP7_75t_L U26529 (.Y(n20085),
	.A1(n20084),
	.A2(n21932),
	.B(n26315),
	.C(FE_OCPN27780_n20083));
   O2A1O1Ixp5_ASAP7_75t_L U26530 (.Y(n20087),
	.A1(n27071),
	.A2(n20086),
	.B(n26942),
	.C(n20085));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26531 (.Y(n20090),
	.A1(n26407),
	.A2(n25510),
	.B(FE_OCPN8218_n25507),
	.C(w2_5_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26532 (.Y(n306),
	.A1(n26407),
	.A2(n25510),
	.B(n20091),
	.C(n20090));
   NAND3xp33_ASAP7_75t_SRAM U26533 (.Y(n20097),
	.A(n20094),
	.B(n20093),
	.C(n20092));
   NOR3xp33_ASAP7_75t_SRAM U26534 (.Y(n20099),
	.A(n20097),
	.B(n20096),
	.C(n20095));
   NAND3xp33_ASAP7_75t_L U26535 (.Y(n20101),
	.A(n20100),
	.B(n20099),
	.C(n20098));
   NAND3xp33_ASAP7_75t_R U26536 (.Y(n20110),
	.A(n20116),
	.B(n20109),
	.C(n20108));
   NOR3xp33_ASAP7_75t_L U26537 (.Y(n20115),
	.A(n20113),
	.B(n22370),
	.C(n20112));
   NAND3xp33_ASAP7_75t_R U26538 (.Y(n20119),
	.A(n22390),
	.B(n20117),
	.C(n22378));
   NOR3xp33_ASAP7_75t_SRAM U26539 (.Y(n20120),
	.A(n20119),
	.B(n20118),
	.C(n22369));
   NAND2xp33_ASAP7_75t_SRAM U26540 (.Y(n20126),
	.A(FE_OCPN29539_n24927),
	.B(FE_OFN25896_w3_4));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26541 (.Y(n20125),
	.A1(n22405),
	.A2(n24930),
	.B(FE_OCPN29538_n24927),
	.C(FE_OFN25899_w3_4));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26542 (.Y(n312),
	.A1(n22405),
	.A2(n24930),
	.B(n20126),
	.C(n20125));
   NOR2xp33_ASAP7_75t_R U26543 (.Y(n20996),
	.A(n20962),
	.B(FE_OCPN29545_n22529));
   NOR3xp33_ASAP7_75t_SRAM U26544 (.Y(n20128),
	.A(n25523),
	.B(n22872),
	.C(n22871));
   NAND3xp33_ASAP7_75t_SRAM U26545 (.Y(n20131),
	.A(n20128),
	.B(n20127),
	.C(n22059));
   NOR2xp33_ASAP7_75t_SRAM U26546 (.Y(n20146),
	.A(n20170),
	.B(n20144));
   NOR2xp33_ASAP7_75t_SRAM U26547 (.Y(n20149),
	.A(n17757),
	.B(n25296));
   NOR3xp33_ASAP7_75t_SL U26548 (.Y(n20154),
	.A(n22562),
	.B(n20194),
	.C(n22873));
   OAI21xp5_ASAP7_75t_SL U26549 (.Y(n20175),
	.A1(FE_OCPN27919_n20155),
	.A2(FE_OCPN27503_n20195),
	.B(n20154));
   OA21x2_ASAP7_75t_SRAM U26550 (.Y(n20157),
	.A1(FE_OCPN29545_n22529),
	.A2(FE_OCPN7645_n20962),
	.B(n22069));
   NAND3xp33_ASAP7_75t_SL U26551 (.Y(n20163),
	.A(n20955),
	.B(n20954),
	.C(n22070));
   A2O1A1Ixp33_ASAP7_75t_SL U26552 (.Y(n22112),
	.A1(FE_OFN108_n26971),
	.A2(FE_OCPN27634_n20169),
	.B(n20161),
	.C(FE_OFN26159_n22080));
   NOR3x1_ASAP7_75t_SL U26553 (.Y(n25299),
	.A(n20165),
	.B(n22561),
	.C(FE_OCPN27424_n22560));
   A2O1A1Ixp33_ASAP7_75t_L U26554 (.Y(n20171),
	.A1(n20170),
	.A2(FE_OCPN27634_n20169),
	.B(n20168),
	.C(FE_OFN26159_n22080));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26555 (.Y(n20184),
	.A1(n27216),
	.A2(n26494),
	.B(FE_OCPN28307_n26491),
	.C(w2_28_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26556 (.Y(n288),
	.A1(n27216),
	.A2(n26494),
	.B(n20185),
	.C(n20184));
   NOR3xp33_ASAP7_75t_L U26557 (.Y(n20188),
	.A(n25525),
	.B(n20186),
	.C(n20995));
   NOR3xp33_ASAP7_75t_SL U26558 (.Y(n20187),
	.A(n20994),
	.B(n22060),
	.C(n20194));
   NAND3xp33_ASAP7_75t_SRAM U26559 (.Y(n20192),
	.A(n17775),
	.B(n25302),
	.C(n25299));
   NOR3xp33_ASAP7_75t_SRAM U26560 (.Y(n20193),
	.A(n20192),
	.B(n25298),
	.C(n20191));
   A2O1A1Ixp33_ASAP7_75t_L U26561 (.Y(n22901),
	.A1(FE_OCPN27574_n20196),
	.A2(FE_OCPN27503_n20195),
	.B(FE_OCPN29545_n22529),
	.C(n22058));
   NOR2x1_ASAP7_75t_L U26562 (.Y(n22073),
	.A(n25912),
	.B(FE_OFN26033_n20197));
   NAND3xp33_ASAP7_75t_SL U26563 (.Y(n20199),
	.A(n20198),
	.B(n25914),
	.C(n22073));
   NAND3xp33_ASAP7_75t_SRAM U26564 (.Y(n20201),
	.A(n20200),
	.B(n22069),
	.C(n20969));
   NAND3xp33_ASAP7_75t_L U26565 (.Y(n20211),
	.A(n22534),
	.B(n22554),
	.C(n20210));
   O2A1O1Ixp33_ASAP7_75t_SRAM U26566 (.Y(n20217),
	.A1(n25310),
	.A2(n25309),
	.B(n27183),
	.C(n25626));
   A2O1A1Ixp33_ASAP7_75t_R U26567 (.Y(n20219),
	.A1(n25307),
	.A2(n25306),
	.B(n26976),
	.C(n20217));
   A2O1A1Ixp33_ASAP7_75t_R U26568 (.Y(n20220),
	.A1(n27216),
	.A2(n20222),
	.B(n20219),
	.C(w2_25_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26569 (.Y(n327),
	.A1(n27216),
	.A2(n20222),
	.B(n20221),
	.C(n20220));
   NAND2xp5_ASAP7_75t_SL U26570 (.Y(n22992),
	.A(n20223),
	.B(n22941));
   NOR3xp33_ASAP7_75t_SRAM U26571 (.Y(n24774),
	.A(FE_OCPN8241_n22041),
	.B(n20224),
	.C(n22992));
   O2A1O1Ixp5_ASAP7_75t_SRAM U26572 (.Y(n20225),
	.A1(FE_OFN28752_n),
	.A2(FE_OFN28787_n19000),
	.B(FE_OFN16248_n20235),
	.C(n22930));
   NAND3xp33_ASAP7_75t_L U26573 (.Y(n20229),
	.A(n24774),
	.B(n24775),
	.C(n20226));
   NAND3xp33_ASAP7_75t_R U26574 (.Y(n20236),
	.A(n22984),
	.B(n22038),
	.C(n20234));
   OAI21xp33_ASAP7_75t_R U26575 (.Y(n22929),
	.A1(FE_OFN29187_FE_OCPN27571_n20235),
	.A2(n22010),
	.B(FE_OCPN29548_n25717));
   NOR2xp33_ASAP7_75t_L U26576 (.Y(n20254),
	.A(n20240),
	.B(n20239));
   A2O1A1Ixp33_ASAP7_75t_L U26577 (.Y(n20248),
	.A1(n20241),
	.A2(n20920),
	.B(FE_OCPN28363_n22979),
	.C(n23002));
   NAND3xp33_ASAP7_75t_SL U26578 (.Y(n20252),
	.A(n25097),
	.B(n20250),
	.C(n20249));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26579 (.Y(n20267),
	.A1(n20256),
	.A2(FE_OCPN27743_n22009),
	.B(n20255),
	.C(FE_OFN27126_sa23_3));
   NAND3xp33_ASAP7_75t_R U26580 (.Y(n20271),
	.A(n26556),
	.B(n26162),
	.C(n26163));
   NOR2xp33_ASAP7_75t_SRAM U26581 (.Y(n20273),
	.A(FE_OFN16272_n24767),
	.B(n26149));
   NOR2xp33_ASAP7_75t_SRAM U26582 (.Y(n20275),
	.A(n18971),
	.B(n26149));
   A2O1A1Ixp33_ASAP7_75t_SL U26583 (.Y(n25695),
	.A1(FE_OFN26032_n20230),
	.A2(n20283),
	.B(n26571),
	.C(n20282));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26584 (.Y(n20284),
	.A1(FE_OFN16169_n26567),
	.A2(n20286),
	.B(FE_OCPN27507_n25695),
	.C(w1_8_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26585 (.Y(n387),
	.A1(FE_OFN16169_n26567),
	.A2(n20286),
	.B(n20285),
	.C(n20284));
   NOR2xp33_ASAP7_75t_SRAM U26586 (.Y(n20290),
	.A(FE_OCPN28299_n),
	.B(n22331));
   NOR2xp33_ASAP7_75t_L U26587 (.Y(n22344),
	.A(FE_OFN28820_n),
	.B(n20289));
   NOR2xp33_ASAP7_75t_SRAM U26588 (.Y(n20292),
	.A(FE_OCPN27690_n16757),
	.B(n22331));
   NAND3xp33_ASAP7_75t_SRAM U26589 (.Y(n20297),
	.A(n25350),
	.B(n25355),
	.C(FE_OCPN27774_n25351));
   NAND3xp33_ASAP7_75t_SL U26590 (.Y(n20302),
	.A(n20300),
	.B(n20299),
	.C(n20298));
   NOR2xp33_ASAP7_75t_SRAM U26591 (.Y(n20317),
	.A(FE_OCPN27616_n16760),
	.B(n20318));
   NOR2xp33_ASAP7_75t_L U26592 (.Y(n20316),
	.A(FE_OFN27163_n20304),
	.B(n22677));
   NOR2xp33_ASAP7_75t_SRAM U26593 (.Y(n20320),
	.A(FE_OCPN28298_n),
	.B(n20318));
   NAND3xp33_ASAP7_75t_SL U26594 (.Y(n20328),
	.A(n20327),
	.B(n20332),
	.C(n20326));
   NOR3xp33_ASAP7_75t_SL U26595 (.Y(n20330),
	.A(n20328),
	.B(n22679),
	.C(n25578));
   NAND3xp33_ASAP7_75t_SL U26596 (.Y(n20352),
	.A(n20331),
	.B(n20330),
	.C(n22352));
   NOR2xp33_ASAP7_75t_SRAM U26597 (.Y(n20338),
	.A(FE_OCPN27642_n16758),
	.B(FE_OCPN27508_n20339));
   NOR2xp33_ASAP7_75t_SRAM U26598 (.Y(n20341),
	.A(FE_OFN16447_n16749),
	.B(FE_OCPN27508_n20339));
   NOR2xp33_ASAP7_75t_R U26599 (.Y(n22682),
	.A(FE_OFN29023_n16750),
	.B(n20345));
   NOR2xp33_ASAP7_75t_R U26600 (.Y(n22681),
	.A(FE_OFN28981_n16767),
	.B(n20345));
   O2A1O1Ixp33_ASAP7_75t_SL U26601 (.Y(n20353),
	.A1(n22688),
	.A2(n20352),
	.B(n25575),
	.C(n20351));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26602 (.Y(n20356),
	.A1(n26829),
	.A2(n20358),
	.B(FE_OCPN29342_n25357),
	.C(FE_OFN26164_w3_13));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26603 (.Y(n307),
	.A1(n26829),
	.A2(n20358),
	.B(n20357),
	.C(n20356));
   NOR2xp33_ASAP7_75t_L U26604 (.Y(n20359),
	.A(n17329),
	.B(n20360));
   NOR2xp33_ASAP7_75t_L U26605 (.Y(n20362),
	.A(FE_OCPN29388_n22461),
	.B(n20360));
   NOR2xp33_ASAP7_75t_SRAM U26606 (.Y(n20379),
	.A(n26456),
	.B(n20380));
   NOR2xp33_ASAP7_75t_SL U26607 (.Y(n20370),
	.A(FE_OFN29254_n),
	.B(n21569));
   NAND3xp33_ASAP7_75t_SRAM U26608 (.Y(n20386),
	.A(n17326),
	.B(FE_OCPN29408_n22461),
	.C(FE_OFN26054_sa01_3));
   NOR2xp33_ASAP7_75t_R U26609 (.Y(n20390),
	.A(FE_OCPN29408_n22461),
	.B(FE_OCPN28301_n22448));
   NOR2xp33_ASAP7_75t_R U26610 (.Y(n20392),
	.A(n17382),
	.B(FE_OCPN28301_n22448));
   NOR3xp33_ASAP7_75t_SL U26611 (.Y(n20400),
	.A(n20399),
	.B(FE_OCPN8236_n22438),
	.C(n22216));
   NOR3xp33_ASAP7_75t_SL U26613 (.Y(n20402),
	.A(n23092),
	.B(n21560),
	.C(n20401));
   NAND3xp33_ASAP7_75t_SRAM U26614 (.Y(n20407),
	.A(n22422),
	.B(n22469),
	.C(n20402));
   NOR3xp33_ASAP7_75t_SL U26615 (.Y(n20403),
	.A(n21549),
	.B(FE_OCPN28301_n22448),
	.C(n22582));
   NAND2x1_ASAP7_75t_SL U26616 (.Y(n22463),
	.A(n25064),
	.B(n20403));
   NAND3x1_ASAP7_75t_SL U26617 (.Y(n22206),
	.A(n24389),
	.B(n20406),
	.C(n20405));
   NOR2xp33_ASAP7_75t_SRAM U26618 (.Y(n20408),
	.A(n26456),
	.B(n20409));
   NOR2xp33_ASAP7_75t_SRAM U26619 (.Y(n20411),
	.A(FE_OCPN27988_n26454),
	.B(n20409));
   NAND2x1p5_ASAP7_75t_SL U26620 (.Y(n26461),
	.A(n20415),
	.B(n25063));
   NOR3x1_ASAP7_75t_SL U26622 (.Y(n24138),
	.A(n25066),
	.B(n25071),
	.C(n20417));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26623 (.Y(n20418),
	.A1(n26282),
	.A2(n24142),
	.B(n24139),
	.C(w1_28_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26624 (.Y(n305),
	.A1(n26282),
	.A2(n24142),
	.B(n20419),
	.C(n20418));
   NOR2xp33_ASAP7_75t_SRAM U26625 (.Y(n20422),
	.A(FE_OFN28895_sa30_2),
	.B(n17603));
   NOR2xp33_ASAP7_75t_SRAM U26626 (.Y(n20424),
	.A(n20422),
	.B(n20421));
   NOR2xp33_ASAP7_75t_R U26627 (.Y(n20432),
	.A(n21602),
	.B(n20430));
   NOR2xp33_ASAP7_75t_R U26628 (.Y(n20444),
	.A(n21590),
	.B(n20438));
   NOR2xp33_ASAP7_75t_L U26629 (.Y(n20442),
	.A(n22624),
	.B(n20439));
   NAND3xp33_ASAP7_75t_L U26630 (.Y(n20445),
	.A(n24131),
	.B(n20444),
	.C(n25086));
   NOR2xp33_ASAP7_75t_SRAM U26632 (.Y(n20452),
	.A(n26028),
	.B(n20451));
   NOR2xp33_ASAP7_75t_SRAM U26633 (.Y(n20461),
	.A(n25108),
	.B(n22139));
   NOR2xp33_ASAP7_75t_SRAM U26634 (.Y(n20463),
	.A(FE_OCPN29467_n25102),
	.B(n22139));
   NAND3xp33_ASAP7_75t_R U26635 (.Y(n20482),
	.A(n21596),
	.B(n22621),
	.C(n20469));
   NAND3xp33_ASAP7_75t_SRAM U26636 (.Y(n20479),
	.A(n20478),
	.B(n20477),
	.C(n20476));
   NOR3xp33_ASAP7_75t_R U26637 (.Y(n20483),
	.A(n20482),
	.B(n20481),
	.C(FE_OFN28563_n20480));
   O2A1O1Ixp33_ASAP7_75t_SL U26638 (.Y(n20486),
	.A1(n25087),
	.A2(n20485),
	.B(n25081),
	.C(n20484));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26639 (.Y(n20488),
	.A1(FE_OFN16163_n26584),
	.A2(FE_OCPN7638_n26183),
	.B(n26180),
	.C(w1_1_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26640 (.Y(n348),
	.A1(FE_OFN16163_n26584),
	.A2(n26183),
	.B(n20489),
	.C(n20488));
   NOR3xp33_ASAP7_75t_L U26641 (.Y(n20493),
	.A(n25281),
	.B(FE_OCPN28189_n20491),
	.C(n20490));
   NAND2xp33_ASAP7_75t_L U26642 (.Y(n20503),
	.A(n20500),
	.B(n25222));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26643 (.Y(n20501),
	.A1(FE_OCPN8242_n20527),
	.A2(FE_OCPN27836_n16976),
	.B(FE_OFN28738_n16989),
	.C(n25286));
   NOR2xp33_ASAP7_75t_SRAM U26645 (.Y(n20512),
	.A(FE_OFN16319_n20527),
	.B(n20513));
   AND3x1_ASAP7_75t_SRAM U26646 (.Y(n20515),
	.A(FE_OFN26572_n19405),
	.B(n20510),
	.C(n20509));
   NOR2xp33_ASAP7_75t_SRAM U26647 (.Y(n20516),
	.A(FE_OCPN27902_n20514),
	.B(n20513));
   NOR3xp33_ASAP7_75t_SRAM U26648 (.Y(n20524),
	.A(n20523),
	.B(n20522),
	.C(n20521));
   NAND3xp33_ASAP7_75t_R U26649 (.Y(n20530),
	.A(n25551),
	.B(n20525),
	.C(n20524));
   NOR2xp33_ASAP7_75t_SRAM U26650 (.Y(n20528),
	.A(n20527),
	.B(FE_OCPN28204_n20526));
   NOR3x1_ASAP7_75t_SL U26651 (.Y(n26748),
	.A(n20536),
	.B(n20535),
	.C(n20534));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26652 (.Y(n20538),
	.A1(n26915),
	.A2(n26753),
	.B(FE_OFN28573_n26748),
	.C(w2_16_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26653 (.Y(n333),
	.A1(n26915),
	.A2(n26753),
	.B(n20539),
	.C(n20538));
   NOR3xp33_ASAP7_75t_SRAM U26654 (.Y(n24047),
	.A(n20540),
	.B(n23214),
	.C(n20591));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26655 (.Y(n20541),
	.A1(FE_OCPN29485_sa12_3),
	.A2(n17906),
	.B(n23587),
	.C(n22745));
   NAND3xp33_ASAP7_75t_L U26656 (.Y(n20551),
	.A(n20543),
	.B(n20542),
	.C(n20541));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26657 (.Y(n24048),
	.A1(n17906),
	.A2(FE_OCPN29559_n17900),
	.B(n20556),
	.C(FE_OCPN27429_sa12_3));
   NAND3xp33_ASAP7_75t_SRAM U26658 (.Y(n20612),
	.A(n24047),
	.B(n20553),
	.C(n24048));
   OAI22xp5_ASAP7_75t_L U26659 (.Y(n23234),
	.A1(n25741),
	.A2(n20556),
	.B1(FE_OFN29211_n23587),
	.B2(n20556));
   NOR3xp33_ASAP7_75t_SRAM U26660 (.Y(n20607),
	.A(n24053),
	.B(n24052),
	.C(FE_PSN8296_FE_OFN26588_n24062));
   OAI21xp33_ASAP7_75t_L U26661 (.Y(n22239),
	.A1(FE_OCPN27804_sa12_1),
	.A2(n22226),
	.B(n20561));
   NAND3xp33_ASAP7_75t_SL U26662 (.Y(n24381),
	.A(n23596),
	.B(n20565),
	.C(n20564));
   NOR2xp33_ASAP7_75t_SRAM U26663 (.Y(n20567),
	.A(FE_OCPN28386_n17899),
	.B(n24381));
   NOR2xp33_ASAP7_75t_SRAM U26664 (.Y(n20574),
	.A(FE_OCPN5137_n23600),
	.B(FE_OFN26556_n23236));
   OAI22xp33_ASAP7_75t_L U26665 (.Y(n20573),
	.A1(FE_OFN29211_n23587),
	.A2(n20571),
	.B1(n25741),
	.B2(n20571));
   NAND3xp33_ASAP7_75t_SL U26666 (.Y(n23225),
	.A(n20573),
	.B(n24592),
	.C(n20572));
   NOR2xp33_ASAP7_75t_SRAM U26667 (.Y(n20576),
	.A(n23603),
	.B(FE_OFN26556_n23236));
   AND3x1_ASAP7_75t_SRAM U26668 (.Y(n20580),
	.A(n23617),
	.B(n20595),
	.C(n20579));
   NOR3xp33_ASAP7_75t_SRAM U26669 (.Y(n20590),
	.A(n20583),
	.B(n22718),
	.C(n20784));
   NAND3xp33_ASAP7_75t_SRAM U26670 (.Y(n20601),
	.A(n20595),
	.B(n20594),
	.C(n23617));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26671 (.Y(n20610),
	.A1(n26139),
	.A2(n20612),
	.B(n20609),
	.C(w1_21_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26672 (.Y(n298),
	.A1(n26139),
	.A2(n20612),
	.B(n20611),
	.C(n20610));
   NOR2xp33_ASAP7_75t_SRAM U26673 (.Y(n20613),
	.A(FE_OFN28729_n20617),
	.B(n23840));
   NOR2xp33_ASAP7_75t_R U26674 (.Y(n20614),
	.A(n18583),
	.B(n23840));
   NOR2x1_ASAP7_75t_SL U26675 (.Y(n23806),
	.A(n23838),
	.B(n23711));
   NOR2xp33_ASAP7_75t_SRAM U26676 (.Y(n20625),
	.A(n20685),
	.B(n21193));
   NAND3xp33_ASAP7_75t_SL U26677 (.Y(n23853),
	.A(n21195),
	.B(n23869),
	.C(FE_OFN29150_sa20_5));
   NOR2xp33_ASAP7_75t_R U26678 (.Y(n20637),
	.A(FE_OFN27083_n),
	.B(n20678));
   NOR2xp33_ASAP7_75t_SRAM U26679 (.Y(n20639),
	.A(FE_OFN29112_FE_OCPN27870_n18527),
	.B(n20678));
   NOR2xp33_ASAP7_75t_SRAM U26680 (.Y(n20648),
	.A(FE_OFN28729_n20617),
	.B(n23763));
   OAI22xp33_ASAP7_75t_SRAM U26681 (.Y(n20647),
	.A1(FE_OFN28869_FE_OCPN27715_n23875),
	.A2(n23831),
	.B1(n18529),
	.B2(n23831));
   A2O1A1Ixp33_ASAP7_75t_R U26682 (.Y(n20659),
	.A1(n18521),
	.A2(n23869),
	.B(n23866),
	.C(FE_OFN29251_n18536));
   NOR2xp33_ASAP7_75t_SL U26683 (.Y(n20656),
	.A(FE_OFN28652_n21642),
	.B(n21658));
   NOR3xp33_ASAP7_75t_R U26684 (.Y(n20655),
	.A(n20654),
	.B(n20653),
	.C(n23792));
   NAND3xp33_ASAP7_75t_L U26685 (.Y(n20657),
	.A(n20656),
	.B(n23699),
	.C(n20655));
   OAI22xp33_ASAP7_75t_SRAM U26686 (.Y(n23870),
	.A1(FE_OFN28986_n18597),
	.A2(n23814),
	.B1(FE_OCPN27896_n18583),
	.B2(n23814));
   NOR2xp33_ASAP7_75t_SRAM U26687 (.Y(n20663),
	.A(n18583),
	.B(n23775));
   NOR2xp33_ASAP7_75t_L U26688 (.Y(n20671),
	.A(FE_OFN27083_n),
	.B(n20669));
   NAND3xp33_ASAP7_75t_L U26689 (.Y(n20675),
	.A(n23833),
	.B(n21665),
	.C(n20674));
   A2O1A1Ixp33_ASAP7_75t_L U26690 (.Y(n21683),
	.A1(FE_OFN29076_n18540),
	.A2(FE_OFN28776_n18532),
	.B(FE_OCPN28017_n18548),
	.C(FE_OCPN7660_FE_OFN28720_sa20_1));
   NAND3xp33_ASAP7_75t_L U26691 (.Y(n20692),
	.A(n23871),
	.B(n21239),
	.C(n21683));
   OAI21xp5_ASAP7_75t_L U26692 (.Y(n21650),
	.A1(FE_OFN28815_n18523),
	.A2(n21639),
	.B(FE_OCPN27591_n23742));
   NAND2xp5_ASAP7_75t_SL U26693 (.Y(n20684),
	.A(n20683),
	.B(n20682));
   NAND3x1_ASAP7_75t_SL U26694 (.Y(n26900),
	.A(n20684),
	.B(n23709),
	.C(n18579));
   NOR2xp33_ASAP7_75t_R U26695 (.Y(n20687),
	.A(FE_OFN28988_n18597),
	.B(n23792));
   NOR2x1_ASAP7_75t_L U26696 (.Y(n23829),
	.A(n20670),
	.B(n21639));
   NOR3x1_ASAP7_75t_L U26697 (.Y(n20690),
	.A(n21241),
	.B(FE_OCPN28432_n23829),
	.C(n23791));
   NAND3x1_ASAP7_75t_SL U26698 (.Y(n23885),
	.A(n20691),
	.B(n20690),
	.C(n23731));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26699 (.Y(n20700),
	.A1(FE_OFN16176_n27207),
	.A2(n26196),
	.B(FE_OCPN27583_n26193),
	.C(w2_12_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26700 (.Y(n292),
	.A1(FE_OFN16176_n27207),
	.A2(n26196),
	.B(n20701),
	.C(n20700));
   NAND3xp33_ASAP7_75t_SRAM U26701 (.Y(n20705),
	.A(n22311),
	.B(n23191),
	.C(n21126));
   NOR3xp33_ASAP7_75t_SRAM U26702 (.Y(n20704),
	.A(n23162),
	.B(FE_OFN29195_n22850),
	.C(FE_OCPN27933_n23328));
   NOR3xp33_ASAP7_75t_SRAM U26703 (.Y(n20713),
	.A(n20705),
	.B(n22305),
	.C(n21766));
   NOR2xp33_ASAP7_75t_R U26704 (.Y(n20708),
	.A(n18159),
	.B(n21764));
   NOR2xp33_ASAP7_75t_SRAM U26706 (.Y(n20715),
	.A(FE_PSN8320_n18176),
	.B(n22796));
   NOR2xp33_ASAP7_75t_SRAM U26707 (.Y(n20717),
	.A(FE_OCPN27722_n23336),
	.B(n22796));
   NAND3xp33_ASAP7_75t_SRAM U26708 (.Y(n20736),
	.A(n21105),
	.B(n23172),
	.C(n20759));
   NAND2xp5_ASAP7_75t_SL U26709 (.Y(n21133),
	.A(n18161),
	.B(n23315));
   NOR2xp33_ASAP7_75t_SL U26710 (.Y(n20728),
	.A(n23315),
	.B(n20726));
   NAND3xp33_ASAP7_75t_SL U26711 (.Y(n20734),
	.A(n20766),
	.B(FE_OCPN28016_n21124),
	.C(n20732));
   NOR2xp33_ASAP7_75t_SRAM U26712 (.Y(n20738),
	.A(n18159),
	.B(n23323));
   A2O1A1Ixp33_ASAP7_75t_L U26713 (.Y(n20737),
	.A1(FE_OCPN27719_n23306),
	.A2(n18178),
	.B(n20753),
	.C(n22295));
   NOR2xp33_ASAP7_75t_SRAM U26714 (.Y(n20741),
	.A(n20739),
	.B(n23323));
   NAND2x1_ASAP7_75t_SL U26715 (.Y(n22856),
	.A(n20745),
	.B(n22271));
   NAND2x1_ASAP7_75t_SL U26716 (.Y(n22852),
	.A(n20764),
	.B(n20763));
   NOR2xp33_ASAP7_75t_SRAM U26717 (.Y(n20767),
	.A(n23315),
	.B(FE_OFN29241_n22811));
   NOR2xp33_ASAP7_75t_SL U26718 (.Y(n20765),
	.A(n24694),
	.B(n22838));
   AND3x1_ASAP7_75t_SRAM U26719 (.Y(n20768),
	.A(n20766),
	.B(n22272),
	.C(n20765));
   NAND3xp33_ASAP7_75t_SRAM U26720 (.Y(n20775),
	.A(n22311),
	.B(n20773),
	.C(n20772));
   NOR3x1_ASAP7_75t_SL U26721 (.Y(n20774),
	.A(FE_OFN26009_n18213),
	.B(n23297),
	.C(n21130));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26722 (.Y(n20782),
	.A1(n27117),
	.A2(n27116),
	.B(FE_OFN29010_n27113),
	.C(w0_13_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26723 (.Y(n365),
	.A1(n27117),
	.A2(n27116),
	.B(n20783),
	.C(n20782));
   NOR2xp33_ASAP7_75t_SRAM U26724 (.Y(n20788),
	.A(n25439),
	.B(n25438));
   OAI21xp33_ASAP7_75t_SRAM U26725 (.Y(n20786),
	.A1(FE_OFN26125_n22742),
	.A2(n20796),
	.B(FE_OFN28834_FE_OCPN28371_n17900));
   NAND3xp33_ASAP7_75t_R U26726 (.Y(n25440),
	.A(n20786),
	.B(n20785),
	.C(n22225));
   NOR2xp33_ASAP7_75t_SRAM U26727 (.Y(n20787),
	.A(n26599),
	.B(n25440));
   NAND3xp33_ASAP7_75t_L U26728 (.Y(n20794),
	.A(n20791),
	.B(n20790),
	.C(n20789));
   NOR2xp33_ASAP7_75t_SRAM U26729 (.Y(n20798),
	.A(n20796),
	.B(n20799));
   AND2x2_ASAP7_75t_SL U26730 (.Y(n20800),
	.A(n20797),
	.B(n24056));
   NOR2xp33_ASAP7_75t_SRAM U26731 (.Y(n20801),
	.A(FE_OCPN29559_n17900),
	.B(n20799));
   NAND3xp33_ASAP7_75t_SL U26732 (.Y(n20811),
	.A(n22227),
	.B(n20805),
	.C(n20804));
   NOR3x1_ASAP7_75t_SL U26733 (.Y(n20823),
	.A(n20811),
	.B(n24589),
	.C(n20810));
   NAND3xp33_ASAP7_75t_SRAM U26734 (.Y(n20816),
	.A(n20812),
	.B(n22778),
	.C(n23609));
   OAI21xp33_ASAP7_75t_SRAM U26735 (.Y(n20820),
	.A1(FE_OCPN28346_n24051),
	.A2(n20826),
	.B(n25682));
   A2O1A1Ixp33_ASAP7_75t_L U26736 (.Y(n26597),
	.A1(n20824),
	.A2(n20823),
	.B(n24377),
	.C(n20820));
   A2O1A1Ixp33_ASAP7_75t_SL U26737 (.Y(n25443),
	.A1(n20828),
	.A2(n26594),
	.B(n26607),
	.C(n20827));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26738 (.Y(n20829),
	.A1(n26139),
	.A2(n20831),
	.B(FE_OCPN5116_n25443),
	.C(w1_16_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26739 (.Y(n407),
	.A1(n26139),
	.A2(n20831),
	.B(n20830),
	.C(n20829));
   OAI21xp33_ASAP7_75t_SRAM U26740 (.Y(n20834),
	.A1(n20853),
	.A2(n20854),
	.B(n20832));
   NOR3xp33_ASAP7_75t_L U26741 (.Y(n20835),
	.A(n20834),
	.B(n24184),
	.C(n20833));
   NOR2xp33_ASAP7_75t_SRAM U26742 (.Y(n20839),
	.A(n21963),
	.B(n25319));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26743 (.Y(n21966),
	.A1(n20868),
	.A2(n16300),
	.B(n20837),
	.C(FE_OFN26060_sa31_4));
   NAND3xp33_ASAP7_75t_R U26744 (.Y(n20844),
	.A(n20839),
	.B(n20838),
	.C(n21966));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26745 (.Y(n21992),
	.A1(FE_OFN28710_n20841),
	.A2(FE_OFN28753_sa31_2),
	.B(n20840),
	.C(n16295));
   NOR3xp33_ASAP7_75t_R U26746 (.Y(n20845),
	.A(n20844),
	.B(FE_OCPN27316_n25849),
	.C(n20843));
   NAND3xp33_ASAP7_75t_SRAM U26747 (.Y(n20852),
	.A(n20882),
	.B(n20856),
	.C(n20849));
   AND2x2_ASAP7_75t_SRAM U26748 (.Y(n20859),
	.A(n20855),
	.B(n20856));
   A2O1A1Ixp33_ASAP7_75t_SL U26750 (.Y(n26198),
	.A1(n20896),
	.A2(n20895),
	.B(n26315),
	.C(n20894));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26752 (.Y(n20897),
	.A1(n26942),
	.A2(n26201),
	.B(FE_OCPN8220_n26198),
	.C(w2_3_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26753 (.Y(n437),
	.A1(n26942),
	.A2(n26201),
	.B(n20898),
	.C(n20897));
   NAND3xp33_ASAP7_75t_L U26754 (.Y(n20902),
	.A(n20930),
	.B(n26160),
	.C(n26147));
   NOR2xp33_ASAP7_75t_SRAM U26755 (.Y(n20905),
	.A(n22048),
	.B(n23496));
   NAND3xp33_ASAP7_75t_SRAM U26756 (.Y(n20910),
	.A(n20905),
	.B(n20904),
	.C(n20924));
   NAND3xp33_ASAP7_75t_SRAM U26757 (.Y(n20908),
	.A(FE_OCPN28098_n20907),
	.B(FE_OFN26557_n19302),
	.C(n22987));
   NOR2xp33_ASAP7_75t_R U26758 (.Y(n26663),
	.A(n20911),
	.B(FE_OCPN27803_sa23_4));
   NAND3xp33_ASAP7_75t_L U26759 (.Y(n20918),
	.A(n20914),
	.B(n24216),
	.C(n20915));
   NOR2xp33_ASAP7_75t_R U26760 (.Y(n20936),
	.A(n23500),
	.B(n20931));
   NAND3xp33_ASAP7_75t_SL U26761 (.Y(n23479),
	.A(n20941),
	.B(n20940),
	.C(n23002));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26764 (.Y(n20950),
	.A1(n24038),
	.A2(n24037),
	.B(FE_OCPN27772_n24234),
	.C(w1_14_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26765 (.Y(n286),
	.A1(n24038),
	.A2(n24037),
	.B(n20951),
	.C(n20950));
   NAND3xp33_ASAP7_75t_SRAM U26766 (.Y(n20958),
	.A(n20953),
	.B(n22902),
	.C(n22107));
   NAND3xp33_ASAP7_75t_SRAM U26767 (.Y(n20956),
	.A(n20955),
	.B(n20954),
	.C(n22058));
   NOR2xp33_ASAP7_75t_SRAM U26768 (.Y(n20972),
	.A(FE_OCPN29546_n),
	.B(n20973));
   NOR2xp33_ASAP7_75t_SRAM U26769 (.Y(n20975),
	.A(FE_OCPN29469_n17747),
	.B(n20973));
   NOR2xp33_ASAP7_75t_SRAM U26770 (.Y(n20980),
	.A(n22060),
	.B(FE_OCPN27972_n20988));
   NOR2xp33_ASAP7_75t_SRAM U26771 (.Y(n20979),
	.A(n20978),
	.B(n25297));
   NAND3xp33_ASAP7_75t_R U26772 (.Y(n20984),
	.A(n20980),
	.B(n22534),
	.C(n20979));
   NOR3xp33_ASAP7_75t_SRAM U26773 (.Y(n21008),
	.A(n20984),
	.B(FE_OCPN28196_n22547),
	.C(n22109));
   OAI22xp33_ASAP7_75t_L U26774 (.Y(n20999),
	.A1(FE_OFN25998_n17781),
	.A2(n20994),
	.B1(FE_OCPN8230_n20993),
	.B2(n20994));
   NOR3xp33_ASAP7_75t_SL U26775 (.Y(n20998),
	.A(n20996),
	.B(n20995),
	.C(n22540));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26776 (.Y(n21010),
	.A1(n27216),
	.A2(n25860),
	.B(FE_OCPN7610_n25861),
	.C(w2_27_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26777 (.Y(n326),
	.A1(n27216),
	.A2(n25860),
	.B(n21011),
	.C(n21010));
   NOR2xp33_ASAP7_75t_R U26778 (.Y(n21016),
	.A(n21708),
	.B(n21017));
   NAND3xp33_ASAP7_75t_R U26779 (.Y(n21709),
	.A(FE_OCPN27617_n18016),
	.B(FE_OCPN28214_n21500),
	.C(FE_OFN29109_n));
   NOR2xp33_ASAP7_75t_L U26780 (.Y(n21030),
	.A(n23431),
	.B(n23443));
   OAI21xp33_ASAP7_75t_L U26782 (.Y(n21520),
	.A1(FE_OFN28948_n18011),
	.A2(FE_OFN26581_n21317),
	.B(n21035));
   NOR2xp33_ASAP7_75t_R U26783 (.Y(n21050),
	.A(FE_OFN29122_n),
	.B(n21051));
   NOR3xp33_ASAP7_75t_SRAM U26785 (.Y(n21527),
	.A(FE_OCPN27675_n17986),
	.B(FE_OCPN29314_n),
	.C(FE_OFN27125_n21057));
   NOR3xp33_ASAP7_75t_R U26786 (.Y(n21061),
	.A(n21527),
	.B(n21740),
	.C(n21058));
   NAND3xp33_ASAP7_75t_R U26787 (.Y(n21062),
	.A(n21061),
	.B(n21060),
	.C(n21059));
   NOR2xp33_ASAP7_75t_SRAM U26788 (.Y(n21073),
	.A(n18045),
	.B(n21066));
   NOR2xp33_ASAP7_75t_SRAM U26789 (.Y(n21072),
	.A(FE_OCPN27285_n18011),
	.B(n21066));
   AND3x2_ASAP7_75t_SL U26790 (.Y(n21742),
	.A(n21071),
	.B(n21070),
	.C(n21069));
   NAND2xp33_ASAP7_75t_SRAM U26792 (.Y(n21082),
	.A(FE_OFN16271_n26814),
	.B(n26355));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26793 (.Y(n21081),
	.A1(n26819),
	.A2(n26818),
	.B(n26815),
	.C(FE_OCPN28096_w3_31));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26794 (.Y(n301),
	.A1(n26819),
	.A2(n26818),
	.B(n21082),
	.C(n21081));
   NAND3xp33_ASAP7_75t_SRAM U26795 (.Y(n21083),
	.A(n22801),
	.B(FE_OCPN28016_n21124),
	.C(n21120));
   NOR3xp33_ASAP7_75t_SRAM U26796 (.Y(n21089),
	.A(n21083),
	.B(n21122),
	.C(n22309));
   INVxp33_ASAP7_75t_SRAM U26797 (.Y(n21086),
	.A(n21084));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26798 (.Y(n21087),
	.A1(n18166),
	.A2(n21086),
	.B(n18186),
	.C(n21085));
   NAND3xp33_ASAP7_75t_SL U26799 (.Y(n21092),
	.A(n21091),
	.B(FE_OCPN28016_n21124),
	.C(n20747));
   NOR2xp33_ASAP7_75t_L U26800 (.Y(n21100),
	.A(n23322),
	.B(n23323));
   NOR2xp33_ASAP7_75t_SRAM U26801 (.Y(n21106),
	.A(FE_OFN28798_FE_OCPN27947_n18177),
	.B(n21107));
   NOR3xp33_ASAP7_75t_SRAM U26802 (.Y(n21116),
	.A(n21115),
	.B(n21114),
	.C(FE_OFN16304_n22808));
   OAI22xp5_ASAP7_75t_L U26803 (.Y(n22797),
	.A1(n23315),
	.A2(n22278),
	.B1(n18177),
	.B2(n22278));
   NAND3xp33_ASAP7_75t_SL U26804 (.Y(n21128),
	.A(n21127),
	.B(n21126),
	.C(n23324));
   NOR2x1_ASAP7_75t_SL U26805 (.Y(n23340),
	.A(n23168),
	.B(n21128));
   NAND3xp33_ASAP7_75t_SL U26806 (.Y(n21131),
	.A(n22797),
	.B(n23340),
	.C(n22819));
   NAND3x1_ASAP7_75t_SL U26807 (.Y(n23194),
	.A(n21133),
	.B(n23325),
	.C(n21132));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26809 (.Y(n21145),
	.A1(n27117),
	.A2(FE_PSN8331_n24113),
	.B(n24114),
	.C(FE_OFN43_w0_10));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26810 (.Y(n366),
	.A1(n27117),
	.A2(FE_PSN8331_n24113),
	.B(n21146),
	.C(n21145));
   NOR2xp33_ASAP7_75t_SL U26811 (.Y(n21149),
	.A(n24348),
	.B(n24344));
   A2O1A1Ixp33_ASAP7_75t_R U26812 (.Y(n21451),
	.A1(FE_OCPN29542_n21151),
	.A2(n21154),
	.B(n21150),
	.C(FE_OCPN29396_n19149));
   NAND3xp33_ASAP7_75t_SRAM U26813 (.Y(n21161),
	.A(n21157),
	.B(n21156),
	.C(n21155));
   NOR2xp33_ASAP7_75t_R U26814 (.Y(n21169),
	.A(n21166),
	.B(n21444));
   AND2x2_ASAP7_75t_L U26815 (.Y(n21170),
	.A(n21168),
	.B(n21167));
   NOR2xp33_ASAP7_75t_SRAM U26816 (.Y(n21171),
	.A(n12998),
	.B(n21444));
   O2A1O1Ixp33_ASAP7_75t_SL U26817 (.Y(n21187),
	.A1(n21186),
	.A2(n21185),
	.B(n27127),
	.C(n21184));
   A2O1A1Ixp33_ASAP7_75t_SL U26818 (.Y(n26633),
	.A1(n21189),
	.A2(n21188),
	.B(n26777),
	.C(n21187));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26820 (.Y(n21190),
	.A1(FE_OFN16170_n26637),
	.A2(n26636),
	.B(FE_OCPN7662_n26633),
	.C(w0_29_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26821 (.Y(n321),
	.A1(FE_OFN16170_n26637),
	.A2(n26636),
	.B(n21191),
	.C(n21190));
   O2A1O1Ixp33_ASAP7_75t_R U26822 (.Y(n21194),
	.A1(n21669),
	.A2(n20617),
	.B(FE_OCPN27715_n23875),
	.C(n21192));
   NOR2xp33_ASAP7_75t_SL U26824 (.Y(n21199),
	.A(FE_OFN28986_n18597),
	.B(n23864));
   NOR2xp33_ASAP7_75t_R U26825 (.Y(n21198),
	.A(FE_OFN29140_n18527),
	.B(n23864));
   NAND3xp33_ASAP7_75t_SRAM U26826 (.Y(n21196),
	.A(FE_OFN29178_sa20_4),
	.B(n23869),
	.C(FE_OFN29251_n18536));
   OA21x2_ASAP7_75t_L U26827 (.Y(n21201),
	.A1(n21199),
	.A2(n21198),
	.B(n21197));
   NAND3xp33_ASAP7_75t_SL U26828 (.Y(n25905),
	.A(n23800),
	.B(n21201),
	.C(n21200));
   NOR3xp33_ASAP7_75t_SRAM U26829 (.Y(n21207),
	.A(n21203),
	.B(FE_OFN16301_n25905),
	.C(n21202));
   NAND3xp33_ASAP7_75t_SRAM U26830 (.Y(n21267),
	.A(n25902),
	.B(n21207),
	.C(n25899));
   NOR2xp33_ASAP7_75t_R U26831 (.Y(n21210),
	.A(FE_OFN16295_n23837),
	.B(FE_OFN27088_n23754));
   NAND3xp33_ASAP7_75t_SL U26832 (.Y(n21208),
	.A(n21665),
	.B(n21637),
	.C(n25328));
   NOR2xp33_ASAP7_75t_SRAM U26833 (.Y(n21212),
	.A(n18532),
	.B(FE_OFN27088_n23754));
   NAND2xp5_ASAP7_75t_L U26834 (.Y(n21636),
	.A(n21221),
	.B(n21220));
   NAND3xp33_ASAP7_75t_R U26835 (.Y(n21236),
	.A(n21235),
	.B(FE_OFN16221_n21234),
	.C(n23777));
   INVxp33_ASAP7_75t_L U26836 (.Y(n21242),
	.A(FE_OFN29112_FE_OCPN27870_n18527));
   NOR2xp33_ASAP7_75t_SL U26837 (.Y(n21243),
	.A(FE_OFN28729_n20617),
	.B(n23739));
   O2A1O1Ixp5_ASAP7_75t_SRAM U26838 (.Y(n21254),
	.A1(n21669),
	.A2(n18529),
	.B(FE_OFN29076_n18540),
	.C(FE_OFN26150_n21253));
   O2A1O1Ixp5_ASAP7_75t_SL U26839 (.Y(n21262),
	.A1(n21698),
	.A2(n21261),
	.B(n27207),
	.C(n21260));
   OAI21xp5_ASAP7_75t_SL U26840 (.Y(n25921),
	.A1(n21263),
	.A2(n26517),
	.B(n21262));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26842 (.Y(n21265),
	.A1(n26323),
	.A2(n21267),
	.B(FE_OCPN27522_n25921),
	.C(w2_8_));
   NAND3xp33_ASAP7_75t_L U26843 (.Y(n21274),
	.A(n21271),
	.B(n23419),
	.C(n21270));
   NOR3xp33_ASAP7_75t_R U26844 (.Y(n21281),
	.A(n21279),
	.B(n21524),
	.C(n21278));
   NOR2xp33_ASAP7_75t_SRAM U26845 (.Y(n21303),
	.A(n21295),
	.B(n17989));
   A2O1A1Ixp33_ASAP7_75t_R U26846 (.Y(n21300),
	.A1(n21708),
	.A2(FE_OFN21730_sa03_3),
	.B(n21296),
	.C(n21327));
   NOR3x1_ASAP7_75t_L U26847 (.Y(n24245),
	.A(n21302),
	.B(FE_OCPN7584_n23447),
	.C(n21301));
   NOR2xp33_ASAP7_75t_SRAM U26848 (.Y(n21305),
	.A(n21304),
	.B(n17989));
   NOR2xp33_ASAP7_75t_SRAM U26849 (.Y(n21312),
	.A(FE_OCPN28001_n21310),
	.B(n18008));
   NOR2xp33_ASAP7_75t_SRAM U26850 (.Y(n21326),
	.A(FE_OCPN4680_n21317),
	.B(FE_OCPN27628_n23455));
   A2O1A1Ixp33_ASAP7_75t_L U26851 (.Y(n21325),
	.A1(FE_OCPN29283_n23439),
	.A2(n17996),
	.B(FE_OCPN27675_n17986),
	.C(n21324));
   NOR3x1_ASAP7_75t_SL U26852 (.Y(n25946),
	.A(n21337),
	.B(n21336),
	.C(n21335));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26853 (.Y(n21338),
	.A1(n26819),
	.A2(FE_OCPN8227_n25950),
	.B(n25947),
	.C(FE_OFN28452_w3_29));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26854 (.Y(n316),
	.A1(n26819),
	.A2(FE_OCPN8227_n25950),
	.B(n21339),
	.C(n21338));
   NOR2xp33_ASAP7_75t_SRAM U26855 (.Y(n26066),
	.A(n21365),
	.B(n22501));
   NAND2xp33_ASAP7_75t_SRAM U26856 (.Y(n21343),
	.A(n26066),
	.B(n26065));
   NAND2xp33_ASAP7_75t_SRAM U26858 (.Y(n21342),
	.A(n26068),
	.B(n26065));
   NOR2xp33_ASAP7_75t_L U26859 (.Y(n21345),
	.A(n21344),
	.B(n21406));
   NAND3xp33_ASAP7_75t_SRAM U26860 (.Y(n21347),
	.A(n24710),
	.B(n26064),
	.C(n26073));
   NOR2xp33_ASAP7_75t_SRAM U26861 (.Y(n21348),
	.A(n26076),
	.B(n21347));
   NAND3xp33_ASAP7_75t_SL U26862 (.Y(n21350),
	.A(n21362),
	.B(n21411),
	.C(n21847));
   NOR2xp33_ASAP7_75t_SRAM U26863 (.Y(n21357),
	.A(n22501),
	.B(n22500));
   OAI22xp5_ASAP7_75t_SL U26864 (.Y(n23389),
	.A1(n17445),
	.A2(n21860),
	.B1(FE_OCPN27730_n17464),
	.B2(n21860));
   NAND3xp33_ASAP7_75t_R U26865 (.Y(n21361),
	.A(n21357),
	.B(n22510),
	.C(n23389));
   NOR2xp33_ASAP7_75t_SRAM U26866 (.Y(n23258),
	.A(n21358),
	.B(n21395));
   NAND3xp33_ASAP7_75t_R U26867 (.Y(n21359),
	.A(n23378),
	.B(FE_OCPN27605_n23357),
	.C(n23258));
   NAND2x1_ASAP7_75t_L U26868 (.Y(n23383),
	.A(n22487),
	.B(n21362));
   NOR3xp33_ASAP7_75t_L U26869 (.Y(n21370),
	.A(n17477),
	.B(n23394),
	.C(n21368));
   NAND3xp33_ASAP7_75t_L U26870 (.Y(n21386),
	.A(n21375),
	.B(n23380),
	.C(n23365));
   NOR2xp33_ASAP7_75t_SRAM U26871 (.Y(n21376),
	.A(n17447),
	.B(n21377));
   NOR2xp33_ASAP7_75t_SRAM U26872 (.Y(n21379),
	.A(n22505),
	.B(n21377));
   NAND3xp33_ASAP7_75t_SL U26873 (.Y(n21842),
	.A(n21384),
	.B(n21383),
	.C(n21382));
   O2A1O1Ixp33_ASAP7_75t_SL U26874 (.Y(n21388),
	.A1(n21417),
	.A2(n26083),
	.B(n26082),
	.C(n26074));
   A2O1A1Ixp33_ASAP7_75t_L U26875 (.Y(n24713),
	.A1(n26080),
	.A2(n26079),
	.B(n26078),
	.C(n21388));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26876 (.Y(n21389),
	.A1(n27062),
	.A2(n21391),
	.B(n24713),
	.C(FE_OFN40_w0_19));
   OAI22xp33_ASAP7_75t_SL U26877 (.Y(n21855),
	.A1(FE_OCPN29513_n17447),
	.A2(n25786),
	.B1(FE_OCPN29435_n17445),
	.B2(n25786));
   NAND3xp33_ASAP7_75t_SRAM U26878 (.Y(n21402),
	.A(n25792),
	.B(n21855),
	.C(n25787));
   NAND3xp33_ASAP7_75t_SRAM U26879 (.Y(n21399),
	.A(n21394),
	.B(n23390),
	.C(n21393));
   NOR3xp33_ASAP7_75t_SL U26880 (.Y(n21397),
	.A(n22504),
	.B(FE_OCPN27584_n22497),
	.C(FE_OCPN27496_n21820));
   NOR2xp33_ASAP7_75t_SRAM U26881 (.Y(n21405),
	.A(FE_OCPN5021_n17446),
	.B(n21406));
   NOR2xp33_ASAP7_75t_SRAM U26882 (.Y(n21407),
	.A(n19162),
	.B(n21406));
   NAND3xp33_ASAP7_75t_R U26883 (.Y(n21432),
	.A(FE_OFN65_n21412),
	.B(n21411),
	.C(n21410));
   NOR3xp33_ASAP7_75t_R U26884 (.Y(n21424),
	.A(FE_OFN29041_n21415),
	.B(n23267),
	.C(n21854));
   NAND3xp33_ASAP7_75t_SRAM U26885 (.Y(n21427),
	.A(n24567),
	.B(n23372),
	.C(n21425));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26886 (.Y(n21436),
	.A1(n27062),
	.A2(n26372),
	.B(FE_OCPN27357_n26369),
	.C(w0_20_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26887 (.Y(n357),
	.A1(n27062),
	.A2(n26372),
	.B(n21437),
	.C(n21436));
   NOR2xp33_ASAP7_75t_SRAM U26888 (.Y(n21443),
	.A(FE_OCPN27819_n17245),
	.B(n21444));
   NOR2xp33_ASAP7_75t_SRAM U26889 (.Y(n21440),
	.A(FE_PSN8290_n21439),
	.B(n21438));
   NAND3xp33_ASAP7_75t_R U26890 (.Y(n24474),
	.A(n21442),
	.B(n21441),
	.C(n21440));
   NAND2xp33_ASAP7_75t_SRAM U26891 (.Y(n21449),
	.A(n21443),
	.B(n21446));
   NOR2xp33_ASAP7_75t_SRAM U26892 (.Y(n21447),
	.A(FE_OCPN28021_n21445),
	.B(n21444));
   NAND2xp33_ASAP7_75t_SRAM U26893 (.Y(n21448),
	.A(n21447),
	.B(n21446));
   NOR2xp33_ASAP7_75t_SRAM U26894 (.Y(n21458),
	.A(FE_OFN28942_n21456),
	.B(n21455));
   NAND3xp33_ASAP7_75t_SRAM U26895 (.Y(n21499),
	.A(n21460),
	.B(n21459),
	.C(FE_OFN27069_n24478));
   NAND3xp33_ASAP7_75t_SRAM U26896 (.Y(n21466),
	.A(n21463),
	.B(FE_OFN28534_n21462),
	.C(n21461));
   NAND2xp33_ASAP7_75t_SRAM U26897 (.Y(n21469),
	.A(n21468),
	.B(n21467));
   NOR3xp33_ASAP7_75t_SRAM U26898 (.Y(n21471),
	.A(n21469),
	.B(n17297),
	.C(FE_OFN28556_n24516));
   NOR2xp33_ASAP7_75t_SRAM U26899 (.Y(n21480),
	.A(FE_OCPN28389_n21479),
	.B(FE_PSN8273_n24087));
   NOR2xp33_ASAP7_75t_SRAM U26900 (.Y(n21483),
	.A(FE_OFN16216_n19573),
	.B(n24087));
   O2A1O1Ixp33_ASAP7_75t_L U26901 (.Y(n21492),
	.A1(FE_OFN28566_n21491),
	.A2(n21490),
	.B(n27127),
	.C(n21489));
   A2O1A1Ixp33_ASAP7_75t_SL U26902 (.Y(n26535),
	.A1(n21495),
	.A2(n21494),
	.B(n21493),
	.C(n21492));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26903 (.Y(n21497),
	.A1(FE_OFN16170_n26637),
	.A2(n21499),
	.B(n26535),
	.C(w0_30_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26904 (.Y(n322),
	.A1(FE_OFN16170_n26637),
	.A2(n21499),
	.B(n21498),
	.C(n21497));
   NOR3xp33_ASAP7_75t_SRAM U26905 (.Y(n21501),
	.A(FE_OFN28956_n18011),
	.B(FE_OFN29109_n),
	.C(FE_OCPN28214_n21500));
   NOR3xp33_ASAP7_75t_SL U26906 (.Y(n24247),
	.A(n21503),
	.B(n21502),
	.C(n21501));
   NOR3xp33_ASAP7_75t_SRAM U26907 (.Y(n21517),
	.A(n21509),
	.B(n21747),
	.C(n21728));
   A2O1A1Ixp33_ASAP7_75t_L U26908 (.Y(n21514),
	.A1(FE_OCPN28184_n18020),
	.A2(FE_OCPN27948_FE_OFN26173_n21511),
	.B(FE_OCPN27998_n18019),
	.C(n21510));
   NOR3xp33_ASAP7_75t_SL U26909 (.Y(n21516),
	.A(n21514),
	.B(n21513),
	.C(n23423));
   OAI22xp33_ASAP7_75t_SRAM U26911 (.Y(n21519),
	.A1(FE_OFN27133_n21725),
	.A2(FE_OFN28677_n17998),
	.B1(n17996),
	.B2(FE_OFN28677_n17998));
   NOR3xp33_ASAP7_75t_SL U26912 (.Y(n21522),
	.A(n21520),
	.B(n21519),
	.C(n21518));
   NOR3xp33_ASAP7_75t_L U26913 (.Y(n21530),
	.A(n21528),
	.B(n23425),
	.C(n21527));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26915 (.Y(n21532),
	.A1(n26819),
	.A2(n24844),
	.B(FE_OFN28578_FE_OFN16316_n24840),
	.C(FE_OCPN27664_w3_25));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26916 (.Y(n336),
	.A1(n26819),
	.A2(n24844),
	.B(n21533),
	.C(n21532));
   NOR3xp33_ASAP7_75t_SL U26917 (.Y(n21536),
	.A(n22436),
	.B(n23076),
	.C(FE_OCPN28301_n22448));
   NAND3x1_ASAP7_75t_SL U26918 (.Y(n27001),
	.A(FE_OCPN29309_n26452),
	.B(n22422),
	.C(n21536));
   NOR3xp33_ASAP7_75t_SL U26919 (.Y(n24205),
	.A(n21538),
	.B(n27001),
	.C(n21537));
   NAND3xp33_ASAP7_75t_L U26920 (.Y(n21543),
	.A(n21539),
	.B(n25060),
	.C(n22456));
   OAI21xp33_ASAP7_75t_R U26921 (.Y(n22187),
	.A1(n17318),
	.A2(n23107),
	.B(n22467));
   NOR3xp33_ASAP7_75t_SRAM U26922 (.Y(n21547),
	.A(n21544),
	.B(n23075),
	.C(n23092));
   NAND3xp33_ASAP7_75t_R U26923 (.Y(n21550),
	.A(n21547),
	.B(n22422),
	.C(n22184));
   NOR2xp33_ASAP7_75t_L U26924 (.Y(n22176),
	.A(FE_OFN27072_n18671),
	.B(FE_OCPN29333_n17330));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26925 (.Y(n21579),
	.A1(n26679),
	.A2(n26678),
	.B(FE_OCPN28279_n),
	.C(w1_30_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26926 (.Y(n294),
	.A1(n26679),
	.A2(n26678),
	.B(n21580),
	.C(n21579));
   NOR2xp33_ASAP7_75t_L U26927 (.Y(n24790),
	.A(FE_OCPN27829_n25102),
	.B(n21604));
   OAI22xp33_ASAP7_75t_SRAM U26928 (.Y(n21581),
	.A1(FE_OCPN28057_n17603),
	.A2(n24790),
	.B1(FE_OFN29094_n21607),
	.B2(n24790));
   NAND3xp33_ASAP7_75t_SRAM U26929 (.Y(n21582),
	.A(n25103),
	.B(n25104),
	.C(n21581));
   NOR3xp33_ASAP7_75t_SRAM U26930 (.Y(n21583),
	.A(n21582),
	.B(FE_PSN8281_n25118),
	.C(n25107));
   NAND3xp33_ASAP7_75t_SRAM U26931 (.Y(n21635),
	.A(n25115),
	.B(n21583),
	.C(n25113));
   NOR2xp33_ASAP7_75t_SRAM U26932 (.Y(n21589),
	.A(n17602),
	.B(n21590));
   NOR2xp33_ASAP7_75t_SRAM U26933 (.Y(n21593),
	.A(FE_OFN25917_n21591),
	.B(n21590));
   NAND2xp5_ASAP7_75t_SL U26934 (.Y(n25121),
	.A(n21595),
	.B(n21594));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26935 (.Y(n21598),
	.A1(FE_OCPN27971_n21627),
	.A2(n21626),
	.B(n21625),
	.C(n21596));
   NOR3xp33_ASAP7_75t_SRAM U26936 (.Y(n21600),
	.A(n21598),
	.B(n21628),
	.C(n21597));
   OAI21xp33_ASAP7_75t_L U26937 (.Y(n21606),
	.A1(FE_OCPN27829_n25102),
	.A2(n21604),
	.B(n21603));
   NOR2xp33_ASAP7_75t_SRAM U26939 (.Y(n21618),
	.A(FE_PSN8335_n17606),
	.B(n21619));
   NOR2xp33_ASAP7_75t_SRAM U26940 (.Y(n21621),
	.A(n17602),
	.B(n21619));
   A2O1A1Ixp33_ASAP7_75t_L U26941 (.Y(n21629),
	.A1(FE_OCPN27971_n21627),
	.A2(n21626),
	.B(n21625),
	.C(n21624));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26942 (.Y(n21632),
	.A1(FE_OCPN28169_n25121),
	.A2(n25120),
	.B(n26926),
	.C(n21631));
   NOR2xp33_ASAP7_75t_SRAM U26943 (.Y(n21645),
	.A(FE_OCPN27532_n21643),
	.B(n21642));
   NOR2xp33_ASAP7_75t_SRAM U26944 (.Y(n21657),
	.A(FE_OFN28776_n18532),
	.B(n21658));
   NOR3xp33_ASAP7_75t_SRAM U26945 (.Y(n21656),
	.A(n23691),
	.B(n23863),
	.C(n21648));
   NOR3xp33_ASAP7_75t_SRAM U26946 (.Y(n21651),
	.A(n21650),
	.B(n23864),
	.C(n21649));
   NAND3xp33_ASAP7_75t_L U26947 (.Y(n21653),
	.A(n21652),
	.B(n21663),
	.C(n21651));
   AND3x1_ASAP7_75t_SRAM U26948 (.Y(n21672),
	.A(n21664),
	.B(n21663),
	.C(n23810));
   NAND3xp33_ASAP7_75t_L U26949 (.Y(n21666),
	.A(FE_OCPN5110_n23721),
	.B(n21665),
	.C(n23787));
   NAND3xp33_ASAP7_75t_R U26950 (.Y(n21668),
	.A(n21667),
	.B(FE_OFN28477_n23853),
	.C(n21690));
   NAND3xp33_ASAP7_75t_L U26951 (.Y(n21697),
	.A(n21672),
	.B(n21671),
	.C(n21670));
   OAI22xp5_ASAP7_75t_L U26952 (.Y(n25327),
	.A1(FE_OFN28868_FE_OCPN27715_n23875),
	.A2(n21682),
	.B1(FE_OFN28986_n18597),
	.B2(n21682));
   AND3x1_ASAP7_75t_L U26953 (.Y(n21686),
	.A(n25327),
	.B(n21684),
	.C(n21683));
   NAND3x1_ASAP7_75t_SL U26954 (.Y(n21693),
	.A(n21691),
	.B(n23767),
	.C(n21690));
   A2O1A1Ixp33_ASAP7_75t_SL U26955 (.Y(n25832),
	.A1(n21701),
	.A2(n21700),
	.B(n26517),
	.C(n21699));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26957 (.Y(n21703),
	.A1(FE_OFN16176_n27207),
	.A2(n21705),
	.B(FE_OCPN5053_n25832),
	.C(w2_13_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26958 (.Y(n372),
	.A1(FE_OFN16176_n27207),
	.A2(n21705),
	.B(n21704),
	.C(n21703));
   OAI22xp33_ASAP7_75t_SRAM U26959 (.Y(n21713),
	.A1(n21708),
	.A2(n21707),
	.B1(FE_OFN28656_FE_OFN25986_n21012),
	.B2(n21707));
   OAI21xp33_ASAP7_75t_L U26960 (.Y(n21710),
	.A1(FE_OFN28677_n17998),
	.A2(FE_OFN27133_n21725),
	.B(n21709));
   NOR3xp33_ASAP7_75t_SRAM U26961 (.Y(n21712),
	.A(n21710),
	.B(n21740),
	.C(n21733));
   NAND3xp33_ASAP7_75t_SRAM U26962 (.Y(n21720),
	.A(n21713),
	.B(n21712),
	.C(n21711));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26963 (.Y(n21732),
	.A1(FE_OCPN27998_n18019),
	.A2(FE_OFN27133_n21725),
	.B(FE_OCPN27675_n17986),
	.C(n21724));
   NOR2xp33_ASAP7_75t_SRAM U26964 (.Y(n21739),
	.A(n21738),
	.B(n21740));
   NOR2xp33_ASAP7_75t_R U26965 (.Y(n21743),
	.A(FE_OCPN27617_n18016),
	.B(n21740));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26966 (.Y(n21762),
	.A1(n26819),
	.A2(n26725),
	.B(n26722),
	.C(FE_OFN27130_w3_28));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26967 (.Y(n303),
	.A1(n26819),
	.A2(n26725),
	.B(n21763),
	.C(n21762));
   O2A1O1Ixp5_ASAP7_75t_SRAM U26968 (.Y(n21765),
	.A1(FE_OFN26141_n23307),
	.A2(n22795),
	.B(FE_OCPN27947_n18177),
	.C(n21764));
   NAND3xp33_ASAP7_75t_L U26969 (.Y(n21784),
	.A(n22848),
	.B(n21780),
	.C(FE_PSN8301_n23197));
   NAND3xp33_ASAP7_75t_SRAM U26970 (.Y(n21783),
	.A(n21782),
	.B(n21781),
	.C(FE_OFN28966_n23329));
   NAND3xp33_ASAP7_75t_SL U26971 (.Y(n21809),
	.A(n23333),
	.B(n21792),
	.C(n23334));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26974 (.Y(n21812),
	.A1(n27117),
	.A2(n26531),
	.B(FE_OCPN29389_n26528),
	.C(w0_15_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26975 (.Y(n369),
	.A1(n27117),
	.A2(n26531),
	.B(n21813),
	.C(n21812));
   OAI21xp33_ASAP7_75t_SRAM U26976 (.Y(n21816),
	.A1(FE_OFN28570_n19172),
	.A2(n21814),
	.B(n19174));
   NOR3xp33_ASAP7_75t_R U26977 (.Y(n24077),
	.A(n21816),
	.B(n22511),
	.C(n22502));
   NAND3xp33_ASAP7_75t_R U26978 (.Y(n21832),
	.A(n24081),
	.B(n24077),
	.C(n24083));
   NOR2xp33_ASAP7_75t_R U26979 (.Y(n21826),
	.A(FE_OCPN5021_n17446),
	.B(n21827));
   NAND3xp33_ASAP7_75t_SRAM U26980 (.Y(n21843),
	.A(n26064),
	.B(n23249),
	.C(n21833));
   NAND2xp5_ASAP7_75t_SL U26981 (.Y(n21835),
	.A(n17473),
	.B(n21834));
   NOR3xp33_ASAP7_75t_SL U26982 (.Y(n21840),
	.A(n21839),
	.B(n21838),
	.C(n21837));
   NAND3xp33_ASAP7_75t_SRAM U26983 (.Y(n21853),
	.A(FE_OCPN27605_n23357),
	.B(n21847),
	.C(n22486));
   NOR2xp33_ASAP7_75t_SL U26984 (.Y(n21849),
	.A(n23267),
	.B(n21848));
   A2O1A1Ixp33_ASAP7_75t_SL U26985 (.Y(n24552),
	.A1(n21868),
	.A2(n21867),
	.B(n17506),
	.C(n21866));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26986 (.Y(n21869),
	.A1(n23400),
	.A2(FE_RN_278_0),
	.B(FE_OFN28934_n24552),
	.C(FE_OFN38_w0_17));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26987 (.Y(n353),
	.A1(n23400),
	.A2(FE_RN_278_0),
	.B(n21870),
	.C(n21869));
   NOR3xp33_ASAP7_75t_L U26988 (.Y(n21878),
	.A(FE_OFN28554_n21876),
	.B(n21875),
	.C(n21874));
   NOR3xp33_ASAP7_75t_SRAM U26989 (.Y(n21883),
	.A(n23043),
	.B(n21894),
	.C(n21906));
   NAND3xp33_ASAP7_75t_SRAM U26990 (.Y(n21889),
	.A(n21884),
	.B(n21883),
	.C(n21882));
   NOR3xp33_ASAP7_75t_R U26991 (.Y(n21917),
	.A(n21889),
	.B(n21888),
	.C(n21887));
   NOR3xp33_ASAP7_75t_L U26992 (.Y(n21898),
	.A(n21891),
	.B(n24460),
	.C(n21890));
   NAND3xp33_ASAP7_75t_L U26993 (.Y(n21895),
	.A(n23127),
	.B(n23950),
	.C(n23034));
   NOR3xp33_ASAP7_75t_L U26994 (.Y(n21897),
	.A(n21895),
	.B(n21894),
	.C(n21893));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26995 (.Y(n21919),
	.A1(n26857),
	.A2(n26793),
	.B(n26787),
	.C(FE_OFN16432_w3_16));
   A2O1A1Ixp33_ASAP7_75t_SRAM U26996 (.Y(n341),
	.A1(n26857),
	.A2(n26793),
	.B(n21920),
	.C(n21919));
   NOR3xp33_ASAP7_75t_SRAM U26997 (.Y(n21923),
	.A(n25318),
	.B(FE_OFN26533_n21922),
	.C(FE_OCPN27817_n21921));
   NAND3xp33_ASAP7_75t_SRAM U26998 (.Y(n21926),
	.A(FE_PSN8293_n25317),
	.B(n25316),
	.C(n21923));
   NOR3xp33_ASAP7_75t_SRAM U26999 (.Y(n21927),
	.A(n21926),
	.B(n25319),
	.C(n25325));
   NOR3xp33_ASAP7_75t_SRAM U27000 (.Y(n21931),
	.A(n21930),
	.B(n21929),
	.C(n21928));
   NOR2xp33_ASAP7_75t_SRAM U27001 (.Y(n21937),
	.A(FE_OFN28549_n21934),
	.B(n21972));
   NAND3xp33_ASAP7_75t_L U27002 (.Y(n21943),
	.A(n21937),
	.B(n21936),
	.C(n21935));
   NOR3xp33_ASAP7_75t_SL U27003 (.Y(n21949),
	.A(n26304),
	.B(n21945),
	.C(n21944));
   O2A1O1Ixp5_ASAP7_75t_SL U27004 (.Y(n27164),
	.A1(n21956),
	.A2(n21955),
	.B(n26942),
	.C(n21954));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27005 (.Y(n21958),
	.A1(n21961),
	.A2(n21960),
	.B(FE_OFN26650_n27164),
	.C(w2_0_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27006 (.Y(n436),
	.A1(n21961),
	.A2(n21960),
	.B(n21959),
	.C(n21958));
   NOR3xp33_ASAP7_75t_SRAM U27007 (.Y(n21971),
	.A(n21964),
	.B(n21963),
	.C(n21962));
   NOR3xp33_ASAP7_75t_L U27008 (.Y(n21970),
	.A(n21969),
	.B(n21968),
	.C(n25325));
   NOR2xp33_ASAP7_75t_SRAM U27009 (.Y(n21987),
	.A(FE_OFN28753_sa31_2),
	.B(n16295));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27011 (.Y(n22000),
	.A1(n26942),
	.A2(n26941),
	.B(FE_OCPN27809_n26938),
	.C(w2_1_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27012 (.Y(n435),
	.A1(n26942),
	.A2(n26941),
	.B(n22001),
	.C(n22000));
   NOR2xp33_ASAP7_75t_SRAM U27013 (.Y(n22005),
	.A(n22004),
	.B(n23499));
   NAND3xp33_ASAP7_75t_SRAM U27014 (.Y(n22014),
	.A(n22007),
	.B(n22006),
	.C(n22005));
   OAI22xp33_ASAP7_75t_L U27015 (.Y(n22011),
	.A1(FE_OFN16272_n24767),
	.A2(n22998),
	.B1(FE_OCPN27743_n22009),
	.B2(n22998));
   A2O1A1Ixp33_ASAP7_75t_L U27016 (.Y(n22982),
	.A1(n18970),
	.A2(FE_OCPN28381_n26660),
	.B(n22930),
	.C(FE_OCPN29373_FE_OFN29191_sa23_2));
   NAND3xp33_ASAP7_75t_SRAM U27017 (.Y(n22032),
	.A(n22019),
	.B(n22968),
	.C(n22018));
   NOR2xp33_ASAP7_75t_SL U27018 (.Y(n22026),
	.A(FE_OCPN28112_n26664),
	.B(FE_OFN27046_n22024));
   NAND2xp5_ASAP7_75t_SL U27019 (.Y(n22029),
	.A(n22028),
	.B(n22027));
   NAND3x1_ASAP7_75t_SL U27020 (.Y(n26659),
	.A(n22030),
	.B(n26556),
	.C(n22029));
   NOR3xp33_ASAP7_75t_SL U27021 (.Y(n22044),
	.A(n22042),
	.B(FE_OCPN8241_n22041),
	.C(n22040));
   NAND2xp33_ASAP7_75t_SRAM U27022 (.Y(n22057),
	.A(n27023),
	.B(n24821));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27023 (.Y(n22056),
	.A1(FE_OFN16169_n26567),
	.A2(FE_OFN28506_n26996),
	.B(FE_OFN28512_n27020),
	.C(w1_9_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27024 (.Y(n388),
	.A1(FE_OFN16169_n26567),
	.A2(FE_OFN28506_n26996),
	.B(n22057),
	.C(n22056));
   NAND3xp33_ASAP7_75t_SRAM U27025 (.Y(n22061),
	.A(n22059),
	.B(n22085),
	.C(n22058));
   NOR3xp33_ASAP7_75t_SL U27026 (.Y(n25915),
	.A(n22061),
	.B(n22060),
	.C(n25536));
   NAND2x1_ASAP7_75t_SL U27027 (.Y(n22911),
	.A(n22066),
	.B(n22065));
   NOR3xp33_ASAP7_75t_SL U27028 (.Y(n22068),
	.A(n22911),
	.B(n25528),
	.C(n22871));
   NAND2xp5_ASAP7_75t_SL U27029 (.Y(n26980),
	.A(n22068),
	.B(n22067));
   NOR3xp33_ASAP7_75t_SRAM U27030 (.Y(n22072),
	.A(n22071),
	.B(FE_OCPN28316_n26980),
	.C(n25911));
   NOR2xp33_ASAP7_75t_R U27031 (.Y(n22079),
	.A(FE_OFN108_n26971),
	.B(FE_OCPN27685_n26968));
   AND2x2_ASAP7_75t_L U27032 (.Y(n22078),
	.A(n22077),
	.B(FE_OCPN29423_n26970));
   NOR2xp33_ASAP7_75t_L U27033 (.Y(n22087),
	.A(FE_OCPN27771_n19275),
	.B(n22088));
   NOR2xp33_ASAP7_75t_SRAM U27034 (.Y(n22096),
	.A(FE_OFN25998_n17781),
	.B(FE_OCPN29318_n25524));
   NOR2xp33_ASAP7_75t_SRAM U27035 (.Y(n22099),
	.A(FE_OFN108_n26971),
	.B(FE_OCPN29318_n25524));
   O2A1O1Ixp5_ASAP7_75t_SL U27037 (.Y(n26983),
	.A1(n22115),
	.A2(n22114),
	.B(n27183),
	.C(n22113));
   A2O1A1Ixp33_ASAP7_75t_SL U27038 (.Y(n25916),
	.A1(n22117),
	.A2(n22116),
	.B(n26976),
	.C(n26983));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27039 (.Y(n22119),
	.A1(n27216),
	.A2(n22121),
	.B(FE_OCPN5131_n25916),
	.C(w2_24_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27040 (.Y(n328),
	.A1(n27216),
	.A2(n22121),
	.B(n22120),
	.C(n22119));
   NOR2xp33_ASAP7_75t_L U27041 (.Y(n22123),
	.A(FE_PSN8335_n17606),
	.B(n22124));
   NAND3xp33_ASAP7_75t_SL U27042 (.Y(n22150),
	.A(FE_OCPN28241_n22142),
	.B(n22141),
	.C(n22140));
   NOR2xp33_ASAP7_75t_R U27044 (.Y(n22158),
	.A(n17616),
	.B(n22156));
   NAND2xp33_ASAP7_75t_L U27045 (.Y(n22622),
	.A(n17602),
	.B(n22157));
   NOR3xp33_ASAP7_75t_SRAM U27046 (.Y(n22170),
	.A(n22169),
	.B(n22168),
	.C(n26029));
   NOR3x1_ASAP7_75t_SL U27047 (.Y(n26579),
	.A(n26031),
	.B(n26036),
	.C(n22172));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27049 (.Y(n22173),
	.A1(FE_OFN16163_n26584),
	.A2(n26583),
	.B(FE_OCPN29473_n26579),
	.C(FE_OFN47_w1_2));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27050 (.Y(n347),
	.A1(FE_OFN16163_n26584),
	.A2(n26583),
	.B(n22174),
	.C(n22173));
   NOR2xp33_ASAP7_75t_SRAM U27051 (.Y(n22180),
	.A(n22189),
	.B(n22176));
   A2O1A1Ixp33_ASAP7_75t_L U27052 (.Y(n22178),
	.A1(FE_OCPN29333_n17330),
	.A2(FE_OFN27052_n21551),
	.B(FE_OFN26648_n22197),
	.C(n26999));
   NAND3xp33_ASAP7_75t_SL U27053 (.Y(n25172),
	.A(n23113),
	.B(n22181),
	.C(n22182));
   NOR2xp33_ASAP7_75t_SRAM U27054 (.Y(n22195),
	.A(n17321),
	.B(n22196));
   NOR2xp33_ASAP7_75t_SRAM U27055 (.Y(n22199),
	.A(FE_OCPN29461_n22197),
	.B(n22196));
   NOR2xp33_ASAP7_75t_SRAM U27056 (.Y(n22207),
	.A(FE_OFN16208_n23101),
	.B(n22597));
   A2O1A1Ixp33_ASAP7_75t_SL U27057 (.Y(n25169),
	.A1(n22219),
	.A2(n22218),
	.B(n26464),
	.C(n22217));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27058 (.Y(n22220),
	.A1(n26679),
	.A2(n25172),
	.B(FE_OCPN27825_n25169),
	.C(w1_31_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27059 (.Y(n293),
	.A1(n26679),
	.A2(n25172),
	.B(n22221),
	.C(n22220));
   OAI21xp5_ASAP7_75t_SL U27060 (.Y(n22765),
	.A1(FE_OFN26158_n22224),
	.A2(n22223),
	.B(n22222));
   NAND3xp33_ASAP7_75t_SL U27061 (.Y(n22231),
	.A(n24591),
	.B(n24592),
	.C(n24587));
   NAND3xp33_ASAP7_75t_SRAM U27062 (.Y(n22243),
	.A(n22234),
	.B(n22778),
	.C(FE_OCPN28309_n22779));
   NOR3xp33_ASAP7_75t_SL U27063 (.Y(n22249),
	.A(n22248),
	.B(FE_OFN28475_n23573),
	.C(n22247));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27065 (.Y(n22267),
	.A1(n26139),
	.A2(n24214),
	.B(n25485),
	.C(w1_22_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27066 (.Y(n404),
	.A1(n26139),
	.A2(n24214),
	.B(n22268),
	.C(n22267));
   NAND3xp33_ASAP7_75t_SL U27067 (.Y(n22274),
	.A(n23165),
	.B(n22270),
	.C(n22269));
   NOR2xp33_ASAP7_75t_L U27068 (.Y(n22279),
	.A(n22278),
	.B(n22277));
   NAND3xp33_ASAP7_75t_L U27069 (.Y(n22298),
	.A(n24701),
	.B(FE_PSN8301_n23197),
	.C(n22291));
   OAI22xp33_ASAP7_75t_SRAM U27070 (.Y(n22322),
	.A1(FE_OFN28798_FE_OCPN27947_n18177),
	.A2(n22321),
	.B1(FE_RN_0_0),
	.B2(n22321));
   NOR3x1_ASAP7_75t_SL U27071 (.Y(n26362),
	.A(n22326),
	.B(n22325),
	.C(n22324));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27073 (.Y(n22327),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(FE_OCPN27744_n26362),
	.C(FE_OFN46_w0_12));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27074 (.Y(n290),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(n22328),
	.C(n22327));
   OAI21xp33_ASAP7_75t_SRAM U27075 (.Y(n22332),
	.A1(n22662),
	.A2(n22329),
	.B(n22669));
   NOR3xp33_ASAP7_75t_SRAM U27076 (.Y(n22338),
	.A(n22332),
	.B(n22331),
	.C(n22330));
   NOR3xp33_ASAP7_75t_SRAM U27077 (.Y(n22337),
	.A(n22334),
	.B(FE_OCPN8250_n22692),
	.C(n24278));
   NAND2xp33_ASAP7_75t_SRAM U27078 (.Y(n22365),
	.A(n25000),
	.B(FE_OFN27111_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27079 (.Y(n22364),
	.A1(n26829),
	.A2(n25005),
	.B(n25002),
	.C(FE_OFN16448_n));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27080 (.Y(n422),
	.A1(n26829),
	.A2(n25005),
	.B(n22365),
	.C(n22364));
   NOR3xp33_ASAP7_75t_SRAM U27081 (.Y(n22373),
	.A(n24991),
	.B(n22367),
	.C(n22366));
   NOR3xp33_ASAP7_75t_SRAM U27082 (.Y(n22371),
	.A(n22370),
	.B(n22369),
	.C(n22368));
   NAND3xp33_ASAP7_75t_SRAM U27083 (.Y(n22376),
	.A(n22373),
	.B(n22372),
	.C(n22371));
   NAND3xp33_ASAP7_75t_SRAM U27084 (.Y(n22382),
	.A(n22379),
	.B(n22378),
	.C(n22377));
   NAND3xp33_ASAP7_75t_R U27085 (.Y(n22406),
	.A(n22395),
	.B(n22394),
	.C(n22393));
   NAND3xp33_ASAP7_75t_SRAM U27086 (.Y(n22400),
	.A(n22397),
	.B(n24866),
	.C(n22396));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27090 (.Y(n22411),
	.A1(n25367),
	.A2(FE_OFN16189_n25672),
	.B(n25667),
	.C(FE_OFN26591_w3_3));
   NOR2xp33_ASAP7_75t_SRAM U27091 (.Y(n22423),
	.A(FE_OCPN27887_n17331),
	.B(n24392));
   NOR2xp33_ASAP7_75t_R U27092 (.Y(n22425),
	.A(n17321),
	.B(n24392));
   NAND3xp33_ASAP7_75t_SRAM U27093 (.Y(n22434),
	.A(n22432),
	.B(n22469),
	.C(n22431));
   NOR2x1_ASAP7_75t_R U27094 (.Y(n26453),
	.A(n23087),
	.B(n22435));
   NOR3xp33_ASAP7_75t_SL U27095 (.Y(n22446),
	.A(n22437),
	.B(n22436),
	.C(n24225));
   NOR2xp33_ASAP7_75t_R U27096 (.Y(n22439),
	.A(n17382),
	.B(n23093));
   NOR2xp33_ASAP7_75t_R U27098 (.Y(n22442),
	.A(FE_OCPN29408_n22461),
	.B(n23093));
   NOR3xp33_ASAP7_75t_SRAM U27099 (.Y(n22449),
	.A(n23092),
	.B(FE_OCPN28301_n22448),
	.C(n22447));
   NAND3xp33_ASAP7_75t_L U27100 (.Y(n22464),
	.A(n22458),
	.B(FE_OCPN29505_n22457),
	.C(n25062));
   A2O1A1Ixp33_ASAP7_75t_R U27101 (.Y(n22460),
	.A1(FE_OFN26054_sa01_3),
	.A2(FE_OFN28594_n26454),
	.B(n22459),
	.C(FE_OCPN27871_n17317));
   A2O1A1Ixp33_ASAP7_75t_L U27102 (.Y(n27008),
	.A1(n17382),
	.A2(FE_OFN27152_n17315),
	.B(n22591),
	.C(FE_OCPN27887_n17331));
   NAND3xp33_ASAP7_75t_R U27103 (.Y(n22471),
	.A(n22470),
	.B(n23078),
	.C(n22469));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27105 (.Y(n22478),
	.A1(n26282),
	.A2(n26250),
	.B(n26251),
	.C(w1_27_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27106 (.Y(n398),
	.A1(n26282),
	.A2(n26250),
	.B(n22479),
	.C(n22478));
   NOR2xp33_ASAP7_75t_SRAM U27107 (.Y(n22481),
	.A(n23247),
	.B(n23374));
   NAND3xp33_ASAP7_75t_SRAM U27108 (.Y(n22488),
	.A(n24547),
	.B(n24548),
	.C(n22485));
   NAND3x1_ASAP7_75t_SL U27109 (.Y(n24545),
	.A(n22487),
	.B(n22486),
	.C(n26080));
   NOR2xp33_ASAP7_75t_SRAM U27110 (.Y(n22491),
	.A(n22489),
	.B(n23375));
   NAND3xp33_ASAP7_75t_R U27111 (.Y(n22496),
	.A(n22495),
	.B(FE_OCPN27848_n23255),
	.C(n22494));
   NOR3xp33_ASAP7_75t_R U27112 (.Y(n22503),
	.A(n22502),
	.B(n22501),
	.C(n22500));
   A2O1A1Ixp33_ASAP7_75t_SL U27113 (.Y(n26735),
	.A1(n22522),
	.A2(n22521),
	.B(n26078),
	.C(n22520));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27114 (.Y(n22523),
	.A1(n27062),
	.A2(FE_OFN171_n26739),
	.B(FE_OFN28474_FE_OCPN5038_n26735),
	.C(w0_16_));
   NOR2xp33_ASAP7_75t_SL U27115 (.Y(n22548),
	.A(FE_OCPN27384_n22888),
	.B(FE_OCPN27424_n22560));
   NOR2xp33_ASAP7_75t_R U27116 (.Y(n22550),
	.A(FE_OCPN29469_n17747),
	.B(FE_OCPN27424_n22560));
   NOR3xp33_ASAP7_75t_SL U27117 (.Y(n22558),
	.A(n22556),
	.B(n22565),
	.C(n26980));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27119 (.Y(n22574),
	.A1(n27183),
	.A2(n27182),
	.B(n27177),
	.C(w2_31_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27120 (.Y(n289),
	.A1(n27183),
	.A2(n27182),
	.B(n22575),
	.C(n22574));
   NOR2xp33_ASAP7_75t_SRAM U27121 (.Y(n22576),
	.A(n22597),
	.B(n27006));
   NOR3xp33_ASAP7_75t_SRAM U27122 (.Y(n22586),
	.A(n18698),
	.B(n22584),
	.C(n22597));
   NAND3xp33_ASAP7_75t_SRAM U27123 (.Y(n22587),
	.A(n27002),
	.B(FE_OFN28576_n27003),
	.C(n22586));
   NOR3xp33_ASAP7_75t_SRAM U27124 (.Y(n22594),
	.A(n22592),
	.B(n22603),
	.C(n22591));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27125 (.Y(n22600),
	.A1(FE_OCPN27399_n22598),
	.A2(FE_OFN60_n27007),
	.B(FE_OFN27152_n17315),
	.C(n22596));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27126 (.Y(n22611),
	.A1(n26679),
	.A2(n25694),
	.B(n25444),
	.C(w1_24_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27127 (.Y(n397),
	.A1(n26679),
	.A2(n25694),
	.B(n22612),
	.C(n22611));
   NOR2xp33_ASAP7_75t_SRAM U27128 (.Y(n22616),
	.A(n22614),
	.B(n22613));
   NAND3xp33_ASAP7_75t_R U27129 (.Y(n22618),
	.A(n22617),
	.B(n22616),
	.C(n22615));
   NOR2xp33_ASAP7_75t_SRAM U27130 (.Y(n22627),
	.A(FE_PSN8308_n22624),
	.B(n22623));
   NOR3xp33_ASAP7_75t_R U27131 (.Y(n22638),
	.A(n22637),
	.B(n22636),
	.C(n22635));
   NAND3xp33_ASAP7_75t_L U27132 (.Y(n22644),
	.A(n24127),
	.B(n22643),
	.C(n25115));
   A2O1A1Ixp33_ASAP7_75t_SL U27133 (.Y(n24421),
	.A1(n22654),
	.A2(n22653),
	.B(n26926),
	.C(n22652));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27134 (.Y(n22655),
	.A1(FE_OFN16164_n25081),
	.A2(n24422),
	.B(n24421),
	.C(w1_5_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27135 (.Y(n277),
	.A1(FE_OFN16164_n25081),
	.A2(n24422),
	.B(n22656),
	.C(n22655));
   OAI21xp33_ASAP7_75t_R U27136 (.Y(n22664),
	.A1(FE_OCPN27246_n22663),
	.A2(n22662),
	.B(n22661));
   NOR3xp33_ASAP7_75t_SRAM U27137 (.Y(n22674),
	.A(n22664),
	.B(FE_OCPN27458_n24891),
	.C(FE_OFN28920_n24254));
   NAND3xp33_ASAP7_75t_SRAM U27138 (.Y(n22673),
	.A(n22667),
	.B(n22666),
	.C(n22665));
   NOR3xp33_ASAP7_75t_SRAM U27139 (.Y(n22687),
	.A(n22677),
	.B(n22676),
	.C(n22675));
   NOR3xp33_ASAP7_75t_SRAM U27140 (.Y(n22686),
	.A(n24256),
	.B(n22679),
	.C(n22678));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27141 (.Y(n24917),
	.A1(FE_OCPN5126_sa21_2),
	.A2(FE_OFN16153_n16747),
	.B(FE_OFN28981_n16767),
	.C(FE_OFN28529_n16774));
   NOR3xp33_ASAP7_75t_SRAM U27142 (.Y(n22714),
	.A(n22688),
	.B(n23638),
	.C(n23671));
   NOR2xp33_ASAP7_75t_SRAM U27143 (.Y(n22695),
	.A(n22694),
	.B(n22696));
   NOR2xp33_ASAP7_75t_SRAM U27144 (.Y(n22698),
	.A(FE_OFN28698_sa21_1),
	.B(n22696));
   NOR3xp33_ASAP7_75t_L U27145 (.Y(n22710),
	.A(n22709),
	.B(n23652),
	.C(n22708));
   NAND2xp33_ASAP7_75t_SRAM U27146 (.Y(n22717),
	.A(n26824),
	.B(FE_OFN26639_w3_14));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27147 (.Y(n22716),
	.A1(n26829),
	.A2(n26828),
	.B(FE_OCPN8221_n26825),
	.C(FE_OCPN29536_FE_OFN8_w3_14));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27148 (.Y(n279),
	.A1(n26829),
	.A2(n26828),
	.B(n22717),
	.C(n22716));
   NOR3xp33_ASAP7_75t_SRAM U27149 (.Y(n22733),
	.A(n22719),
	.B(n22718),
	.C(n24370));
   NAND3xp33_ASAP7_75t_SRAM U27150 (.Y(n22727),
	.A(n25398),
	.B(n23235),
	.C(n22720));
   NOR3xp33_ASAP7_75t_R U27151 (.Y(n22732),
	.A(n22727),
	.B(n22726),
	.C(n22756));
   NOR3x1_ASAP7_75t_SL U27152 (.Y(n23599),
	.A(n22731),
	.B(n22730),
	.C(FE_OFN26588_n24062));
   NOR2xp33_ASAP7_75t_SL U27153 (.Y(n22736),
	.A(n24364),
	.B(n22734));
   NOR2xp33_ASAP7_75t_L U27154 (.Y(n22768),
	.A(FE_OCPN5137_n23600),
	.B(n23581));
   NAND3xp33_ASAP7_75t_SL U27155 (.Y(n22757),
	.A(n23616),
	.B(n22741),
	.C(n22740));
   NOR2xp33_ASAP7_75t_L U27156 (.Y(n22744),
	.A(FE_OFN26125_n22742),
	.B(n25439));
   NAND3xp33_ASAP7_75t_SRAM U27157 (.Y(n22761),
	.A(n22759),
	.B(n25398),
	.C(n22758));
   NOR2xp33_ASAP7_75t_R U27158 (.Y(n22766),
	.A(n24364),
	.B(n23581));
   NAND3x1_ASAP7_75t_SL U27159 (.Y(n22775),
	.A(n22773),
	.B(n22772),
	.C(n22771));
   NOR2xp33_ASAP7_75t_SRAM U27161 (.Y(n22780),
	.A(n25741),
	.B(n22781));
   AND3x1_ASAP7_75t_SRAM U27162 (.Y(n22782),
	.A(FE_OCPN28309_n22779),
	.B(n22778),
	.C(n22777));
   NOR2xp33_ASAP7_75t_SRAM U27163 (.Y(n22783),
	.A(n17898),
	.B(n22781));
   INVxp67_ASAP7_75t_SL U27164 (.Y(n26134),
	.A(n26135));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27165 (.Y(n22793),
	.A1(n26139),
	.A2(n26138),
	.B(n26135),
	.C(w1_20_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27166 (.Y(n403),
	.A1(n26139),
	.A2(n26138),
	.B(n22794),
	.C(n22793));
   OAI22xp33_ASAP7_75t_SRAM U27167 (.Y(n22799),
	.A1(FE_OCPN27722_n23336),
	.A2(n22796),
	.B1(n22795),
	.B2(n22796));
   NAND3xp33_ASAP7_75t_SRAM U27168 (.Y(n22804),
	.A(n22799),
	.B(n22798),
	.C(n22797));
   NAND3xp33_ASAP7_75t_SRAM U27169 (.Y(n22803),
	.A(n22802),
	.B(n22801),
	.C(n22800));
   NOR3xp33_ASAP7_75t_SRAM U27170 (.Y(n22809),
	.A(FE_OCPN8257_n18178),
	.B(FE_OCPN27979_FE_OFN16147_sa22_1),
	.C(n24691));
   NOR3xp33_ASAP7_75t_R U27171 (.Y(n22817),
	.A(n22809),
	.B(FE_OFN16304_n22808),
	.C(n22807));
   NOR2xp33_ASAP7_75t_R U27172 (.Y(n22810),
	.A(FE_OFN26141_n23307),
	.B(FE_OFN29241_n22811));
   NOR2xp33_ASAP7_75t_R U27173 (.Y(n22813),
	.A(FE_OCPN27947_n18177),
	.B(FE_OFN29241_n22811));
   NOR2xp33_ASAP7_75t_SL U27174 (.Y(n22820),
	.A(FE_OFN26528_n23302),
	.B(n22821));
   NOR2xp33_ASAP7_75t_L U27175 (.Y(n22822),
	.A(n18176),
	.B(n22821));
   NOR2xp33_ASAP7_75t_R U27176 (.Y(n22826),
	.A(n23315),
	.B(n22827));
   NOR2xp33_ASAP7_75t_SRAM U27177 (.Y(n22830),
	.A(n22828),
	.B(n22827));
   NAND3xp33_ASAP7_75t_L U27178 (.Y(n22835),
	.A(n22834),
	.B(n23312),
	.C(n22833));
   NOR2xp33_ASAP7_75t_SRAM U27179 (.Y(n22837),
	.A(FE_OCPN27721_n23336),
	.B(n22838));
   NOR2xp33_ASAP7_75t_SRAM U27180 (.Y(n22840),
	.A(FE_RN_0_0),
	.B(n22838));
   NOR2xp33_ASAP7_75t_SRAM U27181 (.Y(n22844),
	.A(FE_OCPN27722_n23336),
	.B(n23169));
   NOR2xp33_ASAP7_75t_SRAM U27182 (.Y(n22845),
	.A(n18159),
	.B(n23169));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27183 (.Y(n22858),
	.A1(n18166),
	.A2(FE_OCPN8257_n18178),
	.B(FE_OFN16450_n23315),
	.C(n22854));
   A2O1A1Ixp33_ASAP7_75t_SL U27184 (.Y(n26479),
	.A1(n22868),
	.A2(n22867),
	.B(n23345),
	.C(n22866));
   INVx2_ASAP7_75t_SL U27185 (.Y(n26477),
	.A(FE_OCPN27494_n26479));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27186 (.Y(n22869),
	.A1(n27117),
	.A2(FE_PSN8300_n26482),
	.B(FE_OCPN27494_n26479),
	.C(FE_OFN53_w0_8));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27187 (.Y(n367),
	.A1(n27117),
	.A2(FE_PSN8300_n26482),
	.B(n22870),
	.C(n22869));
   NOR2xp33_ASAP7_75t_SRAM U27188 (.Y(n22880),
	.A(FE_PSN8313_FE_OCPN29469_n17747),
	.B(n22881));
   NAND3xp33_ASAP7_75t_L U27189 (.Y(n22879),
	.A(n22878),
	.B(n22877),
	.C(n22876));
   NOR2xp33_ASAP7_75t_SRAM U27190 (.Y(n22884),
	.A(n22882),
	.B(n22881));
   AND3x1_ASAP7_75t_SRAM U27191 (.Y(n22889),
	.A(FE_OCPN27384_n22888),
	.B(FE_OCPN27579_FE_OFN16138_sa02_5),
	.C(FE_OFN28730_FE_OCPN28416_sa02_3));
   NOR3xp33_ASAP7_75t_SRAM U27192 (.Y(n22898),
	.A(n22889),
	.B(n22900),
	.C(n22899));
   NAND3xp33_ASAP7_75t_SRAM U27193 (.Y(n22895),
	.A(n22892),
	.B(n22891),
	.C(n22890));
   NOR3xp33_ASAP7_75t_L U27194 (.Y(n22897),
	.A(n22895),
	.B(n22894),
	.C(n22893));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27196 (.Y(n22914),
	.A1(n27183),
	.A2(n24178),
	.B(n24175),
	.C(w2_29_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27197 (.Y(n319),
	.A1(n27183),
	.A2(n24178),
	.B(n22915),
	.C(n22914));
   NOR2xp33_ASAP7_75t_SRAM U27198 (.Y(n22918),
	.A(FE_OFN29003_n23491),
	.B(n22998));
   NAND3xp33_ASAP7_75t_R U27199 (.Y(n22924),
	.A(n26163),
	.B(n26162),
	.C(n22921));
   OAI21xp33_ASAP7_75t_L U27200 (.Y(n22933),
	.A1(n22010),
	.A2(FE_OCPN28363_n22979),
	.B(n22932));
   NOR2xp33_ASAP7_75t_SRAM U27201 (.Y(n22937),
	.A(n19000),
	.B(n22935));
   OAI22xp33_ASAP7_75t_SL U27203 (.Y(n22960),
	.A1(n22967),
	.A2(n26571),
	.B1(n22949),
	.B2(n26571));
   OAI21xp33_ASAP7_75t_L U27204 (.Y(n22956),
	.A1(FE_OCPN27803_sa23_4),
	.A2(n22990),
	.B(n19010));
   NOR3xp33_ASAP7_75t_R U27205 (.Y(n24765),
	.A(n22952),
	.B(n22951),
	.C(n22950));
   NAND3xp33_ASAP7_75t_SL U27206 (.Y(n22955),
	.A(n22954),
	.B(n22953),
	.C(n26152));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27208 (.Y(n22962),
	.A1(n26249),
	.A2(n25736),
	.B(n26178),
	.C(w1_10_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27209 (.Y(n385),
	.A1(n26249),
	.A2(n25736),
	.B(n22963),
	.C(n22962));
   O2A1O1Ixp5_ASAP7_75t_SRAM U27210 (.Y(n26669),
	.A1(FE_OFN29026_n20911),
	.A2(FE_OFN16248_n20235),
	.B(FE_OFN29001_n23491),
	.C(n26154));
   NAND3xp33_ASAP7_75t_SRAM U27211 (.Y(n22965),
	.A(FE_OCPN29548_n25717),
	.B(n25716),
	.C(n26669));
   NOR3xp33_ASAP7_75t_SRAM U27212 (.Y(n22972),
	.A(n22971),
	.B(FE_OCPN27916_n),
	.C(n22970));
   NAND3xp33_ASAP7_75t_SL U27213 (.Y(n22989),
	.A(n22987),
	.B(n22986),
	.C(n22985));
   NOR2xp33_ASAP7_75t_L U27214 (.Y(n22993),
	.A(FE_OCPN27577_sa23_4),
	.B(n22990));
   NAND3xp33_ASAP7_75t_SL U27215 (.Y(n23001),
	.A(n19010),
	.B(n23000),
	.C(n24041));
   O2A1O1Ixp5_ASAP7_75t_SL U27217 (.Y(n23007),
	.A1(n23515),
	.A2(n23006),
	.B(n26249),
	.C(n23005));
   OAI21x1_ASAP7_75t_SL U27218 (.Y(n26683),
	.A1(n23008),
	.A2(n26571),
	.B(n23007));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27220 (.Y(n23009),
	.A1(FE_OFN16169_n26567),
	.A2(n24812),
	.B(FE_OCPN28383_n24808),
	.C(w1_15_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27221 (.Y(n389),
	.A1(FE_OFN16169_n26567),
	.A2(n24812),
	.B(n23010),
	.C(n23009));
   NAND3xp33_ASAP7_75t_SRAM U27222 (.Y(n23017),
	.A(n23980),
	.B(FE_OFN25959_n23011),
	.C(FE_OFN28722_sa10_3));
   NOR2xp33_ASAP7_75t_SRAM U27223 (.Y(n23984),
	.A(n24944),
	.B(n23141));
   OR2x2_ASAP7_75t_SRAM U27224 (.Y(n23990),
	.A(n16533),
	.B(n23012));
   NAND2xp33_ASAP7_75t_SRAM U27225 (.Y(n23014),
	.A(n23984),
	.B(n23990));
   NOR2xp33_ASAP7_75t_SRAM U27226 (.Y(n23986),
	.A(FE_OFN28912_n16534),
	.B(n23141));
   NAND2xp33_ASAP7_75t_SRAM U27227 (.Y(n23013),
	.A(n23986),
	.B(n23990));
   NAND2xp33_ASAP7_75t_SRAM U27228 (.Y(n23016),
	.A(n23014),
	.B(n23013));
   NAND3xp33_ASAP7_75t_SRAM U27229 (.Y(n23020),
	.A(n23017),
	.B(n23016),
	.C(n23979));
   NOR3xp33_ASAP7_75t_SRAM U27230 (.Y(n23021),
	.A(n23020),
	.B(FE_OFN169_n23992),
	.C(n23018));
   NAND3xp33_ASAP7_75t_SRAM U27231 (.Y(n23058),
	.A(n23993),
	.B(n23021),
	.C(n23994));
   NOR3xp33_ASAP7_75t_SRAM U27232 (.Y(n23053),
	.A(n23999),
	.B(n23997),
	.C(n23022));
   NAND3xp33_ASAP7_75t_SL U27234 (.Y(n23032),
	.A(n23029),
	.B(n23028),
	.C(n24949));
   NOR3xp33_ASAP7_75t_L U27235 (.Y(n23033),
	.A(n23032),
	.B(FE_OCPN5015_n23031),
	.C(FE_OFN16378_n23030));
   OA21x2_ASAP7_75t_SRAM U27236 (.Y(n23039),
	.A1(n23036),
	.A2(n23982),
	.B(n23950));
   NOR2xp33_ASAP7_75t_L U27237 (.Y(n23040),
	.A(FE_OCPN28157_n16534),
	.B(n23038));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27238 (.Y(n23055),
	.A1(n23053),
	.A2(n23052),
	.B(n24978),
	.C(FE_OCPN8260_n26335));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27239 (.Y(n23056),
	.A1(n24974),
	.A2(n23058),
	.B(n23055),
	.C(FE_OFN16441_w3_21));
   NOR2xp33_ASAP7_75t_SRAM U27240 (.Y(n23061),
	.A(n23059),
	.B(n23062));
   NOR2xp33_ASAP7_75t_SRAM U27241 (.Y(n23063),
	.A(FE_OFN27152_n17315),
	.B(n17331));
   NOR2xp33_ASAP7_75t_SRAM U27242 (.Y(n23065),
	.A(n23063),
	.B(n23062));
   NOR2xp33_ASAP7_75t_SRAM U27243 (.Y(n23077),
	.A(n23076),
	.B(n23075));
   NAND3xp33_ASAP7_75t_R U27244 (.Y(n23080),
	.A(n23079),
	.B(n23078),
	.C(n23077));
   NOR2xp33_ASAP7_75t_SRAM U27245 (.Y(n23089),
	.A(n17329),
	.B(n23087));
   NOR3xp33_ASAP7_75t_SRAM U27246 (.Y(n23095),
	.A(n23094),
	.B(n23093),
	.C(n23092));
   NOR2xp33_ASAP7_75t_SRAM U27247 (.Y(n23100),
	.A(n23099),
	.B(FE_OFN78_n22457));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27248 (.Y(n23117),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(FE_OFN27123_n26275),
	.C(w1_25_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27249 (.Y(n395),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(n23118),
	.C(n23117));
   NOR3xp33_ASAP7_75t_SRAM U27250 (.Y(n23124),
	.A(FE_OFN27094_n24956),
	.B(n23119),
	.C(FE_OFN28586_n24736));
   NOR3xp33_ASAP7_75t_SRAM U27251 (.Y(n23123),
	.A(n24735),
	.B(n24734),
	.C(FE_OCPN5158_n24742));
   NAND3xp33_ASAP7_75t_SRAM U27252 (.Y(n23130),
	.A(FE_OCPN5153_n23127),
	.B(n23126),
	.C(FE_OCPN29529_n23125));
   NOR3xp33_ASAP7_75t_SRAM U27253 (.Y(n23136),
	.A(n23133),
	.B(n23132),
	.C(n23131));
   OR2x2_ASAP7_75t_SRAM U27254 (.Y(n23147),
	.A(FE_OCPN29407_FE_OFN142_sa10_0),
	.B(FE_OCPN29424_FE_OFN26039_sa10_2));
   NOR2xp33_ASAP7_75t_SRAM U27255 (.Y(n23150),
	.A(n23148),
	.B(n23948));
   O2A1O1Ixp33_ASAP7_75t_L U27256 (.Y(n23156),
	.A1(n24732),
	.A2(n24731),
	.B(n26857),
	.C(n24740));
   A2O1A1Ixp33_ASAP7_75t_SL U27257 (.Y(n24936),
	.A1(n24964),
	.A2(n23157),
	.B(n25139),
	.C(n23156));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27258 (.Y(n23158),
	.A1(n24974),
	.A2(n24939),
	.B(n24936),
	.C(FE_OFN26072_n26720));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27259 (.Y(n342),
	.A1(n24974),
	.A2(n24939),
	.B(n23159),
	.C(n23158));
   NOR3xp33_ASAP7_75t_SRAM U27260 (.Y(n23166),
	.A(n23164),
	.B(FE_OFN26009_n18213),
	.C(n23162));
   NAND3xp33_ASAP7_75t_R U27261 (.Y(n23167),
	.A(n23190),
	.B(n23166),
	.C(n23165));
   NOR3xp33_ASAP7_75t_SRAM U27262 (.Y(n23171),
	.A(n23170),
	.B(n23169),
	.C(n23168));
   NOR2xp33_ASAP7_75t_SRAM U27263 (.Y(n23177),
	.A(FE_OCPN27722_n23336),
	.B(n23297));
   NOR2xp33_ASAP7_75t_SRAM U27264 (.Y(n23179),
	.A(FE_OFN16407_n23322),
	.B(n23297));
   OAI21xp33_ASAP7_75t_SRAM U27265 (.Y(n23186),
	.A1(n18186),
	.A2(n18166),
	.B(n23182));
   NOR3xp33_ASAP7_75t_R U27266 (.Y(n23188),
	.A(n23186),
	.B(n23185),
	.C(n23184));
   NAND3xp33_ASAP7_75t_R U27267 (.Y(n23199),
	.A(n23189),
	.B(n23188),
	.C(n23187));
   NAND3xp33_ASAP7_75t_R U27268 (.Y(n23193),
	.A(n23192),
	.B(n23191),
	.C(n23190));
   A2O1A1Ixp33_ASAP7_75t_SL U27269 (.Y(n25976),
	.A1(n23203),
	.A2(n23202),
	.B(n26889),
	.C(n23201));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27271 (.Y(n23204),
	.A1(n27117),
	.A2(FE_OFN28690_n25979),
	.B(n25974),
	.C(FE_OFN44_w0_9));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27272 (.Y(n364),
	.A1(n27117),
	.A2(FE_OFN28690_n25979),
	.B(n23205),
	.C(n23204));
   NOR2xp33_ASAP7_75t_SRAM U27273 (.Y(n23207),
	.A(n25741),
	.B(n23208));
   NOR2xp33_ASAP7_75t_SRAM U27274 (.Y(n23210),
	.A(FE_OFN29211_n23587),
	.B(n23208));
   NOR2xp33_ASAP7_75t_SRAM U27275 (.Y(n23219),
	.A(n25741),
	.B(n23214));
   A2O1A1Ixp33_ASAP7_75t_SL U27276 (.Y(n23218),
	.A1(n23217),
	.A2(FE_OCPN29324_n23216),
	.B(n23215),
	.C(n24378));
   NAND2xp5_ASAP7_75t_SL U27277 (.Y(n25162),
	.A(n23223),
	.B(n23222));
   NAND3xp33_ASAP7_75t_SRAM U27278 (.Y(n23239),
	.A(n23236),
	.B(n23235),
	.C(n23234));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27279 (.Y(n23244),
	.A1(n26139),
	.A2(n25725),
	.B(n25722),
	.C(w1_23_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27280 (.Y(n274),
	.A1(n26139),
	.A2(n25725),
	.B(n23245),
	.C(n23244));
   NAND3xp33_ASAP7_75t_SL U27281 (.Y(n23263),
	.A(n23258),
	.B(n23257),
	.C(n23256));
   NAND3xp33_ASAP7_75t_SRAM U27282 (.Y(n23271),
	.A(n23269),
	.B(n23391),
	.C(n23268));
   INVxp33_ASAP7_75t_SRAM U27283 (.Y(n23279),
	.A(n25786));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27284 (.Y(n23294),
	.A1(n27062),
	.A2(n27061),
	.B(n27058),
	.C(w0_22_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27285 (.Y(n276),
	.A1(n27062),
	.A2(n27061),
	.B(n23295),
	.C(n23294));
   NOR3xp33_ASAP7_75t_SRAM U27286 (.Y(n23314),
	.A(FE_OCPN27719_n23306),
	.B(FE_OFN28688_sa22_2),
	.C(FE_OFN29152_sa22_0));
   NOR2xp33_ASAP7_75t_SRAM U27287 (.Y(n23317),
	.A(n23315),
	.B(n23314));
   OAI22xp33_ASAP7_75t_SRAM U27288 (.Y(n23326),
	.A1(n23336),
	.A2(n23323),
	.B1(n23322),
	.B2(n23323));
   NAND3xp33_ASAP7_75t_R U27289 (.Y(n23332),
	.A(n23326),
	.B(n23325),
	.C(n23324));
   NAND3xp33_ASAP7_75t_SRAM U27290 (.Y(n23330),
	.A(FE_OFN28966_n23329),
	.B(n20733),
	.C(n23327));
   A2O1A1Ixp33_ASAP7_75t_SL U27291 (.Y(n27049),
	.A1(n23352),
	.A2(n23351),
	.B(n26889),
	.C(n23350));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27293 (.Y(n23353),
	.A1(n27117),
	.A2(n27052),
	.B(FE_OCPN28073_n27049),
	.C(w0_14_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27294 (.Y(n278),
	.A1(n27117),
	.A2(n27052),
	.B(n23354),
	.C(n23353));
   NOR2xp33_ASAP7_75t_SRAM U27295 (.Y(n23358),
	.A(n23355),
	.B(n25786));
   AND2x2_ASAP7_75t_R U27296 (.Y(n23360),
	.A(FE_OCPN27605_n23357),
	.B(n23356));
   NOR2xp33_ASAP7_75t_SRAM U27297 (.Y(n23361),
	.A(FE_OCPN27414_n23359),
	.B(n25786));
   NOR2xp33_ASAP7_75t_SRAM U27298 (.Y(n23379),
	.A(n23375),
	.B(n23374));
   NAND3xp33_ASAP7_75t_L U27299 (.Y(n23396),
	.A(n23391),
	.B(n23390),
	.C(n23389));
   NOR2xp33_ASAP7_75t_SRAM U27300 (.Y(n23395),
	.A(n23393),
	.B(FE_OCPN28447_n23392));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27301 (.Y(n23410),
	.A1(n26082),
	.A2(n25605),
	.B(n25606),
	.C(FE_OFN39_w0_21));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27302 (.Y(n358),
	.A1(n26082),
	.A2(FE_PSN8278_n25605),
	.B(n23411),
	.C(n23410));
   NAND3xp33_ASAP7_75t_SRAM U27303 (.Y(n23424),
	.A(n23416),
	.B(n23415),
	.C(n23414));
   NOR2xp33_ASAP7_75t_SRAM U27304 (.Y(n23427),
	.A(FE_OCPN27611_n23426),
	.B(n23425));
   NOR2xp33_ASAP7_75t_SRAM U27305 (.Y(n23433),
	.A(n23431),
	.B(n23430));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27306 (.Y(n23440),
	.A1(FE_OCPN29283_n23439),
	.A2(FE_OCPN27733_n17996),
	.B(FE_OCPN27675_n17986),
	.C(n23438));
   NOR3xp33_ASAP7_75t_SRAM U27307 (.Y(n23468),
	.A(n23442),
	.B(n23441),
	.C(n23440));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27308 (.Y(n23470),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(FE_OCPN28106_FE_OFN25876_n25462),
	.C(FE_OFN27206_w3_30));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27309 (.Y(n302),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(n23471),
	.C(n23470));
   NOR3xp33_ASAP7_75t_R U27310 (.Y(n23477),
	.A(n23474),
	.B(n23473),
	.C(n23472));
   NOR2xp33_ASAP7_75t_SRAM U27311 (.Y(n23489),
	.A(FE_OFN29026_n20911),
	.B(n23490));
   NOR2xp33_ASAP7_75t_SRAM U27312 (.Y(n23493),
	.A(FE_OFN28580_n23491),
	.B(n23490));
   NOR3xp33_ASAP7_75t_SRAM U27313 (.Y(n23509),
	.A(n23498),
	.B(FE_OFN25890_n23497),
	.C(n23496));
   NOR2xp33_ASAP7_75t_SRAM U27314 (.Y(n23503),
	.A(n23500),
	.B(n23499));
   INVxp33_ASAP7_75t_SRAM U27315 (.Y(n23505),
	.A(FE_OCPN28107_n23504));
   NAND3xp33_ASAP7_75t_SRAM U27316 (.Y(n23512),
	.A(FE_OFN29003_n23491),
	.B(n23510),
	.C(FE_OCPN29373_FE_OFN29191_sa23_2));
   NAND3xp33_ASAP7_75t_R U27317 (.Y(n23516),
	.A(n23513),
	.B(n23512),
	.C(n23511));
   NOR3xp33_ASAP7_75t_SL U27318 (.Y(n23518),
	.A(n23516),
	.B(n23515),
	.C(n23514));
   O2A1O1Ixp5_ASAP7_75t_SL U27319 (.Y(n23523),
	.A1(n23522),
	.A2(n23521),
	.B(n24038),
	.C(n23520));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27320 (.Y(n23526),
	.A1(n26249),
	.A2(n26248),
	.B(FE_OFN26149_n26245),
	.C(w1_12_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27321 (.Y(n304),
	.A1(n26249),
	.A2(n26248),
	.B(n23527),
	.C(n23526));
   NAND3xp33_ASAP7_75t_SRAM U27322 (.Y(n23570),
	.A(n26358),
	.B(n26359),
	.C(n26360));
   NOR2xp33_ASAP7_75t_SRAM U27323 (.Y(n23567),
	.A(FE_OFN29005_n23558),
	.B(n23530));
   NAND3xp33_ASAP7_75t_SRAM U27324 (.Y(n23536),
	.A(n23533),
	.B(FE_OCPN29561_n23532),
	.C(n23531));
   NOR3xp33_ASAP7_75t_SRAM U27325 (.Y(n23541),
	.A(n23538),
	.B(n26122),
	.C(n23537));
   NOR2xp33_ASAP7_75t_SRAM U27326 (.Y(n23540),
	.A(FE_OCPN7607_n23539),
	.B(n24300));
   NAND3xp33_ASAP7_75t_R U27327 (.Y(n23545),
	.A(n23542),
	.B(n23541),
	.C(n23540));
   NAND3xp33_ASAP7_75t_R U27328 (.Y(n23563),
	.A(n23562),
	.B(n23561),
	.C(n23560));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27329 (.Y(n23568),
	.A1(n23571),
	.A2(n23570),
	.B(FE_OCPN27641_n27121),
	.C(w0_4_));
   NOR3xp33_ASAP7_75t_L U27330 (.Y(n24375),
	.A(n23583),
	.B(n23582),
	.C(n23581));
   NOR2xp33_ASAP7_75t_SRAM U27331 (.Y(n23589),
	.A(n23587),
	.B(n23590));
   NOR2xp33_ASAP7_75t_SRAM U27332 (.Y(n23592),
	.A(n23603),
	.B(n23590));
   NAND3xp33_ASAP7_75t_SL U27333 (.Y(n23620),
	.A(n24046),
	.B(n23599),
	.C(n23598));
   NAND3xp33_ASAP7_75t_SL U27334 (.Y(n23614),
	.A(n23613),
	.B(n23612),
	.C(n23611));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27335 (.Y(n23623),
	.A1(n26139),
	.A2(n25455),
	.B(n25452),
	.C(w1_17_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27336 (.Y(n406),
	.A1(n26139),
	.A2(n25455),
	.B(n23624),
	.C(n23623));
   NAND3xp33_ASAP7_75t_SRAM U27337 (.Y(n23632),
	.A(n23626),
	.B(n23625),
	.C(n24919));
   O2A1O1Ixp5_ASAP7_75t_SRAM U27338 (.Y(n23627),
	.A1(FE_OFN28779_n24257),
	.A2(FE_OFN16447_n16749),
	.B(FE_OCPN27690_n16757),
	.C(n25353));
   NOR2xp33_ASAP7_75t_SRAM U27339 (.Y(n23634),
	.A(FE_OFN27157_n23928),
	.B(n23632));
   NOR2xp33_ASAP7_75t_SRAM U27340 (.Y(n23646),
	.A(FE_OCPN28299_n),
	.B(n23643));
   NAND3xp33_ASAP7_75t_R U27341 (.Y(n23653),
	.A(FE_OCPN27774_n25351),
	.B(n23650),
	.C(n23649));
   NOR3xp33_ASAP7_75t_L U27342 (.Y(n23655),
	.A(n23653),
	.B(n23652),
	.C(n23651));
   NOR2xp33_ASAP7_75t_SRAM U27343 (.Y(n23660),
	.A(FE_OFN28778_FE_OCPN28352_n16748),
	.B(n23661));
   NOR2xp33_ASAP7_75t_R U27344 (.Y(n23663),
	.A(FE_OFN29023_n16750),
	.B(n23661));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27345 (.Y(n23675),
	.A1(n26829),
	.A2(n25959),
	.B(FE_OFN16249_n25956),
	.C(FE_OFN102_w3_12));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27346 (.Y(n423),
	.A1(n26829),
	.A2(n25959),
	.B(n23676),
	.C(n23675));
   NOR2xp33_ASAP7_75t_SRAM U27347 (.Y(n23679),
	.A(FE_OFN16295_n23837),
	.B(n23680));
   AND3x1_ASAP7_75t_SRAM U27348 (.Y(n23681),
	.A(n23678),
	.B(FE_OFN29096_n25188),
	.C(n23752));
   NOR2xp33_ASAP7_75t_SRAM U27349 (.Y(n23682),
	.A(FE_OFN29081_n18526),
	.B(n23680));
   NOR2xp33_ASAP7_75t_L U27350 (.Y(n23690),
	.A(FE_OCPN28257_n23689),
	.B(n23688));
   NOR2xp33_ASAP7_75t_SL U27351 (.Y(n23692),
	.A(FE_OFN29081_n18526),
	.B(n23693));
   NOR2xp33_ASAP7_75t_L U27352 (.Y(n23695),
	.A(FE_OFN29140_n18527),
	.B(n23693));
   A2O1A1Ixp33_ASAP7_75t_SL U27353 (.Y(n23700),
	.A1(FE_OFN29139_n18527),
	.A2(FE_OFN29091_n),
	.B(n23698),
	.C(n18522));
   NOR3x1_ASAP7_75t_SL U27354 (.Y(n23781),
	.A(n23701),
	.B(n23719),
	.C(n23741));
   NAND2x1p5_ASAP7_75t_SL U27355 (.Y(n25628),
	.A(n23708),
	.B(n23707));
   OAI21xp33_ASAP7_75t_R U27356 (.Y(n23712),
	.A1(n18530),
	.A2(n23711),
	.B(n23710));
   OAI22xp33_ASAP7_75t_SRAM U27357 (.Y(n23722),
	.A1(n23869),
	.A2(n23719),
	.B1(FE_OFN29076_n18540),
	.B2(n23719));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27358 (.Y(n23737),
	.A1(FE_OFN16177_n27207),
	.A2(n27206),
	.B(FE_OCPN5166_n27203),
	.C(w2_9_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27359 (.Y(n373),
	.A1(FE_OFN16177_n27207),
	.A2(n27206),
	.B(n23738),
	.C(n23737));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27360 (.Y(n23743),
	.A1(n23838),
	.A2(n20670),
	.B(n23677),
	.C(FE_OCPN28246_n));
   NAND3xp33_ASAP7_75t_SRAM U27361 (.Y(n23751),
	.A(n18532),
	.B(FE_OFN29200_n18521),
	.C(FE_OCPN27542_sa20_3));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27364 (.Y(n23789),
	.A1(FE_OFN16176_n27207),
	.A2(n27192),
	.B(n27188),
	.C(w2_14_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27365 (.Y(n281),
	.A1(FE_OFN16176_n27207),
	.A2(n27192),
	.B(n23790),
	.C(n23789));
   NOR2xp33_ASAP7_75t_SRAM U27366 (.Y(n23794),
	.A(n23792),
	.B(n23791));
   NOR3xp33_ASAP7_75t_SRAM U27367 (.Y(n23796),
	.A(n25634),
	.B(n26900),
	.C(n23795));
   NAND3xp33_ASAP7_75t_R U27368 (.Y(n23807),
	.A(n23802),
	.B(n23801),
	.C(n23800));
   NOR2xp33_ASAP7_75t_SRAM U27369 (.Y(n23816),
	.A(FE_OFN29081_n18526),
	.B(n23814));
   NOR2xp33_ASAP7_75t_SRAM U27370 (.Y(n23822),
	.A(FE_OCPN27896_n18583),
	.B(n23823));
   NOR2xp33_ASAP7_75t_SRAM U27371 (.Y(n23824),
	.A(FE_OFN28776_n18532),
	.B(n23823));
   NOR3xp33_ASAP7_75t_R U27372 (.Y(n23834),
	.A(n23831),
	.B(n23830),
	.C(FE_OCPN28432_n23829));
   NOR2xp33_ASAP7_75t_L U27373 (.Y(n23836),
	.A(n23863),
	.B(n23835));
   OAI21xp33_ASAP7_75t_L U27374 (.Y(n25631),
	.A1(n23838),
	.A2(n23677),
	.B(n23836));
   NAND2xp5_ASAP7_75t_SL U27375 (.Y(n26898),
	.A(n23808),
	.B(n23847));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27376 (.Y(n23849),
	.A1(n27207),
	.A2(n23851),
	.B(FE_OCPN7621_n26898),
	.C(w2_10_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27377 (.Y(n297),
	.A1(n27207),
	.A2(n23851),
	.B(n23850),
	.C(n23849));
   NOR2xp33_ASAP7_75t_SRAM U27378 (.Y(n23854),
	.A(n18540),
	.B(n23855));
   NOR2xp33_ASAP7_75t_SRAM U27379 (.Y(n23858),
	.A(n23856),
	.B(n23855));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27381 (.Y(n23896),
	.A1(FE_OFN16177_n27207),
	.A2(n26057),
	.B(n26054),
	.C(w2_15_));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27382 (.Y(n374),
	.A1(FE_OFN16177_n27207),
	.A2(n26057),
	.B(n23897),
	.C(n23896));
   OAI22xp33_ASAP7_75t_SRAM U27383 (.Y(n23901),
	.A1(n23900),
	.A2(n23899),
	.B1(n23898),
	.B2(n23899));
   OAI22xp33_ASAP7_75t_R U27384 (.Y(n23923),
	.A1(n22405),
	.A2(n23903),
	.B1(n24289),
	.B2(n23903));
   NOR2xp33_ASAP7_75t_L U27385 (.Y(n23908),
	.A(n24844),
	.B(n23906));
   A2O1A1Ixp33_ASAP7_75t_L U27386 (.Y(n23914),
	.A1(n23916),
	.A2(FE_OFN16148_n25466),
	.B(n23913),
	.C(n23937));
   A2O1A1Ixp33_ASAP7_75t_L U27387 (.Y(n23918),
	.A1(FE_OFN16148_n25466),
	.A2(n23916),
	.B(n23915),
	.C(n23914));
   NAND3xp33_ASAP7_75t_L U27388 (.Y(n23917),
	.A(n23918),
	.B(n23920),
	.C(n23919));
   A2O1A1Ixp33_ASAP7_75t_SL U27389 (.Y(n23922),
	.A1(n23920),
	.A2(n23919),
	.B(n23918),
	.C(n23917));
   NAND3xp33_ASAP7_75t_L U27390 (.Y(n23921),
	.A(n23923),
	.B(n23924),
	.C(n23922));
   A2O1A1Ixp33_ASAP7_75t_SL U27391 (.Y(n23940),
	.A1(n23924),
	.A2(n23923),
	.B(n23922),
	.C(n23921));
   NOR3xp33_ASAP7_75t_SRAM U27392 (.Y(n23927),
	.A(n23926),
	.B(FE_OCPN29294_n23925),
	.C(n24881));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27393 (.Y(n23931),
	.A1(n23633),
	.A2(FE_OFN28820_n),
	.B(n16762),
	.C(n23927));
   O2A1O1Ixp5_ASAP7_75t_SL U27394 (.Y(n23932),
	.A1(n23931),
	.A2(n23930),
	.B(n26829),
	.C(n23968));
   A2O1A1Ixp33_ASAP7_75t_SL U27395 (.Y(n23934),
	.A1(n25044),
	.A2(FE_OCPN29586_n26857),
	.B(FE_OCPN29433_n25040),
	.C(FE_OCPN28437_n23932));
   A2O1A1Ixp33_ASAP7_75t_SL U27396 (.Y(n477),
	.A1(n23940),
	.A2(n25423),
	.B(n23939),
	.C(n23938));
   O2A1O1Ixp5_ASAP7_75t_SL U27397 (.Y(n23944),
	.A1(FE_OFN25937_n23943),
	.A2(n23942),
	.B(n25466),
	.C(n23941));
   NOR3xp33_ASAP7_75t_SRAM U27398 (.Y(n23964),
	.A(FE_OFN28971_n23947),
	.B(sa03_6_),
	.C(sa03_7_));
   NAND3xp33_ASAP7_75t_SRAM U27399 (.Y(n23957),
	.A(n23954),
	.B(n23956),
	.C(n23955));
   O2A1O1Ixp5_ASAP7_75t_SL U27400 (.Y(n23960),
	.A1(FE_OCPN5156_n23958),
	.A2(n23957),
	.B(n26857),
	.C(n25011));
   O2A1O1Ixp5_ASAP7_75t_SL U27401 (.Y(n23978),
	.A1(FE_OCPN5178_n25039),
	.A2(n23964),
	.B(FE_OCPN27446_n24847),
	.C(n23963));
   INVx1_ASAP7_75t_SL U27402 (.Y(n23967),
	.A(n23966));
   A2O1A1Ixp33_ASAP7_75t_L U27403 (.Y(n23969),
	.A1(n26829),
	.A2(n23971),
	.B(n23968),
	.C(n23967));
   A2O1A1Ixp33_ASAP7_75t_SL U27404 (.Y(n25437),
	.A1(n26829),
	.A2(n23971),
	.B(n23970),
	.C(n23969));
   AOI22xp33_ASAP7_75t_SL U27406 (.Y(n23977),
	.A1(FE_OCPN27282_n25437),
	.A2(FE_OFN16421_n23974),
	.B1(FE_OFN51_w3_18),
	.B2(n23972));
   A2O1A1Ixp33_ASAP7_75t_SL U27407 (.Y(n428),
	.A1(n23978),
	.A2(n23977),
	.B(n23976),
	.C(n23975));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27408 (.Y(n23983),
	.A1(n23982),
	.A2(n23981),
	.B(FE_OFN25956_n16575),
	.C(n23979));
   NAND3xp33_ASAP7_75t_SRAM U27409 (.Y(n24004),
	.A(n23994),
	.B(n23993),
	.C(n23992));
   O2A1O1Ixp33_ASAP7_75t_SL U27410 (.Y(n26336),
	.A1(n24005),
	.A2(n24004),
	.B(n24974),
	.C(n24003));
   NOR2xp33_ASAP7_75t_SRAM U27411 (.Y(n24013),
	.A(n25354),
	.B(sa21_6_));
   NOR2xp33_ASAP7_75t_L U27412 (.Y(n24015),
	.A(n24014),
	.B(sa21_6_));
   A2O1A1Ixp33_ASAP7_75t_L U27413 (.Y(n24018),
	.A1(n26819),
	.A2(n26725),
	.B(n26722),
	.C(FE_OFN16278_w3_5));
   O2A1O1Ixp5_ASAP7_75t_SL U27414 (.Y(n24023),
	.A1(FE_OCPN27226_n25357),
	.A2(n24659),
	.B(n24021),
	.C(n24020));
   A2O1A1Ixp33_ASAP7_75t_SL U27415 (.Y(n24029),
	.A1(FE_OCPN29539_n24927),
	.A2(n24024),
	.B(n24023),
	.C(n24022));
   A2O1A1Ixp33_ASAP7_75t_SL U27416 (.Y(n457),
	.A1(FE_OCPN27505_n24684),
	.A2(n24029),
	.B(n24028),
	.C(n24027));
   A2O1A1Ixp33_ASAP7_75t_L U27417 (.Y(n24035),
	.A1(n24038),
	.A2(n24037),
	.B(FE_OCPN27772_n24234),
	.C(n24034));
   NAND3xp33_ASAP7_75t_SL U27419 (.Y(n24043),
	.A(n24041),
	.B(n24040),
	.C(FE_OFN26032_n20230));
   NAND3xp33_ASAP7_75t_SRAM U27420 (.Y(n24050),
	.A(n24048),
	.B(n24047),
	.C(n24046));
   NOR2xp33_ASAP7_75t_SRAM U27421 (.Y(n24054),
	.A(FE_OCPN28386_n17899),
	.B(n24055));
   A2O1A1Ixp33_ASAP7_75t_L U27422 (.Y(n24066),
	.A1(n26679),
	.A2(n26678),
	.B(FE_OCPN28279_n),
	.C(w1_22_));
   A2O1A1Ixp33_ASAP7_75t_SL U27423 (.Y(n24071),
	.A1(FE_OCPN28023_n25770),
	.A2(FE_OCPN27815_n25769),
	.B(n24069),
	.C(n24068));
   A2O1A1Ixp33_ASAP7_75t_L U27424 (.Y(n24076),
	.A1(FE_OCPN5107_n24418),
	.A2(n24147),
	.B(n24071),
	.C(n24070));
   OAI21xp5_ASAP7_75t_L U27425 (.Y(n24075),
	.A1(n24076),
	.A2(FE_OCPN28077_n),
	.B(FE_OFN28486_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27426 (.Y(n489),
	.A1(FE_OCPN28077_n),
	.A2(n24076),
	.B(n24075),
	.C(n24074));
   NOR3xp33_ASAP7_75t_SRAM U27428 (.Y(n24082),
	.A(n24080),
	.B(n24079),
	.C(n24078));
   NAND3xp33_ASAP7_75t_SRAM U27429 (.Y(n24088),
	.A(n24085),
	.B(FE_OFN28767_n26103),
	.C(n24084));
   NOR3xp33_ASAP7_75t_L U27430 (.Y(n24091),
	.A(n24088),
	.B(FE_PSN8273_n24087),
	.C(n24086));
   NAND3xp33_ASAP7_75t_SL U27432 (.Y(n24095),
	.A(n24092),
	.B(n24091),
	.C(n24090));
   NOR2xp33_ASAP7_75t_SRAM U27433 (.Y(n24098),
	.A(n24097),
	.B(n24096));
   NAND3xp33_ASAP7_75t_SL U27434 (.Y(n24104),
	.A(FE_OFN16392_n24102),
	.B(n24101),
	.C(n25258));
   NOR2xp67_ASAP7_75t_SL U27435 (.Y(n24106),
	.A(w0_18_),
	.B(n26771));
   A2O1A1Ixp33_ASAP7_75t_SL U27436 (.Y(n24111),
	.A1(FE_OFN16263_n25976),
	.A2(n24109),
	.B(n24108),
	.C(n24107));
   A2O1A1Ixp33_ASAP7_75t_L U27437 (.Y(n26093),
	.A1(n26770),
	.A2(n26769),
	.B(n24116),
	.C(n24115));
   OAI22xp33_ASAP7_75t_SRAM U27438 (.Y(n24117),
	.A1(text_in_r_114_),
	.A2(FE_OFN28484_ld_r),
	.B1(n24118),
	.B2(FE_OFN28484_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27439 (.Y(n391),
	.A1(n24121),
	.A2(FE_OCPN27941_n),
	.B(n24120),
	.C(n24119));
   NAND2x1p5_ASAP7_75t_SL U27440 (.Y(n26467),
	.A(n25769),
	.B(n25770));
   A2O1A1Ixp33_ASAP7_75t_L U27441 (.Y(n24124),
	.A1(n26282),
	.A2(n24126),
	.B(n24123),
	.C(n26466));
   A2O1A1Ixp33_ASAP7_75t_SL U27442 (.Y(n25483),
	.A1(n26282),
	.A2(n24126),
	.B(n24125),
	.C(n24124));
   NOR3xp33_ASAP7_75t_SL U27443 (.Y(n24143),
	.A(FE_OCPN7620_n25761),
	.B(n24144),
	.C(FE_OCPN5119_n25762));
   O2A1O1Ixp5_ASAP7_75t_SL U27444 (.Y(n24146),
	.A1(FE_OCPN7620_n25761),
	.A2(FE_OCPN5119_n25762),
	.B(n24144),
	.C(n24143));
   NAND3xp33_ASAP7_75t_SL U27445 (.Y(n24145),
	.A(n24146),
	.B(FE_OCPN5107_n24418),
	.C(n24147));
   A2O1A1Ixp33_ASAP7_75t_SL U27446 (.Y(n24152),
	.A1(FE_OCPN5107_n24418),
	.A2(n24147),
	.B(n24146),
	.C(n24145));
   OAI21xp5_ASAP7_75t_SL U27447 (.Y(n24151),
	.A1(n24152),
	.A2(FE_OCPN27467_n25483),
	.B(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27448 (.Y(n492),
	.A1(FE_OCPN27467_n25483),
	.A2(n24152),
	.B(n24151),
	.C(n24150));
   NOR2xp33_ASAP7_75t_SRAM U27449 (.Y(n24158),
	.A(n24156),
	.B(FE_OFN28919_n24155));
   NAND3xp33_ASAP7_75t_SL U27450 (.Y(n24168),
	.A(n24166),
	.B(n24165),
	.C(n24164));
   O2A1O1Ixp5_ASAP7_75t_SL U27451 (.Y(n24170),
	.A1(n24169),
	.A2(n24168),
	.B(n26915),
	.C(n24167));
   NOR2x1_ASAP7_75t_SL U27453 (.Y(n24174),
	.A(n26235),
	.B(n26236));
   A2O1A1Ixp33_ASAP7_75t_SL U27454 (.Y(n24176),
	.A1(n27183),
	.A2(n24178),
	.B(n24175),
	.C(n24174));
   NOR3xp33_ASAP7_75t_R U27455 (.Y(n24179),
	.A(FE_OCPN5053_n25832),
	.B(FE_OCPN7589_n26420),
	.C(n25831));
   NOR2xp33_ASAP7_75t_SRAM U27456 (.Y(n24183),
	.A(n24181),
	.B(n24184));
   NOR2xp33_ASAP7_75t_SRAM U27457 (.Y(n24186),
	.A(FE_OFN27043_n),
	.B(n24184));
   NAND2xp5_ASAP7_75t_R U27458 (.Y(n24196),
	.A(FE_OFN25911_n26491),
	.B(n24200));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27459 (.Y(n24195),
	.A1(n27216),
	.A2(n26494),
	.B(FE_OCPN28307_n26491),
	.C(w2_5_));
   A2O1A1Ixp33_ASAP7_75t_L U27460 (.Y(n24198),
	.A1(n27216),
	.A2(n26494),
	.B(n24196),
	.C(n24195));
   O2A1O1Ixp33_ASAP7_75t_L U27461 (.Y(n24203),
	.A1(FE_OCPN5077_n25855),
	.A2(n25856),
	.B(n24198),
	.C(n24197));
   A2O1A1Ixp33_ASAP7_75t_SL U27462 (.Y(n475),
	.A1(n24204),
	.A2(n24203),
	.B(n24202),
	.C(n24201));
   A2O1A1Ixp33_ASAP7_75t_SL U27463 (.Y(n24212),
	.A1(n26139),
	.A2(n24214),
	.B(n25485),
	.C(n24211));
   OAI22xp5_ASAP7_75t_L U27464 (.Y(n24223),
	.A1(n24222),
	.A2(n27004),
	.B1(n24221),
	.B2(n27004));
   O2A1O1Ixp5_ASAP7_75t_SL U27465 (.Y(n24433),
	.A1(n24228),
	.A2(n24227),
	.B(n26679),
	.C(n24226));
   A2O1A1Ixp33_ASAP7_75t_L U27466 (.Y(n24231),
	.A1(FE_OFN16164_n25081),
	.A2(n24422),
	.B(n24421),
	.C(n24230));
   A2O1A1Ixp33_ASAP7_75t_SL U27467 (.Y(n25768),
	.A1(FE_OFN16164_n25081),
	.A2(n24422),
	.B(n24232),
	.C(n24231));
   NOR3xp33_ASAP7_75t_R U27468 (.Y(n24233),
	.A(FE_OCPN27772_n24234),
	.B(FE_OCPN27421_n25768),
	.C(FE_OFN28495_n24584));
   O2A1O1Ixp5_ASAP7_75t_SL U27469 (.Y(n24239),
	.A1(FE_OCPN27772_n24234),
	.A2(FE_OFN28495_n24584),
	.B(FE_OCPN27421_n25768),
	.C(n24233));
   A2O1A1Ixp33_ASAP7_75t_L U27470 (.Y(n511),
	.A1(n24240),
	.A2(n24239),
	.B(n24238),
	.C(n24237));
   NOR3xp33_ASAP7_75t_SRAM U27472 (.Y(n24246),
	.A(n24244),
	.B(n24243),
	.C(FE_OFN16398_n24241));
   NAND3xp33_ASAP7_75t_R U27473 (.Y(n24248),
	.A(n24247),
	.B(n24246),
	.C(n24245));
   O2A1O1Ixp33_ASAP7_75t_SL U27474 (.Y(n25383),
	.A1(FE_OFN28922_n24249),
	.A2(n24248),
	.B(n26819),
	.C(FE_OFN16316_n24840));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27475 (.Y(n24250),
	.A1(n26857),
	.A2(n19640),
	.B(FE_OCPN27478_n25011),
	.C(FE_OCPN27538_n25383));
   O2A1O1Ixp33_ASAP7_75t_SL U27476 (.Y(n24274),
	.A1(n24267),
	.A2(n24266),
	.B(n26829),
	.C(n24265));
   NOR3xp33_ASAP7_75t_SRAM U27477 (.Y(n24280),
	.A(n24279),
	.B(n24278),
	.C(n24277));
   A2O1A1Ixp33_ASAP7_75t_SL U27478 (.Y(n24284),
	.A1(n22405),
	.A2(n26842),
	.B(n26839),
	.C(n24283));
   A2O1A1Ixp33_ASAP7_75t_SL U27479 (.Y(n26796),
	.A1(n22405),
	.A2(FE_OCPN27940_n26842),
	.B(n24285),
	.C(n24284));
   A2O1A1Ixp33_ASAP7_75t_R U27480 (.Y(n24287),
	.A1(n24289),
	.A2(n22405),
	.B(FE_OCPN5073_n24996),
	.C(FE_OFN27111_n));
   A2O1A1Ixp33_ASAP7_75t_L U27481 (.Y(n24290),
	.A1(n22405),
	.A2(n24289),
	.B(n24288),
	.C(n24287));
   OAI22xp33_ASAP7_75t_SRAM U27482 (.Y(n24291),
	.A1(text_in_r_9_),
	.A2(FE_OFN28489_ld_r),
	.B1(FE_OFN27111_n),
	.B2(FE_OFN28489_ld_r));
   NOR2xp33_ASAP7_75t_SRAM U27483 (.Y(n24308),
	.A(FE_OFN44_w0_9),
	.B(FE_OCPN28024_n26427));
   A2O1A1Ixp33_ASAP7_75t_L U27484 (.Y(n24313),
	.A1(n27117),
	.A2(FE_PSN8300_n26482),
	.B(n24312),
	.C(n24311));
   FAx1_ASAP7_75t_SL U27485 (.SN(n24323),
	.A(FE_OCPN28123_n27047),
	.B(n24314),
	.CI(n24313));
   NOR2x1_ASAP7_75t_SL U27486 (.Y(n24318),
	.A(n24315),
	.B(FE_OFN28934_n24552));
   OAI22xp33_ASAP7_75t_SRAM U27487 (.Y(n24319),
	.A1(text_in_r_105_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(n24320),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27488 (.Y(n456),
	.A1(n24323),
	.A2(FE_OCPN27310_n26389),
	.B(n24322),
	.C(n24321));
   O2A1O1Ixp5_ASAP7_75t_SL U27489 (.Y(n27152),
	.A1(n24335),
	.A2(n24334),
	.B(n26770),
	.C(n24333));
   O2A1O1Ixp5_ASAP7_75t_SL U27490 (.Y(n27153),
	.A1(n24339),
	.A2(n24338),
	.B(n24610),
	.C(n24337));
   A2O1A1Ixp33_ASAP7_75t_L U27491 (.Y(n24342),
	.A1(n27117),
	.A2(n27116),
	.B(FE_OFN29010_n27113),
	.C(n24341));
   A2O1A1Ixp33_ASAP7_75t_SL U27492 (.Y(n24491),
	.A1(n27117),
	.A2(n27116),
	.B(n24343),
	.C(n24342));
   OAI222xp33_ASAP7_75t_R U27493 (.Y(n24354),
	.A1(n25795),
	.A2(n17506),
	.B1(n24349),
	.B2(n17506),
	.C1(n25794),
	.C2(n17506));
   A2O1A1Ixp33_ASAP7_75t_SL U27494 (.Y(n24350),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(FE_OCPN27744_n26362),
	.C(FE_OFN39_w0_21));
   O2A1O1Ixp5_ASAP7_75t_SL U27495 (.Y(n24356),
	.A1(FE_OCPN27357_n26369),
	.A2(n24354),
	.B(n24353),
	.C(n24352));
   A2O1A1Ixp33_ASAP7_75t_SL U27496 (.Y(n24361),
	.A1(FE_OCPN28235_n26631),
	.A2(n24502),
	.B(n24356),
	.C(n24355));
   OAI22xp33_ASAP7_75t_SRAM U27497 (.Y(n24357),
	.A1(text_in_r_117_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(n24358),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27498 (.Y(n458),
	.A1(FE_OCPN27412_n24491),
	.A2(n24361),
	.B(n24360),
	.C(n24359));
   OAI22xp33_ASAP7_75t_SRAM U27499 (.Y(n24366),
	.A1(n24364),
	.A2(n24363),
	.B1(FE_OCPN27729_n24362),
	.B2(n24363));
   NOR2xp33_ASAP7_75t_SRAM U27500 (.Y(n24369),
	.A(n24367),
	.B(n24370));
   NOR2xp33_ASAP7_75t_R U27501 (.Y(n24372),
	.A(n17906),
	.B(n24370));
   O2A1O1Ixp33_ASAP7_75t_SRAM U27502 (.Y(n24388),
	.A1(n24381),
	.A2(n24380),
	.B(n26139),
	.C(n24379));
   A2O1A1Ixp33_ASAP7_75t_SL U27504 (.Y(n26285),
	.A1(n24388),
	.A2(n24387),
	.B(n25688),
	.C(n24386));
   NAND3xp33_ASAP7_75t_SRAM U27505 (.Y(n24394),
	.A(FE_OFN28590_n24391),
	.B(n24390),
	.C(n24389));
   NOR3xp33_ASAP7_75t_SRAM U27506 (.Y(n24397),
	.A(n24394),
	.B(n24393),
	.C(n24392));
   OA222x2_ASAP7_75t_SRAM U27507 (.Y(n24400),
	.A1(n24397),
	.A2(n27015),
	.B1(n24396),
	.B2(n27015),
	.C1(n24395),
	.C2(n27015));
   NOR2xp33_ASAP7_75t_SRAM U27508 (.Y(n24401),
	.A(FE_OCPN29352_n25173),
	.B(n24399));
   NAND2xp33_ASAP7_75t_SRAM U27509 (.Y(n24407),
	.A(w1_18_),
	.B(n27023));
   A2O1A1Ixp33_ASAP7_75t_R U27510 (.Y(n24406),
	.A1(FE_OFN28506_n26996),
	.A2(FE_OFN16169_n26567),
	.B(FE_OFN28512_n27020),
	.C(n24412));
   A2O1A1Ixp33_ASAP7_75t_SL U27511 (.Y(n24415),
	.A1(n24410),
	.A2(n24405),
	.B(n24409),
	.C(n24408));
   OAI22xp33_ASAP7_75t_SRAM U27512 (.Y(n24411),
	.A1(text_in_r_82_),
	.A2(FE_OFN28487_ld_r),
	.B1(n24412),
	.B2(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27513 (.Y(n393),
	.A1(n26285),
	.A2(n24415),
	.B(n24414),
	.C(n24413));
   NAND2xp33_ASAP7_75t_SRAM U27515 (.Y(n24429),
	.A(w1_21_),
	.B(FE_OFN26148_n26245));
   A2O1A1Ixp33_ASAP7_75t_R U27516 (.Y(n24428),
	.A1(n26248),
	.A2(n26249),
	.B(FE_OFN26149_n26245),
	.C(n24435));
   A2O1A1Ixp33_ASAP7_75t_L U27517 (.Y(n24431),
	.A1(n26249),
	.A2(n26248),
	.B(n24429),
	.C(n24428));
   A2O1A1Ixp33_ASAP7_75t_L U27518 (.Y(n24438),
	.A1(n24433),
	.A2(n24432),
	.B(n24431),
	.C(n24430));
   OAI21xp5_ASAP7_75t_R U27519 (.Y(n24437),
	.A1(n24438),
	.A2(n26472),
	.B(FE_OFN28487_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U27520 (.Y(n24434),
	.A1(text_in_r_85_),
	.A2(FE_OFN28487_ld_r),
	.B1(n24435),
	.B2(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27521 (.Y(n483),
	.A1(FE_OCPN8238_n26472),
	.A2(n24438),
	.B(n24437),
	.C(n24436));
   NOR2xp33_ASAP7_75t_SRAM U27522 (.Y(n24439),
	.A(n24834),
	.B(sa03_6_));
   NOR3xp33_ASAP7_75t_SRAM U27523 (.Y(n24442),
	.A(n24441),
	.B(n24440),
	.C(n24839));
   NOR2xp33_ASAP7_75t_SL U27524 (.Y(n24444),
	.A(n24442),
	.B(sa03_6_));
   NOR3xp33_ASAP7_75t_SL U27525 (.Y(n24447),
	.A(n24837),
	.B(FE_OCPN28131_n26796),
	.C(n24448));
   A2O1A1Ixp33_ASAP7_75t_L U27526 (.Y(n24451),
	.A1(FE_OCPN29587_n26857),
	.A2(FE_OFN29242_n26856),
	.B(FE_OCPN27377_n26853),
	.C(n24450));
   NAND3xp33_ASAP7_75t_SL U27527 (.Y(n24453),
	.A(FE_OFN28489_ld_r),
	.B(n24454),
	.C(n25390));
   NOR3xp33_ASAP7_75t_SRAM U27529 (.Y(n24462),
	.A(n24460),
	.B(n24459),
	.C(n24458));
   NAND3xp33_ASAP7_75t_SRAM U27530 (.Y(n24463),
	.A(n24964),
	.B(n24462),
	.C(n24461));
   OAI21xp33_ASAP7_75t_SRAM U27531 (.Y(n24465),
	.A1(n24901),
	.A2(n24463),
	.B(n26857));
   NAND3xp33_ASAP7_75t_SL U27532 (.Y(n24464),
	.A(n25041),
	.B(n24465),
	.C(FE_OCPN27282_n25437));
   A2O1A1Ixp33_ASAP7_75t_SL U27533 (.Y(n24467),
	.A1(n24465),
	.A2(n25041),
	.B(FE_OCPN27282_n25437),
	.C(n24464));
   A2O1A1Ixp33_ASAP7_75t_SL U27534 (.Y(n24472),
	.A1(n24468),
	.A2(FE_OFN28490_ld_r),
	.B(n24467),
	.C(n24466));
   NAND3xp33_ASAP7_75t_SL U27535 (.Y(n24469),
	.A(n24470),
	.B(n24472),
	.C(n24471));
   A2O1A1Ixp33_ASAP7_75t_SL U27536 (.Y(n411),
	.A1(n24472),
	.A2(n24471),
	.B(n24470),
	.C(n24469));
   A2O1A1Ixp33_ASAP7_75t_L U27537 (.Y(n24481),
	.A1(n27062),
	.A2(n27061),
	.B(n27058),
	.C(FE_OFN28963_n24480));
   O2A1O1Ixp5_ASAP7_75t_SL U27538 (.Y(n24493),
	.A1(FE_OCPN29481_n26537),
	.A2(n25610),
	.B(FE_OCPN27412_n24491),
	.C(n24490));
   A2O1A1Ixp33_ASAP7_75t_L U27539 (.Y(n24498),
	.A1(n27117),
	.A2(n27052),
	.B(FE_OFN29142_n27049),
	.C(w0_6_));
   A2O1A1Ixp33_ASAP7_75t_L U27540 (.Y(n24504),
	.A1(n24502),
	.A2(FE_OCPN28235_n26631),
	.B(n24501),
	.C(n24500));
   A2O1A1Ixp33_ASAP7_75t_SL U27541 (.Y(n24509),
	.A1(FE_OCPN28173_n27153),
	.A2(FE_OCPN28150_n27152),
	.B(n24504),
	.C(n24503));
   A2O1A1Ixp33_ASAP7_75t_SL U27542 (.Y(n521),
	.A1(FE_OCPN27379_n26809),
	.A2(n24509),
	.B(n24508),
	.C(n24507));
   A2O1A1Ixp33_ASAP7_75t_SL U27543 (.Y(n24512),
	.A1(n26082),
	.A2(n24633),
	.B(n24630),
	.C(n24511));
   NOR3xp33_ASAP7_75t_SRAM U27544 (.Y(n24519),
	.A(n24518),
	.B(n24517),
	.C(FE_OFN28556_n24516));
   NOR2xp33_ASAP7_75t_R U27545 (.Y(n24520),
	.A(n24519),
	.B(FE_OFN28499_sa00_6));
   A2O1A1Ixp33_ASAP7_75t_SL U27546 (.Y(n24524),
	.A1(n27127),
	.A2(FE_OCPN7622_n24526),
	.B(FE_OCPN27402_n24523),
	.C(n24537));
   NOR3xp33_ASAP7_75t_R U27547 (.Y(n24527),
	.A(n24529),
	.B(FE_OCPN27514_n25981),
	.C(n24528));
   A2O1A1Ixp33_ASAP7_75t_SL U27548 (.Y(n479),
	.A1(n24535),
	.A2(n24534),
	.B(n24533),
	.C(n24532));
   A2O1A1Ixp33_ASAP7_75t_L U27549 (.Y(n24538),
	.A1(n27117),
	.A2(FE_OFN28690_n25979),
	.B(n25974),
	.C(FE_OCPN29263_n24537));
   A2O1A1Ixp33_ASAP7_75t_L U27550 (.Y(n24639),
	.A1(n27117),
	.A2(FE_OFN28690_n25979),
	.B(n24539),
	.C(n24538));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27551 (.Y(n24541),
	.A1(n24543),
	.A2(n27127),
	.B(FE_OCPN27314_n26113),
	.C(n24575));
   O2A1O1Ixp5_ASAP7_75t_SL U27552 (.Y(n25971),
	.A1(n24551),
	.A2(n24550),
	.B(n27062),
	.C(n26735));
   FAx1_ASAP7_75t_SL U27553 (.SN(n24578),
	.A(FE_OCPN29365_n24639),
	.B(n24558),
	.CI(n24557));
   NAND3xp33_ASAP7_75t_R U27554 (.Y(n24563),
	.A(n25787),
	.B(n24560),
	.C(n24559));
   NOR2x1p5_ASAP7_75t_L U27556 (.Y(n25967),
	.A(n26267),
	.B(n26268));
   A2O1A1Ixp33_ASAP7_75t_SL U27557 (.Y(n24572),
	.A1(n27127),
	.A2(n25255),
	.B(n27056),
	.C(n25967));
   A2O1A1Ixp33_ASAP7_75t_SL U27558 (.Y(n352),
	.A1(n24578),
	.A2(FE_OCPN29540_FE_OFN25927_n26527),
	.B(n24577),
	.C(n24576));
   A2O1A1Ixp33_ASAP7_75t_SL U27559 (.Y(n24582),
	.A1(n26679),
	.A2(n25172),
	.B(FE_OCPN27825_n25169),
	.C(n24809));
   NAND3xp33_ASAP7_75t_SRAM U27560 (.Y(n24588),
	.A(n24587),
	.B(n24586),
	.C(n24585));
   A2O1A1Ixp33_ASAP7_75t_SL U27561 (.Y(n24595),
	.A1(FE_OFN16169_n26567),
	.A2(n24812),
	.B(n26683),
	.C(w1_23_));
   O2A1O1Ixp33_ASAP7_75t_SL U27562 (.Y(n24600),
	.A1(FE_OCPN27723_n),
	.A2(n25484),
	.B(n24598),
	.C(n24597));
   A2O1A1Ixp33_ASAP7_75t_SL U27563 (.Y(n24605),
	.A1(n24602),
	.A2(n24601),
	.B(n24600),
	.C(n24599));
   NOR2x1p5_ASAP7_75t_L U27564 (.Y(n27031),
	.A(FE_OFN16213_ld_r),
	.B(n25407));
   A2O1A1Ixp33_ASAP7_75t_L U27566 (.Y(n24606),
	.A1(n27034),
	.A2(FE_OFN28486_ld_r),
	.B(n24605),
	.C(n24604));
   A2O1A1Ixp33_ASAP7_75t_SL U27567 (.Y(n486),
	.A1(text_in_r_87_),
	.A2(n24608),
	.B(n24607),
	.C(n24606));
   O2A1O1Ixp5_ASAP7_75t_SRAM U27568 (.Y(n24636),
	.A1(n24612),
	.A2(n24611),
	.B(n24610),
	.C(n24609));
   OAI22xp33_ASAP7_75t_SRAM U27569 (.Y(n24615),
	.A1(FE_OCPN27555_n16422),
	.A2(n24613),
	.B1(FE_OFN28592_n16427),
	.B2(n24613));
   NAND2xp33_ASAP7_75t_SRAM U27570 (.Y(n24616),
	.A(n24615),
	.B(n24614));
   NOR3xp33_ASAP7_75t_R U27571 (.Y(n24620),
	.A(n24618),
	.B(n24617),
	.C(n24616));
   NAND3xp33_ASAP7_75t_SRAM U27572 (.Y(n24623),
	.A(FE_OFN25940_n24621),
	.B(n24620),
	.C(n24619));
   A2O1A1Ixp33_ASAP7_75t_SL U27573 (.Y(n24719),
	.A1(n26082),
	.A2(n24633),
	.B(n24632),
	.C(n24631));
   NAND3xp33_ASAP7_75t_SRAM U27574 (.Y(n24650),
	.A(n24646),
	.B(FE_OFN26553_n24644),
	.C(n24645));
   O2A1O1Ixp5_ASAP7_75t_SL U27575 (.Y(n24652),
	.A1(n24650),
	.A2(n24649),
	.B(n22405),
	.C(n25470));
   A2O1A1Ixp33_ASAP7_75t_SL U27576 (.Y(n24655),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(FE_OCPN28106_FE_OFN25876_n25462),
	.C(FE_OFN34_w3_22));
   A2O1A1Ixp33_ASAP7_75t_SL U27577 (.Y(n24658),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(n24656),
	.C(n24655));
   O2A1O1Ixp33_ASAP7_75t_SL U27578 (.Y(n24661),
	.A1(FE_OCPN27226_n25357),
	.A2(n24659),
	.B(n24658),
	.C(n24657));
   A2O1A1Ixp33_ASAP7_75t_SL U27579 (.Y(n24666),
	.A1(FE_OCPN27991_n26336),
	.A2(FE_OCPN28110_n),
	.B(n24661),
	.C(n24660));
   OAI22xp33_ASAP7_75t_SRAM U27580 (.Y(n24662),
	.A1(text_in_r_22_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(FE_OFN7_w3_22),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U27581 (.Y(n24668),
	.A1(n24729),
	.A2(n25139),
	.B1(n24667),
	.B2(n25139));
   NOR2xp33_ASAP7_75t_SRAM U27582 (.Y(n24670),
	.A(n24669),
	.B(FE_OFN59_sa10_7));
   AND2x2_ASAP7_75t_SRAM U27583 (.Y(n24679),
	.A(n24675),
	.B(n24674));
   NAND3xp33_ASAP7_75t_SL U27584 (.Y(n24683),
	.A(n26822),
	.B(n26823),
	.C(n24684));
   NOR2xp33_ASAP7_75t_SRAM U27585 (.Y(n24693),
	.A(n24691),
	.B(n24694));
   NOR2xp33_ASAP7_75t_SRAM U27586 (.Y(n24696),
	.A(n18162),
	.B(n24694));
   NAND2xp33_ASAP7_75t_SRAM U27587 (.Y(n24703),
	.A(n26872),
	.B(n24702));
   NOR2xp33_ASAP7_75t_SL U27589 (.Y(n24709),
	.A(n26765),
	.B(FE_OFN25973_n26087));
   O2A1O1Ixp33_ASAP7_75t_SL U27590 (.Y(n24708),
	.A1(n26542),
	.A2(n18158),
	.B(n26088),
	.C(FE_OFN29039_n26763));
   O2A1O1Ixp33_ASAP7_75t_SL U27591 (.Y(n26227),
	.A1(FE_OFN16180_n26542),
	.A2(n18158),
	.B(n24709),
	.C(n24708));
   NAND3xp33_ASAP7_75t_SRAM U27592 (.Y(n24712),
	.A(n24710),
	.B(n26064),
	.C(n26071));
   NOR3xp33_ASAP7_75t_R U27593 (.Y(n24717),
	.A(n24712),
	.B(n24711),
	.C(n26076));
   O2A1O1Ixp5_ASAP7_75t_SL U27594 (.Y(n24718),
	.A1(n17506),
	.A2(n24717),
	.B(n24716),
	.C(n24715));
   FAx1_ASAP7_75t_SL U27595 (.SN(n24724),
	.A(FE_OCPN27361_n24719),
	.B(FE_OCPN29460_n26227),
	.CI(n24718));
   A2O1A1Ixp33_ASAP7_75t_SL U27596 (.Y(n451),
	.A1(n24724),
	.A2(FE_OCPN29540_FE_OFN25927_n26527),
	.B(n24723),
	.C(n24722));
   O2A1O1Ixp33_ASAP7_75t_L U27597 (.Y(n25953),
	.A1(n24732),
	.A2(n24731),
	.B(n26857),
	.C(n24730));
   O2A1O1Ixp33_ASAP7_75t_SL U27598 (.Y(n25954),
	.A1(FE_OCPN5158_n24742),
	.A2(n24741),
	.B(n24974),
	.C(n24740));
   NAND2xp33_ASAP7_75t_SRAM U27599 (.Y(n24748),
	.A(n24925),
	.B(FE_OCPN29520_n24755));
   A2O1A1Ixp33_ASAP7_75t_L U27600 (.Y(n24747),
	.A1(n22405),
	.A2(n24930),
	.B(FE_OCPN29538_n24927),
	.C(FE_OFN102_w3_12));
   NOR2xp33_ASAP7_75t_L U27601 (.Y(n24752),
	.A(n25133),
	.B(n25667));
   O2A1O1Ixp33_ASAP7_75t_SL U27602 (.Y(n24751),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25669),
	.C(n25134));
   O2A1O1Ixp5_ASAP7_75t_SL U27603 (.Y(n25422),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n24752),
	.C(n24751));
   OAI22xp33_ASAP7_75t_SRAM U27605 (.Y(n24754),
	.A1(text_in_r_12_),
	.A2(FE_OFN28489_ld_r),
	.B1(FE_OCPN29520_n24755),
	.B2(FE_OFN28489_ld_r));
   NAND3xp33_ASAP7_75t_SRAM U27606 (.Y(n24763),
	.A(n24760),
	.B(n25104),
	.C(n24759));
   OA21x2_ASAP7_75t_SRAM U27607 (.Y(n24770),
	.A1(n22010),
	.A2(FE_OCPN27288_n25091),
	.B(n24766));
   NOR2xp33_ASAP7_75t_L U27608 (.Y(n24771),
	.A(FE_OFN28787_n19000),
	.B(n24769));
   NOR2xp33_ASAP7_75t_SRAM U27609 (.Y(n24778),
	.A(n25108),
	.B(n24779));
   NAND3xp33_ASAP7_75t_SRAM U27610 (.Y(n24788),
	.A(n24787),
	.B(n24786),
	.C(n24785));
   NOR2x1_ASAP7_75t_R U27611 (.Y(n24806),
	.A(n24803),
	.B(FE_OFN28451_n26990));
   A2O1A1Ixp33_ASAP7_75t_SL U27615 (.Y(n24810),
	.A1(FE_OFN16169_n26567),
	.A2(n24812),
	.B(n26683),
	.C(n24809));
   A2O1A1Ixp33_ASAP7_75t_R U27616 (.Y(n24813),
	.A1(FE_OFN16163_n26584),
	.A2(n26183),
	.B(n26180),
	.C(w1_9_));
   A2O1A1Ixp33_ASAP7_75t_SL U27617 (.Y(n24815),
	.A1(FE_OFN16163_n26584),
	.A2(n26183),
	.B(n24814),
	.C(n24813));
   FAx1_ASAP7_75t_SL U27618 (.SN(n24824),
	.A(FE_OFN16227_n26602),
	.B(FE_OCPN29531_FE_OFN25926_n26922),
	.CI(n24815));
   A2O1A1Ixp33_ASAP7_75t_SL U27619 (.Y(n27030),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(n24819),
	.C(n24818));
   A2O1A1Ixp33_ASAP7_75t_L U27620 (.Y(n433),
	.A1(n24824),
	.A2(FE_OCPN27439_n27030),
	.B(n24823),
	.C(n24822));
   OAI22xp33_ASAP7_75t_SRAM U27621 (.Y(n24851),
	.A1(FE_OCPN27985_n24831),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_1_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27622 (.Y(n24828),
	.A1(n17580),
	.A2(n24830),
	.B(FE_OCPN27491_n26351),
	.C(n24827));
   A2O1A1Ixp33_ASAP7_75t_L U27623 (.Y(n24832),
	.A1(n22405),
	.A2(FE_OCPN27940_n26842),
	.B(n26839),
	.C(FE_OFN16423_n24831));
   NAND3xp33_ASAP7_75t_SL U27624 (.Y(n24838),
	.A(FE_OFN26001_n24836),
	.B(n24835),
	.C(n24834));
   O2A1O1Ixp5_ASAP7_75t_SL U27625 (.Y(n25007),
	.A1(n24839),
	.A2(n24838),
	.B(n26819),
	.C(FE_OFN95_n19498));
   A2O1A1Ixp33_ASAP7_75t_SL U27626 (.Y(n24842),
	.A1(n24844),
	.A2(n26819),
	.B(FE_OFN28578_FE_OFN16316_n24840),
	.C(n25006));
   A2O1A1Ixp33_ASAP7_75t_SL U27627 (.Y(n24845),
	.A1(n26819),
	.A2(FE_OCPN8239_n24844),
	.B(n24843),
	.C(n24842));
   NAND3xp33_ASAP7_75t_SRAM U27629 (.Y(n24875),
	.A(n24854),
	.B(n24853),
	.C(n24852));
   NOR3xp33_ASAP7_75t_R U27631 (.Y(n24865),
	.A(n24864),
	.B(n24863),
	.C(n24862));
   NAND3xp33_ASAP7_75t_R U27632 (.Y(n24870),
	.A(n24867),
	.B(n24866),
	.C(n24865));
   NAND3xp33_ASAP7_75t_R U27633 (.Y(n24874),
	.A(n24873),
	.B(n24872),
	.C(n24871));
   NOR2xp33_ASAP7_75t_SRAM U27635 (.Y(n24880),
	.A(FE_OCPN27690_n16757),
	.B(n24881));
   NAND2xp33_ASAP7_75t_SRAM U27636 (.Y(n24886),
	.A(n24880),
	.B(n24883));
   NOR2xp33_ASAP7_75t_SRAM U27637 (.Y(n24884),
	.A(FE_OFN28836_FE_OCPN27631_n16774),
	.B(n24881));
   NAND2xp33_ASAP7_75t_SRAM U27638 (.Y(n24885),
	.A(n24884),
	.B(n24883));
   NAND2xp33_ASAP7_75t_SRAM U27639 (.Y(n24889),
	.A(n24886),
	.B(n24885));
   NAND3xp33_ASAP7_75t_SRAM U27640 (.Y(n24890),
	.A(n24889),
	.B(n24888),
	.C(n24887));
   NOR3xp33_ASAP7_75t_SRAM U27641 (.Y(n24897),
	.A(n24895),
	.B(n24894),
	.C(n24893));
   A2O1A1Ixp33_ASAP7_75t_SL U27642 (.Y(n24905),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(n25462),
	.C(n24904));
   A2O1A1Ixp33_ASAP7_75t_SL U27644 (.Y(n24916),
	.A1(n26824),
	.A2(n24911),
	.B(n24910),
	.C(n24909));
   OAI22xp33_ASAP7_75t_SRAM U27645 (.Y(n24912),
	.A1(text_in_r_6_),
	.A2(FE_OFN28490_ld_r),
	.B1(n24913),
	.B2(FE_OFN28490_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27646 (.Y(n505),
	.A1(FE_OCPN7641_n25778),
	.A2(n24916),
	.B(n24915),
	.C(n24914));
   NAND3xp33_ASAP7_75t_R U27647 (.Y(n24923),
	.A(n24919),
	.B(n24918),
	.C(n24917));
   O2A1O1Ixp33_ASAP7_75t_SL U27648 (.Y(n24926),
	.A1(n24923),
	.A2(n24922),
	.B(n26829),
	.C(n25956));
   A2O1A1Ixp33_ASAP7_75t_SL U27649 (.Y(n24928),
	.A1(n22405),
	.A2(n24930),
	.B(FE_OCPN29538_n24927),
	.C(n24926));
   A2O1A1Ixp33_ASAP7_75t_L U27650 (.Y(n24937),
	.A1(n24974),
	.A2(n24939),
	.B(n24936),
	.C(FE_OFN27130_w3_28));
   NOR2xp33_ASAP7_75t_SRAM U27651 (.Y(n24942),
	.A(FE_OCPN28157_n16534),
	.B(n24943));
   NAND3xp33_ASAP7_75t_L U27652 (.Y(n24954),
	.A(n24951),
	.B(n24950),
	.C(n24949));
   NOR2xp33_ASAP7_75t_SRAM U27653 (.Y(n24957),
	.A(n24955),
	.B(n24958));
   NAND2xp33_ASAP7_75t_R U27654 (.Y(n24963),
	.A(n24957),
	.B(n24960));
   NOR2xp33_ASAP7_75t_SRAM U27655 (.Y(n24961),
	.A(n24959),
	.B(n24958));
   NAND3xp33_ASAP7_75t_L U27656 (.Y(n24975),
	.A(n24966),
	.B(n24965),
	.C(n24964));
   OAI21x1_ASAP7_75t_SL U27657 (.Y(n25132),
	.A1(n24979),
	.A2(n24978),
	.B(n24977));
   O2A1O1Ixp33_ASAP7_75t_R U27658 (.Y(n24980),
	.A1(n25139),
	.A2(FE_OCPN29562_n25138),
	.B(FE_OCPN5112_n25135),
	.C(n25657));
   A2O1A1Ixp33_ASAP7_75t_SL U27659 (.Y(n429),
	.A1(FE_OCPN27787_n26728),
	.A2(n24987),
	.B(n24986),
	.C(n24985));
   OAI21xp33_ASAP7_75t_SRAM U27660 (.Y(n24989),
	.A1(FE_OFN28686_FE_OCPN27812),
	.A2(FE_OFN26035_n),
	.B(FE_OCPN28434_n17546));
   OAI21xp33_ASAP7_75t_SRAM U27661 (.Y(n24993),
	.A1(FE_OFN28893_n),
	.A2(n24989),
	.B(n24988));
   O2A1O1Ixp5_ASAP7_75t_SL U27662 (.Y(n25001),
	.A1(n24998),
	.A2(n24997),
	.B(n22405),
	.C(n24996));
   A2O1A1Ixp33_ASAP7_75t_L U27663 (.Y(n25389),
	.A1(n26829),
	.A2(n25005),
	.B(n25004),
	.C(n25003));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27664 (.Y(n25012),
	.A1(n19640),
	.A2(n26857),
	.B(FE_OCPN27478_n25011),
	.C(FE_OCPN27659_w3_25));
   FAx1_ASAP7_75t_SL U27665 (.SN(n25019),
	.A(FE_OFN28565_n26845),
	.B(FE_OFN154_n26788),
	.CI(n25014));
   OAI21xp5_ASAP7_75t_L U27666 (.Y(n25018),
	.A1(n25019),
	.A2(FE_PSN8279_FE_OCPN27292_n25389),
	.B(FE_OFN28490_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27667 (.Y(n337),
	.A1(FE_PSN8279_FE_OCPN27292_n25389),
	.A2(n25019),
	.B(n25018),
	.C(n25017));
   NAND3xp33_ASAP7_75t_SRAM U27669 (.Y(n25032),
	.A(n25026),
	.B(n25025),
	.C(n25024));
   OAI21xp33_ASAP7_75t_SRAM U27670 (.Y(n25030),
	.A1(n19920),
	.A2(FE_OCPN29298_n25028),
	.B(n25027));
   NOR3xp33_ASAP7_75t_SRAM U27671 (.Y(n25033),
	.A(n25032),
	.B(FE_OFN28557_n25031),
	.C(n25030));
   NOR2xp33_ASAP7_75t_R U27672 (.Y(n25035),
	.A(n25033),
	.B(n17732));
   NOR3xp33_ASAP7_75t_L U27673 (.Y(n25045),
	.A(n25047),
	.B(n25679),
	.C(n25046));
   O2A1O1Ixp5_ASAP7_75t_SL U27674 (.Y(n25049),
	.A1(n25047),
	.A2(n25046),
	.B(FE_OCPN27362_n25679),
	.C(n25045));
   NOR2xp33_ASAP7_75t_SRAM U27675 (.Y(n25056),
	.A(n27007),
	.B(n25055));
   A2O1A1Ixp33_ASAP7_75t_L U27676 (.Y(n25070),
	.A1(n26457),
	.A2(n25069),
	.B(n27004),
	.C(n26463));
   A2O1A1Ixp33_ASAP7_75t_L U27677 (.Y(n25074),
	.A1(n26139),
	.A2(n26138),
	.B(n26135),
	.C(n25073));
   NAND3xp33_ASAP7_75t_SRAM U27678 (.Y(n25089),
	.A(n25086),
	.B(n25085),
	.C(n25084));
   OAI21xp5_ASAP7_75t_L U27679 (.Y(n25094),
	.A1(FE_OCPN28071_n25092),
	.A2(FE_OCPN27288_n25091),
	.B(n25090));
   NOR3xp33_ASAP7_75t_L U27680 (.Y(n26555),
	.A(n25094),
	.B(FE_OFN26542_n26155),
	.C(n25093));
   NOR3xp33_ASAP7_75t_SRAM U27681 (.Y(n25098),
	.A(n25096),
	.B(n25095),
	.C(n26559));
   NAND3xp33_ASAP7_75t_SRAM U27682 (.Y(n25101),
	.A(n26555),
	.B(n25098),
	.C(n25097));
   O2A1O1Ixp5_ASAP7_75t_SL U27683 (.Y(n25122),
	.A1(n25101),
	.A2(n25100),
	.B(n26249),
	.C(n25099));
   AND3x1_ASAP7_75t_SRAM U27684 (.Y(n25109),
	.A(n25105),
	.B(n25104),
	.C(n25103));
   O2A1O1Ixp33_ASAP7_75t_SL U27685 (.Y(n25119),
	.A1(FE_PSN8281_n25118),
	.A2(n25117),
	.B(n26584),
	.C(n25116));
   A2O1A1Ixp33_ASAP7_75t_SL U27686 (.Y(n26252),
	.A1(FE_OCPN28169_n25121),
	.A2(n25120),
	.B(n26926),
	.C(n25119));
   NOR2xp33_ASAP7_75t_SL U27687 (.Y(n25125),
	.A(FE_OFN25955_n25122),
	.B(FE_OFN16311_n26252));
   FAx1_ASAP7_75t_SL U27688 (.SN(n25131),
	.A(FE_OCPN29531_FE_OFN25926_n26922),
	.B(n25126),
	.CI(FE_OCPN27322_n25755));
   OAI22xp33_ASAP7_75t_SRAM U27689 (.Y(n25156),
	.A1(FE_OCPN8254_w3_3),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_3_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL U27690 (.Y(n25137),
	.A(n25133),
	.B(n25132));
   NAND3xp33_ASAP7_75t_SL U27692 (.Y(n25159),
	.A(FE_OFN16375_n25750),
	.B(n25397),
	.C(n25395));
   O2A1O1Ixp5_ASAP7_75t_SL U27693 (.Y(n25161),
	.A1(n25160),
	.A2(n25159),
	.B(n26139),
	.C(n25158));
   A2O1A1Ixp33_ASAP7_75t_SL U27694 (.Y(n25170),
	.A1(n26679),
	.A2(n25172),
	.B(FE_OCPN27825_n25169),
	.C(n25168));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27695 (.Y(n25180),
	.A1(n25682),
	.A2(n25680),
	.B(n25681),
	.C(w1_27_));
   A2O1A1Ixp33_ASAP7_75t_L U27696 (.Y(n25182),
	.A1(n25682),
	.A2(n25680),
	.B(n25181),
	.C(n25180));
   FAx1_ASAP7_75t_SL U27697 (.SN(n25187),
	.A(FE_OCPN29383_n26674),
	.B(n26171),
	.CI(n25182));
   OAI22xp33_ASAP7_75t_SRAM U27698 (.Y(n25183),
	.A1(text_in_r_91_),
	.A2(FE_OFN28487_ld_r),
	.B1(n25184),
	.B2(FE_OFN28487_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27699 (.Y(n399),
	.A1(n25187),
	.A2(FE_OCPN27560_n25755),
	.B(n25186),
	.C(n25185));
   NOR3xp33_ASAP7_75t_L U27700 (.Y(n25205),
	.A(n25203),
	.B(n25202),
	.C(n25201));
   OAI222xp33_ASAP7_75t_L U27701 (.Y(n25207),
	.A1(n25206),
	.A2(n26976),
	.B1(n25205),
	.B2(n26976),
	.C1(n25204),
	.C2(n26976));
   O2A1O1Ixp33_ASAP7_75t_SL U27702 (.Y(n26620),
	.A1(FE_OCPN29387_n25273),
	.A2(n25208),
	.B(n27183),
	.C(n25207));
   NOR3xp33_ASAP7_75t_SL U27703 (.Y(n25214),
	.A(n25212),
	.B(n25211),
	.C(n25210));
   O2A1O1Ixp5_ASAP7_75t_SL U27704 (.Y(n26621),
	.A1(n25217),
	.A2(n25216),
	.B(n27216),
	.C(n25215));
   NOR2xp33_ASAP7_75t_SL U27706 (.Y(n25239),
	.A(n25235),
	.B(n25237));
   OAI22xp33_ASAP7_75t_SRAM U27707 (.Y(n25272),
	.A1(w0_1_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_97_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27708 (.Y(n25253),
	.A1(n27127),
	.A2(n25255),
	.B(FE_OCPN28442_n27056),
	.C(n25252));
   A2O1A1Ixp33_ASAP7_75t_SL U27709 (.Y(n26115),
	.A1(n27127),
	.A2(n25255),
	.B(n25254),
	.C(n25253));
   NOR3xp33_ASAP7_75t_SRAM U27711 (.Y(n25259),
	.A(n25257),
	.B(n26100),
	.C(FE_OFN28783_n26099));
   O2A1O1Ixp5_ASAP7_75t_SL U27712 (.Y(n25261),
	.A1(n26106),
	.A2(n25260),
	.B(n27127),
	.C(n26113));
   NOR2xp33_ASAP7_75t_SL U27713 (.Y(n25264),
	.A(n25261),
	.B(n26427));
   NOR2x1p5_ASAP7_75t_SL U27715 (.Y(n26781),
	.A(FE_OFN2_ld_r),
	.B(n26784));
   NAND3xp33_ASAP7_75t_SRAM U27716 (.Y(n25288),
	.A(n25286),
	.B(n25285),
	.C(FE_OFN27147_n25284));
   NOR3xp33_ASAP7_75t_R U27717 (.Y(n25300),
	.A(n25298),
	.B(n25297),
	.C(n25296));
   NAND3xp33_ASAP7_75t_SL U27718 (.Y(n25304),
	.A(n25301),
	.B(n25300),
	.C(n25299));
   NAND3xp33_ASAP7_75t_SL U27719 (.Y(n25303),
	.A(n17775),
	.B(n25302),
	.C(n25504));
   A2O1A1Ixp33_ASAP7_75t_L U27720 (.Y(n25308),
	.A1(n25307),
	.A2(n25306),
	.B(n26976),
	.C(n25305));
   O2A1O1Ixp5_ASAP7_75t_SL U27721 (.Y(n26910),
	.A1(n27140),
	.A2(n27139),
	.B(n25313),
	.C(n25312));
   NAND3xp33_ASAP7_75t_R U27723 (.Y(n25324),
	.A(n25323),
	.B(FE_OFN28618_n25322),
	.C(n25321));
   NAND3xp33_ASAP7_75t_SRAM U27724 (.Y(n25331),
	.A(n25901),
	.B(n25328),
	.C(n25327));
   O2A1O1Ixp5_ASAP7_75t_SL U27725 (.Y(n26982),
	.A1(n27168),
	.A2(n27167),
	.B(n25333),
	.C(n25332));
   A2O1A1Ixp33_ASAP7_75t_L U27726 (.Y(n25334),
	.A1(n26941),
	.A2(n26942),
	.B(FE_OCPN27809_n26938),
	.C(n25346));
   A2O1A1Ixp33_ASAP7_75t_SL U27727 (.Y(n25336),
	.A1(n26942),
	.A2(n26941),
	.B(n25335),
	.C(n25334));
   FAx1_ASAP7_75t_SL U27728 (.SN(n25349),
	.A(FE_OCPN27741_n),
	.B(FE_OCPN27354_n26982),
	.CI(n25336));
   OAI22xp33_ASAP7_75t_SRAM U27729 (.Y(n25345),
	.A1(text_in_r_41_),
	.A2(FE_OFN16215_ld_r),
	.B1(n25346),
	.B2(FE_OFN16215_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27730 (.Y(n370),
	.A1(n25349),
	.A2(FE_OCPN7629_FE_OFN105_n27178),
	.B(n25348),
	.C(n25347));
   NOR2xp33_ASAP7_75t_SRAM U27731 (.Y(n25356),
	.A(n25353),
	.B(n25352));
   NAND3xp33_ASAP7_75t_L U27732 (.Y(n25358),
	.A(n25356),
	.B(n25355),
	.C(n25354));
   A2O1A1Ixp33_ASAP7_75t_SL U27734 (.Y(n25364),
	.A1(n25367),
	.A2(n25366),
	.B(n25363),
	.C(n25362));
   NOR3xp33_ASAP7_75t_SL U27735 (.Y(n25370),
	.A(FE_OCPN28100_n25470),
	.B(n26349),
	.C(n25469));
   OAI21xp5_ASAP7_75t_L U27736 (.Y(n25371),
	.A1(FE_OFN16214_ld_r),
	.A2(FE_OCPN27534_n),
	.B(n25372));
   A2O1A1Ixp33_ASAP7_75t_SL U27737 (.Y(n25376),
	.A1(FE_OCPN27534_n),
	.A2(FE_OFN28489_ld_r),
	.B(n25372),
	.C(n25371));
   A2O1A1Ixp33_ASAP7_75t_L U27738 (.Y(n499),
	.A1(n25376),
	.A2(n25375),
	.B(FE_OFN26640_w3_14),
	.C(n25373));
   OAI22xp33_ASAP7_75t_SRAM U27739 (.Y(n25394),
	.A1(n25377),
	.A2(FE_OFN28489_ld_r),
	.B1(text_in_r_17_),
	.B2(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_R U27740 (.Y(n25380),
	.A1(n25575),
	.A2(n25382),
	.B(FE_OFN28960_n25379),
	.C(n25377));
   A2O1A1Ixp33_ASAP7_75t_L U27741 (.Y(n25385),
	.A1(n26793),
	.A2(n26857),
	.B(n26787),
	.C(n25384));
   O2A1O1Ixp5_ASAP7_75t_SL U27743 (.Y(n410),
	.A1(n25377),
	.A2(text_in_r_17_),
	.B(n25394),
	.C(n25393));
   NAND3xp33_ASAP7_75t_SRAM U27744 (.Y(n25400),
	.A(n25399),
	.B(n25398),
	.C(n25397));
   NOR2xp33_ASAP7_75t_SRAM U27745 (.Y(n25401),
	.A(FE_OCPN8229_n25750),
	.B(n25400));
   NOR2xp33_ASAP7_75t_R U27746 (.Y(n25402),
	.A(n25401),
	.B(FE_OFN165_sa12_7));
   O2A1O1Ixp33_ASAP7_75t_SL U27747 (.Y(n25417),
	.A1(n25420),
	.A2(FE_OFN28561_n25419),
	.B(FE_OCPN27682_n25414),
	.C(FE_OFN29087_n));
   NOR2x1_ASAP7_75t_SL U27749 (.Y(n25424),
	.A(n26729),
	.B(n25425));
   O2A1O1Ixp5_ASAP7_75t_SL U27750 (.Y(n418),
	.A1(FE_OFN16179_w3_19),
	.A2(text_in_r_19_),
	.B(n25427),
	.C(n25426));
   O2A1O1Ixp33_ASAP7_75t_SRAM U27752 (.Y(n25428),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25669),
	.C(FE_OFN28853_FE_OCPN28408));
   OAI22xp33_ASAP7_75t_SRAM U27753 (.Y(n25432),
	.A1(text_in_r_11_),
	.A2(FE_OFN28489_ld_r),
	.B1(FE_OFN28853_FE_OCPN28408),
	.B2(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27754 (.Y(n442),
	.A1(FE_OCPN27282_n25437),
	.A2(n25436),
	.B(n25435),
	.C(n25434));
   NOR3xp33_ASAP7_75t_SRAM U27755 (.Y(n25441),
	.A(n25440),
	.B(n25439),
	.C(n25438));
   O2A1O1Ixp5_ASAP7_75t_SL U27756 (.Y(n25696),
	.A1(n26599),
	.A2(n26598),
	.B(n26139),
	.C(n25443));
   A2O1A1Ixp33_ASAP7_75t_L U27757 (.Y(n25445),
	.A1(n26679),
	.A2(n25694),
	.B(n25444),
	.C(FE_OCPN29361_n25696));
   A2O1A1Ixp33_ASAP7_75t_L U27758 (.Y(n26930),
	.A1(n26679),
	.A2(n25694),
	.B(n25446),
	.C(n25445));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27759 (.Y(n25453),
	.A1(n25455),
	.A2(n26139),
	.B(n25452),
	.C(FE_OFN66_w1_25));
   FAx1_ASAP7_75t_SL U27760 (.SN(n25461),
	.A(FE_OCPN29576_n26930),
	.B(FE_OCPN27462_n26215),
	.CI(n25456));
   A2O1A1Ixp33_ASAP7_75t_SL U27761 (.Y(n405),
	.A1(FE_OCPN29382_n26674),
	.A2(n25461),
	.B(n25460),
	.C(n25459));
   OR2x2_ASAP7_75t_SL U27762 (.Y(n25464),
	.A(FE_OCPN28106_FE_OFN25876_n25462),
	.B(FE_OFN16283_n26788));
   A2O1A1Ixp33_ASAP7_75t_L U27763 (.Y(n25463),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(FE_OCPN28106_FE_OFN25876_n25462),
	.C(FE_OFN16283_n26788));
   A2O1A1Ixp33_ASAP7_75t_SL U27764 (.Y(n25468),
	.A1(FE_OFN16148_n25466),
	.A2(FE_OFN29051_n25465),
	.B(n25464),
	.C(n25463));
   NOR3xp33_ASAP7_75t_SL U27765 (.Y(n25467),
	.A(FE_OCPN28100_n25470),
	.B(n25468),
	.C(n25469));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27766 (.Y(n25473),
	.A1(n25475),
	.A2(n25575),
	.B(n25472),
	.C(FE_OCPN29501_FE_OFN28662_w3_7));
   OAI21xp5_ASAP7_75t_SL U27767 (.Y(n25479),
	.A1(n25480),
	.A2(n25481),
	.B(FE_OFN28489_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U27768 (.Y(n25476),
	.A1(text_in_r_7_),
	.A2(FE_OFN28489_ld_r),
	.B1(FE_OCPN29501_FE_OFN28662_w3_7),
	.B2(FE_OFN28489_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U27769 (.Y(n25487),
	.A1(FE_OCPN27723_n),
	.A2(n25484),
	.B(FE_OCPN27467_n25483),
	.C(n25482));
   A2O1A1Ixp33_ASAP7_75t_SL U27770 (.Y(n25492),
	.A1(FE_OCPN28077_n),
	.A2(FE_OFN28487_ld_r),
	.B(n25487),
	.C(n25486));
   NOR3xp33_ASAP7_75t_SL U27771 (.Y(n25493),
	.A(FE_OCPN27753_n26685),
	.B(FE_OFN160_n26440),
	.C(n25494));
   A2O1A1Ixp33_ASAP7_75t_SL U27772 (.Y(n25501),
	.A1(FE_OCPN4698_n25497),
	.A2(FE_OFN28487_ld_r),
	.B(n25496),
	.C(n25495));
   NAND3xp33_ASAP7_75t_SL U27773 (.Y(n25498),
	.A(n25499),
	.B(n25501),
	.C(n25500));
   A2O1A1Ixp33_ASAP7_75t_SL U27774 (.Y(n496),
	.A1(n25501),
	.A2(n25500),
	.B(n25499),
	.C(n25498));
   NAND3xp33_ASAP7_75t_SRAM U27775 (.Y(n25505),
	.A(n25504),
	.B(n25503),
	.C(n25502));
   A2O1A1Ixp33_ASAP7_75t_SL U27776 (.Y(n25512),
	.A1(n26407),
	.A2(n25510),
	.B(n25509),
	.C(n25508));
   A2O1A1Ixp33_ASAP7_75t_SL U27778 (.Y(n25520),
	.A1(n26651),
	.A2(FE_OCPN29471_n24175),
	.B(n25512),
	.C(n25511));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27779 (.Y(n25513),
	.A1(n27192),
	.A2(FE_OFN16176_n27207),
	.B(n27188),
	.C(n25516));
   OAI22xp33_ASAP7_75t_SRAM U27780 (.Y(n25515),
	.A1(text_in_r_38_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(n25516),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27781 (.Y(n503),
	.A1(n25520),
	.A2(n25519),
	.B(n25518),
	.C(n25517));
   A2O1A1Ixp33_ASAP7_75t_SL U27782 (.Y(n25521),
	.A1(n26942),
	.A2(n26201),
	.B(n26198),
	.C(n26495));
   NOR3xp33_ASAP7_75t_SRAM U27783 (.Y(n25534),
	.A(n25525),
	.B(FE_OCPN29318_n25524),
	.C(n25523));
   NOR3xp33_ASAP7_75t_L U27784 (.Y(n25533),
	.A(n25529),
	.B(n25528),
	.C(n25527));
   NOR3xp33_ASAP7_75t_SRAM U27785 (.Y(n25532),
	.A(n26967),
	.B(n25531),
	.C(n25530));
   NAND3xp33_ASAP7_75t_SL U27786 (.Y(n25535),
	.A(n25534),
	.B(n25533),
	.C(n25532));
   A2O1A1Ixp33_ASAP7_75t_SL U27787 (.Y(n25537),
	.A1(n26915),
	.A2(n26914),
	.B(FE_OFN28473_n26911),
	.C(n26317));
   NAND3xp33_ASAP7_75t_R U27789 (.Y(n25542),
	.A(n25541),
	.B(n25540),
	.C(n25562));
   NOR2xp33_ASAP7_75t_L U27790 (.Y(n25546),
	.A(n25545),
	.B(n25544));
   NOR2x1_ASAP7_75t_SL U27791 (.Y(n26955),
	.A(n25557),
	.B(n25556));
   FAx1_ASAP7_75t_SL U27792 (.SN(n25573),
	.A(n26520),
	.B(n25621),
	.CI(n25560));
   NAND2xp5_ASAP7_75t_L U27793 (.Y(n25568),
	.A(FE_OFN104_n27179),
	.B(n26051));
   OAI22xp33_ASAP7_75t_SRAM U27794 (.Y(n25569),
	.A1(text_in_r_59_),
	.A2(FE_OFN16215_ld_r),
	.B1(n25570),
	.B2(FE_OFN16215_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27795 (.Y(n417),
	.A1(n25573),
	.A2(FE_OCPN29356_n27110),
	.B(n25572),
	.C(n25571));
   NOR3xp33_ASAP7_75t_SRAM U27796 (.Y(n25584),
	.A(n25581),
	.B(n25580),
	.C(n25579));
   O2A1O1Ixp5_ASAP7_75t_SRAM U27797 (.Y(n25591),
	.A1(FE_OCPN27629_n25589),
	.A2(n25588),
	.B(n26829),
	.C(n25587));
   A2O1A1Ixp33_ASAP7_75t_SL U27798 (.Y(n25594),
	.A1(n25592),
	.A2(n25591),
	.B(n26852),
	.C(n25590));
   A2O1A1Ixp33_ASAP7_75t_SL U27799 (.Y(n25598),
	.A1(FE_OFN28565_n26845),
	.A2(FE_OFN28489_ld_r),
	.B(n25594),
	.C(n25593));
   NAND2xp33_ASAP7_75t_R U27800 (.Y(n25597),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_0_));
   NAND3xp33_ASAP7_75t_SL U27801 (.Y(n25595),
	.A(n25596),
	.B(n25598),
	.C(n25597));
   A2O1A1Ixp33_ASAP7_75t_SL U27802 (.Y(n383),
	.A1(n25598),
	.A2(n25597),
	.B(n25596),
	.C(n25595));
   NOR2xp33_ASAP7_75t_SRAM U27803 (.Y(n25600),
	.A(FE_OFN27069_n24478),
	.B(sa00_7_));
   NOR2xp33_ASAP7_75t_SRAM U27804 (.Y(n25602),
	.A(n25601),
	.B(sa00_7_));
   A2O1A1Ixp33_ASAP7_75t_R U27805 (.Y(n25607),
	.A1(n27117),
	.A2(n27116),
	.B(FE_OFN29010_n27113),
	.C(FE_OCPN8268_n26632));
   A2O1A1Ixp33_ASAP7_75t_SL U27806 (.Y(n25613),
	.A1(n27117),
	.A2(n27052),
	.B(FE_OFN29142_n27049),
	.C(n25612));
   A2O1A1Ixp33_ASAP7_75t_SL U27808 (.Y(n446),
	.A1(n25620),
	.A2(n25619),
	.B(n25618),
	.C(n25617));
   A2O1A1Ixp33_ASAP7_75t_L U27809 (.Y(n25622),
	.A1(n26942),
	.A2(n26941),
	.B(FE_OCPN27809_n26938),
	.C(n26944));
   A2O1A1Ixp33_ASAP7_75t_SL U27810 (.Y(n25625),
	.A1(n26942),
	.A2(n26941),
	.B(n25623),
	.C(n25622));
   NOR3xp33_ASAP7_75t_SL U27811 (.Y(n25624),
	.A(FE_OCPN29515_n27136),
	.B(n25625),
	.C(n25626));
   NAND3xp33_ASAP7_75t_SRAM U27812 (.Y(n25633),
	.A(n25630),
	.B(n25629),
	.C(n25628));
   OAI21xp5_ASAP7_75t_SL U27813 (.Y(n25640),
	.A1(n25639),
	.A2(n25638),
	.B(n26323));
   O2A1O1Ixp5_ASAP7_75t_SL U27814 (.Y(n26513),
	.A1(n26900),
	.A2(n26899),
	.B(n27207),
	.C(n25644));
   OAI22xp33_ASAP7_75t_SRAM U27815 (.Y(n25647),
	.A1(text_in_r_34_),
	.A2(FE_OFN16215_ld_r),
	.B1(n25648),
	.B2(FE_OFN16215_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U27816 (.Y(n25666),
	.A1(FE_OFN25897_w3_4),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_4_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SRAM U27818 (.Y(n25670),
	.A1(n17584),
	.A2(FE_OFN16353_n25672),
	.B(n25669),
	.C(FE_OFN26120_n));
   FAx1_ASAP7_75t_SL U27819 (.SN(n25678),
	.A(FE_OFN155_n26788),
	.B(FE_OCPN27359_n26726),
	.CI(n25673));
   OAI22xp33_ASAP7_75t_SRAM U27820 (.Y(n25674),
	.A1(text_in_r_27_),
	.A2(FE_OFN28490_ld_r),
	.B1(FE_OFN26120_n),
	.B2(FE_OFN28490_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27821 (.Y(n25683),
	.A1(n26282),
	.A2(n26250),
	.B(n26251),
	.C(n26704));
   O2A1O1Ixp33_ASAP7_75t_R U27822 (.Y(n25685),
	.A1(FE_OFN16413_n26687),
	.A2(n26258),
	.B(n26255),
	.C(n25690));
   FAx1_ASAP7_75t_SL U27823 (.SN(n25693),
	.A(FE_OCPN29353_n26586),
	.B(FE_OCPN27441_n25688),
	.CI(n25687));
   OAI22xp33_ASAP7_75t_SRAM U27825 (.Y(n25689),
	.A1(text_in_r_75_),
	.A2(FE_OFN28486_ld_r),
	.B1(n25690),
	.B2(FE_OFN28486_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27826 (.Y(n463),
	.A1(n25693),
	.A2(FE_OCPN7585_FE_OFN25926_n26922),
	.B(n25692),
	.C(n25691));
   NAND3xp33_ASAP7_75t_SL U27827 (.Y(n25702),
	.A(n26213),
	.B(n25710),
	.C(n25709));
   A2O1A1Ixp33_ASAP7_75t_SL U27828 (.Y(n25704),
	.A1(n25710),
	.A2(n25709),
	.B(n26213),
	.C(n25702));
   O2A1O1Ixp33_ASAP7_75t_SL U27829 (.Y(n448),
	.A1(n25707),
	.A2(n25706),
	.B(w1_0_),
	.C(n25705));
   A2O1A1Ixp33_ASAP7_75t_SL U27830 (.Y(n25727),
	.A1(n25710),
	.A2(n25709),
	.B(FE_OCPN29335_n),
	.C(n25708));
   A2O1A1Ixp33_ASAP7_75t_SL U27831 (.Y(n25723),
	.A1(n26139),
	.A2(n25725),
	.B(n25722),
	.C(n25721));
   A2O1A1Ixp33_ASAP7_75t_SL U27832 (.Y(n26717),
	.A1(n26139),
	.A2(n25725),
	.B(n25724),
	.C(n25723));
   NOR3xp33_ASAP7_75t_SL U27833 (.Y(n25726),
	.A(n25727),
	.B(FE_OFN16214_ld_r),
	.C(FE_OCPN27884_n26717));
   A2O1A1Ixp33_ASAP7_75t_L U27835 (.Y(n25734),
	.A1(n26249),
	.A2(n25736),
	.B(n26178),
	.C(w1_19_));
   NOR2xp33_ASAP7_75t_SRAM U27836 (.Y(n25739),
	.A(FE_OFN28739_n17898),
	.B(n25740));
   O2A1O1Ixp33_ASAP7_75t_SL U27837 (.Y(n26276),
	.A1(FE_OCPN8229_n25750),
	.A2(n25749),
	.B(n26139),
	.C(n25748));
   NAND2x1p5_ASAP7_75t_L U27838 (.Y(n26443),
	.A(FE_OCPN27884_n26717),
	.B(FE_OFN28486_ld_r));
   NOR2xp33_ASAP7_75t_SRAM U27839 (.Y(n25785),
	.A(FE_OCPN29513_n17447),
	.B(n25786));
   NOR2xp33_ASAP7_75t_SRAM U27840 (.Y(n25788),
	.A(FE_OCPN29435_n17445),
	.B(n25786));
   NAND3xp33_ASAP7_75t_R U27841 (.Y(n25797),
	.A(n25792),
	.B(n25791),
	.C(n26073));
   O2A1O1Ixp5_ASAP7_75t_SL U27842 (.Y(n25799),
	.A1(n25797),
	.A2(n25796),
	.B(n27062),
	.C(n26369));
   A2O1A1Ixp33_ASAP7_75t_SL U27843 (.Y(n25800),
	.A1(n27127),
	.A2(n27126),
	.B(n27122),
	.C(n25799));
   A2O1A1Ixp33_ASAP7_75t_SL U27844 (.Y(n26380),
	.A1(n27127),
	.A2(n27126),
	.B(n25801),
	.C(n25800));
   A2O1A1Ixp33_ASAP7_75t_SL U27845 (.Y(n25810),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(n25804),
	.C(n25803));
   O2A1O1Ixp5_ASAP7_75t_SL U27847 (.Y(n25822),
	.A1(n25821),
	.A2(n25820),
	.B(n26942),
	.C(n25819));
   NAND2xp5_ASAP7_75t_SL U27848 (.Y(n25829),
	.A(FE_OCPN27456_n27189),
	.B(n25826));
   A2O1A1Ixp33_ASAP7_75t_SL U27849 (.Y(n25828),
	.A1(FE_OFN16176_n27207),
	.A2(n27192),
	.B(FE_OCPN29447_n27189),
	.C(n25827));
   O2A1O1Ixp33_ASAP7_75t_L U27850 (.Y(n25845),
	.A1(FE_OCPN5053_n25832),
	.A2(n25831),
	.B(FE_OCPN5020_n27079),
	.C(n25830));
   O2A1O1Ixp33_ASAP7_75t_SL U27851 (.Y(n25844),
	.A1(FE_OCPN27451_n26236),
	.A2(n26235),
	.B(n25839),
	.C(n25838));
   OAI22xp33_ASAP7_75t_SRAM U27852 (.Y(n25840),
	.A1(text_in_r_54_),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B1(n25841),
	.B2(FE_OFN16_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27853 (.Y(n510),
	.A1(n25845),
	.A2(n25844),
	.B(n25843),
	.C(n25842));
   A2O1A1Ixp33_ASAP7_75t_SL U27854 (.Y(n25854),
	.A1(FE_OFN28521_n26007),
	.A2(n25853),
	.B(n26315),
	.C(n26012));
   A2O1A1Ixp33_ASAP7_75t_SL U27855 (.Y(n26501),
	.A1(FE_OFN16176_n27207),
	.A2(n26196),
	.B(n25859),
	.C(n25858));
   O2A1O1Ixp33_ASAP7_75t_L U27856 (.Y(n25862),
	.A1(FE_OFN16158_n26959),
	.A2(n26958),
	.B(FE_OCPN28119_n26955),
	.C(n26507));
   NAND3xp33_ASAP7_75t_SRAM U27857 (.Y(n25867),
	.A(n26001),
	.B(FE_OFN28502_n25865),
	.C(n25997));
   NOR3xp33_ASAP7_75t_SRAM U27858 (.Y(n25892),
	.A(n25867),
	.B(FE_OCPN29525_n18947),
	.C(n25866));
   NOR2xp33_ASAP7_75t_SRAM U27859 (.Y(n25874),
	.A(FE_OCPN27859_n25868),
	.B(n25875));
   OAI21xp33_ASAP7_75t_SRAM U27860 (.Y(n25873),
	.A1(FE_OFN16396_n25869),
	.A2(FE_OCPN27761_n16977),
	.B(FE_OCPN8213_FE_OFN29234_n16996));
   AND3x1_ASAP7_75t_SRAM U27862 (.Y(n25876),
	.A(n25873),
	.B(n25872),
	.C(FE_OFN28994_FE_OCPN5176_n25870));
   NAND2xp33_ASAP7_75t_R U27863 (.Y(n25879),
	.A(n25874),
	.B(n25876));
   NOR2xp33_ASAP7_75t_SRAM U27864 (.Y(n25877),
	.A(FE_OFN28584_n17001),
	.B(n25875));
   NAND2xp33_ASAP7_75t_R U27865 (.Y(n25878),
	.A(n25877),
	.B(n25876));
   A2O1A1Ixp33_ASAP7_75t_L U27866 (.Y(n25888),
	.A1(n25887),
	.A2(n25886),
	.B(n27102),
	.C(FE_OCPN5106_n25999));
   A2O1A1Ixp33_ASAP7_75t_SL U27867 (.Y(n468),
	.A1(n25898),
	.A2(FE_OCPN29356_n27110),
	.B(n25897),
	.C(n25896));
   NOR2xp33_ASAP7_75t_SRAM U27868 (.Y(n25900),
	.A(n25899),
	.B(sa20_6_));
   NAND3xp33_ASAP7_75t_SRAM U27869 (.Y(n25904),
	.A(n25903),
	.B(n25902),
	.C(n25901));
   NOR2xp33_ASAP7_75t_R U27870 (.Y(n25906),
	.A(FE_OFN16301_n25905),
	.B(n25904));
   NOR2xp33_ASAP7_75t_SRAM U27871 (.Y(n25913),
	.A(FE_OFN28924_n25912),
	.B(n25911));
   O2A1O1Ixp5_ASAP7_75t_SL U27872 (.Y(n25934),
	.A1(FE_OCPN28316_n26980),
	.A2(n26979),
	.B(n27216),
	.C(n25916));
   O2A1O1Ixp5_ASAP7_75t_SL U27873 (.Y(n25927),
	.A1(FE_OCPN27522_n25921),
	.A2(n25920),
	.B(n27171),
	.C(n25919));
   A2O1A1Ixp33_ASAP7_75t_L U27874 (.Y(n25924),
	.A1(n27183),
	.A2(n27182),
	.B(n27177),
	.C(n25923));
   NAND3xp33_ASAP7_75t_SL U27875 (.Y(n25926),
	.A(FE_DBTN0_ld_r),
	.B(n25927),
	.C(FE_OCPN7636_n25940));
   O2A1O1Ixp33_ASAP7_75t_SL U27876 (.Y(n426),
	.A1(n25930),
	.A2(n25929),
	.B(w2_0_),
	.C(n25928));
   OAI22xp33_ASAP7_75t_SRAM U27877 (.Y(n25944),
	.A1(w2_1_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_33_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_SL U27878 (.Y(n25932),
	.A1(n27168),
	.A2(n27167),
	.B(n27163),
	.C(n25931));
   O2A1O1Ixp33_ASAP7_75t_SL U27879 (.Y(n25939),
	.A1(n27168),
	.A2(n27167),
	.B(n25933),
	.C(n25932));
   A2O1A1Ixp33_ASAP7_75t_SL U27880 (.Y(n25938),
	.A1(FE_OFN16177_n27207),
	.A2(n27206),
	.B(n25937),
	.C(n25936));
   NOR2x1_ASAP7_75t_L U27882 (.Y(n26327),
	.A(FE_OFN1_ld_r),
	.B(FE_OCPN7636_n25940));
   A2O1A1Ixp33_ASAP7_75t_SL U27884 (.Y(n25948),
	.A1(n26819),
	.A2(FE_OCPN8227_n25950),
	.B(n25947),
	.C(n26339));
   A2O1A1Ixp33_ASAP7_75t_SL U27886 (.Y(n25965),
	.A1(FE_OCPN28320_n25954),
	.A2(FE_OCPN28328_n25953),
	.B(n25952),
	.C(n25951));
   NAND2xp33_ASAP7_75t_SRAM U27887 (.Y(n25958),
	.A(FE_OFN16441_w3_21),
	.B(FE_OFN28504_n25956));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27888 (.Y(n25957),
	.A1(n25959),
	.A2(n26829),
	.B(FE_OFN16249_n25956),
	.C(n25961));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27889 (.Y(n25964),
	.A1(n26829),
	.A2(n25959),
	.B(n25958),
	.C(n25957));
   OAI21xp5_ASAP7_75t_SL U27890 (.Y(n25963),
	.A1(n25965),
	.A2(n25964),
	.B(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27891 (.Y(n25968),
	.A1(n27117),
	.A2(n26531),
	.B(FE_OCPN29389_n26528),
	.C(n25967));
   NAND2xp33_ASAP7_75t_SRAM U27893 (.Y(n25992),
	.A(n25989),
	.B(n25988));
   NOR3xp33_ASAP7_75t_SL U27894 (.Y(n25993),
	.A(n25992),
	.B(FE_OCPN29525_n18947),
	.C(n25990));
   NAND3xp33_ASAP7_75t_SRAM U27895 (.Y(n25998),
	.A(n25995),
	.B(n25994),
	.C(n25993));
   A2O1A1Ixp33_ASAP7_75t_L U27896 (.Y(n26004),
	.A1(n27216),
	.A2(n26494),
	.B(FE_OCPN28307_n26491),
	.C(n26192));
   A2O1A1Ixp33_ASAP7_75t_SL U27897 (.Y(n26234),
	.A1(n27216),
	.A2(n26494),
	.B(n26005),
	.C(n26004));
   NOR2xp33_ASAP7_75t_SRAM U27898 (.Y(n26014),
	.A(w2_12_),
	.B(FE_OFN16281_n26011));
   O2A1O1Ixp33_ASAP7_75t_SRAM U27899 (.Y(n26013),
	.A1(n26315),
	.A2(n26015),
	.B(n26012),
	.C(n26018));
   FAx1_ASAP7_75t_SL U27900 (.SN(n26021),
	.A(n27176),
	.B(FE_PSN8321_n26520),
	.CI(n26016));
   OAI22xp33_ASAP7_75t_SRAM U27901 (.Y(n26017),
	.A1(text_in_r_44_),
	.A2(FE_OFN16215_ld_r),
	.B1(n26018),
	.B2(FE_OFN16215_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27902 (.Y(n514),
	.A1(FE_OCPN7605_n26234),
	.A2(n26021),
	.B(n26020),
	.C(n26019));
   NOR3xp33_ASAP7_75t_SRAM U27903 (.Y(n26034),
	.A(n26024),
	.B(n26023),
	.C(n26022));
   OAI21xp33_ASAP7_75t_SRAM U27904 (.Y(n26030),
	.A1(FE_OCPN27428_n26027),
	.A2(FE_OFN29121_n26026),
	.B(n26025));
   NOR3xp33_ASAP7_75t_SRAM U27905 (.Y(n26033),
	.A(n26030),
	.B(n26029),
	.C(n26028));
   OAI22xp33_ASAP7_75t_L U27906 (.Y(n26032),
	.A1(FE_OFN16163_n26584),
	.A2(n26031),
	.B1(n26583),
	.B2(n26031));
   OAI22xp33_ASAP7_75t_L U27908 (.Y(n26047),
	.A1(n26045),
	.A2(n27168),
	.B1(n26044),
	.B2(n27168));
   A2O1A1Ixp33_ASAP7_75t_L U27909 (.Y(n26059),
	.A1(FE_OCPN5086_n26050),
	.A2(n27074),
	.B(n25506),
	.C(n26048));
   A2O1A1Ixp33_ASAP7_75t_L U27910 (.Y(n26502),
	.A1(FE_OFN16177_n27207),
	.A2(n26057),
	.B(n26056),
	.C(n26055));
   O2A1O1Ixp5_ASAP7_75t_SL U27911 (.Y(n26077),
	.A1(n26076),
	.A2(n26075),
	.B(n27062),
	.C(n26074));
   A2O1A1Ixp33_ASAP7_75t_SL U27912 (.Y(n26081),
	.A1(n26080),
	.A2(n26079),
	.B(n26078),
	.C(n26077));
   A2O1A1Ixp33_ASAP7_75t_L U27913 (.Y(n26085),
	.A1(FE_OFN16170_n26637),
	.A2(n26226),
	.B(n26222),
	.C(FE_OCPN27283_n26867));
   A2O1A1Ixp33_ASAP7_75t_SL U27914 (.Y(n450),
	.A1(FE_OCPN5045_n26098),
	.A2(FE_OCPN28140_FE_OFN133_n24306),
	.B(n26097),
	.C(n26096));
   NOR3xp33_ASAP7_75t_SRAM U27915 (.Y(n26102),
	.A(FE_OFN28625_n26101),
	.B(n26100),
	.C(FE_OFN28783_n26099));
   NAND3xp33_ASAP7_75t_SRAM U27916 (.Y(n26105),
	.A(n26104),
	.B(FE_OFN28767_n26103),
	.C(n26102));
   NOR2xp33_ASAP7_75t_SRAM U27917 (.Y(n26107),
	.A(n26106),
	.B(n26105));
   NOR2xp33_ASAP7_75t_SRAM U27918 (.Y(n26108),
	.A(n26107),
	.B(FE_OFN28499_sa00_6));
   NOR3xp33_ASAP7_75t_SL U27919 (.Y(n26111),
	.A(FE_OCPN27314_n26113),
	.B(FE_OCPN27525_n26434),
	.C(n26112));
   O2A1O1Ixp5_ASAP7_75t_SL U27920 (.Y(n26116),
	.A1(FE_OCPN27314_n26113),
	.A2(n26112),
	.B(FE_OCPN27525_n26434),
	.C(n26111));
   NAND3xp33_ASAP7_75t_SRAM U27921 (.Y(n26123),
	.A(n26120),
	.B(n26358),
	.C(n26360));
   NOR3xp33_ASAP7_75t_SRAM U27922 (.Y(n26127),
	.A(n26123),
	.B(n26122),
	.C(n26121));
   OAI22xp33_ASAP7_75t_SRAM U27924 (.Y(n26129),
	.A1(text_in_r_108_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(n26130),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27925 (.Y(n515),
	.A1(FE_OCPN27321_n26380),
	.A2(n26133),
	.B(n26132),
	.C(n26131));
   A2O1A1Ixp33_ASAP7_75t_L U27926 (.Y(n26136),
	.A1(n26138),
	.A2(n26139),
	.B(n26135),
	.C(n26142));
   FAx1_ASAP7_75t_SL U27927 (.SN(n26145),
	.A(FE_OCPN29277_n26713),
	.B(FE_OCPN29359_n26586),
	.CI(n26140));
   A2O1A1Ixp33_ASAP7_75t_SL U27928 (.Y(n441),
	.A1(FE_OCPN29382_n26674),
	.A2(FE_OCPN7609_n26145),
	.B(n26144),
	.C(n26143));
   NAND2xp33_ASAP7_75t_SRAM U27929 (.Y(n26150),
	.A(n26147),
	.B(n26146));
   NOR3xp33_ASAP7_75t_SRAM U27930 (.Y(n26153),
	.A(n26150),
	.B(n26149),
	.C(n26148));
   NAND3xp33_ASAP7_75t_SRAM U27931 (.Y(n26156),
	.A(n26153),
	.B(n26152),
	.C(n26151));
   NOR3xp33_ASAP7_75t_SRAM U27932 (.Y(n26157),
	.A(n26156),
	.B(FE_OFN26542_n26155),
	.C(n26154));
   NOR2xp33_ASAP7_75t_SRAM U27933 (.Y(n26158),
	.A(n26157),
	.B(sa23_7_));
   NAND3xp33_ASAP7_75t_SRAM U27934 (.Y(n26166),
	.A(n26161),
	.B(n26160),
	.C(n26159));
   NAND3xp33_ASAP7_75t_SRAM U27935 (.Y(n26164),
	.A(n26163),
	.B(n26162),
	.C(n20914));
   NOR2xp33_ASAP7_75t_SRAM U27936 (.Y(n26168),
	.A(n26167),
	.B(sa23_7_));
   A2O1A1Ixp33_ASAP7_75t_L U27937 (.Y(n26173),
	.A1(n26282),
	.A2(FE_OCPN5172_n26281),
	.B(FE_OFN27123_n26275),
	.C(FE_OCPN27373_n26172));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27939 (.Y(n26181),
	.A1(FE_OCPN7638_n26183),
	.A2(FE_OFN16163_n26584),
	.B(n26180),
	.C(n26185));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27940 (.Y(n26188),
	.A1(FE_OFN16163_n26584),
	.A2(FE_OCPN7638_n26183),
	.B(n26182),
	.C(n26181));
   OAI22xp33_ASAP7_75t_SRAM U27941 (.Y(n26184),
	.A1(text_in_r_66_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(n26185),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U27942 (.Y(n26199),
	.A1(n26942),
	.A2(n26201),
	.B(n26198),
	.C(n26508));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27943 (.Y(n26203),
	.A1(n26494),
	.A2(n27216),
	.B(FE_OCPN28307_n26491),
	.C(n26202));
   OAI22xp33_ASAP7_75t_SRAM U27944 (.Y(n26220),
	.A1(w1_17_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_81_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL U27946 (.Y(n26446),
	.A(FE_OFN16213_ld_r),
	.B(FE_OCPN27884_n26717));
   NOR2xp67_ASAP7_75t_SL U27947 (.Y(n26216),
	.A(n26446),
	.B(n26217));
   OAI22xp33_ASAP7_75t_SRAM U27948 (.Y(n26232),
	.A1(FE_OFN40_w0_19),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_115_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U27949 (.Y(n26224),
	.A1(FE_OFN16170_n26637),
	.A2(n26226),
	.B(n26222),
	.C(FE_OFN40_w0_19));
   O2A1O1Ixp33_ASAP7_75t_SL U27950 (.Y(n26238),
	.A1(FE_OCPN27451_n26236),
	.A2(n26235),
	.B(n26234),
	.C(n26233));
   OAI22xp33_ASAP7_75t_SRAM U27951 (.Y(n26265),
	.A1(w1_4_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_68_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   NAND2xp33_ASAP7_75t_SRAM U27952 (.Y(n26247),
	.A(FE_OFN26148_n26245),
	.B(n26243));
   A2O1A1Ixp33_ASAP7_75t_L U27953 (.Y(n26246),
	.A1(n26249),
	.A2(n26248),
	.B(FE_OFN26149_n26245),
	.C(FE_OFN58_w1_4));
   A2O1A1Ixp33_ASAP7_75t_SL U27954 (.Y(n26260),
	.A1(n26249),
	.A2(n26248),
	.B(n26247),
	.C(n26246));
   NOR2xp33_ASAP7_75t_L U27955 (.Y(n26257),
	.A(n26253),
	.B(FE_OFN16311_n26252));
   O2A1O1Ixp33_ASAP7_75t_L U27956 (.Y(n26256),
	.A1(FE_OFN16413_n26687),
	.A2(n26258),
	.B(n26255),
	.C(n26254));
   NOR2xp67_ASAP7_75t_SL U27958 (.Y(n26262),
	.A(n27031),
	.B(n26263));
   O2A1O1Ixp5_ASAP7_75t_SL U27959 (.Y(n508),
	.A1(w1_4_),
	.A2(text_in_r_68_),
	.B(n26265),
	.C(n26264));
   O2A1O1Ixp33_ASAP7_75t_SL U27960 (.Y(n26270),
	.A1(n26268),
	.A2(n26267),
	.B(FE_OCPN27447_n26638),
	.C(n26266));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27961 (.Y(n26279),
	.A1(FE_OCPN5172_n26281),
	.A2(n26282),
	.B(FE_OFN27123_n26275),
	.C(n26277));
   O2A1O1Ixp5_ASAP7_75t_SRAM U27962 (.Y(n26295),
	.A1(FE_OFN27043_n),
	.A2(FE_OCPN27516_n26292),
	.B(FE_OFN28808_n26291),
	.C(n26290));
   NAND3xp33_ASAP7_75t_SRAM U27963 (.Y(n26299),
	.A(n26296),
	.B(n26295),
	.C(n26294));
   NOR3xp33_ASAP7_75t_SRAM U27964 (.Y(n26314),
	.A(n26299),
	.B(n26298),
	.C(n26297));
   OAI21xp5_ASAP7_75t_L U27965 (.Y(n26305),
	.A1(FE_OCPN28156_n26304),
	.A2(n26303),
	.B(n26407));
   A2O1A1Ixp33_ASAP7_75t_SRAM U27966 (.Y(n26320),
	.A1(n26322),
	.A2(n26323),
	.B(n26319),
	.C(FE_OFN16340_n26317));
   A2O1A1Ixp33_ASAP7_75t_L U27967 (.Y(n26324),
	.A1(n26323),
	.A2(n26322),
	.B(n26321),
	.C(n26320));
   O2A1O1Ixp33_ASAP7_75t_SL U27968 (.Y(n26331),
	.A1(FE_OFN1_ld_r),
	.A2(n26330),
	.B(n26329),
	.C(n26328));
   O2A1O1Ixp5_ASAP7_75t_SL U27969 (.Y(n471),
	.A1(w2_3_),
	.A2(text_in_r_35_),
	.B(n26332),
	.C(n26331));
   NAND3xp33_ASAP7_75t_SL U27970 (.Y(n26333),
	.A(FE_OCPN28110_n),
	.B(FE_OCPN27991_n26336),
	.C(n26334));
   A2O1A1Ixp33_ASAP7_75t_SL U27971 (.Y(n26338),
	.A1(FE_OCPN27991_n26336),
	.A2(FE_OCPN28110_n),
	.B(n26334),
	.C(n26333));
   A2O1A1Ixp33_ASAP7_75t_SL U27972 (.Y(n26343),
	.A1(FE_OCPN27534_n),
	.A2(FE_OFN28490_ld_r),
	.B(n26338),
	.C(n26337));
   NOR3xp33_ASAP7_75t_SL U27973 (.Y(n26352),
	.A(n26353),
	.B(FE_OFN16214_ld_r),
	.C(n26732));
   A2O1A1Ixp33_ASAP7_75t_SL U27974 (.Y(n460),
	.A1(n26357),
	.A2(n26356),
	.B(n26355),
	.C(n26354));
   A2O1A1Ixp33_ASAP7_75t_L U27975 (.Y(n26365),
	.A1(n27117),
	.A2(FE_OFN28846_n26367),
	.B(FE_OCPN27744_n26362),
	.C(n26363));
   A2O1A1Ixp33_ASAP7_75t_SL U27976 (.Y(n26370),
	.A1(n26372),
	.A2(n27062),
	.B(FE_OCPN27357_n26369),
	.C(n26375));
   FAx1_ASAP7_75t_SL U27977 (.SN(n26378),
	.A(FE_OCPN27765_FE_OFN16265_n26527),
	.B(FE_OFN28968_n26780),
	.CI(n26373));
   NAND3xp33_ASAP7_75t_SL U27978 (.Y(n26379),
	.A(FE_OCPN28150_n27152),
	.B(FE_OCPN28173_n27153),
	.C(n26380));
   A2O1A1Ixp33_ASAP7_75t_SL U27979 (.Y(n26382),
	.A1(n27153),
	.A2(FE_OCPN28150_n27152),
	.B(n26380),
	.C(n26379));
   A2O1A1Ixp33_ASAP7_75t_SL U27980 (.Y(n26387),
	.A1(n26383),
	.A2(FE_OFN28483_ld_r),
	.B(n26382),
	.C(n26381));
   NAND2xp33_ASAP7_75t_R U27981 (.Y(n26386),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_125_));
   NAND3xp33_ASAP7_75t_SL U27982 (.Y(n26384),
	.A(n26385),
	.B(n26387),
	.C(n26386));
   A2O1A1Ixp33_ASAP7_75t_SL U27983 (.Y(n392),
	.A1(n26387),
	.A2(n26386),
	.B(n26385),
	.C(n26384));
   NAND2xp33_ASAP7_75t_SRAM U27984 (.Y(n26403),
	.A(FE_OFN26584_n20059),
	.B(n26399));
   NOR3xp33_ASAP7_75t_SRAM U27985 (.Y(n26405),
	.A(n26403),
	.B(n26402),
	.C(n26401));
   NAND3xp33_ASAP7_75t_SRAM U27986 (.Y(n26408),
	.A(n26406),
	.B(n26405),
	.C(FE_PSN8291_n26404));
   OAI21xp5_ASAP7_75t_SRAM U27987 (.Y(n26412),
	.A1(n26409),
	.A2(n26408),
	.B(n26407));
   NOR3xp33_ASAP7_75t_SL U27988 (.Y(n26419),
	.A(FE_OFN116_n27187),
	.B(FE_OCPN7589_n26420),
	.C(n27186));
   A2O1A1Ixp33_ASAP7_75t_SL U27989 (.Y(n26426),
	.A1(FE_OCPN5088_n27079),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B(n26422),
	.C(n26421));
   NAND2xp33_ASAP7_75t_R U27990 (.Y(n26425),
	.A(FE_OFN1_ld_r),
	.B(text_in_r_62_));
   NAND3xp33_ASAP7_75t_SL U27991 (.Y(n26423),
	.A(n26424),
	.B(n26426),
	.C(n26425));
   A2O1A1Ixp33_ASAP7_75t_SL U27992 (.Y(n473),
	.A1(n26426),
	.A2(n26425),
	.B(n26424),
	.C(n26423));
   A2O1A1Ixp33_ASAP7_75t_SL U27993 (.Y(n26438),
	.A1(FE_OCPN27525_n26434),
	.A2(FE_OFN28484_ld_r),
	.B(n26433),
	.C(n26432));
   NAND2xp33_ASAP7_75t_R U27994 (.Y(n26437),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_120_));
   O2A1O1Ixp5_ASAP7_75t_SL U27995 (.Y(n26445),
	.A1(FE_OCPN29458_n26442),
	.A2(n26441),
	.B(FE_OFN160_n26440),
	.C(n26439));
   NAND3xp33_ASAP7_75t_SL U27996 (.Y(n26447),
	.A(n26448),
	.B(n26450),
	.C(n26449));
   NAND3xp33_ASAP7_75t_SRAM U27997 (.Y(n26455),
	.A(n26453),
	.B(FE_OCPN29309_n26452),
	.C(FE_OCPN28305_n26451));
   OAI22xp33_ASAP7_75t_L U27998 (.Y(n26458),
	.A1(n26456),
	.A2(n26455),
	.B1(FE_OCPN27988_n26454),
	.B2(n26455));
   A2O1A1Ixp33_ASAP7_75t_L U28000 (.Y(n26480),
	.A1(FE_PSN8300_n26482),
	.A2(n27117),
	.B(FE_OCPN27494_n26479),
	.C(FE_OCPN29274_n26478));
   NOR3x1_ASAP7_75t_SL U28002 (.Y(n26483),
	.A(n26484),
	.B(FE_OFN2_ld_r),
	.C(n26895));
   NAND3x1_ASAP7_75t_L U28003 (.Y(n26485),
	.A(n26486),
	.B(n26488),
	.C(n26487));
   A2O1A1Ixp33_ASAP7_75t_SL U28004 (.Y(n350),
	.A1(n26488),
	.A2(n26487),
	.B(n26486),
	.C(n26485));
   A2O1A1Ixp33_ASAP7_75t_SL U28005 (.Y(n26500),
	.A1(n27216),
	.A2(n26494),
	.B(n26493),
	.C(n26492));
   FAx1_ASAP7_75t_SL U28006 (.SN(n26504),
	.A(FE_OCPN28054_n26501),
	.B(n26500),
	.CI(n26499));
   NOR2x1_ASAP7_75t_L U28007 (.Y(n27144),
	.A(FE_OFN12_FE_DBTN0_ld_r),
	.B(FE_OCPN29397_n26502));
   O2A1O1Ixp5_ASAP7_75t_SL U28008 (.Y(n494),
	.A1(w2_20_),
	.A2(text_in_r_52_),
	.B(n26506),
	.C(n26505));
   A2O1A1Ixp33_ASAP7_75t_L U28009 (.Y(n26509),
	.A1(n26915),
	.A2(n26914),
	.B(FE_OFN28473_n26911),
	.C(n26508));
   A2O1A1Ixp33_ASAP7_75t_L U28010 (.Y(n26519),
	.A1(n26915),
	.A2(n26914),
	.B(n26510),
	.C(n26509));
   O2A1O1Ixp5_ASAP7_75t_L U28012 (.Y(n455),
	.A1(w2_19_),
	.A2(text_in_r_51_),
	.B(n26524),
	.C(n26523));
   A2O1A1Ixp33_ASAP7_75t_L U28013 (.Y(n26529),
	.A1(n27117),
	.A2(n26531),
	.B(FE_OCPN29389_n26528),
	.C(FE_OFN16265_n26527));
   NOR3xp33_ASAP7_75t_SL U28014 (.Y(n26532),
	.A(FE_OCPN5056_n26535),
	.B(n26533),
	.C(n26534));
   OAI22xp33_ASAP7_75t_SRAM U28015 (.Y(n26543),
	.A1(text_in_r_103_),
	.A2(FE_OFN28484_ld_r),
	.B1(n26544),
	.B2(FE_OFN28484_ld_r));
   OAI22xp33_ASAP7_75t_SRAM U28016 (.Y(n26593),
	.A1(w1_3_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(text_in_r_67_),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   NOR2xp33_ASAP7_75t_SL U28017 (.Y(n26554),
	.A(n26553),
	.B(sa23_7_));
   NAND3xp33_ASAP7_75t_L U28018 (.Y(n26560),
	.A(n26557),
	.B(n26556),
	.C(n26555));
   NOR3xp33_ASAP7_75t_L U28019 (.Y(n26561),
	.A(n26560),
	.B(n26559),
	.C(n26558));
   A2O1A1Ixp33_ASAP7_75t_SL U28020 (.Y(n26703),
	.A1(n26573),
	.A2(FE_OCPN8258_n26572),
	.B(n26571),
	.C(n26570));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28021 (.Y(n26581),
	.A1(FE_OFN16163_n26584),
	.A2(n26583),
	.B(FE_OFN29029_n26579),
	.C(w1_3_));
   A2O1A1Ixp33_ASAP7_75t_L U28022 (.Y(n26585),
	.A1(FE_OFN16163_n26584),
	.A2(n26583),
	.B(n26582),
	.C(n26581));
   XOR2xp5_ASAP7_75t_SL U28023 (.Y(n26588),
	.A(n26587),
	.B(FE_OCPN27358_n26586));
   XOR2xp5_ASAP7_75t_SL U28024 (.Y(n26591),
	.A(n26589),
	.B(n26588));
   O2A1O1Ixp33_ASAP7_75t_SRAM U28025 (.Y(n26603),
	.A1(n26599),
	.A2(n26598),
	.B(n26139),
	.C(n26597));
   NOR2xp67_ASAP7_75t_SL U28026 (.Y(n26605),
	.A(n26601),
	.B(n26600));
   O2A1O1Ixp33_ASAP7_75t_SL U28027 (.Y(n26604),
	.A1(n26607),
	.A2(n26606),
	.B(n26603),
	.C(FE_OCPN29335_n));
   O2A1O1Ixp5_ASAP7_75t_SL U28028 (.Y(n26609),
	.A1(n26607),
	.A2(n26606),
	.B(n26605),
	.C(n26604));
   A2O1A1Ixp33_ASAP7_75t_SL U28029 (.Y(n26613),
	.A1(FE_OCPN29382_n26674),
	.A2(FE_OFN28487_ld_r),
	.B(n26609),
	.C(n26608));
   NAND2xp5_ASAP7_75t_L U28030 (.Y(n26617),
	.A(FE_OFN104_n27179),
	.B(n26615));
   A2O1A1Ixp33_ASAP7_75t_SL U28031 (.Y(n26619),
	.A1(n27183),
	.A2(n27182),
	.B(n26617),
	.C(n26616));
   A2O1A1Ixp33_ASAP7_75t_SL U28033 (.Y(n26627),
	.A1(n26625),
	.A2(n26624),
	.B(n26623),
	.C(n26622));
   NAND2xp5_ASAP7_75t_SL U28034 (.Y(n26635),
	.A(n26631),
	.B(n26630));
   A2O1A1Ixp33_ASAP7_75t_SL U28035 (.Y(n26634),
	.A1(FE_OFN16170_n26637),
	.A2(n26636),
	.B(FE_OCPN27284_n26633),
	.C(n26632));
   A2O1A1Ixp33_ASAP7_75t_SL U28036 (.Y(n27151),
	.A1(FE_OFN16170_n26637),
	.A2(n26636),
	.B(n26635),
	.C(n26634));
   NAND2xp5_ASAP7_75t_SL U28037 (.Y(n26641),
	.A(FE_OCPN27447_n26638),
	.B(n27057));
   A2O1A1Ixp33_ASAP7_75t_L U28038 (.Y(n26640),
	.A1(n27061),
	.A2(n27062),
	.B(n27058),
	.C(n26639));
   A2O1A1Ixp33_ASAP7_75t_SL U28039 (.Y(n26643),
	.A1(n27062),
	.A2(n27061),
	.B(n26641),
	.C(n26640));
   NOR2xp33_ASAP7_75t_SRAM U28041 (.Y(n26662),
	.A(n26660),
	.B(n26663));
   NOR2xp33_ASAP7_75t_SRAM U28042 (.Y(n26666),
	.A(FE_OCPN28112_n26664),
	.B(n26663));
   A2O1A1Ixp33_ASAP7_75t_SL U28043 (.Y(n26681),
	.A1(n26679),
	.A2(n26678),
	.B(n26677),
	.C(n26676));
   NOR3xp33_ASAP7_75t_SL U28044 (.Y(n26680),
	.A(FE_OCPN28383_n24808),
	.B(n26681),
	.C(n26682));
   O2A1O1Ixp5_ASAP7_75t_SL U28045 (.Y(n26696),
	.A1(FE_OCPN28383_n24808),
	.A2(n26682),
	.B(n26681),
	.C(n26680));
   OAI22xp33_ASAP7_75t_SRAM U28046 (.Y(n26691),
	.A1(text_in_r_71_),
	.A2(FE_OFN14_FE_DBTN0_ld_r),
	.B1(n26692),
	.B2(FE_OFN14_FE_DBTN0_ld_r));
   O2A1O1Ixp5_ASAP7_75t_SL U28047 (.Y(n498),
	.A1(w1_20_),
	.A2(text_in_r_84_),
	.B(n26719),
	.C(n26718));
   OAI22xp33_ASAP7_75t_SRAM U28048 (.Y(n26734),
	.A1(FE_OFN26072_n26720),
	.A2(FE_OFN28489_ld_r),
	.B1(text_in_r_20_),
	.B2(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U28049 (.Y(n26723),
	.A1(n26819),
	.A2(n26725),
	.B(n26722),
	.C(FE_OFN26072_n26720));
   NOR2xp33_ASAP7_75t_L U28050 (.Y(n26738),
	.A(n24306),
	.B(FE_OCPN5038_n26735));
   O2A1O1Ixp5_ASAP7_75t_L U28051 (.Y(n26737),
	.A1(n17506),
	.A2(n26739),
	.B(n26736),
	.C(FE_OFN133_n24306));
   A2O1A1Ixp33_ASAP7_75t_SL U28052 (.Y(n26746),
	.A1(n26742),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B(n26741),
	.C(n26740));
   A2O1A1Ixp33_ASAP7_75t_SL U28053 (.Y(n375),
	.A1(n26746),
	.A2(n26745),
	.B(n26744),
	.C(n26743));
   A2O1A1Ixp33_ASAP7_75t_R U28054 (.Y(n26751),
	.A1(n26915),
	.A2(n26753),
	.B(n26750),
	.C(n26749));
   A2O1A1Ixp33_ASAP7_75t_L U28055 (.Y(n27142),
	.A1(n26915),
	.A2(n26753),
	.B(n26752),
	.C(n26751));
   NOR2xp33_ASAP7_75t_SL U28056 (.Y(n26756),
	.A(n27110),
	.B(FE_OFN26650_n27164));
   O2A1O1Ixp5_ASAP7_75t_L U28057 (.Y(n26755),
	.A1(n27168),
	.A2(n27167),
	.B(n27163),
	.C(n26754));
   O2A1O1Ixp33_ASAP7_75t_SL U28058 (.Y(n26758),
	.A1(n27168),
	.A2(n27167),
	.B(n26756),
	.C(n26755));
   A2O1A1Ixp33_ASAP7_75t_SL U28059 (.Y(n26762),
	.A1(n27142),
	.A2(FE_OFN16215_ld_r),
	.B(n26758),
	.C(n26757));
   NAND2xp33_ASAP7_75t_R U28060 (.Y(n26761),
	.A(FE_OFN1_ld_r),
	.B(text_in_r_56_));
   A2O1A1Ixp33_ASAP7_75t_SL U28061 (.Y(n332),
	.A1(n26762),
	.A2(n26761),
	.B(n26760),
	.C(n26759));
   A2O1A1Ixp33_ASAP7_75t_SL U28062 (.Y(n26767),
	.A1(n26770),
	.A2(n26769),
	.B(n26766),
	.C(n26765));
   NOR2x1_ASAP7_75t_SL U28065 (.Y(n26782),
	.A(n26781),
	.B(n26783));
   O2A1O1Ixp5_ASAP7_75t_SL U28066 (.Y(n484),
	.A1(w0_3_),
	.A2(text_in_r_99_),
	.B(n26786),
	.C(n26785));
   NOR2xp33_ASAP7_75t_L U28067 (.Y(n26805),
	.A(n24306),
	.B(n26802));
   O2A1O1Ixp5_ASAP7_75t_L U28068 (.Y(n26804),
	.A1(n17463),
	.A2(n26806),
	.B(n26803),
	.C(FE_OFN133_n24306));
   O2A1O1Ixp5_ASAP7_75t_SL U28069 (.Y(n26808),
	.A1(n17463),
	.A2(n26806),
	.B(n26805),
	.C(n26804));
   A2O1A1Ixp33_ASAP7_75t_SL U28070 (.Y(n526),
	.A1(n26813),
	.A2(n26812),
	.B(n26811),
	.C(n26810));
   A2O1A1Ixp33_ASAP7_75t_SL U28071 (.Y(n26821),
	.A1(n26819),
	.A2(n26818),
	.B(n26817),
	.C(n26816));
   A2O1A1Ixp33_ASAP7_75t_SL U28072 (.Y(n26835),
	.A1(n26823),
	.A2(n26822),
	.B(n26821),
	.C(n26820));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28073 (.Y(n26826),
	.A1(n26828),
	.A2(n26829),
	.B(n26825),
	.C(FE_OCPN29502_w3_23));
   OAI22xp33_ASAP7_75t_SRAM U28074 (.Y(n26830),
	.A1(text_in_r_23_),
	.A2(FE_OFN28489_ld_r),
	.B1(FE_OCPN29502_w3_23),
	.B2(FE_OFN28489_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U28075 (.Y(n26854),
	.A1(FE_OFN29242_n26856),
	.A2(FE_OCPN29587_n26857),
	.B(FE_OCPN27377_n26853),
	.C(FE_OCPN27295_n26851));
   A2O1A1Ixp33_ASAP7_75t_SL U28076 (.Y(n26864),
	.A1(FE_OCPN27375_n26860),
	.A2(FE_OFN28489_ld_r),
	.B(n26859),
	.C(n26858));
   NAND3xp33_ASAP7_75t_SL U28077 (.Y(n26861),
	.A(FE_OFN26129_w3_15),
	.B(n26864),
	.C(n26863));
   A2O1A1Ixp33_ASAP7_75t_SL U28078 (.Y(n512),
	.A1(n26864),
	.A2(n26863),
	.B(FE_OFN26129_w3_15),
	.C(n26861));
   OAI22xp33_ASAP7_75t_SRAM U28079 (.Y(n26897),
	.A1(w0_20_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(text_in_r_116_),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_L U28080 (.Y(n26868),
	.A1(n27127),
	.A2(n27126),
	.B(n27122),
	.C(FE_OCPN27283_n26867));
   NOR2xp33_ASAP7_75t_SRAM U28081 (.Y(n26873),
	.A(n26871),
	.B(n26870));
   NAND3xp33_ASAP7_75t_SRAM U28082 (.Y(n26877),
	.A(n26874),
	.B(n26873),
	.C(n26872));
   NOR3xp33_ASAP7_75t_SRAM U28083 (.Y(n26888),
	.A(n26877),
	.B(n26876),
	.C(n26875));
   O2A1O1Ixp5_ASAP7_75t_SL U28084 (.Y(n513),
	.A1(w0_20_),
	.A2(text_in_r_116_),
	.B(n26897),
	.C(n26896));
   A2O1A1Ixp33_ASAP7_75t_SL U28085 (.Y(n26905),
	.A1(n26942),
	.A2(n26907),
	.B(n26904),
	.C(n26903));
   NAND2xp5_ASAP7_75t_L U28086 (.Y(n26913),
	.A(FE_OCPN27302_n26910),
	.B(FE_OFN26558_n26911));
   A2O1A1Ixp33_ASAP7_75t_SL U28087 (.Y(n26912),
	.A1(n26914),
	.A2(n26915),
	.B(FE_OFN28473_n26911),
	.C(n26910));
   A2O1A1Ixp33_ASAP7_75t_SL U28088 (.Y(n26917),
	.A1(n26915),
	.A2(n26914),
	.B(n26913),
	.C(n26912));
   NOR2xp33_ASAP7_75t_SL U28090 (.Y(n26925),
	.A(n26923),
	.B(FE_OFN28451_n26990));
   O2A1O1Ixp33_ASAP7_75t_SL U28091 (.Y(n26929),
	.A1(n26926),
	.A2(n26995),
	.B(n26925),
	.C(n26924));
   A2O1A1Ixp33_ASAP7_75t_SL U28092 (.Y(n26934),
	.A1(FE_OFN28487_ld_r),
	.A2(FE_OCPN29576_n26930),
	.B(n26929),
	.C(n26928));
   NAND2xp33_ASAP7_75t_R U28093 (.Y(n26933),
	.A(FE_OFN16214_ld_r),
	.B(text_in_r_72_));
   A2O1A1Ixp33_ASAP7_75t_L U28095 (.Y(n26939),
	.A1(n26942),
	.A2(n26941),
	.B(n26938),
	.C(n26937));
   NOR3xp33_ASAP7_75t_L U28096 (.Y(n26943),
	.A(n26946),
	.B(n26944),
	.C(n26945));
   O2A1O1Ixp33_ASAP7_75t_L U28097 (.Y(n26948),
	.A1(n26946),
	.A2(n26945),
	.B(FE_OCPN8249_n26944),
	.C(n26943));
   A2O1A1Ixp33_ASAP7_75t_L U28098 (.Y(n26953),
	.A1(FE_OCPN8246_n27143),
	.A2(FE_OFN16215_ld_r),
	.B(n26948),
	.C(n26947));
   FAx1_ASAP7_75t_SL U28099 (.SN(n26966),
	.A(FE_OCPN27442_n27202),
	.B(FE_OCPN27271_n26961),
	.CI(n26960));
   OAI22xp33_ASAP7_75t_SRAM U28100 (.Y(n26962),
	.A1(text_in_r_43_),
	.A2(FE_OFN16215_ld_r),
	.B1(n26963),
	.B2(FE_OFN16215_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U28101 (.Y(n467),
	.A1(n27176),
	.A2(n26966),
	.B(n26965),
	.C(n26964));
   NOR3xp33_ASAP7_75t_SRAM U28102 (.Y(n26975),
	.A(n26969),
	.B(FE_OCPN27685_n26968),
	.C(n26967));
   OAI21xp33_ASAP7_75t_SRAM U28103 (.Y(n26973),
	.A1(FE_OFN28941_sa02_2),
	.A2(FE_OCPN29533_n26971),
	.B(FE_OCPN29423_n26970));
   O2A1O1Ixp5_ASAP7_75t_SRAM U28104 (.Y(n26984),
	.A1(FE_OCPN28316_n26980),
	.A2(n26979),
	.B(n27216),
	.C(n26978));
   NAND3xp33_ASAP7_75t_SL U28105 (.Y(n26981),
	.A(n26982),
	.B(n26984),
	.C(FE_OCPN7583_n26983));
   A2O1A1Ixp33_ASAP7_75t_SL U28106 (.Y(n26986),
	.A1(n26984),
	.A2(FE_OCPN7583_n26983),
	.B(n26982),
	.C(n26981));
   O2A1O1Ixp33_ASAP7_75t_SL U28107 (.Y(n408),
	.A1(n26989),
	.A2(n26988),
	.B(w2_16_),
	.C(n26987));
   NAND3xp33_ASAP7_75t_SL U28108 (.Y(n27000),
	.A(n26999),
	.B(n26998),
	.C(n26997));
   NAND3xp33_ASAP7_75t_SL U28110 (.Y(n27013),
	.A(FE_OFN16307_n27010),
	.B(n27009),
	.C(n27008));
   NOR3xp33_ASAP7_75t_L U28111 (.Y(n27016),
	.A(n27013),
	.B(n27012),
	.C(n27011));
   A2O1A1Ixp33_ASAP7_75t_SL U28112 (.Y(n27018),
	.A1(n27017),
	.A2(n27016),
	.B(n27015),
	.C(n27014));
   FAx1_ASAP7_75t_SL U28113 (.SN(n27033),
	.A(FE_OCPN27439_n27030),
	.B(n27029),
	.CI(n27028));
   NOR2xp33_ASAP7_75t_SRAM U28115 (.Y(n27038),
	.A(n27037),
	.B(FE_OFN28499_sa00_6));
   NOR3xp33_ASAP7_75t_SRAM U28116 (.Y(n27042),
	.A(FE_OFN26147_n27041),
	.B(n27040),
	.C(n27039));
   NOR2xp33_ASAP7_75t_SRAM U28117 (.Y(n27044),
	.A(n27042),
	.B(FE_OFN28499_sa00_6));
   A2O1A1Ixp33_ASAP7_75t_SL U28118 (.Y(n27054),
	.A1(n27117),
	.A2(n27052),
	.B(n27051),
	.C(n27050));
   NOR3xp33_ASAP7_75t_SL U28119 (.Y(n27053),
	.A(FE_OCPN28442_n27056),
	.B(n27054),
	.C(n27055));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28120 (.Y(n27059),
	.A1(n27061),
	.A2(n27062),
	.B(n27058),
	.C(n27064));
   OAI22xp33_ASAP7_75t_SRAM U28121 (.Y(n27063),
	.A1(text_in_r_119_),
	.A2(FE_OFN15_FE_DBTN0_ld_r),
	.B1(n27064),
	.B2(FE_OFN15_FE_DBTN0_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U28122 (.Y(n506),
	.A1(n27068),
	.A2(n27067),
	.B(n27066),
	.C(n27065));
   NOR2xp33_ASAP7_75t_SRAM U28123 (.Y(n27077),
	.A(n27070),
	.B(n27069));
   NOR3xp33_ASAP7_75t_SRAM U28124 (.Y(n27076),
	.A(n27073),
	.B(n27072),
	.C(n27071));
   A2O1A1Ixp33_ASAP7_75t_L U28125 (.Y(n27081),
	.A1(n27077),
	.A2(n27076),
	.B(n27075),
	.C(n27074));
   A2O1A1Ixp33_ASAP7_75t_SL U28127 (.Y(n27087),
	.A1(FE_OCPN7650_n27110),
	.A2(FE_OFN16215_ld_r),
	.B(n27083),
	.C(n27082));
   NAND3xp33_ASAP7_75t_SRAM U28128 (.Y(n27093),
	.A(n27090),
	.B(n27089),
	.C(n27088));
   NOR3xp33_ASAP7_75t_SRAM U28129 (.Y(n27096),
	.A(n27093),
	.B(FE_OFN28548_n27092),
	.C(n27091));
   O2A1O1Ixp33_ASAP7_75t_R U28130 (.Y(n27099),
	.A1(n27102),
	.A2(n27101),
	.B(n27098),
	.C(n27106));
   O2A1O1Ixp33_ASAP7_75t_L U28131 (.Y(n27103),
	.A1(n27102),
	.A2(n27101),
	.B(n27100),
	.C(n27099));
   OAI22xp33_ASAP7_75t_SRAM U28132 (.Y(n27105),
	.A1(text_in_r_57_),
	.A2(FE_OFN16215_ld_r),
	.B1(n27106),
	.B2(FE_OFN16215_ld_r));
   A2O1A1Ixp33_ASAP7_75t_SL U28133 (.Y(n409),
	.A1(FE_OFN26559_n26754),
	.A2(n27109),
	.B(n27108),
	.C(n27107));
   A2O1A1Ixp33_ASAP7_75t_SL U28134 (.Y(n27114),
	.A1(n27117),
	.A2(n27116),
	.B(FE_OFN29010_n27113),
	.C(n27151));
   A2O1A1Ixp33_ASAP7_75t_SL U28135 (.Y(n27119),
	.A1(n27117),
	.A2(n27116),
	.B(n27115),
	.C(n27114));
   NOR3xp33_ASAP7_75t_SL U28136 (.Y(n27118),
	.A(FE_OCPN27641_n27121),
	.B(n27119),
	.C(n27120));
   O2A1O1Ixp33_ASAP7_75t_SL U28137 (.Y(n27133),
	.A1(FE_OCPN27641_n27121),
	.A2(n27120),
	.B(n27119),
	.C(n27118));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28138 (.Y(n27124),
	.A1(n27126),
	.A2(n27127),
	.B(n27122),
	.C(n27129));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28139 (.Y(n27132),
	.A1(n27127),
	.A2(n27126),
	.B(n27125),
	.C(n27124));
   OAI22xp33_ASAP7_75t_SRAM U28140 (.Y(n27149),
	.A1(w2_17_),
	.A2(FE_OFN16_FE_DBTN0_ld_r),
	.B1(text_in_r_49_),
	.B2(FE_OFN16_FE_DBTN0_ld_r));
   O2A1O1Ixp33_ASAP7_75t_R U28141 (.Y(n27137),
	.A1(n27140),
	.A2(n27139),
	.B(n27136),
	.C(n27135));
   O2A1O1Ixp33_ASAP7_75t_L U28142 (.Y(n27141),
	.A1(n27140),
	.A2(n27139),
	.B(n27138),
	.C(n27137));
   NAND3xp33_ASAP7_75t_L U28143 (.Y(n27150),
	.A(FE_OCPN28150_n27152),
	.B(FE_OCPN28173_n27153),
	.C(FE_OFN16329_n27151));
   A2O1A1Ixp33_ASAP7_75t_L U28144 (.Y(n27156),
	.A1(FE_OCPN28173_n27153),
	.A2(FE_OCPN28150_n27152),
	.B(FE_OFN16329_n27151),
	.C(n27150));
   NAND2xp33_ASAP7_75t_R U28145 (.Y(n27161),
	.A(FE_OFN2_ld_r),
	.B(text_in_r_109_));
   NAND3xp33_ASAP7_75t_SL U28146 (.Y(n27159),
	.A(n27160),
	.B(n27162),
	.C(n27161));
   NAND2xp33_ASAP7_75t_SL U28147 (.Y(n27181),
	.A(FE_OFN104_n27179),
	.B(FE_OFN105_n27178));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28149 (.Y(n27190),
	.A1(n27192),
	.A2(FE_OFN16176_n27207),
	.B(n27188),
	.C(n27195));
   A2O1A1Ixp33_ASAP7_75t_SL U28150 (.Y(n27204),
	.A1(FE_OFN16177_n27207),
	.A2(n27206),
	.B(FE_OCPN29445_n27203),
	.C(n27202));
   A2O1A1Ixp33_ASAP7_75t_SRAM U28151 (.Y(n27213),
	.A1(n27215),
	.A2(n27216),
	.B(n27212),
	.C(n27219));
   A2O1A1Ixp33_ASAP7_75t_R U28152 (.Y(n27222),
	.A1(n27216),
	.A2(n27215),
	.B(n27214),
	.C(n27213));
endmodule

