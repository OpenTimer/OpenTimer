module ac97_ctrl (
x1542,
x1203,
x806,
x1557,
x130646,
x1390,
x1424,
x1564,
x1511,
x1006,
x1486,
x1398,
x1459,
x130629,
x130652,
x130647,
x1572,
x130631,
x1587,
x130641,
x1322,
x130638,
x1501,
x1209,
x1432,
x1215,
x130633,
x1155,
x130637,
x1451,
x1519,
x1062,
x1358,
x1261,
x940,
x130632,
x906,
x1417,
x1034,
x130648,
x1101,
x130649,
x1580,
x130636,
x130644,
x1406,
x821,
x1822,
x1494,
x977,
x1286,
x1126,
x130654,
x130657,
x1231,
x837,
x130645,
x1550,
x130656,
x130651,
x130655,
x1345,
x1479,
x130635,
x1527,
x130640,
x1351,
x130634,
x1374,
x1382,
x130639,
x1467,
x130630,
x130642,
x130643,
x1193,
x1366,
x868,
x889,
x1534,
x130650,
x130653,
x1595,
x1443,
x718,
x124,
x30,
x589,
x397,
x84,
x217,
x765,
x361,
x149,
x138,
x315,
x522,
x172,
x786,
x131,
x681,
x476,
x145,
x638,
x390,
x63,
x379,
x447,
x96,
x179,
x699,
x195,
x0,
x106,
x420,
x101,
x620,
x187,
x538,
x264,
x744,
x234,
x114,
x77,
x657,
x342,
x494,
x14,
x287,
x561,
x249,
x38);

// Start PIs
input x1542;
input x1203;
input x806;
input x1557;
input x130646;
input x1390;
input x1424;
input x1564;
input x1511;
input x1006;
input x1486;
input x1398;
input x1459;
input x130629;
input x130652;
input x130647;
input x1572;
input x130631;
input x1587;
input x130641;
input x1322;
input x130638;
input x1501;
input x1209;
input x1432;
input x1215;
input x130633;
input x1155;
input x130637;
input x1451;
input x1519;
input x1062;
input x1358;
input x1261;
input x940;
input x130632;
input x906;
input x1417;
input x1034;
input x130648;
input x1101;
input x130649;
input x1580;
input x130636;
input x130644;
input x1406;
input x821;
input x1822;
input x1494;
input x977;
input x1286;
input x1126;
input x130654;
input x130657;
input x1231;
input x837;
input x130645;
input x1550;
input x130656;
input x130651;
input x130655;
input x1345;
input x1479;
input x130635;
input x1527;
input x130640;
input x1351;
input x130634;
input x1374;
input x1382;
input x130639;
input x1467;
input x130630;
input x130642;
input x130643;
input x1193;
input x1366;
input x868;
input x889;
input x1534;
input x130650;
input x130653;
input x1595;
input x1443;

// Start POs
output x718;
output x124;
output x30;
output x589;
output x397;
output x84;
output x217;
output x765;
output x361;
output x149;
output x138;
output x315;
output x522;
output x172;
output x786;
output x131;
output x681;
output x476;
output x145;
output x638;
output x390;
output x63;
output x379;
output x447;
output x96;
output x179;
output x699;
output x195;
output x0;
output x106;
output x420;
output x101;
output x620;
output x187;
output x538;
output x264;
output x744;
output x234;
output x114;
output x77;
output x657;
output x342;
output x494;
output x14;
output x287;
output x561;
output x249;
output x38;

// Start wires
wire net_8298;
wire net_8631;
wire net_4065;
wire net_11968;
wire net_4854;
wire net_2418;
wire net_14199;
wire net_7279;
wire net_943;
wire net_11788;
wire net_10413;
wire net_4598;
wire net_4392;
wire net_11330;
wire net_12833;
wire net_1897;
wire net_9435;
wire net_980;
wire net_13088;
wire net_5499;
wire net_9803;
wire net_2542;
wire net_12029;
wire net_7081;
wire net_10629;
wire net_11370;
wire net_5515;
wire net_3996;
wire net_11996;
wire net_7594;
wire net_6241;
wire net_7298;
wire net_4382;
wire net_13988;
wire net_12537;
wire net_13226;
wire net_12501;
wire net_8105;
wire net_4934;
wire net_2256;
wire net_4306;
wire net_264;
wire net_12959;
wire net_11178;
wire net_12809;
wire net_3904;
wire net_4122;
wire net_4315;
wire net_8914;
wire net_11757;
wire net_9072;
wire net_2769;
wire net_8503;
wire net_11190;
wire net_4996;
wire net_14016;
wire net_3707;
wire net_1064;
wire net_14405;
wire net_2082;
wire net_10165;
wire net_6227;
wire net_7173;
wire net_5035;
wire net_12907;
wire net_4832;
wire net_4464;
wire net_8577;
wire net_9784;
wire net_12704;
wire net_13544;
wire net_10988;
wire net_7191;
wire net_703;
wire net_5330;
wire net_193;
wire net_11377;
wire net_9989;
wire net_12447;
wire net_6037;
wire net_14381;
wire net_10554;
wire net_6773;
wire net_5273;
wire net_12413;
wire net_7283;
wire net_5627;
wire net_2942;
wire net_3817;
wire net_9441;
wire net_13993;
wire net_3281;
wire net_13916;
wire net_10659;
wire net_4442;
wire net_3949;
wire net_3134;
wire net_13458;
wire net_8185;
wire net_10215;
wire net_5523;
wire net_1720;
wire net_14164;
wire net_13885;
wire net_8191;
wire net_6231;
wire net_3818;
wire net_3434;
wire net_6104;
wire net_2060;
wire net_2051;
wire net_6087;
wire net_4535;
wire net_9464;
wire net_3756;
wire net_6426;
wire net_593;
wire net_5563;
wire net_10156;
wire net_6238;
wire net_4169;
wire net_2765;
wire net_13451;
wire net_7845;
wire net_9957;
wire net_11979;
wire net_742;
wire net_8341;
wire net_5139;
wire net_6384;
wire net_11044;
wire net_12976;
wire net_9597;
wire net_7092;
wire net_10343;
wire net_2830;
wire net_10320;
wire net_4509;
wire net_1198;
wire net_3975;
wire net_2862;
wire net_8100;
wire net_2457;
wire net_8260;
wire net_883;
wire net_13476;
wire net_11605;
wire net_8124;
wire net_4108;
wire net_9970;
wire net_5533;
wire net_2957;
wire net_446;
wire net_1516;
wire net_1712;
wire net_6782;
wire net_6473;
wire net_3063;
wire net_1083;
wire net_3423;
wire net_1499;
wire net_964;
wire net_2913;
wire net_8242;
wire net_3295;
wire net_13729;
wire net_6402;
wire net_11003;
wire net_4379;
wire net_2268;
wire net_10000;
wire net_6114;
wire net_14352;
wire net_2846;
wire net_2303;
wire net_13331;
wire net_11685;
wire net_9479;
wire net_4369;
wire net_1735;
wire net_2210;
wire net_8249;
wire net_2176;
wire net_13191;
wire net_11933;
wire net_8563;
wire net_997;
wire net_12243;
wire net_10837;
wire net_6401;
wire net_11060;
wire net_10007;
wire net_256;
wire net_8762;
wire net_4929;
wire net_3959;
wire net_4309;
wire net_8873;
wire net_12393;
wire net_11226;
wire net_6573;
wire net_1140;
wire net_2764;
wire net_1464;
wire net_7490;
wire net_10931;
wire net_5797;
wire net_11985;
wire net_4973;
wire net_12891;
wire net_3196;
wire net_5962;
wire net_515;
wire net_4835;
wire net_10620;
wire net_5342;
wire net_13216;
wire net_11124;
wire net_7463;
wire net_6806;
wire net_5121;
wire net_3987;
wire net_223;
wire net_6557;
wire net_7146;
wire net_2077;
wire net_8468;
wire net_7496;
wire net_2219;
wire net_2745;
wire net_7343;
wire net_11166;
wire net_5680;
wire net_13973;
wire net_5084;
wire net_3965;
wire net_13827;
wire net_7483;
wire net_1876;
wire net_13130;
wire net_6706;
wire net_130;
wire net_7212;
wire net_572;
wire net_9810;
wire net_5289;
wire net_10955;
wire net_9614;
wire net_5116;
wire net_369;
wire net_12709;
wire net_12051;
wire net_7850;
wire net_1662;
wire net_10396;
wire net_4358;
wire net_7543;
wire net_9835;
wire net_1079;
wire net_10495;
wire net_7959;
wire net_3935;
wire net_11290;
wire net_10148;
wire net_6760;
wire net_5198;
wire net_2809;
wire net_14318;
wire net_3235;
wire net_780;
wire net_4938;
wire net_3586;
wire net_3184;
wire net_7099;
wire net_6812;
wire net_12226;
wire net_13261;
wire net_9272;
wire net_2391;
wire net_10095;
wire net_5263;
wire net_2802;
wire net_11350;
wire net_7965;
wire net_4614;
wire net_2906;
wire net_456;
wire net_155;
wire net_12555;
wire net_11357;
wire net_9301;
wire net_11299;
wire net_10636;
wire net_7238;
wire net_3850;
wire net_9153;
wire net_9023;
wire net_8222;
wire net_349;
wire net_12923;
wire net_8533;
wire net_14367;
wire net_8547;
wire net_3428;
wire net_1409;
wire net_12576;
wire net_2977;
wire net_493;
wire net_6374;
wire net_6080;
wire net_14306;
wire net_13140;
wire net_6506;
wire net_13679;
wire net_1428;
wire net_987;
wire net_13137;
wire net_6167;
wire net_5222;
wire net_3620;
wire net_10510;
wire net_14340;
wire net_7781;
wire net_13824;
wire net_4238;
wire net_5844;
wire net_8475;
wire net_2350;
wire net_6293;
wire x1366;
wire net_3271;
wire net_13183;
wire net_11197;
wire net_10675;
wire net_13098;
wire net_12568;
wire net_10506;
wire net_5740;
wire net_12276;
wire net_12418;
wire net_721;
wire net_12366;
wire net_9033;
wire net_8950;
wire net_7779;
wire net_3226;
wire net_3143;
wire net_8164;
wire net_12127;
wire net_9819;
wire net_2757;
wire net_13634;
wire net_12776;
wire net_9531;
wire net_1018;
wire net_11085;
wire net_3629;
wire net_7315;
wire net_11701;
wire net_2369;
wire net_2038;
wire net_13289;
wire net_6591;
wire net_823;
wire net_9067;
wire net_12878;
wire net_9269;
wire net_1676;
wire net_7271;
wire net_4788;
wire net_14230;
wire net_698;
wire net_12969;
wire net_11774;
wire net_9541;
wire net_7892;
wire net_14374;
wire net_11028;
wire net_5428;
wire net_1191;
wire net_13688;
wire net_5259;
wire net_8515;
wire net_2255;
wire net_4649;
wire net_4754;
wire net_2485;
wire net_13906;
wire net_6967;
wire net_3857;
wire net_8970;
wire net_7471;
wire net_12918;
wire net_749;
wire net_11729;
wire net_1019;
wire net_1948;
wire net_1616;
wire net_11500;
wire net_11898;
wire net_6180;
wire net_10348;
wire net_1006;
wire net_2781;
wire net_9415;
wire net_6767;
wire net_14181;
wire net_4342;
wire net_9724;
wire net_12863;
wire net_2969;
wire net_7839;
wire net_7518;
wire net_12522;
wire net_12351;
wire net_5490;
wire net_12960;
wire net_13167;
wire net_7544;
wire net_11406;
wire net_8886;
wire net_2985;
wire net_11551;
wire net_537;
wire net_3056;
wire net_14050;
wire net_12943;
wire net_11310;
wire net_10893;
wire net_8710;
wire net_12477;
wire net_3614;
wire net_7624;
wire net_13446;
wire net_13007;
wire net_5501;
wire net_12294;
wire net_3252;
wire net_6792;
wire net_5790;
wire net_5891;
wire net_513;
wire net_12020;
wire net_7950;
wire net_1576;
wire net_1421;
wire net_14282;
wire net_12462;
wire net_9525;
wire net_4496;
wire net_8737;
wire net_6067;
wire net_3407;
wire net_2736;
wire net_2127;
wire net_1280;
wire net_459;
wire net_12616;
wire net_9239;
wire net_8720;
wire net_13569;
wire net_3656;
wire net_737;
wire net_6590;
wire net_2284;
wire net_3412;
wire net_2113;
wire net_13305;
wire net_9397;
wire net_4793;
wire net_5865;
wire net_13372;
wire x1390;
wire net_4760;
wire net_3915;
wire net_12737;
wire net_5957;
wire net_5606;
wire net_11722;
wire net_11541;
wire net_12375;
wire net_5201;
wire net_8063;
wire net_8353;
wire net_1156;
wire net_14127;
wire net_5150;
wire net_13641;
wire net_1966;
wire net_13049;
wire net_14299;
wire net_12188;
wire net_11718;
wire net_4571;
wire net_9212;
wire net_12713;
wire net_8176;
wire net_12873;
wire net_5977;
wire net_11493;
wire net_7709;
wire net_12672;
wire net_1659;
wire net_326;
wire net_2381;
wire net_589;
wire net_11012;
wire net_10286;
wire net_9504;
wire net_1814;
wire net_5403;
wire net_11610;
wire net_5981;
wire net_10242;
wire net_6735;
wire net_6668;
wire net_3175;
wire net_10186;
wire net_10076;
wire net_7319;
wire net_2829;
wire net_10288;
wire net_8698;
wire net_724;
wire net_9826;
wire net_9123;
wire net_4815;
wire net_4099;
wire net_3142;
wire net_1219;
wire net_12826;
wire net_14410;
wire net_8058;
wire net_10886;
wire net_10871;
wire net_13815;
wire net_2384;
wire net_3884;
wire net_7760;
wire net_8745;
wire net_3736;
wire net_2877;
wire net_5889;
wire net_2480;
wire net_9943;
wire net_12181;
wire net_9868;
wire net_9352;
wire net_874;
wire net_8334;
wire net_13706;
wire net_1632;
wire net_3796;
wire net_1661;
wire net_11399;
wire net_1236;
wire net_13627;
wire net_4277;
wire net_13771;
wire net_8987;
wire net_7907;
wire net_12107;
wire net_3674;
wire net_7555;
wire net_2700;
wire net_7996;
wire net_7868;
wire net_10307;
wire net_9548;
wire net_6841;
wire net_6273;
wire net_1488;
wire net_6187;
wire net_4966;
wire net_2812;
wire net_5244;
wire net_12721;
wire net_10178;
wire net_5691;
wire net_352;
wire net_11182;
wire net_9320;
wire net_12857;
wire net_3920;
wire net_436;
wire net_2837;
wire net_7963;
wire net_7181;
wire net_5641;
wire net_11157;
wire net_2824;
wire net_6342;
wire net_1777;
wire net_12983;
wire net_8263;
wire net_7373;
wire net_13647;
wire net_7903;
wire net_1641;
wire net_7511;
wire net_12325;
wire net_7246;
wire net_12153;
wire net_12134;
wire net_5556;
wire net_4919;
wire net_1702;
wire net_1103;
wire net_4403;
wire net_767;
wire net_7974;
wire net_6358;
wire net_1838;
wire net_4557;
wire net_11365;
wire net_10857;
wire net_131;
wire net_9754;
wire net_5488;
wire net_358;
wire net_1973;
wire net_8693;
wire net_8748;
wire net_7564;
wire net_4292;
wire net_2016;
wire net_14169;
wire net_2934;
wire net_7702;
wire net_10486;
wire x84;
wire net_11427;
wire net_3125;
wire x1126;
wire net_1285;
wire net_10364;
wire net_5912;
wire net_3112;
wire net_13952;
wire net_1175;
wire net_13207;
wire net_13118;
wire net_12544;
wire net_10962;
wire net_9453;
wire net_6550;
wire x476;
wire net_9101;
wire net_9934;
wire net_5722;
wire net_13021;
wire net_9312;
wire net_9191;
wire net_2922;
wire net_9022;
wire net_10043;
wire net_1742;
wire net_13321;
wire net_11884;
wire net_7526;
wire net_7641;
wire net_11823;
wire net_468;
wire net_9308;
wire net_6890;
wire net_9372;
wire net_9257;
wire net_11654;
wire net_9738;
wire net_8011;
wire net_13734;
wire net_3370;
wire net_7025;
wire net_13040;
wire net_9497;
wire net_3947;
wire net_3441;
wire net_179;
wire net_9665;
wire net_4947;
wire net_4015;
wire net_3662;
wire net_10171;
wire net_12730;
wire net_8677;
wire net_8729;
wire net_3261;
wire net_9187;
wire net_13441;
wire net_6349;
wire net_2289;
wire net_10756;
wire x1587;
wire net_7300;
wire net_11244;
wire net_6759;
wire net_5919;
wire net_3539;
wire net_2031;
wire net_1868;
wire net_1560;
wire net_13942;
wire net_4414;
wire net_12451;
wire net_4409;
wire net_10110;
wire net_7205;
wire net_12160;
wire net_10453;
wire net_6754;
wire net_13690;
wire net_12684;
wire net_3863;
wire net_10538;
wire net_9856;
wire net_8538;
wire net_9684;
wire net_8715;
wire net_14227;
wire net_13111;
wire net_5778;
wire net_7724;
wire net_6489;
wire net_3382;
wire net_4257;
wire net_1545;
wire net_13756;
wire net_4662;
wire net_4872;
wire net_8204;
wire net_990;
wire net_10798;
wire net_13838;
wire net_11728;
wire net_11485;
wire net_7423;
wire net_10428;
wire net_10473;
wire net_11763;
wire net_2332;
wire net_3774;
wire net_12491;
wire net_2715;
wire net_1803;
wire net_13803;
wire net_1941;
wire net_8031;
wire net_13074;
wire net_1134;
wire net_13968;
wire net_14276;
wire net_3899;
wire net_363;
wire net_1319;
wire net_8757;
wire net_776;
wire net_4550;
wire net_3080;
wire net_11075;
wire net_2508;
wire net_12118;
wire net_9624;
wire net_10353;
wire net_8451;
wire net_1650;
wire net_1582;
wire net_13574;
wire net_12696;
wire net_10717;
wire net_3149;
wire net_11253;
wire net_6454;
wire net_1675;
wire net_4016;
wire net_2247;
wire net_6028;
wire net_13747;
wire net_2333;
wire net_6544;
wire net_6464;
wire net_8115;
wire net_1368;
wire net_1248;
wire net_6525;
wire net_2291;
wire net_11108;
wire net_10531;
wire net_2238;
wire net_845;
wire net_10745;
wire x287;
wire net_8003;
wire net_10973;
wire net_11096;
wire net_9081;
wire net_8414;
wire net_695;
wire net_12404;
wire net_7692;
wire net_2525;
wire net_1201;
wire net_14086;
wire net_12073;
wire net_2671;
wire net_9701;
wire net_6787;
wire net_6569;
wire net_14331;
wire net_5106;
wire net_8074;
wire net_13852;
wire net_12761;
wire net_859;
wire net_7259;
wire net_1167;
wire net_5896;
wire net_12788;
wire net_8636;
wire net_12610;
wire net_2198;
wire net_9043;
wire net_1044;
wire net_5250;
wire net_6435;
wire net_6661;
wire net_4322;
wire net_10948;
wire net_2940;
wire net_10617;
wire net_8672;
wire net_2043;
wire net_6775;
wire net_5583;
wire net_2095;
wire net_4681;
wire net_6955;
wire net_5231;
wire net_10662;
wire net_9726;
wire net_2314;
wire net_9905;
wire net_5454;
wire net_2613;
wire net_9995;
wire net_3605;
wire net_14336;
wire net_12174;
wire net_10865;
wire net_6635;
wire net_9010;
wire net_8849;
wire net_11055;
wire net_7250;
wire net_4114;
wire net_14220;
wire net_11479;
wire net_10330;
wire net_865;
wire net_13500;
wire net_9896;
wire net_231;
wire net_10197;
wire net_13326;
wire net_2621;
wire net_13832;
wire net_3024;
wire net_1223;
wire net_4691;
wire net_2750;
wire net_5816;
wire net_11961;
wire net_926;
wire net_4623;
wire net_12381;
wire net_7264;
wire net_7403;
wire net_4223;
wire net_6153;
wire net_11321;
wire net_8642;
wire net_2297;
wire net_13052;
wire net_9439;
wire net_7188;
wire net_3325;
wire net_12868;
wire net_10595;
wire net_9185;
wire net_6466;
wire net_6171;
wire net_2048;
wire net_582;
wire net_12485;
wire net_4481;
wire net_7419;
wire net_2341;
wire net_661;
wire net_3633;
wire net_3360;
wire net_13537;
wire net_11854;
wire net_7337;
wire net_7036;
wire net_9086;
wire net_3561;
wire net_1543;
wire net_1295;
wire net_10006;
wire net_13692;
wire net_10993;
wire net_9429;
wire net_5661;
wire net_9460;
wire net_2071;
wire net_1923;
wire net_1275;
wire net_210;
wire net_13481;
wire net_11031;
wire net_916;
wire net_13463;
wire net_3395;
wire net_11641;
wire net_940;
wire net_4335;
wire net_851;
wire net_9924;
wire net_4411;
wire net_4857;
wire net_3719;
wire net_10572;
wire net_13247;
wire net_2426;
wire net_6061;
wire net_8311;
wire net_5350;
wire net_7405;
wire net_14329;
wire net_12330;
wire net_12237;
wire net_9627;
wire net_3310;
wire net_671;
wire net_8817;
wire net_8846;
wire net_13631;
wire net_12849;
wire net_5335;
wire net_12431;
wire net_6830;
wire net_6965;
wire net_12438;
wire net_10133;
wire net_8734;
wire net_9485;
wire net_12978;
wire net_9054;
wire net_1454;
wire net_307;
wire net_6949;
wire net_3342;
wire net_13938;
wire net_3547;
wire net_1550;
wire net_3543;
wire net_11470;
wire net_10069;
wire net_9642;
wire net_5104;
wire net_6069;
wire net_233;
wire net_5138;
wire net_3459;
wire net_2656;
wire net_13411;
wire net_1268;
wire net_11127;
wire net_6326;
wire net_3922;
wire net_3212;
wire net_13783;
wire net_3780;
wire net_6530;
wire net_4051;
wire net_1115;
wire net_11465;
wire net_9632;
wire net_1764;
wire net_6641;
wire net_14067;
wire net_961;
wire net_9643;
wire net_3513;
wire net_9968;
wire net_13290;
wire net_4042;
wire net_2106;
wire net_9691;
wire net_3335;
wire net_5377;
wire net_3682;
wire net_6456;
wire net_5175;
wire net_14196;
wire net_11909;
wire net_4894;
wire net_12245;
wire net_5655;
wire net_9424;
wire net_7856;
wire net_9480;
wire net_3327;
wire net_5091;
wire net_13719;
wire net_2667;
wire net_13700;
wire net_3456;
wire net_12818;
wire net_7627;
wire net_13220;
wire net_12453;
wire net_12250;
wire net_5431;
wire net_9907;
wire net_4407;
wire net_13713;
wire net_8443;
wire net_1586;
wire net_14113;
wire net_5354;
wire net_480;
wire net_7662;
wire net_13284;
wire net_216;
wire net_4507;
wire net_10727;
wire net_4986;
wire net_2897;
wire net_5810;
wire net_2881;
wire net_836;
wire net_13817;
wire net_12630;
wire net_2161;
wire net_4602;
wire net_12075;
wire net_12057;
wire net_10671;
wire net_5635;
wire net_9495;
wire net_6568;
wire net_8408;
wire net_6059;
wire net_370;
wire net_8806;
wire net_8379;
wire net_11237;
wire net_13429;
wire net_12520;
wire net_9097;
wire net_6443;
wire net_5881;
wire net_1120;
wire net_2848;
wire net_7126;
wire net_1169;
wire net_973;
wire net_11832;
wire net_13416;
wire net_1139;
wire net_7057;
wire net_6998;
wire net_7013;
wire net_9337;
wire net_7394;
wire net_13677;
wire net_9238;
wire net_7389;
wire net_3902;
wire net_2206;
wire net_11206;
wire net_1392;
wire net_1574;
wire net_9008;
wire net_4842;
wire net_11576;
wire net_6121;
wire net_311;
wire net_2479;
wire net_10132;
wire net_8016;
wire net_154;
wire net_3699;
wire net_11119;
wire net_4469;
wire net_11452;
wire net_13847;
wire net_12527;
wire net_12056;
wire net_9986;
wire net_14075;
wire net_13210;
wire net_2520;
wire net_1478;
wire net_10166;
wire net_2179;
wire net_1696;
wire net_587;
wire net_1262;
wire net_10768;
wire net_9163;
wire net_10704;
wire net_4027;
wire net_14106;
wire net_6676;
wire net_8750;
wire net_4505;
wire net_4213;
wire net_2197;
wire net_10521;
wire net_5399;
wire net_10220;
wire net_4131;
wire net_12089;
wire net_10779;
wire net_9473;
wire net_7396;
wire net_11323;
wire net_2905;
wire net_1907;
wire net_10372;
wire net_200;
wire net_4435;
wire net_8612;
wire net_5220;
wire net_4164;
wire net_6312;
wire net_195;
wire net_5995;
wire net_10200;
wire net_1853;
wire net_9741;
wire net_10247;
wire net_10119;
wire net_10240;
wire net_2170;
wire net_6851;
wire net_10104;
wire net_8980;
wire net_2678;
wire net_11036;
wire net_8346;
wire net_13999;
wire net_9119;
wire net_9042;
wire net_8323;
wire net_7002;
wire net_10256;
wire net_9196;
wire net_8906;
wire net_3761;
wire net_6698;
wire net_13722;
wire net_11267;
wire net_242;
wire net_7722;
wire net_7719;
wire net_7076;
wire net_10381;
wire net_7717;
wire net_6988;
wire x1519;
wire net_9543;
wire net_6281;
wire net_6209;
wire net_2864;
wire net_8938;
wire net_1998;
wire net_11384;
wire net_9341;
wire net_13621;
wire net_11656;
wire net_8336;
wire net_13514;
wire net_2795;
wire net_1311;
wire net_13587;
wire net_5939;
wire net_5540;
wire net_13307;
wire net_11230;
wire net_7068;
wire net_1918;
wire net_12790;
wire net_10207;
wire net_10549;
wire net_5870;
wire net_11911;
wire net_7894;
wire net_5937;
wire net_8208;
wire net_3236;
wire net_5837;
wire net_12314;
wire net_3201;
wire net_11812;
wire net_11169;
wire net_9678;
wire net_3558;
wire net_8147;
wire net_8096;
wire net_5613;
wire net_555;
wire net_9560;
wire net_8966;
wire net_13016;
wire net_7758;
wire net_7163;
wire net_1613;
wire net_8024;
wire net_6897;
wire net_12912;
wire net_11938;
wire net_790;
wire net_5300;
wire net_12359;
wire net_8926;
wire net_11466;
wire net_1417;
wire net_11520;
wire net_13423;
wire x0;
wire net_11063;
wire net_2386;
wire net_2166;
wire net_5803;
wire net_5410;
wire net_3650;
wire net_8359;
wire net_2465;
wire net_5078;
wire net_11588;
wire net_5447;
wire net_12830;
wire net_12043;
wire net_10650;
wire net_8485;
wire net_10388;
wire net_7150;
wire net_13699;
wire net_7462;
wire net_9900;
wire net_6023;
wire net_13862;
wire net_898;
wire net_6136;
wire net_10416;
wire net_6537;
wire net_13023;
wire net_8364;
wire net_7229;
wire net_7045;
wire net_4416;
wire net_5015;
wire net_714;
wire net_8640;
wire net_2999;
wire net_1309;
wire net_9567;
wire net_683;
wire net_1771;
wire net_148;
wire net_1376;
wire net_12136;
wire net_5005;
wire net_4493;
wire net_13555;
wire net_13409;
wire net_8810;
wire net_6885;
wire net_7220;
wire net_6701;
wire net_1980;
wire net_13793;
wire net_9171;
wire net_10362;
wire net_9303;
wire net_7751;
wire net_7449;
wire net_1302;
wire net_244;
wire net_7341;
wire net_5547;
wire net_9361;
wire net_9149;
wire net_8687;
wire net_2395;
wire net_6012;
wire net_7353;
wire net_5616;
wire net_5347;
wire net_12117;
wire net_7113;
wire net_5439;
wire net_4002;
wire net_1989;
wire net_2855;
wire net_1795;
wire net_13310;
wire net_9247;
wire net_8588;
wire net_12186;
wire net_7740;
wire net_2403;
wire net_1539;
wire net_9626;
wire net_14147;
wire net_4261;
wire net_7913;
wire net_10123;
wire net_3490;
wire net_3035;
wire net_7646;
wire net_8550;
wire x522;
wire net_11483;
wire net_1548;
wire net_394;
wire net_810;
wire net_13434;
wire net_3778;
wire net_1189;
wire net_6359;
wire net_12082;
wire net_11131;
wire net_7430;
wire net_409;
wire net_7183;
wire net_7437;
wire net_1469;
wire net_3470;
wire net_11908;
wire net_11626;
wire net_4081;
wire net_13354;
wire net_2436;
wire net_8036;
wire net_11509;
wire net_10754;
wire net_3419;
wire net_10793;
wire net_1254;
wire net_10733;
wire net_14176;
wire net_11417;
wire net_11878;
wire net_621;
wire net_12793;
wire net_10018;
wire net_5153;
wire net_13316;
wire net_10375;
wire net_13171;
wire net_10533;
wire net_11862;
wire net_7240;
wire net_12586;
wire net_7365;
wire net_7729;
wire net_5361;
wire net_8703;
wire net_5598;
wire net_12591;
wire net_11276;
wire net_3985;
wire net_12390;
wire net_9792;
wire net_9383;
wire net_9552;
wire net_10229;
wire net_9689;
wire x1432;
wire net_12663;
wire net_9841;
wire net_4675;
wire net_8378;
wire net_327;
wire net_13032;
wire net_3877;
wire net_999;
wire net_8549;
wire net_353;
wire net_13799;
wire net_8052;
wire net_11730;
wire net_12322;
wire net_10888;
wire net_8838;
wire net_13924;
wire net_9584;
wire net_9752;
wire net_8552;
wire net_5730;
wire net_14209;
wire net_4994;
wire net_3588;
wire net_14140;
wire net_9151;
wire net_8770;
wire net_1480;
wire net_6927;
wire net_12628;
wire net_3046;
wire net_7700;
wire net_6019;
wire net_4952;
wire net_164;
wire net_377;
wire net_8836;
wire net_4702;
wire net_288;
wire net_7632;
wire net_2649;
wire net_3096;
wire net_8947;
wire net_1629;
wire net_1459;
wire net_12252;
wire net_7290;
wire net_5265;
wire net_11650;
wire net_11387;
wire net_3277;
wire net_805;
wire net_12032;
wire net_12093;
wire net_7749;
wire net_6740;
wire net_3741;
wire net_3590;
wire net_13257;
wire net_4470;
wire net_9168;
wire net_2151;
wire net_540;
wire net_8521;
wire net_2688;
wire net_2642;
wire net_14304;
wire net_6650;
wire net_1622;
wire net_891;
wire net_12899;
wire net_9388;
wire net_5224;
wire net_3065;
wire net_13392;
wire net_11664;
wire net_6299;
wire net_5149;
wire net_5821;
wire net_4167;
wire net_7796;
wire net_6746;
wire net_4711;
wire net_10236;
wire net_5868;
wire net_10358;
wire net_7815;
wire net_7453;
wire net_4802;
wire net_12998;
wire net_13420;
wire net_11744;
wire net_618;
wire net_12825;
wire net_2244;
wire net_9075;
wire net_3688;
wire net_5759;
wire net_12001;
wire net_11737;
wire net_7826;
wire net_12399;
wire net_8256;
wire net_783;
wire net_11955;
wire net_6970;
wire net_14255;
wire net_5945;
wire net_13686;
wire net_6148;
wire net_754;
wire net_10785;
wire net_9211;
wire net_11703;
wire net_6305;
wire net_9469;
wire net_2605;
wire net_7193;
wire net_921;
wire net_9875;
wire net_9113;
wire net_550;
wire net_7989;
wire net_11581;
wire net_4957;
wire net_10821;
wire net_12292;
wire net_5238;
wire net_3308;
wire net_12607;
wire net_10274;
wire net_9158;
wire net_5086;
wire net_3991;
wire net_2192;
wire net_1533;
wire net_10912;
wire net_8565;
wire net_7999;
wire net_461;
wire net_7681;
wire net_7778;
wire net_6879;
wire net_12962;
wire net_8524;
wire net_6657;
wire net_9284;
wire net_9138;
wire net_14185;
wire net_11158;
wire net_9884;
wire net_3502;
wire net_14014;
wire net_1512;
wire net_4827;
wire net_654;
wire net_330;
wire net_8047;
wire net_5025;
wire net_1330;
wire net_3506;
wire net_8082;
wire net_4275;
wire net_11011;
wire net_3015;
wire net_1785;
wire net_13507;
wire net_11077;
wire net_9116;
wire net_4771;
wire net_570;
wire net_444;
wire net_525;
wire net_10680;
wire net_3829;
wire net_3646;
wire net_1210;
wire net_1067;
wire net_9516;
wire net_6624;
wire net_5058;
wire net_6870;
wire net_5998;
wire net_9655;
wire net_7820;
wire net_5060;
wire net_12596;
wire net_6200;
wire net_5668;
wire net_10408;
wire net_6259;
wire net_4679;
wire net_985;
wire net_6719;
wire net_12190;
wire net_3933;
wire net_7061;
wire net_424;
wire net_11629;
wire net_6837;
wire net_1729;
wire net_12623;
wire net_3353;
wire net_9325;
wire net_4247;
wire net_4820;
wire net_5719;
wire net_13486;
wire net_10055;
wire net_7577;
wire net_14404;
wire net_3639;
wire net_8065;
wire net_12311;
wire net_12148;
wire net_11992;
wire net_3086;
wire net_4585;
wire net_11110;
wire net_9409;
wire net_2058;
wire net_12206;
wire net_9404;
wire net_3045;
wire net_1178;
wire net_9722;
wire net_5573;
wire net_4875;
wire net_7098;
wire net_2018;
wire net_13100;
wire net_11731;
wire net_3825;
wire net_11142;
wire net_6218;
wire net_12380;
wire net_340;
wire net_6039;
wire net_2510;
wire net_9952;
wire net_2634;
wire net_434;
wire net_7881;
wire net_3808;
wire net_12941;
wire net_6915;
wire net_8434;
wire net_7024;
wire net_6936;
wire net_6243;
wire net_14200;
wire net_7882;
wire net_1797;
wire net_6415;
wire net_9443;
wire net_14393;
wire net_11086;
wire net_9201;
wire net_4906;
wire net_4524;
wire net_6302;
wire net_8916;
wire net_339;
wire net_2279;
wire net_7686;
wire net_14048;
wire net_3447;
wire net_13105;
wire net_8401;
wire net_6174;
wire net_3468;
wire net_10443;
wire net_11775;
wire net_12753;
wire net_2710;
wire net_9267;
wire net_2660;
wire net_8624;
wire net_10083;
wire net_13893;
wire net_10826;
wire net_8087;
wire net_5389;
wire net_8497;
wire net_3671;
wire net_8236;
wire net_8651;
wire net_10295;
wire net_3691;
wire net_7801;
wire net_3217;
wire net_6362;
wire net_4387;
wire net_1291;
wire net_1865;
wire net_13896;
wire net_678;
wire net_6076;
wire net_5168;
wire net_5329;
wire net_11631;
wire net_8979;
wire net_10985;
wire net_928;
wire x1534;
wire net_10490;
wire net_8460;
wire net_5459;
wire net_13363;
wire net_2578;
wire net_208;
wire net_9225;
wire net_7878;
wire net_8658;
wire net_8215;
wire net_10462;
wire net_2744;
wire net_2377;
wire net_1433;
wire net_415;
wire net_116;
wire net_3251;
wire net_2786;
wire net_11672;
wire net_347;
wire net_13745;
wire net_13526;
wire net_11059;
wire net_3794;
wire net_12664;
wire net_8606;
wire net_7306;
wire net_5440;
wire net_9425;
wire net_1335;
wire net_5928;
wire net_2574;
wire net_14235;
wire net_3531;
wire net_12210;
wire net_5477;
wire net_3747;
wire net_2212;
wire net_5453;
wire net_11535;
wire net_7730;
wire net_12212;
wire net_5732;
wire net_8593;
wire net_3571;
wire net_4642;
wire x940;
wire net_610;
wire net_1844;
wire net_8130;
wire net_11512;
wire net_7870;
wire net_389;
wire net_902;
wire net_13981;
wire net_2344;
wire net_11287;
wire net_10588;
wire net_1323;
wire net_14130;
wire net_1506;
wire net_10470;
wire net_13386;
wire net_13237;
wire net_6496;
wire net_13193;
wire net_736;
wire net_8771;
wire net_539;
wire net_13068;
wire net_692;
wire net_5462;
wire net_5282;
wire net_4568;
wire net_6498;
wire net_8372;
wire net_10807;
wire net_6262;
wire net_4377;
wire net_14261;
wire net_7704;
wire net_13125;
wire net_10905;
wire net_10311;
wire net_12517;
wire net_1400;
wire net_14092;
wire net_885;
wire net_10034;
wire net_9202;
wire net_7249;
wire net_11698;
wire net_14320;
wire net_9918;
wire net_5717;
wire net_10770;
wire net_869;
wire net_12144;
wire net_6822;
wire net_3714;
wire net_8308;
wire net_11280;
wire net_4077;
wire net_11607;
wire net_2441;
wire net_6594;
wire net_3517;
wire net_496;
wire net_761;
wire net_11396;
wire net_6799;
wire net_5828;
wire net_4749;
wire net_1554;
wire net_7101;
wire net_8775;
wire net_13774;
wire net_12092;
wire net_2459;
wire net_10638;
wire net_4370;
wire net_10394;
wire net_4979;
wire net_12578;
wire net_2249;
wire net_5422;
wire net_6629;
wire net_5686;
wire net_6704;
wire net_739;
wire net_12395;
wire net_8760;
wire net_6508;
wire net_2548;
wire net_2075;
wire net_826;
wire net_1738;
wire net_10384;
wire net_10504;
wire net_3359;
wire net_5848;
wire net_10085;
wire net_12296;
wire net_11644;
wire net_9069;
wire net_6716;
wire net_7548;
wire net_2624;
wire net_12889;
wire net_11761;
wire net_343;
wire net_6165;
wire net_4795;
wire net_511;
wire net_9263;
wire net_12759;
wire net_7313;
wire net_3967;
wire net_9672;
wire net_8456;
wire net_5236;
wire net_4424;
wire net_7541;
wire net_9615;
wire net_2654;
wire net_7451;
wire net_2487;
wire net_11791;
wire net_7803;
wire net_2911;
wire net_1819;
wire net_8258;
wire net_12821;
wire net_8227;
wire net_12763;
wire net_13132;
wire net_2975;
wire net_4625;
wire net_7236;
wire net_5257;
wire net_8220;
wire net_2779;
wire net_14187;
wire net_11552;
wire net_6392;
wire net_13181;
wire net_11379;
wire net_9031;
wire net_9346;
wire net_13661;
wire net_11352;
wire net_8169;
wire x195;
wire net_1490;
wire net_11083;
wire net_9274;
wire net_4282;
wire net_989;
wire net_11806;
wire net_12774;
wire net_8446;
wire net_14342;
wire net_5742;
wire net_458;
wire net_4356;
wire net_11748;
wire net_685;
wire net_8466;
wire net_7442;
wire net_8322;
wire net_10998;
wire net_9030;
wire net_10957;
wire net_12349;
wire net_14183;
wire net_13333;
wire net_11843;
wire net_4052;
wire net_8513;
wire net_4616;
wire net_8681;
wire net_13096;
wire net_11408;
wire net_4786;
wire net_8616;
wire net_7872;
wire net_5893;
wire net_10542;
wire net_13469;
wire net_10891;
wire net_10652;
wire net_7160;
wire net_12876;
wire net_4686;
wire net_3410;
wire net_2111;
wire net_1946;
wire net_2733;
wire net_8162;
wire net_5525;
wire net_12496;
wire net_14280;
wire net_6764;
wire net_13252;
wire net_5610;
wire net_14278;
wire net_6769;
wire net_3612;
wire net_11634;
wire net_1605;
wire net_12795;
wire net_13045;
wire net_2535;
wire net_13165;
wire net_3191;
wire net_5118;
wire net_14396;
wire net_13822;
wire net_747;
wire net_10355;
wire net_2305;
wire net_1653;
wire net_12865;
wire net_14125;
wire net_5842;
wire net_12125;
wire net_9817;
wire net_7377;
wire net_2983;
wire net_12916;
wire net_10024;
wire net_2258;
wire net_198;
wire net_1647;
wire net_12460;
wire net_11168;
wire net_12510;
wire net_14327;
wire net_10058;
wire net_7509;
wire net_4756;
wire net_13280;
wire net_6500;
wire net_5196;
wire net_2367;
wire net_4573;
wire net_4127;
wire net_2892;
wire net_13263;
wire net_2810;
wire net_13546;
wire net_13077;
wire net_1053;
wire net_4444;
wire net_11292;
wire net_1004;
wire net_848;
wire net_4921;
wire net_11716;
wire net_11359;
wire net_9550;
wire net_12022;
wire net_1080;
wire net_10641;
wire net_3232;
wire net_1890;
wire net_13356;
wire net_13648;
wire net_4498;
wire net_11293;
wire net_3228;
wire net_2282;
wire net_10029;
wire net_4501;
wire net_2357;
wire net_13319;
wire net_12449;
wire net_11114;
wire net_1546;
wire net_11772;
wire net_11367;
wire net_8542;
wire net_5492;
wire net_12383;
wire net_6042;
wire net_13654;
wire net_11372;
wire net_10199;
wire net_1046;
wire net_6536;
wire net_11502;
wire net_7417;
wire net_4363;
wire x1424;
wire net_606;
wire net_10332;
wire net_4960;
wire net_3906;
wire net_623;
wire net_12503;
wire net_663;
wire net_1213;
wire net_1891;
wire net_2265;
wire net_8118;
wire net_10163;
wire net_5180;
wire net_3998;
wire net_579;
wire net_9490;
wire net_8597;
wire net_5795;
wire net_12812;
wire net_769;
wire net_1780;
wire net_2062;
wire net_13668;
wire net_13666;
wire net_9828;
wire net_10844;
wire net_6418;
wire net_1025;
wire net_3758;
wire net_7296;
wire net_4834;
wire net_9317;
wire net_8061;
wire net_4067;
wire net_4717;
wire net_13157;
wire net_10403;
wire net_7502;
wire net_1518;
wire net_4618;
wire net_1089;
wire net_12169;
wire net_1194;
wire net_1437;
wire net_11998;
wire net_5517;
wire net_6770;
wire net_11923;
wire net_7587;
wire net_1664;
wire net_13651;
wire net_4528;
wire net_6233;
wire net_5625;
wire net_10326;
wire net_705;
wire net_4141;
wire net_2948;
wire net_10523;
wire net_14094;
wire net_12535;
wire net_10669;
wire net_1036;
wire net_6052;
wire net_5608;
wire net_11966;
wire net_7497;
wire net_5146;
wire net_4537;
wire net_8701;
wire net_1196;
wire net_6331;
wire net_3973;
wire net_5326;
wire net_12921;
wire net_4394;
wire net_9077;
wire net_6762;
wire net_5531;
wire net_5953;
wire net_12442;
wire net_11047;
wire net_12702;
wire net_9433;
wire net_6085;
wire net_10816;
wire net_6598;
wire net_14124;
wire net_13248;
wire net_5701;
wire net_11786;
wire net_3626;
wire net_12095;
wire net_5779;
wire net_3136;
wire net_12553;
wire net_6417;
wire net_4726;
wire net_4090;
wire net_14377;
wire net_13086;
wire net_9588;
wire net_6149;
wire net_10809;
wire net_9178;
wire net_5344;
wire net_3834;
wire net_7492;
wire net_12468;
wire net_5364;
wire x217;
wire net_10300;
wire net_13471;
wire net_8743;
wire net_3152;
wire net_6388;
wire net_14311;
wire net_13478;
wire net_3648;
wire net_740;
wire net_1722;
wire net_4072;
wire net_6395;
wire net_2008;
wire net_11633;
wire net_11090;
wire net_5825;
wire net_3183;
wire net_2808;
wire net_3908;
wire net_8265;
wire net_4837;
wire net_730;
wire net_9055;
wire net_4150;
wire x96;
wire net_14008;
wire net_8049;
wire net_7094;
wire net_5405;
wire net_11931;
wire net_6575;
wire net_2105;
wire net_13918;
wire net_7226;
wire net_6432;
wire net_4707;
wire net_1127;
wire net_6381;
wire net_9458;
wire net_11243;
wire net_12771;
wire net_6420;
wire net_957;
wire net_1287;
wire net_13831;
wire net_10625;
wire net_7465;
wire net_14040;
wire net_9297;
wire net_2726;
wire net_4143;
wire net_12900;
wire net_8679;
wire net_7285;
wire net_1340;
wire net_5140;
wire net_7277;
wire net_3123;
wire net_2955;
wire net_7165;
wire net_9599;
wire net_12363;
wire net_771;
wire net_2844;
wire net_2301;
wire net_12415;
wire net_2978;
wire net_9977;
wire net_5538;
wire net_5185;
wire net_13139;
wire net_9941;
wire net_6804;
wire net_4852;
wire net_10341;
wire net_14361;
wire net_3950;
wire net_10435;
wire net_4437;
wire net_4028;
wire net_2860;
wire net_432;
wire net_6025;
wire net_4927;
wire net_1062;
wire net_6329;
wire net_14395;
wire net_10627;
wire net_4936;
wire net_3293;
wire net_1142;
wire net_4120;
wire net_9246;
wire net_7733;
wire net_3159;
wire net_5644;
wire net_6050;
wire net_2240;
wire net_2416;
wire net_13214;
wire net_12882;
wire net_6404;
wire net_5188;
wire net_4590;
wire net_8727;
wire x889;
wire net_14354;
wire net_6185;
wire net_6116;
wire net_9713;
wire net_1411;
wire net_12549;
wire net_505;
wire net_5383;
wire net_4088;
wire net_10471;
wire net_3723;
wire net_10540;
wire net_7487;
wire net_13520;
wire net_10493;
wire net_10426;
wire net_7152;
wire net_6527;
wire net_4013;
wire net_992;
wire net_11517;
wire net_7485;
wire net_9781;
wire net_6727;
wire net_782;
wire net_2144;
wire net_2236;
wire net_10527;
wire net_13576;
wire net_11106;
wire net_11057;
wire net_3443;
wire net_6291;
wire net_4186;
wire net_13328;
wire net_4738;
wire net_3314;
wire net_7422;
wire net_3945;
wire net_2971;
wire net_5776;
wire net_8824;
wire net_13322;
wire net_11529;
wire net_10339;
wire net_8072;
wire net_8244;
wire net_2836;
wire net_1505;
wire net_10615;
wire net_5689;
wire net_7429;
wire net_1805;
wire net_4667;
wire net_13836;
wire net_11536;
wire net_8279;
wire net_3952;
wire net_3669;
wire net_13448;
wire net_10660;
wire net_1861;
wire net_3635;
wire net_9999;
wire net_4388;
wire net_11852;
wire net_13559;
wire net_5672;
wire net_221;
wire net_1594;
wire net_7120;
wire net_1110;
wire net_442;
wire net_542;
wire net_14218;
wire net_13026;
wire net_13789;
wire net_12483;
wire net_6487;
wire net_7202;
wire net_4562;
wire net_9437;
wire net_3087;
wire net_2376;
wire net_6562;
wire net_1520;
wire net_6713;
wire net_13900;
wire net_1821;
wire net_8579;
wire net_9638;
wire net_11675;
wire net_7480;
wire net_3865;
wire net_1588;
wire net_9029;
wire net_4037;
wire net_8005;
wire net_3937;
wire net_1495;
wire net_2992;
wire net_12974;
wire net_3664;
wire net_5124;
wire net_3233;
wire net_9731;
wire net_3522;
wire net_7178;
wire net_10937;
wire net_668;
wire net_7601;
wire net_11814;
wire net_9649;
wire net_3079;
wire net_1584;
wire net_14203;
wire net_13539;
wire net_12612;
wire net_2330;
wire net_8040;
wire net_5814;
wire net_7890;
wire net_12707;
wire net_3397;
wire net_1070;
wire net_9777;
wire net_8878;
wire net_1225;
wire net_812;
wire net_5898;
wire net_6785;
wire net_7814;
wire net_4391;
wire net_11473;
wire net_13805;
wire net_9045;
wire net_6314;
wire net_12659;
wire net_6875;
wire net_6972;
wire net_2857;
wire net_1107;
wire net_8674;
wire net_2767;
wire net_9594;
wire net_6120;
wire net_11491;
wire net_11053;
wire net_3384;
wire net_12652;
wire net_6604;
wire net_1203;
wire net_13347;
wire net_825;
wire net_309;
wire net_1366;
wire net_13054;
wire net_2615;
wire net_9011;
wire net_12402;
wire net_12176;
wire net_10867;
wire net_10715;
wire net_14268;
wire net_5321;
wire net_11434;
wire net_9290;
wire net_7367;
wire net_12789;
wire net_8158;
wire net_1151;
wire net_5240;
wire net_5318;
wire net_9993;
wire net_11138;
wire net_8291;
wire net_5884;
wire net_3213;
wire net_2818;
wire net_863;
wire net_7131;
wire net_7690;
wire net_6468;
wire net_3164;
wire net_4173;
wire net_580;
wire net_14058;
wire net_13150;
wire net_9805;
wire net_2136;
wire net_904;
wire net_2339;
wire net_8884;
wire net_7699;
wire net_12850;
wire net_14226;
wire net_4157;
wire net_13552;
wire net_1879;
wire net_6777;
wire net_12286;
wire net_6663;
wire net_12122;
wire net_13224;
wire net_8202;
wire net_6633;
wire net_8126;
wire net_4941;
wire net_4221;
wire net_6092;
wire net_6732;
wire net_6559;
wire net_12524;
wire net_11360;
wire net_9183;
wire net_4845;
wire net_1160;
wire net_12683;
wire net_159;
wire net_11147;
wire net_9379;
wire net_3268;
wire net_11022;
wire net_5604;
wire net_11612;
wire net_5863;
wire net_8351;
wire net_11615;
wire net_9523;
wire net_10181;
wire net_4887;
wire net_9354;
wire net_13116;
wire net_2875;
wire net_763;
wire net_13704;
wire net_12952;
wire net_14088;
wire net_10213;
wire net_7762;
wire net_5639;
wire net_1740;
wire net_324;
wire net_6848;
wire net_11724;
wire net_10284;
wire net_10074;
wire net_13397;
wire net_9455;
wire net_5480;
wire net_10309;
wire net_7257;
wire net_872;
wire net_13047;
wire net_9706;
wire net_14248;
wire net_14103;
wire net_9125;
wire net_12647;
wire net_10964;
wire net_10502;
wire net_5046;
wire net_3066;
wire net_8251;
wire net_6270;
wire net_3880;
wire net_6275;
wire net_5581;
wire net_4333;
wire net_4181;
wire net_11285;
wire net_376;
wire net_5558;
wire x131;
wire net_7575;
wire net_2133;
wire net_13643;
wire net_4817;
wire net_4880;
wire net_13374;
wire net_2515;
wire net_1812;
wire net_8174;
wire net_3173;
wire net_12584;
wire net_8038;
wire net_4825;
wire net_10850;
wire net_3738;
wire net_8696;
wire net_7994;
wire net_4138;
wire net_5298;
wire net_5119;
wire net_3203;
wire net_422;
wire net_4290;
wire net_1345;
wire net_12811;
wire net_1450;
wire net_561;
wire net_12694;
wire net_11881;
wire net_4899;
wire net_12670;
wire net_7515;
wire net_2659;
wire net_2589;
wire net_12739;
wire net_591;
wire net_1700;
wire net_12985;
wire net_5955;
wire net_8501;
wire net_4299;
wire net_2290;
wire net_12741;
wire net_10188;
wire net_7557;
wire net_2851;
wire net_178;
wire net_11751;
wire net_8427;
wire net_9074;
wire net_2843;
wire net_14081;
wire net_14019;
wire net_6780;
wire net_7961;
wire net_10191;
wire net_3772;
wire net_7901;
wire net_3807;
wire net_4868;
wire net_10480;
wire net_2698;
wire net_809;
wire net_13995;
wire net_8393;
wire net_6552;
wire net_8453;
wire net_3450;
wire net_635;
wire net_4279;
wire net_266;
wire net_1235;
wire net_14412;
wire net_2691;
wire net_3528;
wire net_8559;
wire net_8610;
wire net_12600;
wire net_8956;
wire net_350;
wire net_6622;
wire net_4270;
wire net_8332;
wire net_6007;
wire net_13205;
wire net_13178;
wire net_10176;
wire net_7606;
wire net_6549;
wire net_13275;
wire net_6542;
wire net_13091;
wire net_3460;
wire net_12859;
wire net_3117;
wire net_14245;
wire net_11816;
wire net_3482;
wire net_6648;
wire net_3198;
wire net_8366;
wire net_5720;
wire net_1626;
wire net_2822;
wire net_7317;
wire net_8413;
wire net_1258;
wire net_7375;
wire net_12041;
wire net_3369;
wire net_9866;
wire net_9020;
wire net_1101;
wire net_994;
wire net_12828;
wire net_12268;
wire net_10231;
wire net_318;
wire net_6685;
wire net_3927;
wire net_11837;
wire net_10859;
wire net_1971;
wire net_8931;
wire net_4166;
wire net_2409;
wire net_4608;
wire net_3192;
wire net_1900;
wire net_1779;
wire net_2647;
wire net_5218;
wire net_3340;
wire net_8492;
wire net_4545;
wire net_3844;
wire net_1849;
wire net_7972;
wire net_10045;
wire net_228;
wire net_5486;
wire net_11886;
wire net_4737;
wire net_2640;
wire net_13011;
wire net_966;
wire net_7083;
wire net_13516;
wire net_4698;
wire net_3372;
wire net_11122;
wire net_6049;
wire net_2201;
wire net_1108;
wire net_2827;
wire net_2025;
wire net_8583;
wire net_7905;
wire net_2936;
wire net_5643;
wire net_9756;
wire net_9936;
wire net_1878;
wire net_13736;
wire net_5728;
wire net_13070;
wire net_9255;
wire net_11446;
wire net_8013;
wire net_3890;
wire net_5975;
wire net_133;
wire net_12425;
wire net_10702;
wire net_10366;
wire net_7528;
wire net_14297;
wire net_4025;
wire net_11414;
wire net_12444;
wire net_11265;
wire net_10920;
wire net_9194;
wire net_7078;
wire net_12529;
wire net_10579;
wire net_7008;
wire net_11957;
wire net_7997;
wire net_4522;
wire net_3882;
wire net_557;
wire net_3043;
wire net_11925;
wire net_8908;
wire net_7860;
wire net_8689;
wire net_6611;
wire net_3652;
wire net_6829;
wire net_2669;
wire net_13891;
wire net_11386;
wire net_4083;
wire net_12316;
wire net_1991;
wire net_1611;
wire net_1173;
wire net_14046;
wire net_1431;
wire net_1754;
wire net_2328;
wire net_7715;
wire net_11401;
wire net_8080;
wire net_1714;
wire net_5571;
wire net_13014;
wire net_11970;
wire net_10205;
wire net_5805;
wire net_8868;
wire net_240;
wire net_12792;
wire net_7254;
wire net_13623;
wire net_7684;
wire net_295;
wire net_8411;
wire net_12991;
wire net_10743;
wire net_13605;
wire net_13565;
wire net_13425;
wire net_9604;
wire net_9241;
wire net_6887;
wire net_9838;
wire net_4462;
wire net_5935;
wire net_11038;
wire net_13490;
wire net_1394;
wire net_7753;
wire net_2963;
wire net_5546;
wire net_5412;
wire net_12115;
wire net_7720;
wire net_6134;
wire net_9395;
wire net_1281;
wire net_2463;
wire net_11239;
wire net_9291;
wire net_12619;
wire net_6691;
wire net_8210;
wire net_12967;
wire net_278;
wire net_6864;
wire net_11258;
wire net_8995;
wire net_8367;
wire net_4058;
wire net_9063;
wire net_8432;
wire net_4874;
wire net_3509;
wire net_1162;
wire net_10090;
wire net_13856;
wire net_13309;
wire net_2443;
wire net_10736;
wire net_2472;
wire net_1307;
wire net_13589;
wire net_4514;
wire net_2790;
wire net_2742;
wire net_13120;
wire net_10738;
wire net_5007;
wire net_10318;
wire net_6940;
wire net_13795;
wire net_10434;
wire net_5591;
wire net_4810;
wire net_11902;
wire net_8360;
wire net_10269;
wire net_6521;
wire net_10561;
wire net_4418;
wire net_3320;
wire net_5221;
wire net_3657;
wire net_5550;
wire net_5385;
wire net_14145;
wire net_6099;
wire net_1353;
wire net_9786;
wire net_11652;
wire net_12679;
wire net_7630;
wire net_5303;
wire net_3581;
wire net_13854;
wire net_13712;
wire net_4049;
wire net_3776;
wire net_1300;
wire net_14322;
wire net_1252;
wire net_12131;
wire x30;
wire net_9173;
wire net_7739;
wire net_9095;
wire net_7784;
wire net_13432;
wire net_14026;
wire net_10941;
wire net_547;
wire net_1098;
wire net_10731;
wire net_507;
wire net_10097;
wire net_10049;
wire net_8981;
wire net_1902;
wire net_6683;
wire net_238;
wire net_3074;
wire net_7111;
wire net_8973;
wire net_5475;
wire net_11354;
wire net_7055;
wire net_7896;
wire net_2438;
wire net_2600;
wire net_1911;
wire net_6906;
wire net_5734;
wire net_3563;
wire net_12224;
wire net_8726;
wire net_6585;
wire net_649;
wire net_9565;
wire net_13597;
wire net_11936;
wire net_4491;
wire net_11543;
wire net_1374;
wire net_13887;
wire net_8282;
wire net_7538;
wire net_4843;
wire net_8959;
wire net_1962;
wire net_291;
wire net_9502;
wire net_7351;
wire net_1964;
wire net_2494;
wire net_857;
wire net_867;
wire net_5964;
wire net_11217;
wire net_6819;
wire net_396;
wire net_12274;
wire net_3700;
wire net_13349;
wire net_10602;
wire x806;
wire net_8851;
wire net_10535;
wire net_530;
wire net_9140;
wire net_1541;
wire net_11839;
wire net_10529;
wire net_14216;
wire net_9748;
wire net_5177;
wire net_271;
wire net_3329;
wire net_10067;
wire net_10004;
wire net_6111;
wire net_673;
wire net_7022;
wire net_4268;
wire net_12247;
wire net_12208;
wire net_7029;
wire net_3611;
wire net_2064;
wire net_9966;
wire net_6256;
wire net_2797;
wire net_3846;
wire net_12261;
wire net_5333;
wire net_1925;
wire net_9790;
wire net_3549;
wire net_1445;
wire net_10227;
wire net_8581;
wire net_1909;
wire net_6729;
wire net_13807;
wire net_9922;
wire net_10126;
wire net_7639;
wire net_1410;
wire net_11454;
wire net_11583;
wire net_365;
wire net_13412;
wire net_5379;
wire net_13340;
wire net_3913;
wire net_11643;
wire net_9988;
wire net_3344;
wire net_12060;
wire net_8374;
wire net_3787;
wire net_10729;
wire net_4413;
wire net_1810;
wire net_10776;
wire net_1118;
wire net_13849;
wire net_8719;
wire net_4313;
wire net_11000;
wire net_12235;
wire net_6858;
wire net_372;
wire net_9882;
wire net_8313;
wire net_7086;
wire net_2990;
wire x977;
wire x1822;
wire net_9339;
wire net_6324;
wire net_7128;
wire net_7915;
wire net_13723;
wire net_11749;
wire net_13730;
wire net_4892;
wire net_803;
wire net_10884;
wire net_3595;
wire net_13787;
wire net_10383;
wire net_8923;
wire net_2788;
wire net_10142;
wire net_6899;
wire net_14111;
wire net_7764;
wire net_6375;
wire net_1476;
wire net_3489;
wire net_1293;
wire net_11098;
wire net_11184;
wire net_13581;
wire net_2883;
wire net_8665;
wire net_563;
wire net_7854;
wire net_13979;
wire net_1147;
wire net_11742;
wire net_13388;
wire net_2681;
wire net_8815;
wire net_13452;
wire net_12159;
wire net_9629;
wire net_2158;
wire net_5136;
wire net_4855;
wire net_4366;
wire net_10234;
wire net_13936;
wire net_10175;
wire net_12254;
wire net_5009;
wire net_1266;
wire net_3684;
wire net_1452;
wire net_8418;
wire net_2773;
wire net_2428;
wire net_909;
wire net_4529;
wire net_10695;
wire net_4898;
wire net_152;
wire net_8652;
wire net_11575;
wire net_10814;
wire net_3105;
wire net_2895;
wire net_13299;
wire net_2138;
wire net_13418;
wire net_8238;
wire net_258;
wire net_12957;
wire net_11192;
wire net_2477;
wire net_10761;
wire net_12935;
wire net_12054;
wire net_9927;
wire net_5653;
wire net_13983;
wire net_13819;
wire net_7664;
wire net_5083;
wire net_2446;
wire net_7171;
wire net_11999;
wire net_4188;
wire net_7605;
wire net_585;
wire net_7611;
wire net_7809;
wire net_6146;
wire net_4040;
wire net_11913;
wire net_11347;
wire net_12766;
wire net_5433;
wire net_12061;
wire net_10593;
wire net_3759;
wire net_3511;
wire net_12839;
wire net_374;
wire net_14069;
wire net_10293;
wire net_8755;
wire net_1987;
wire net_12816;
wire net_12632;
wire net_788;
wire net_12910;
wire net_9090;
wire net_214;
wire net_7011;
wire net_8113;
wire net_3602;
wire net_249;
wire net_13155;
wire net_13028;
wire net_9963;
wire net_8144;
wire net_3578;
wire net_12455;
wire net_5283;
wire net_13903;
wire net_8804;
wire net_9013;
wire net_8871;
wire net_6310;
wire net_6196;
wire net_13488;
wire net_10766;
wire net_4009;
wire net_7648;
wire net_5097;
wire net_13880;
wire net_8508;
wire net_7329;
wire net_5993;
wire net_4259;
wire net_2565;
wire net_8018;
wire net_2632;
wire net_2547;
wire net_8634;
wire net_5076;
wire net_13229;
wire net_9084;
wire net_6783;
wire net_5908;
wire net_2118;
wire net_463;
wire net_2295;
wire net_5831;
wire net_5628;
wire net_9487;
wire net_1817;
wire net_197;
wire net_2560;
wire net_11009;
wire net_9348;
wire net_1381;
wire net_9331;
wire net_6445;
wire net_5017;
wire net_3709;
wire net_202;
wire net_13596;
wire net_3312;
wire net_13085;
wire net_7325;
wire net_1756;
wire net_12803;
wire net_7588;
wire net_11468;
wire net_2208;
wire net_6475;
wire net_5352;
wire net_2595;
wire net_1383;
wire net_7302;
wire net_2751;
wire net_918;
wire net_11204;
wire net_7727;
wire net_9663;
wire net_9165;
wire net_5397;
wire net_9204;
wire net_4446;
wire net_14160;
wire net_10484;
wire net_6269;
wire net_6176;
wire net_5901;
wire net_14170;
wire net_13672;
wire net_13610;
wire net_11116;
wire net_13497;
wire net_1683;
wire net_12515;
wire net_978;
wire net_9356;
wire net_1313;
wire net_10780;
wire net_1129;
wire net_11345;
wire net_7618;
wire net_3331;
wire net_1056;
wire net_4908;
wire net_11994;
wire net_13286;
wire net_10896;
wire net_5712;
wire net_10877;
wire net_8383;
wire net_4781;
wire net_2044;
wire net_9954;
wire net_7402;
wire net_6360;
wire net_2181;
wire net_8626;
wire net_6913;
wire net_1789;
wire net_14035;
wire net_13142;
wire net_13940;
wire net_8406;
wire net_7379;
wire net_4530;
wire net_838;
wire net_3219;
wire net_10441;
wire net_6123;
wire net_7520;
wire net_14316;
wire net_11151;
wire net_14202;
wire net_4587;
wire net_11750;
wire net_5872;
wire net_7107;
wire net_4980;
wire net_2576;
wire net_11270;
wire net_3827;
wire net_2352;
wire net_1038;
wire net_8405;
wire net_12072;
wire net_6931;
wire net_4241;
wire net_9920;
wire net_8168;
wire net_5308;
wire net_5710;
wire net_5369;
wire net_3763;
wire net_3515;
wire net_12747;
wire net_5033;
wire net_8085;
wire net_6333;
wire net_9720;
wire net_11338;
wire net_9223;
wire net_7697;
wire net_3398;
wire net_2277;
wire net_342;
wire net_13400;
wire net_6078;
wire net_975;
wire net_5421;
wire net_612;
wire net_892;
wire net_8098;
wire net_12871;
wire net_4650;
wire net_4198;
wire net_13061;
wire net_10423;
wire net_5434;
wire net_11144;
wire net_6160;
wire net_10848;
wire net_5874;
wire net_2006;
wire net_13570;
wire net_12639;
wire net_8344;
wire net_10060;
wire net_6511;
wire net_1331;
wire net_1537;
wire net_13051;
wire net_11105;
wire net_12307;
wire net_13399;
wire net_5826;
wire net_4074;
wire net_4000;
wire net_13912;
wire net_2214;
wire net_3338;
wire net_5987;
wire net_8604;
wire net_2728;
wire net_13238;
wire net_9929;
wire net_4636;
wire net_417;
wire net_122;
wire net_6264;
wire net_13619;
wire net_12847;
wire net_11514;
wire net_10634;
wire net_10026;
wire net_5387;
wire x1322;
wire net_8217;
wire net_9262;
wire net_7467;
wire net_4092;
wire x447;
wire net_10758;
wire net_12300;
wire net_8595;
wire net_8287;
wire net_3337;
wire net_2662;
wire net_11760;
wire net_10751;
wire net_3752;
wire net_4486;
wire net_9427;
wire net_9131;
wire net_482;
wire net_5144;
wire net_10805;
wire net_3258;
wire net_10942;
wire net_10983;
wire net_7262;
wire net_149;
wire net_387;
wire net_7790;
wire net_3275;
wire net_7447;
wire net_6297;
wire net_13107;
wire net_13127;
wire net_10828;
wire net_5291;
wire net_5160;
wire net_1893;
wire net_14137;
wire net_6494;
wire net_1932;
wire net_9639;
wire net_8896;
wire net_11620;
wire net_8268;
wire net_3836;
wire net_577;
wire net_13245;
wire net_3401;
wire net_10313;
wire net_2550;
wire net_797;
wire net_7747;
wire net_3545;
wire net_1957;
wire net_1799;
wire net_10150;
wire net_11224;
wire net_10102;
wire net_13743;
wire net_13231;
wire net_9368;
wire net_11859;
wire net_12909;
wire net_9218;
wire net_7581;
wire net_2572;
wire net_2414;
wire net_337;
wire net_10581;
wire net_1846;
wire net_13312;
wire net_4476;
wire net_690;
wire net_13381;
wire net_5667;
wire net_11222;
wire net_7933;
wire net_6820;
wire net_9662;
wire net_3743;
wire net_7888;
wire net_12475;
wire net_523;
wire net_11066;
wire net_13984;
wire net_11070;
wire net_4254;
wire net_13760;
wire net_6718;
wire net_3815;
wire net_3555;
wire net_7144;
wire net_5739;
wire net_2371;
wire net_3375;
wire net_6744;
wire net_9620;
wire net_6794;
wire net_14077;
wire net_4926;
wire net_3467;
wire net_9617;
wire net_13368;
wire net_8972;
wire net_11014;
wire net_9760;
wire net_8396;
wire net_12546;
wire net_9640;
wire net_7843;
wire net_7392;
wire net_4467;
wire net_3982;
wire net_1388;
wire net_12129;
wire net_5028;
wire net_4709;
wire net_14409;
wire net_4721;
wire net_5756;
wire net_9858;
wire net_3391;
wire net_2730;
wire net_4426;
wire net_1631;
wire net_1337;
wire net_6835;
wire net_5786;
wire net_14254;
wire net_13553;
wire net_1182;
wire net_4655;
wire net_1624;
wire net_7231;
wire net_6618;
wire net_12332;
wire net_13656;
wire net_1638;
wire net_1950;
wire net_9052;
wire net_7455;
wire net_3875;
wire net_12146;
wire net_9319;
wire net_9280;
wire net_7039;
wire net_10135;
wire net_2421;
wire net_5684;
wire net_5268;
wire net_11389;
wire net_4901;
wire net_4804;
wire net_880;
wire net_1402;
wire net_6335;
wire net_2153;
wire net_1939;
wire net_9582;
wire net_4100;
wire net_8781;
wire net_8474;
wire net_3098;
wire net_7242;
wire net_14190;
wire net_8535;
wire net_6288;
wire net_4673;
wire net_5762;
wire net_9061;
wire net_5151;
wire net_13922;
wire net_10249;
wire net_11876;
wire net_7828;
wire net_2901;
wire net_162;
wire net_8301;
wire net_13255;
wire net_4950;
wire net_7776;
wire net_4944;
wire net_653;
wire net_14301;
wire net_13160;
wire net_5066;
wire net_13919;
wire net_11735;
wire net_12661;
wire net_12030;
wire net_4847;
wire net_3052;
wire net_3145;
wire net_10906;
wire net_6652;
wire net_9558;
wire net_13694;
wire net_3694;
wire net_11554;
wire net_7295;
wire net_10262;
wire net_11592;
wire net_6368;
wire net_3855;
wire net_236;
wire net_12324;
wire net_487;
wire net_9286;
wire net_552;
wire net_10823;
wire net_8861;
wire net_8206;
wire net_7992;
wire net_1787;
wire net_3551;
wire net_6654;
wire net_7440;
wire net_13390;
wire net_5056;
wire net_9518;
wire net_756;
wire net_7067;
wire net_7735;
wire net_13636;
wire net_4765;
wire net_14234;
wire x1398;
wire net_8329;
wire net_12230;
wire net_10101;
wire net_7798;
wire net_14402;
wire net_11301;
wire net_5031;
wire net_3416;
wire net_7198;
wire net_5166;
wire net_11845;
wire net_4886;
wire net_9878;
wire net_3537;
wire net_10914;
wire net_14070;
wire net_12039;
wire net_8522;
wire net_6659;
wire net_12897;
wire net_12192;
wire net_6877;
wire net_711;
wire net_2225;
wire net_7659;
wire net_4741;
wire net_11687;
wire net_8618;
wire net_4700;
wire net_846;
wire net_10469;
wire net_9402;
wire net_12852;
wire net_3017;
wire x1494;
wire net_11864;
wire net_4677;
wire net_11420;
wire net_8033;
wire net_10996;
wire net_10038;
wire net_5768;
wire net_174;
wire net_2607;
wire net_7799;
wire net_7957;
wire net_10971;
wire net_7987;
wire net_7214;
wire net_11691;
wire net_8769;
wire net_6202;
wire net_1831;
wire net_1482;
wire net_13870;
wire net_5023;
wire net_3291;
wire net_2168;
wire net_3306;
wire net_2928;
wire net_7563;
wire net_1030;
wire net_1885;
wire net_4129;
wire net_1485;
wire net_14357;
wire net_10272;
wire net_9236;
wire net_10406;
wire net_10053;
wire net_6929;
wire net_3245;
wire net_13300;
wire net_10682;
wire net_9385;
wire net_7473;
wire net_6920;
wire net_7335;
wire net_7387;
wire net_11987;
wire net_13407;
wire net_12740;
wire net_12711;
wire net_10787;
wire net_11498;
wire net_10031;
wire net_4773;
wire net_4201;
wire net_13929;
wire net_4273;
wire net_1969;
wire net_745;
wire net_9651;
wire net_7991;
wire net_12306;
wire net_8009;
wire net_7064;
wire net_14271;
wire net_933;
wire net_1244;
wire net_12532;
wire net_429;
wire net_12036;
wire net_10966;
wire net_10860;
wire net_3377;
wire net_373;
wire net_12593;
wire net_356;
wire net_13701;
wire net_452;
wire net_11432;
wire net_545;
wire net_3683;
wire net_11700;
wire net_1483;
wire net_2147;
wire net_10361;
wire net_8067;
wire net_560;
wire net_3031;
wire net_9253;
wire net_10098;
wire net_5148;
wire net_4603;
wire net_2645;
wire net_14017;
wire net_10433;
wire net_11951;
wire net_5510;
wire net_5356;
wire net_10500;
wire net_9359;
wire net_6709;
wire net_14386;
wire net_8078;
wire net_7310;
wire net_7674;
wire net_7386;
wire net_6684;
wire net_13151;
wire net_4278;
wire net_7522;
wire net_2674;
wire net_13801;
wire net_2872;
wire net_6833;
wire net_2432;
wire net_12780;
wire net_10193;
wire net_8934;
wire net_7059;
wire net_5401;
wire net_322;
wire net_1671;
wire net_4764;
wire net_420;
wire net_665;
wire net_1746;
wire net_2222;
wire net_8944;
wire net_2322;
wire net_2825;
wire net_7209;
wire net_3670;
wire net_9109;
wire net_5940;
wire net_4344;
wire net_13376;
wire net_3341;
wire net_5985;
wire net_7925;
wire net_1072;
wire net_6606;
wire net_10182;
wire net_10376;
wire net_7136;
wire net_4861;
wire net_13738;
wire net_11666;
wire net_1706;
wire net_4510;
wire net_11113;
wire net_3574;
wire net_6278;
wire net_5994;
wire net_1730;
wire net_10852;
wire net_2921;
wire net_3289;
wire net_8829;
wire net_6311;
wire net_13501;
wire net_4575;
wire net_10225;
wire net_651;
wire net_12097;
wire net_2931;
wire net_3114;
wire net_3415;
wire net_6846;
wire net_10019;
wire net_744;
wire net_8276;
wire net_4967;
wire net_598;
wire net_7985;
wire net_4136;
wire net_2011;
wire net_3455;
wire net_6317;
wire net_12011;
wire net_10068;
wire net_777;
wire net_4806;
wire net_13203;
wire net_7185;
wire net_4818;
wire net_3157;
wire net_8690;
wire net_2820;
wire net_8348;
wire net_7532;
wire net_6091;
wire net_490;
wire net_4404;
wire net_11497;
wire net_3068;
wire net_12677;
wire net_8585;
wire net_5973;
wire net_12130;
wire net_3892;
wire net_13930;
wire net_7921;
wire net_6009;
wire net_3462;
wire net_7080;
wire net_6739;
wire net_5978;
wire net_5670;
wire net_632;
wire net_4439;
wire net_843;
wire net_3860;
wire net_5602;
wire net_12720;
wire net_7638;
wire net_2841;
wire net_10106;
wire net_10063;
wire net_11889;
wire net_5484;
wire net_7255;
wire net_5813;
wire net_1977;
wire net_11959;
wire net_2100;
wire net_2938;
wire net_14009;
wire net_2122;
wire net_12572;
wire net_6617;
wire net_1171;
wire net_10691;
wire net_1540;
wire net_9680;
wire net_248;
wire net_3594;
wire net_6548;
wire net_5341;
wire net_11835;
wire net_9734;
wire net_10393;
wire net_1725;
wire net_14064;
wire net_13583;
wire net_3541;
wire net_5649;
wire net_13718;
wire net_3532;
wire net_12725;
wire net_5112;
wire net_1767;
wire net_4010;
wire net_7333;
wire net_11827;
wire net_1640;
wire net_12956;
wire net_13788;
wire net_10303;
wire net_9750;
wire net_5190;
wire net_2724;
wire net_11916;
wire net_6554;
wire net_12090;
wire net_7504;
wire net_503;
wire net_1741;
wire net_10141;
wire net_13510;
wire net_4227;
wire net_5695;
wire net_11818;
wire net_1672;
wire net_2103;
wire net_996;
wire net_3091;
wire net_7550;
wire net_14165;
wire net_2994;
wire net_11617;
wire net_959;
wire net_5381;
wire net_10838;
wire net_8327;
wire net_11476;
wire net_7911;
wire net_3051;
wire net_8767;
wire net_4004;
wire net_7706;
wire net_2345;
wire net_12342;
wire net_9304;
wire net_2973;
wire net_6981;
wire net_6460;
wire net_3106;
wire net_13792;
wire net_2503;
wire net_9705;
wire net_6660;
wire net_2164;
wire net_11079;
wire net_6646;
wire net_5659;
wire net_11797;
wire net_13578;
wire net_6469;
wire net_3751;
wire net_8330;
wire net_9821;
wire net_6211;
wire net_5311;
wire net_4564;
wire net_13670;
wire net_2338;
wire net_10982;
wire net_10556;
wire net_4606;
wire net_3721;
wire net_2616;
wire net_8200;
wire x1358;
wire net_8894;
wire net_282;
wire net_1596;
wire net_10804;
wire net_6572;
wire net_12397;
wire net_4296;
wire net_11677;
wire net_7416;
wire net_6901;
wire net_11857;
wire net_5051;
wire net_10688;
wire net_10908;
wire net_11693;
wire net_2370;
wire net_2047;
wire net_8320;
wire net_2469;
wire net_11214;
wire net_9647;
wire net_12733;
wire net_2693;
wire net_13115;
wire net_11212;
wire net_10458;
wire net_1012;
wire net_1404;
wire net_12765;
wire net_12185;
wire net_9621;
wire net_907;
wire net_3076;
wire net_8809;
wire net_5807;
wire net_4694;
wire net_395;
wire net_2036;
wire net_12988;
wire net_9182;
wire net_8070;
wire net_2719;
wire net_10219;
wire net_6343;
wire net_8623;
wire net_2323;
wire net_9688;
wire net_3867;
wire net_3677;
wire net_641;
wire net_4811;
wire net_5451;
wire net_2798;
wire net_5071;
wire net_10977;
wire net_10599;
wire net_4972;
wire net_3869;
wire net_14335;
wire net_1152;
wire net_1226;
wire net_10459;
wire net_14212;
wire net_10525;
wire net_8429;
wire net_4890;
wire net_1901;
wire net_3021;
wire net_5315;
wire net_3711;
wire net_10257;
wire net_3805;
wire net_7580;
wire net_3942;
wire net_7836;
wire net_4580;
wire net_602;
wire net_12605;
wire net_8273;
wire net_2379;
wire net_13199;
wire net_1818;
wire net_12783;
wire net_11850;
wire net_13335;
wire net_12288;
wire net_10932;
wire net_8646;
wire net_2918;
wire net_11658;
wire net_9371;
wire net_1497;
wire net_1800;
wire net_4634;
wire net_279;
wire net_1523;
wire net_3347;
wire net_1656;
wire net_6522;
wire net_12281;
wire net_4039;
wire net_11326;
wire net_4030;
wire net_691;
wire net_10212;
wire net_6951;
wire net_10713;
wire net_6337;
wire net_14119;
wire net_5551;
wire net_3178;
wire net_2701;
wire net_14289;
wire net_10422;
wire net_4078;
wire net_1863;
wire net_2833;
wire net_2561;
wire net_12170;
wire net_13775;
wire net_10774;
wire net_8399;
wire net_2519;
wire net_471;
wire net_1055;
wire net_3813;
wire net_878;
wire net_1531;
wire net_3894;
wire net_1159;
wire net_10666;
wire net_518;
wire net_10334;
wire net_861;
wire net_6755;
wire net_7217;
wire net_12645;
wire net_11136;
wire net_10172;
wire net_13533;
wire net_929;
wire net_6696;
wire net_12400;
wire net_11102;
wire net_2523;
wire net_4914;
wire net_11779;
wire net_4210;
wire net_3954;
wire net_12939;
wire net_11811;
wire net_5726;
wire net_1565;
wire net_10882;
wire net_8544;
wire net_5262;
wire net_169;
wire net_12951;
wire net_9948;
wire net_5213;
wire net_7696;
wire net_8567;
wire net_12986;
wire net_2234;
wire net_4552;
wire net_12120;
wire net_6828;
wire net_10481;
wire net_967;
wire net_1527;
wire net_13270;
wire net_13056;
wire net_4420;
wire net_11849;
wire net_8007;
wire net_268;
wire net_13861;
wire net_4318;
wire net_12358;
wire net_11475;
wire net_3386;
wire net_4134;
wire net_4910;
wire net_6631;
wire net_13324;
wire net_1645;
wire net_2962;
wire net_9406;
wire net_4365;
wire net_176;
wire net_3638;
wire net_2570;
wire net_12410;
wire net_5793;
wire net_13195;
wire net_3354;
wire net_9468;
wire net_614;
wire net_2712;
wire net_13976;
wire net_2005;
wire net_12505;
wire net_1123;
wire net_2771;
wire net_8293;
wire net_6040;
wire net_4897;
wire net_3194;
wire net_3572;
wire net_5537;
wire net_13911;
wire net_9343;
wire net_4740;
wire net_9980;
wire net_8338;
wire net_1192;
wire net_11241;
wire net_10697;
wire net_6857;
wire net_4838;
wire net_5958;
wire net_14368;
wire net_4542;
wire net_984;
wire net_3363;
wire net_11894;
wire net_11753;
wire net_11705;
wire net_6407;
wire net_5467;
wire net_10915;
wire net_7263;
wire net_13652;
wire net_8730;
wire net_4061;
wire net_1105;
wire net_12370;
wire net_12201;
wire net_2172;
wire net_3156;
wire net_12109;
wire net_2482;
wire net_13043;
wire net_11448;
wire net_7275;
wire net_707;
wire net_14023;
wire net_6534;
wire net_7491;
wire net_4457;
wire net_5039;
wire net_9519;
wire net_11174;
wire net_6867;
wire net_4850;
wire net_1856;
wire net_830;
wire net_13828;
wire net_4531;
wire net_575;
wire net_1279;
wire net_1047;
wire net_5833;
wire net_13003;
wire net_4715;
wire net_7169;
wire net_9475;
wire net_3697;
wire net_12642;
wire net_11374;
wire net_8439;
wire net_6394;
wire net_12582;
wire net_11425;
wire net_6193;
wire net_4688;
wire net_2631;
wire net_8101;
wire net_12386;
wire net_6431;
wire net_3618;
wire net_12926;
wire net_1467;
wire net_9156;
wire net_7562;
wire net_5623;
wire net_1061;
wire net_3181;
wire net_14012;
wire net_10842;
wire net_5951;
wire net_5512;
wire net_765;
wire net_1342;
wire net_2633;
wire net_1666;
wire net_3837;
wire net_9096;
wire net_4839;
wire net_2288;
wire net_4193;
wire net_8718;
wire net_13752;
wire net_8573;
wire net_8253;
wire net_11189;
wire net_2099;
wire net_5745;
wire net_6750;
wire net_5182;
wire net_7612;
wire net_13454;
wire net_9809;
wire net_10302;
wire net_8195;
wire net_5850;
wire net_5646;
wire net_2021;
wire net_11248;
wire net_1068;
wire net_186;
wire net_14378;
wire net_3983;
wire net_8121;
wire net_2495;
wire net_12823;
wire net_6672;
wire net_3814;
wire net_10534;
wire net_1050;
wire net_6266;
wire net_2072;
wire net_2760;
wire net_5914;
wire net_4751;
wire net_1872;
wire net_2271;
wire net_1716;
wire net_13926;
wire net_5327;
wire net_5003;
wire net_1607;
wire net_14083;
wire net_11768;
wire net_5247;
wire net_12164;
wire net_6125;
wire net_7143;
wire net_13472;
wire net_7983;
wire net_1263;
wire net_12331;
wire net_4591;
wire net_196;
wire net_3452;
wire net_14356;
wire net_11969;
wire net_10324;
wire net_8766;
wire net_2067;
wire net_14243;
wire net_8120;
wire net_3130;
wire net_8881;
wire net_8572;
wire net_5183;
wire net_7200;
wire net_5704;
wire net_1639;
wire net_5267;
wire net_4126;
wire net_4289;
wire net_4549;
wire net_9775;
wire net_7284;
wire net_11431;
wire net_3625;
wire net_9510;
wire net_4145;
wire net_7604;
wire net_13806;
wire net_4712;
wire net_11340;
wire net_260;
wire net_2947;
wire net_12552;
wire net_11784;
wire net_3137;
wire net_11981;
wire net_732;
wire net_2152;
wire net_8649;
wire net_12880;
wire net_12423;
wire net_5286;
wire net_1597;
wire net_8285;
wire net_6105;
wire net_7946;
wire net_2088;
wire net_13083;
wire net_8785;
wire net_7572;
wire net_6423;
wire net_13963;
wire net_10655;
wire net_7593;
wire net_4217;
wire net_2689;
wire net_3988;
wire net_2761;
wire net_6396;
wire net_8422;
wire net_3788;
wire net_4355;
wire net_11678;
wire net_11092;
wire net_10623;
wire net_1503;
wire net_3961;
wire net_13970;
wire net_8430;
wire net_4639;
wire net_8628;
wire net_11089;
wire net_449;
wire net_5494;
wire net_5234;
wire net_9299;
wire net_8225;
wire net_11523;
wire net_11928;
wire net_9574;
wire net_12638;
wire net_1087;
wire net_4234;
wire net_11064;
wire net_3995;
wire net_733;
wire net_8245;
wire net_887;
wire net_5856;
wire net_9606;
wire net_12362;
wire net_11409;
wire net_6098;
wire net_11975;
wire net_7537;
wire net_6595;
wire net_13663;
wire net_11653;
wire net_10491;
wire net_6151;
wire net_13866;
wire net_6301;
wire net_5443;
wire net_2308;
wire net_5211;
wire net_4731;
wire net_2989;
wire net_9105;
wire net_497;
wire net_6720;
wire net_4628;
wire net_12494;
wire net_2770;
wire net_7658;
wire net_1424;
wire net_2636;
wire net_8160;
wire net_1414;
wire net_4375;
wire net_4153;
wire net_4412;
wire net_11307;
wire net_10927;
wire net_9864;
wire net_300;
wire net_9287;
wire net_2652;
wire net_5526;
wire net_10149;
wire net_1233;
wire net_2720;
wire net_8167;
wire net_6351;
wire net_4280;
wire net_12917;
wire net_10347;
wire net_1834;
wire net_9563;
wire net_950;
wire net_6027;
wire net_4925;
wire net_13213;
wire net_13024;
wire net_13313;
wire net_11441;
wire net_11355;
wire net_5474;
wire net_14363;
wire net_9839;
wire net_9745;
wire net_2816;
wire net_6610;
wire net_7651;
wire net_8984;
wire net_14344;
wire net_12565;
wire net_1214;
wire net_9529;
wire net_3641;
wire net_13405;
wire net_12895;
wire net_10203;
wire net_866;
wire net_11946;
wire net_13603;
wire net_12700;
wire net_5194;
wire net_4220;
wire net_12025;
wire net_3150;
wire net_9596;
wire net_10681;
wire net_1032;
wire net_567;
wire net_13985;
wire net_3726;
wire net_3979;
wire net_5255;
wire net_5787;
wire net_272;
wire net_8822;
wire net_13345;
wire net_13384;
wire net_8458;
wire net_3939;
wire net_12712;
wire net_12480;
wire net_1024;
wire net_1590;
wire net_14097;
wire net_1612;
wire net_839;
wire net_11121;
wire net_814;
wire net_13542;
wire net_11778;
wire net_13685;
wire net_7095;
wire net_8128;
wire net_5840;
wire net_6184;
wire net_12705;
wire net_4660;
wire x786;
wire net_12525;
wire net_14003;
wire net_10639;
wire net_4785;
wire net_3930;
wire x1459;
wire net_9815;
wire net_2586;
wire net_3299;
wire net_13013;
wire net_10290;
wire net_1655;
wire net_11294;
wire net_6963;
wire net_7805;
wire net_11313;
wire net_954;
wire net_2365;
wire net_13094;
wire net_4565;
wire net_9051;
wire net_9037;
wire net_4797;
wire net_8796;
wire net_11271;
wire net_8962;
wire net_10897;
wire net_9240;
wire net_10810;
wire net_2361;
wire net_2598;
wire net_11194;
wire net_2879;
wire net_10152;
wire net_1680;
wire net_14219;
wire net_3302;
wire net_13359;
wire net_13265;
wire net_9545;
wire net_10411;
wire net_7540;
wire net_12445;
wire net_11337;
wire net_11989;
wire net_4790;
wire net_3187;
wire net_12048;
wire net_2622;
wire net_5363;
wire net_5966;
wire net_7529;
wire net_10514;
wire net_8294;
wire net_10997;
wire net_8888;
wire net_6665;
wire net_4900;
wire net_9807;
wire net_13222;
wire net_2262;
wire net_7505;
wire net_6502;
wire net_7305;
wire net_6163;
wire net_3011;
wire net_13079;
wire net_10643;
wire net_2087;
wire net_13187;
wire net_10021;
wire net_1002;
wire net_12946;
wire net_6817;
wire net_6000;
wire net_9079;
wire net_8863;
wire net_7620;
wire net_11930;
wire net_7224;
wire net_6118;
wire net_13628;
wire net_3188;
wire net_12466;
wire net_9536;
wire net_13308;
wire net_12887;
wire net_1993;
wire net_8198;
wire net_3010;
wire net_11128;
wire net_881;
wire net_12657;
wire net_8724;
wire net_10544;
wire net_2805;
wire net_8683;
wire net_1397;
wire net_2903;
wire net_14231;
wire net_4474;
wire net_11623;
wire net_8392;
wire net_9556;
wire net_4128;
wire net_4923;
wire net_1954;
wire net_13036;
wire net_11866;
wire net_3873;
wire net_7615;
wire net_6015;
wire net_2155;
wire net_14294;
wire net_6741;
wire net_168;
wire net_2041;
wire net_13090;
wire net_11830;
wire net_10354;
wire net_385;
wire net_13253;
wire net_2609;
wire net_14179;
wire net_5736;
wire net_5365;
wire net_7937;
wire net_7930;
wire net_5404;
wire net_5044;
wire net_10260;
wire net_8657;
wire net_7196;
wire net_8139;
wire net_12197;
wire net_10468;
wire net_11220;
wire net_6236;
wire net_14143;
wire net_2423;
wire net_7660;
wire net_13675;
wire net_7535;
wire net_6723;
wire net_2380;
wire net_3393;
wire net_4548;
wire net_13875;
wire net_8231;
wire net_9323;
wire net_12379;
wire net_11283;
wire net_895;
wire net_10781;
wire net_6412;
wire net_11603;
wire net_5990;
wire net_14358;
wire net_1412;
wire net_12006;
wire net_8240;
wire net_7048;
wire net_9715;
wire net_7767;
wire net_8831;
wire net_12394;
wire net_10683;
wire net_12965;
wire net_12327;
wire net_13357;
wire net_1255;
wire net_7358;
wire net_12603;
wire net_7211;
wire net_1250;
wire net_8247;
wire net_13928;
wire net_207;
wire net_3040;
wire net_13762;
wire net_10825;
wire net_3557;
wire net_10609;
wire net_3643;
wire net_8801;
wire net_3004;
wire net_13639;
wire net_12102;
wire net_8014;
wire net_13382;
wire net_11874;
wire net_1689;
wire net_12624;
wire net_10345;
wire net_10271;
wire net_7244;
wire net_6186;
wire net_7981;
wire net_10315;
wire net_8569;
wire net_9757;
wire net_5698;
wire net_3830;
wire net_8464;
wire net_274;
wire net_13987;
wire net_1075;
wire net_12806;
wire net_12561;
wire net_9387;
wire net_10282;
wire net_13360;
wire net_14044;
wire net_6204;
wire net_833;
wire net_930;
wire net_2387;
wire net_12599;
wire net_12744;
wire net_9316;
wire net_8358;
wire net_6656;
wire net_4723;
wire net_2267;
wire net_4758;
wire net_7323;
wire net_4249;
wire net_4769;
wire net_13590;
wire net_12931;
wire net_13681;
wire net_11349;
wire net_1399;
wire net_8529;
wire net_10016;
wire net_8667;
wire net_4888;
wire net_9539;
wire net_3350;
wire net_3553;
wire net_5161;
wire net_7623;
wire net_3304;
wire net_12751;
wire net_2549;
wire net_11024;
wire net_8654;
wire net_1781;
wire net_14390;
wire net_3465;
wire net_6217;
wire net_7457;
wire net_3049;
wire net_10299;
wire net_6918;
wire net_637;
wire net_13062;
wire net_2514;
wire net_9250;
wire net_2390;
wire net_12183;
wire net_5436;
wire net_4775;
wire net_2686;
wire net_3474;
wire net_5577;
wire net_5472;
wire net_2013;
wire net_1509;
wire net_529;
wire net_7477;
wire net_13503;
wire x1479;
wire net_9447;
wire net_3495;
wire net_11262;
wire net_9887;
wire net_2028;
wire net_2553;
wire net_9758;
wire net_4881;
wire net_1889;
wire net_3766;
wire net_7361;
wire net_12065;
wire net_8717;
wire net_2981;
wire net_8506;
wire net_6477;
wire net_11303;
wire net_1164;
wire net_10817;
wire net_8912;
wire net_6810;
wire net_121;
wire net_5228;
wire net_6923;
wire net_11148;
wire net_7475;
wire net_12500;
wire net_2583;
wire net_9762;
wire x1443;
wire net_5708;
wire net_3820;
wire net_3799;
wire net_8854;
wire net_4175;
wire net_10938;
wire net_5824;
wire net_4665;
wire net_9366;
wire net_2664;
wire net_14206;
wire net_2706;
wire net_11202;
wire net_5163;
wire net_849;
wire net_5580;
wire net_14161;
wire net_11842;
wire net_10577;
wire net_8304;
wire net_7470;
wire net_5294;
wire net_11681;
wire net_2602;
wire net_6366;
wire net_5751;
wire net_401;
wire net_8449;
wire net_8165;
wire net_10720;
wire net_4484;
wire net_3798;
wire net_2714;
wire net_2183;
wire net_2557;
wire net_440;
wire net_14265;
wire net_9229;
wire net_11361;
wire net_8069;
wire net_8048;
wire net_758;
wire net_10866;
wire net_5664;
wire net_13754;
wire net_6874;
wire net_4652;
wire net_718;
wire net_10846;
wire net_7773;
wire net_6178;
wire net_13563;
wire net_7682;
wire net_14193;
wire net_8707;
wire net_5504;
wire net_12995;
wire net_5714;
wire net_13367;
wire net_5838;
wire net_4998;
wire net_3255;
wire net_13946;
wire net_12215;
wire net_12303;
wire net_14078;
wire net_13545;
wire net_9848;
wire net_6564;
wire net_4448;
wire x837;
wire net_9797;
wire net_9419;
wire net_336;
wire net_12973;
wire net_10946;
wire net_5306;
wire net_10404;
wire net_14033;
wire net_9577;
wire net_1578;
wire net_9938;
wire net_11539;
wire net_8417;
wire net_2917;
wire net_8404;
wire net_6711;
wire net_3221;
wire net_697;
wire net_2003;
wire net_7708;
wire net_605;
wire net_3411;
wire net_5053;
wire net_4987;
wire net_10447;
wire net_3426;
wire net_9233;
wire net_13008;
wire net_5095;
wire net_9527;
wire net_924;
wire net_8883;
wire net_12255;
wire net_5469;
wire net_1333;
wire net_5325;
wire net_9205;
wire net_10980;
wire net_7829;
wire net_2348;
wire net_5924;
wire net_489;
wire net_5593;
wire net_5107;
wire net_3082;
wire net_5859;
wire net_11503;
wire net_10802;
wire net_5457;
wire net_13521;
wire net_3676;
wire net_4185;
wire net_6143;
wire net_4646;
wire net_4204;
wire net_5630;
wire net_2748;
wire net_9991;
wire net_11561;
wire net_9611;
wire net_7591;
wire net_6072;
wire net_9135;
wire net_8060;
wire net_251;
wire net_6682;
wire net_2054;
wire net_9880;
wire net_128;
wire net_6295;
wire net_840;
wire net_9206;
wire net_10632;
wire net_9133;
wire net_8086;
wire net_14057;
wire net_10901;
wire net_6933;
wire net_5789;
wire net_13281;
wire net_14133;
wire net_12928;
wire x1261;
wire net_11229;
wire net_2793;
wire net_9914;
wire net_411;
wire net_2137;
wire net_1836;
wire net_10570;
wire net_8783;
wire net_4310;
wire net_11689;
wire net_12220;
wire net_11256;
wire net_12688;
wire net_5922;
wire net_13158;
wire net_7874;
wire net_7293;
wire net_11557;
wire net_8975;
wire net_3430;
wire net_8266;
wire net_1862;
wire net_13889;
wire net_10052;
wire net_2317;
wire net_6795;
wire net_6248;
wire net_8135;
wire net_4244;
wire net_10584;
wire net_7887;
wire net_6035;
wire net_6930;
wire net_6492;
wire net_3583;
wire net_8183;
wire net_4396;
wire net_6158;
wire net_10536;
wire net_8219;
wire net_2373;
wire net_11694;
wire net_14109;
wire net_9273;
wire net_2398;
wire net_4581;
wire net_12140;
wire net_7811;
wire net_4431;
wire net_10943;
wire net_7821;
wire net_7746;
wire net_9282;
wire net_3315;
wire net_2455;
wire net_1609;
wire net_402;
wire net_7847;
wire net_4047;
wire net_3448;
wire net_12732;
wire net_7108;
wire net_3248;
wire net_10753;
wire net_12450;
wire net_2274;
wire net_11597;
wire net_8493;
wire net_8744;
wire net_12681;
wire net_1386;
wire net_11488;
wire net_7841;
wire net_13859;
wire net_10950;
wire net_9431;
wire net_12345;
wire net_2359;
wire net_8949;
wire net_6546;
wire net_6115;
wire net_12805;
wire net_10550;
wire net_13101;
wire net_12574;
wire net_5991;
wire net_10252;
wire net_5101;
wire net_11585;
wire net_10127;
wire net_4102;
wire net_2186;
wire net_3696;
wire net_13551;
wire net_3473;
wire net_6908;
wire net_1430;
wire net_9964;
wire net_12062;
wire net_6892;
wire net_569;
wire net_2478;
wire net_6429;
wire net_2563;
wire net_13877;
wire net_12435;
wire net_9484;
wire net_9243;
wire net_8051;
wire net_5679;
wire net_12767;
wire net_3408;
wire net_4870;
wire net_630;
wire net_12514;
wire net_8857;
wire net_2202;
wire net_2490;
wire net_8841;
wire net_4018;
wire net_4428;
wire net_1791;
wire net_6826;
wire net_4339;
wire net_1471;
wire net_9975;
wire net_8997;
wire net_7667;
wire net_3608;
wire net_13696;
wire net_3124;
wire net_1903;
wire net_2407;
wire net_13467;
wire x130657;
wire net_10600;
wire net_912;
wire net_13162;
wire net_7412;
wire net_13414;
wire net_13562;
wire net_7018;
wire net_4517;
wire net_2078;
wire net_779;
wire net_1928;
wire net_3841;
wire net_12473;
wire net_1328;
wire net_9871;
wire net_234;
wire net_2859;
wire net_12634;
wire net_4151;
wire net_2884;
wire net_3848;
wire net_13258;
wire net_5372;
wire net_5142;
wire net_4942;
wire net_13616;
wire net_3205;
wire net_1094;
wire net_3487;
wire net_2749;
wire net_7390;
wire net_5764;
wire net_855;
wire net_11469;
wire net_674;
wire net_7732;
wire net_11032;
wire net_9506;
wire net_303;
wire net_10041;
wire net_6583;
wire net_9128;
wire net_9982;
wire net_491;
wire net_2475;
wire net_11460;
wire net_9925;
wire net_1299;
wire net_6679;
wire net_948;
wire net_2937;
wire net_7792;
wire net_7657;
wire net_7400;
wire net_6191;
wire net_11573;
wire net_12249;
wire net_12993;
wire net_7865;
wire net_4743;
wire net_13767;
wire net_876;
wire net_2593;
wire net_6479;
wire net_2162;
wire net_10833;
wire net_9478;
wire net_2439;
wire net_13297;
wire net_11048;
wire net_7154;
wire net_172;
wire net_9646;
wire net_4341;
wire net_13460;
wire net_8601;
wire net_11960;
wire net_1458;
wire net_4048;
wire net_5587;
wire net_10749;
wire net_4570;
wire net_10184;
wire net_10244;
wire net_5933;
wire net_6689;
wire x264;
wire net_10591;
wire net_905;
wire net_14122;
wire net_12233;
wire net_13934;
wire net_142;
wire net_7034;
wire net_6446;
wire x1101;
wire net_8029;
wire net_11939;
wire net_9050;
wire net_6198;
wire net_2229;
wire net_13842;
wire net_10613;
wire net_5774;
wire net_158;
wire net_7370;
wire net_3200;
wire net_3733;
wire net_3881;
wire net_12263;
wire net_8598;
wire net_5624;
wire net_11944;
wire net_2504;
wire net_11571;
wire net_5650;
wire net_2175;
wire net_3784;
wire net_10519;
wire net_14136;
wire net_10214;
wire net_8091;
wire net_8057;
wire net_6258;
wire net_8361;
wire net_2116;
wire net_1758;
wire net_4327;
wire net_13840;
wire net_11334;
wire net_8813;
wire net_8035;
wire net_11802;
wire net_9572;
wire net_8090;
wire net_1769;
wire net_9115;
wire net_6694;
wire net_1967;
wire net_11565;
wire net_9333;
wire net_5171;
wire net_1567;
wire net_8020;
wire net_6860;
wire net_6322;
wire net_12087;
wire net_8754;
wire net_465;
wire net_11186;
wire net_8152;
wire net_9520;
wire net_1883;
wire net_11233;
wire net_476;
wire net_2783;
wire net_6055;
wire net_7079;
wire net_382;
wire net_3058;
wire net_11412;
wire net_8484;
wire net_11259;
wire net_5301;
wire net_583;
wire net_1315;
wire net_6994;
wire net_5904;
wire net_7041;
wire net_5358;
wire net_10073;
wire net_9408;
wire net_14173;
wire net_9767;
wire net_5208;
wire net_13144;
wire net_5019;
wire net_9903;
wire net_9376;
wire net_6956;
wire net_13055;
wire net_9695;
wire net_4719;
wire net_10379;
wire net_10138;
wire net_4977;
wire net_9005;
wire net_5075;
wire net_4460;
wire net_11646;
wire net_7327;
wire net_220;
wire net_1465;
wire net_293;
wire net_11153;
wire net_3666;
wire net_13599;
wire net_11890;
wire net_4982;
wire net_13303;
wire net_1938;
wire net_543;
wire net_625;
wire net_3760;
wire net_11411;
wire net_10708;
wire net_1823;
wire net_5081;
wire net_11637;
wire net_13790;
wire net_191;
wire net_3576;
wire net_4331;
wire net_2909;
wire net_4953;
wire net_558;
wire net_2069;
wire net_9607;
wire net_4697;
wire net_5638;
wire net_1618;
wire net_10910;
wire net_14399;
wire net_2497;
wire net_7899;
wire net_11594;
wire net_12157;
wire net_10562;
wire net_7006;
wire net_3562;
wire net_1694;
wire net_12844;
wire net_4991;
wire net_910;
wire net_12356;
wire net_5885;
wire net_7112;
wire x1374;
wire net_11905;
wire net_5394;
wire net_7944;
wire net_2412;
wire net_4023;
wire net_12070;
wire net_4265;
wire net_7755;
wire net_6881;
wire net_4450;
wire net_4158;
wire net_6942;
wire net_13442;
wire net_1984;
wire net_13959;
wire net_13527;
wire net_315;
wire net_1375;
wire net_4670;
wire net_10734;
wire net_1944;
wire net_4006;
wire net_11545;
wire net_8212;
wire net_1351;
wire net_1775;
wire net_10112;
wire net_10158;
wire net_297;
wire net_346;
wire net_1535;
wire net_2400;
wire net_5543;
wire net_10693;
wire net_13725;
wire net_8661;
wire net_10959;
wire net_2034;
wire net_229;
wire net_4360;
wire net_8921;
wire net_4962;
wire net_1808;
wire net_3256;
wire net_687;
wire net_3266;
wire net_13122;
wire net_4160;
wire net_13339;
wire net_3888;
wire net_7072;
wire net_13949;
wire net_13438;
wire net_14303;
wire net_10567;
wire net_3322;
wire net_2533;
wire net_10267;
wire net_3566;
wire net_1913;
wire net_12297;
wire net_3596;
wire net_13243;
wire net_11526;
wire net_7830;
wire net_9673;
wire net_9016;
wire net_7642;
wire net_10143;
wire net_11904;
wire net_5021;
wire net_9732;
wire net_9264;
wire net_6615;
wire net_12279;
wire net_7409;
wire net_13741;
wire net_7671;
wire net_1760;
wire net_9345;
wire net_9296;
wire net_5415;
wire net_13492;
wire net_1184;
wire net_7714;
wire net_4055;
wire x361;
wire net_5339;
wire net_3926;
wire net_6482;
wire net_6961;
wire net_4849;
wire net_7383;
wire net_10722;
wire net_5758;
wire net_5425;
wire net_3403;
wire net_10002;
wire net_1960;
wire net_6977;
wire net_10718;
wire net_9660;
wire net_3093;
wire net_7935;
wire net_12820;
wire net_6886;
wire net_647;
wire net_3247;
wire net_12548;
wire net_7435;
wire net_6452;
wire net_8684;
wire net_2464;
wire net_12272;
wire net_9492;
wire net_9145;
wire net_4256;
wire net_828;
wire net_6222;
wire net_3839;
wire net_6513;
wire net_4490;
wire net_1603;
wire net_14349;
wire net_12222;
wire net_13031;
wire net_2732;
wire net_10009;
wire net_7446;
wire net_10108;
wire net_13483;
wire net_11809;
wire net_11017;
wire net_8368;
wire net_8385;
wire net_7345;
wire net_3521;
wire net_1096;
wire net_795;
wire net_982;
wire net_8153;
wire net_11403;
wire net_9610;
wire net_1580;
wire net_1406;
wire net_9093;
wire net_5287;
wire net_3896;
wire net_4384;
wire net_6462;
wire net_9189;
wire net_8490;
wire net_10463;
wire net_9314;
wire net_1434;
wire net_6996;
wire net_3668;
wire net_6096;
wire net_9576;
wire net_9823;
wire net_4912;
wire net_10012;
wire net_5130;
wire net_11870;
wire net_5617;
wire net_4946;
wire net_6002;
wire net_774;
wire net_10071;
wire net_5748;
wire net_12076;
wire net_8180;
wire net_6958;
wire net_11393;
wire net_10869;
wire net_5049;
wire net_8892;
wire net_13235;
wire net_7221;
wire net_11058;
wire net_501;
wire net_8899;
wire net_3679;
wire net_225;
wire net_4489;
wire net_12344;
wire net_5818;
wire net_3128;
wire net_4733;
wire net_12937;
wire net_6524;
wire net_6213;
wire net_4692;
wire net_9769;
wire net_6644;
wire net_7481;
wire net_9170;
wire net_13327;
wire net_5313;
wire net_447;
wire net_9180;
wire net_871;
wire net_2611;
wire net_11804;
wire net_390;
wire net_13279;
wire net_5772;
wire net_1154;
wire net_6318;
wire net_11789;
wire net_11219;
wire net_6983;
wire net_6593;
wire net_14031;
wire net_10755;
wire net_13371;
wire net_11782;
wire net_9703;
wire net_12368;
wire net_8952;
wire net_13944;
wire net_4294;
wire net_5128;
wire net_10923;
wire net_6062;
wire net_12735;
wire net_7900;
wire net_7494;
wire net_14038;
wire net_4106;
wire net_12798;
wire net_2951;
wire net_8621;
wire net_3631;
wire net_12854;
wire net_2293;
wire net_12132;
wire net_280;
wire net_12027;
wire net_12715;
wire net_495;
wire net_13022;
wire net_10105;
wire net_1802;
wire net_10569;
wire net_7694;
wire net_13180;
wire net_2140;
wire net_5482;
wire net_13975;
wire net_6345;
wire net_10456;
wire net_13211;
wire net_7637;
wire net_2517;
wire net_11318;
wire net_8798;
wire net_2316;
wire net_12105;
wire net_8644;
wire net_6457;
wire net_2755;
wire net_6100;
wire net_12172;
wire net_6356;
wire net_13850;
wire net_1678;
wire net_2703;
wire net_11273;
wire net_13524;
wire net_6638;
wire net_3366;
wire net_14214;
wire net_1441;
wire net_10210;
wire net_969;
wire net_9154;
wire net_8271;
wire net_1525;
wire net_7097;
wire net_12710;
wire net_11458;
wire net_7737;
wire net_7206;
wire net_4003;
wire net_821;
wire net_13444;
wire net_6757;
wire net_4177;
wire net_9350;
wire net_8511;
wire net_7757;
wire net_11726;
wire net_8936;
wire net_10934;
wire net_3436;
wire net_8345;
wire net_2335;
wire net_14159;
wire net_11210;
wire net_3940;
wire net_10812;
wire net_8708;
wire net_7725;
wire net_3911;
wire net_11533;
wire net_13913;
wire net_11161;
wire net_12866;
wire net_5337;
wire net_14153;
wire net_2618;
wire net_8638;
wire net_4316;
wire net_3365;
wire net_10711;
wire net_6045;
wire net_14372;
wire net_14099;
wire net_6540;
wire net_12698;
wire net_8587;
wire net_7952;
wire net_1114;
wire net_12786;
wire net_10619;
wire net_8670;
wire net_13431;
wire net_7090;
wire net_3388;
wire net_5411;
wire net_12691;
wire net_1748;
wire net_10664;
wire net_4116;
wire net_3078;
wire net_3218;
wire net_13005;
wire net_11882;
wire net_4632;
wire net_2964;
wire net_12283;
wire net_9946;
wire net_8171;
wire net_7266;
wire net_6738;
wire net_2232;
wire net_2343;
wire net_726;
wire net_13241;
wire net_6690;
wire net_6565;
wire net_3811;
wire net_1028;
wire net_14287;
wire net_1529;
wire net_600;
wire net_14021;
wire net_3237;
wire net_701;
wire net_397;
wire net_808;
wire net_5553;
wire net_11126;
wire net_7602;
wire net_5595;
wire net_10968;
wire net_9121;
wire net_9894;
wire net_1704;
wire net_12373;
wire net_5026;
wire net_4821;
wire net_1384;
wire net_2738;
wire net_8712;
wire net_3918;
wire net_9107;
wire net_5280;
wire net_320;
wire net_6844;
wire net_4916;
wire net_6902;
wire net_9251;
wire net_2944;
wire net_9103;
wire net_12530;
wire net_7063;
wire net_986;
wire net_12079;
wire net_1242;
wire net_6556;
wire net_14384;
wire net_4346;
wire net_1241;
wire net_13153;
wire net_11953;
wire net_6662;
wire net_3690;
wire net_11176;
wire net_13058;
wire net_9451;
wire net_7927;
wire net_7524;
wire net_11833;
wire net_11019;
wire net_13998;
wire net_13197;
wire net_5654;
wire net_13034;
wire net_8827;
wire net_935;
wire net_3001;
wire net_1511;
wire net_3116;
wire net_645;
wire net_11436;
wire net_3121;
wire net_10368;
wire net_4841;
wire net_4621;
wire net_10289;
wire net_10217;
wire net_4071;
wire net_1634;
wire net_10305;
wire net_6271;
wire net_609;
wire net_12034;
wire net_13343;
wire x1406;
wire net_14242;
wire net_8825;
wire net_10862;
wire net_6155;
wire net_3083;
wire net_5693;
wire net_4533;
wire net_1816;
wire net_9782;
wire net_8076;
wire net_1221;
wire net_7909;
wire net_7158;
wire net_4195;
wire net_14085;
wire net_6911;
wire net_4895;
wire net_9851;
wire net_331;
wire x390;
wire net_12597;
wire net_816;
wire net_9100;
wire net_4644;
wire net_3264;
wire net_7363;
wire net_2092;
wire net_13209;
wire net_8633;
wire net_7134;
wire net_12745;
wire net_8669;
wire net_2220;
wire net_4762;
wire net_2823;
wire net_1217;
wire net_13879;
wire net_7028;
wire net_9719;
wire net_2933;
wire net_3728;
wire net_8141;
wire net_3381;
wire net_10818;
wire net_14156;
wire net_8848;
wire net_5724;
wire net_7138;
wire net_4118;
wire net_4577;
wire net_4970;
wire net_1575;
wire net_4884;
wire net_3279;
wire net_12981;
wire net_657;
wire net_8000;
wire net_8495;
wire net_5042;
wire net_1727;
wire net_12541;
wire net_13808;
wire net_14333;
wire net_12841;
wire net_12199;
wire net_329;
wire net_5809;
wire net_4600;
wire net_4753;
wire net_1259;
wire net_12848;
wire net_11207;
wire net_1924;
wire net_4225;
wire net_2143;
wire net_2839;
wire net_4287;
wire net_1825;
wire net_2196;
wire net_3791;
wire net_7676;
wire net_3168;
wire net_8059;
wire net_10478;
wire net_10078;
wire net_10558;
wire net_11611;
wire net_5275;
wire net_962;
wire net_7914;
wire net_478;
wire net_8695;
wire x179;
wire net_13731;
wire net_7817;
wire net_596;
wire net_11429;
wire net_6608;
wire net_11840;
wire net_1261;
wire net_8733;
wire net_5781;
wire net_4959;
wire net_2120;
wire net_1975;
wire net_4705;
wire net_10430;
wire net_14167;
wire net_8958;
wire net_8375;
wire net_7566;
wire net_13512;
wire net_13067;
wire net_11948;
wire net_13991;
wire net_12893;
wire net_565;
wire net_2569;
wire net_5600;
wire net_7406;
wire net_2832;
wire net_7530;
wire net_4478;
wire net_7253;
wire net_2149;
wire net_3028;
wire net_11281;
wire net_7087;
wire net_1692;
wire net_13174;
wire net_9736;
wire net_12675;
wire net_5079;
wire net_2528;
wire net_2655;
wire net_10611;
wire net_10363;
wire net_5062;
wire net_10854;
wire net_9682;
wire net_6518;
wire net_4236;
wire net_11618;
wire net_1361;
wire net_2450;
wire net_4813;
wire net_9260;
wire net_14118;
wire net_1208;
wire net_10986;
wire net_7948;
wire net_232;
wire net_8920;
wire net_6538;
wire net_14273;
wire net_13201;
wire net_12162;
wire net_13769;
wire net_8560;
wire net_9279;
wire net_12954;
wire net_12778;
wire net_2167;
wire net_2880;
wire net_7923;
wire net_11062;
wire net_13378;
wire net_4710;
wire net_13810;
wire net_4808;
wire net_2996;
wire net_5506;
wire net_2889;
wire net_9537;
wire net_4544;
wire net_7340;
wire net_13901;
wire net_12187;
wire net_137;
wire net_6398;
wire net_3154;
wire net_6386;
wire net_4828;
wire x1511;
wire net_4465;
wire net_532;
wire net_2501;
wire net_3530;
wire net_13179;
wire net_9862;
wire net_13190;
wire net_3622;
wire net_10398;
wire net_9800;
wire net_10389;
wire net_2729;
wire net_4422;
wire net_10116;
wire net_302;
wire net_8223;
wire net_1131;
wire net_889;
wire net_12609;
wire net_1116;
wire net_13018;
wire net_753;
wire net_9034;
wire net_5253;
wire net_5575;
wire net_4373;
wire net_13135;
wire net_9289;
wire net_9710;
wire net_11521;
wire net_2814;
wire x114;
wire net_13609;
wire net_12464;
wire net_689;
wire net_751;
wire net_8084;
wire net_4155;
wire x249;
wire net_13864;
wire net_11297;
wire net_6353;
wire net_6722;
wire net_8288;
wire net_2363;
wire net_14346;
wire net_6283;
wire net_12861;
wire net_3659;
wire net_6578;
wire net_5232;
wire net_5192;
wire net_13708;
wire net_10512;
wire net_3724;
wire net_13129;
wire net_12301;
wire net_13268;
wire net_1228;
wire net_10146;
wire net_7148;
wire net_4593;
wire net_7807;
wire net_13092;
wire net_2722;
wire net_9891;
wire net_12139;
wire net_1426;
wire net_12649;
wire net_9399;
wire net_6504;
wire net_11111;
wire net_12013;
wire net_8531;
wire net_13113;
wire net_9813;
wire net_1407;
wire net_3147;
wire net_4903;
wire net_11548;
wire net_8536;
wire net_11380;
wire net_5409;
wire net_12949;
wire net_13602;
wire net_11795;
wire net_3263;
wire net_10093;
wire net_1057;
wire net_2915;
wire net_14129;
wire net_7235;
wire net_10895;
wire net_5225;
wire net_4931;
wire net_6161;
wire net_6953;
wire net_10647;
wire net_2987;
wire net_10509;
wire net_7261;
wire net_8613;
wire net_8233;
wire net_2253;
wire net_6189;
wire net_1699;
wire net_5114;
wire net_4398;
wire net_9534;
wire net_1042;
wire net_4783;
wire net_4076;
wire net_4792;
wire net_12944;
wire net_7788;
wire net_13267;
wire net_1000;
wire net_11309;
wire net_11133;
wire net_1995;
wire net_2521;
wire net_12915;
wire net_6246;
wire net_11296;
wire net_2545;
wire net_1016;
wire net_6437;
wire net_9035;
wire net_5158;
wire net_11315;
wire net_10017;
wire net_10323;
wire net_3977;
wire net_4567;
wire net_10417;
wire net_10201;
wire net_1744;
wire net_516;
wire net_2870;
wire net_3176;
wire net_3585;
wire net_12655;
wire net_11776;
wire net_12614;
wire net_6182;
wire net_956;
wire net_4320;
wire net_3963;
wire net_11847;
wire net_5799;
wire net_14383;
wire net_2596;
wire net_5496;
wire net_10835;
wire net_2970;
wire net_14388;
wire net_12369;
wire net_438;
wire net_8181;
wire net_8178;
wire net_14001;
wire net_9001;
wire net_2584;
wire net_14052;
wire net_12334;
wire net_2250;
wire net_5278;
wire net_3013;
wire net_5438;
wire net_13826;
wire net_7546;
wire net_11963;
wire net_952;
wire net_3110;
wire net_2967;
wire net_14305;
wire net_4097;
wire net_11743;
wire net_5170;
wire net_3185;
wire net_13821;
wire net_10916;
wire net_8214;
wire net_14290;
wire net_13337;
wire net_9048;
wire net_7598;
wire net_3300;
wire net_6808;
wire net_6438;
wire net_2245;
wire net_10645;
wire net_13185;
wire net_7268;
wire net_12963;
wire net_8187;
wire net_7570;
wire net_13773;
wire net_4231;
wire net_383;
wire net_4068;
wire net_3570;
wire net_14055;
wire net_3140;
wire net_5916;
wire net_6765;
wire net_9773;
wire net_427;
wire net_7823;
wire net_135;
wire net_2785;
wire net_9693;
wire net_10840;
wire net_1121;
wire net_8575;
wire net_13169;
wire net_8274;
wire net_473;
wire net_13687;
wire net_7288;
wire net_13897;
wire net_7559;
wire net_3599;
wire net_7381;
wire net_5099;
wire net_9512;
wire net_8350;
wire net_4329;
wire net_11094;
wire net_6409;
wire net_2777;
wire net_1049;
wire net_13531;
wire net_9440;
wire net_454;
wire net_3901;
wire net_6251;
wire net_5349;
wire net_10674;
wire net_9364;
wire net_6707;
wire net_709;
wire net_2484;
wire net_8437;
wire net_13535;
wire net_9278;
wire net_7582;
wire net_11342;
wire net_6229;
wire net_8608;
wire net_10791;
wire net_5199;
wire net_12905;
wire net_1066;
wire net_5514;
wire net_12388;
wire net_9293;
wire net_9956;
wire net_2591;
wire net_4304;
wire net_10552;
wire net_8985;
wire net_10880;
wire net_5847;
wire net_5189;
wire net_11896;
wire net_4560;
wire net_1344;
wire net_5791;
wire net_1283;
wire net_1084;
wire net_3968;
wire net_12875;
wire net_4554;
wire net_1500;
wire net_354;
wire net_9778;
wire net_11376;
wire net_1136;
wire net_14010;
wire net_12428;
wire net_5418;
wire net_3008;
wire net_11707;
wire net_2763;
wire net_573;
wire net_12099;
wire net_9065;
wire net_3356;
wire net_12412;
wire net_11423;
wire net_7175;
wire net_5465;
wire net_6855;
wire net_13314;
wire net_12640;
wire net_11606;
wire net_3616;
wire net_9494;
wire net_3886;
wire net_7281;
wire net_1592;
wire net_13650;
wire net_2085;
wire net_13352;
wire net_8570;
wire net_5521;
wire net_5037;
wire net_3672;
wire net_11101;
wire net_6089;
wire net_4406;
wire net_9249;
wire net_14371;
wire net_12557;
wire net_5621;
wire net_8764;
wire net_11879;
wire net_10297;
wire net_1637;
wire net_3702;
wire net_9374;
wire net_6480;
wire net_6425;
wire net_5971;
wire net_5811;
wire net_6220;
wire net_8915;
wire net_941;
wire net_7560;
wire net_7629;
wire net_6038;
wire net_11324;
wire net_5854;
wire net_13292;
wire net_14351;
wire net_8129;
wire net_4555;
wire net_2070;
wire net_2311;
wire net_9444;
wire net_11661;
wire net_4611;
wire net_7500;
wire net_10605;
wire net_4124;
wire net_1599;
wire net_6587;
wire net_10575;
wire net_11087;
wire net_12372;
wire net_3828;
wire net_3981;
wire net_13659;
wire net_11504;
wire net_3132;
wire net_3161;
wire net_9973;
wire net_6107;
wire net_4303;
wire net_1290;
wire net_12924;
wire net_4147;
wire net_12240;
wire net_3053;
wire net_9802;
wire net_9579;
wire net_4056;
wire net_7187;
wire net_12589;
wire net_7460;
wire net_3297;
wire net_6601;
wire net_8518;
wire net_2023;
wire net_14028;
wire net_13923;
wire net_4523;
wire net_123;
wire net_11766;
wire net_5249;
wire net_1668;
wire net_527;
wire net_262;
wire net_13474;
wire net_12205;
wire net_3424;
wire net_12151;
wire net_7552;
wire net_6364;
wire net_10169;
wire net_3139;
wire net_5388;
wire net_4063;
wire net_6399;
wire net_5087;
wire net_13218;
wire net_11983;
wire net_1793;
wire net_11714;
wire net_3104;
wire net_3786;
wire net_5508;
wire net_2278;
wire net_8261;
wire net_7161;
wire net_3072;
wire net_6215;
wire net_7286;
wire net_1021;
wire net_10498;
wire net_5269;
wire net_10488;
wire net_1737;
wire net_9979;
wire net_10657;
wire net_5706;
wire net_6801;
wire net_1859;
wire net_12550;
wire net_145;
wire net_3607;
wire net_4654;
wire net_8541;
wire net_4917;
wire net_10699;
wire net_8193;
wire net_1145;
wire net_10431;
wire net_8424;
wire net_4637;
wire net_2804;
wire net_11134;
wire net_9306;
wire net_2261;
wire net_9411;
wire net_5535;
wire net_188;
wire net_3753;
wire net_3061;
wire net_3319;
wire net_4353;
wire net_7414;
wire net_10160;
wire net_7141;
wire net_2958;
wire net_1077;
wire net_14163;
wire net_6520;
wire x1542;
wire net_2924;
wire net_10050;
wire net_8969;
wire net_11328;
wire net_14131;
wire net_12318;
wire net_11825;
wire net_8022;
wire net_5918;
wire net_2410;
wire net_8281;
wire net_10827;
wire net_9208;
wire net_119;
wire net_3108;
wire net_10975;
wire net_10445;
wire net_2185;
wire net_13103;
wire net_6853;
wire net_1321;
wire net_14263;
wire net_13961;
wire net_13624;
wire net_4441;
wire net_6307;
wire net_4192;
wire net_8741;
wire net_5392;
wire net_4949;
wire net_1099;
wire net_11977;
wire net_11733;
wire net_11141;
wire net_11568;
wire net_7106;
wire net_4583;
wire net_7103;
wire net_9885;
wire net_9227;
wire net_12290;
wire net_404;
wire net_11683;
wire net_6033;
wire net_4663;
wire net_14330;
wire net_11624;
wire net_5455;
wire net_9276;
wire net_2666;
wire net_5822;
wire net_4084;
wire net_4500;
wire net_10929;
wire net_8045;
wire net_8402;
wire net_1239;
wire net_10246;
wire net_8663;
wire net_8591;
wire net_5879;
wire net_1463;
wire net_9743;
wire net_14250;
wire net_8793;
wire net_8562;
wire net_12257;
wire net_2056;
wire net_10081;
wire net_5716;
wire net_9266;
wire net_7884;
wire net_3822;
wire net_12217;
wire net_10800;
wire net_9147;
wire net_1628;
wire net_3476;
wire net_13957;
wire net_6872;
wire net_7347;
wire net_484;
wire net_896;
wire net_7655;
wire net_4823;
wire net_12519;
wire net_2512;
wire net_3223;
wire net_12997;
wire net_5894;
wire net_1936;
wire net_11363;
wire net_3802;
wire net_11599;
wire net_10035;
wire net_14339;
wire net_126;
wire net_2708;
wire net_8773;
wire net_8705;
wire net_10088;
wire net_10873;
wire net_9795;
wire net_12971;
wire net_9958;
wire net_2211;
wire net_13106;
wire net_11563;
wire net_7425;
wire net_5479;
wire net_13939;
wire net_11794;
wire net_13001;
wire net_13614;
wire net_11550;
wire net_7917;
wire net_1896;
wire net_14090;
wire net_8388;
wire net_8777;
wire net_9998;
wire net_1732;
wire net_1982;
wire net_13283;
wire net_12687;
wire net_5926;
wire net_8089;
wire net_7866;
wire net_6348;
wire net_12084;
wire net_10014;
wire net_9390;
wire net_11719;
wire net_12149;
wire net_6509;
wire net_12507;
wire net_900;
wire net_3253;
wire net_10630;
wire net_6935;
wire net_13176;
wire net_7597;
wire net_5498;
wire net_1882;
wire net_12347;
wire net_12229;
wire net_12755;
wire net_7744;
wire net_5528;
wire net_413;
wire net_2001;
wire net_11072;
wire net_1491;
wire net_10879;
wire net_9613;
wire net_8306;
wire net_6141;
wire net_10918;
wire net_12666;
wire net_5390;
wire net_7876;
wire net_2419;
wire net_10154;
wire net_1034;
wire net_11559;
wire net_5753;
wire net_7608;
wire net_12203;
wire net_11510;
wire net_14315;
wire net_253;
wire net_11696;
wire net_276;
wire net_9728;
wire net_14229;
wire net_3439;
wire net_12112;
wire net_8470;
wire net_13899;
wire net_13332;
wire net_10586;
wire net_6490;
wire net_13395;
wire net_9799;
wire net_11398;
wire net_1959;
wire net_616;
wire net_1847;
wire net_11506;
wire net_12320;
wire net_2717;
wire net_793;
wire net_9137;
wire net_460;
wire net_7356;
wire net_6797;
wire net_2353;
wire net_6074;
wire net_11919;
wire net_2272;
wire net_9231;
wire net_4206;
wire net_9708;
wire net_1133;
wire net_14222;
wire net_6131;
wire net_4104;
wire net_8133;
wire net_3287;
wire net_11712;
wire net_10724;
wire net_166;
wire net_11305;
wire net_11027;
wire net_2866;
wire net_5866;
wire net_13954;
wire net_5489;
wire net_3025;
wire net_13164;
wire net_3871;
wire net_5407;
wire net_4455;
wire net_7673;
wire net_10995;
wire net_8788;
wire net_3352;
wire net_7507;
wire net_7309;
wire net_10342;
wire net_6071;
wire net_6894;
wire net_3832;
wire net_5663;
wire net_205;
wire net_11702;
wire net_1286;
wire net_6427;
wire net_6017;
wire net_10062;
wire net_11872;
wire net_9764;
wire net_7617;
wire net_7533;
wire net_6925;
wire net_334;
wire net_1952;
wire net_9214;
wire net_10930;
wire net_9846;
wire net_2453;
wire net_3062;
wire net_11495;
wire net_9586;
wire net_5738;
wire net_12512;
wire net_12629;
wire net_4620;
wire net_14141;
wire net_5696;
wire net_380;
wire net_2847;
wire net_10952;
wire net_6515;
wire net_13797;
wire net_7932;
wire net_12626;
wire net_14042;
wire net_12885;
wire net_1556;
wire net_6803;
wire net_5911;
wire net_6790;
wire net_4337;
wire net_13548;
wire net_3768;
wire net_7976;
wire net_4745;
wire x1286;
wire net_1270;
wire net_4905;
wire net_2286;
wire net_14178;
wire net_9717;
wire net_1552;
wire net_13785;
wire net_9380;
wire net_14015;
wire net_6094;
wire net_7712;
wire net_4940;
wire net_3878;
wire net_5674;
wire net_7954;
wire net_8132;
wire net_5585;
wire net_3215;
wire net_1933;
wire net_298;
wire net_3717;
wire net_3241;
wire net_998;
wire net_12620;
wire net_4657;
wire net_2157;
wire net_8945;
wire net_7273;
wire net_2555;
wire net_10317;
wire net_4864;
wire net_11154;
wire net_13148;
wire net_12457;
wire net_9328;
wire net_3504;
wire net_13763;
wire net_14194;
wire net_2405;
wire net_1687;
wire net_835;
wire net_7459;
wire net_5243;
wire net_1762;
wire net_7407;
wire net_13683;
wire net_1181;
wire net_9321;
wire net_10685;
wire net_10466;
wire net_6459;
wire net_638;
wire net_12299;
wire net_7472;
wire net_932;
wire net_313;
wire net_5633;
wire net_6082;
wire net_10028;
wire net_5766;
wire net_11519;
wire net_13403;
wire net_10783;
wire net_12488;
wire net_12801;
wire net_4767;
wire net_1783;
wire net_14257;
wire net_5271;
wire net_12814;
wire net_6771;
wire net_7771;
wire net_1874;
wire net_9554;
wire net_7769;
wire net_972;
wire net_14308;
wire net_9650;
wire net_3499;
wire net_5206;
wire net_4725;
wire net_4777;
wire net_14292;
wire net_13192;
wire net_11669;
wire net_6201;
wire net_14108;
wire net_12808;
wire net_785;
wire net_7047;
wire net_9152;
wire net_1489;
wire net_13665;
wire net_5883;
wire net_4343;
wire net_4215;
wire net_10276;
wire net_9874;
wire net_6677;
wire net_10902;
wire net_13633;
wire net_10409;
wire net_9657;
wire net_7479;
wire net_3746;
wire net_1349;
wire net_7794;
wire net_7194;
wire net_979;
wire net_2392;
wire net_156;
wire net_13251;
wire net_11820;
wire net_10278;
wire net_12563;
wire net_2015;
wire net_8441;
wire net_6658;
wire net_13064;
wire net_10266;
wire net_5947;
wire net_1040;
wire net_9676;
wire net_8978;
wire net_5202;
wire net_4877;
wire net_6781;
wire net_4170;
wire net_3089;
wire net_3101;
wire net_12336;
wire net_6268;
wire net_3037;
wire net_4472;
wire net_12723;
wire net_7331;
wire net_4463;
wire net_3876;
wire net_5982;
wire net_2907;
wire net_3686;
wire net_1887;
wire net_13146;
wire net_7444;
wire net_5470;
wire net_379;
wire net_2243;
wire net_1569;
wire net_4033;
wire net_4245;
wire net_11868;
wire net_9514;
wire net_7795;
wire net_3133;
wire net_5568;
wire net_3047;
wire net_2559;
wire net_8910;
wire net_9532;
wire net_6944;
wire net_6883;
wire net_2657;
wire net_1358;
wire net_8477;
wire net_6815;
wire net_12259;
wire net_11438;
wire net_8415;
wire net_7742;
wire net_2629;
wire net_2486;
wire net_11405;
wire net_6888;
wire net_8927;
wire net_8421;
wire net_7117;
wire net_1206;
wire net_8381;
wire net_3653;
wire net_960;
wire net_13494;
wire net_3704;
wire net_1166;
wire net_10706;
wire net_8155;
wire net_10765;
wire net_801;
wire net_11051;
wire net_2620;
wire net_14062;
wire net_7450;
wire net_1718;
wire net_2581;
wire net_5093;
wire net_12842;
wire net_13365;
wire net_9417;
wire net_7372;
wire net_13996;
wire net_9445;
wire net_6441;
wire net_4348;
wire net_4526;
wire net_11921;
wire net_10391;
wire net_8482;
wire net_2129;
wire net_7832;
wire net_5968;
wire x718;
wire net_6234;
wire net_9909;
wire net_8991;
wire net_581;
wire net_10564;
wire net_13967;
wire net_8799;
wire net_2899;
wire net_9833;
wire net_8856;
wire net_12421;
wire net_9609;
wire net_11382;
wire net_658;
wire net_7115;
wire net_5906;
wire net_7978;
wire net_11391;
wire net_8462;
wire net_13529;
wire net_2090;
wire net_9540;
wire net_7723;
wire net_12509;
wire net_2325;
wire net_8807;
wire net_13715;
wire net_12758;
wire net_806;
wire net_10259;
wire net_11907;
wire net_5801;
wire net_9901;
wire net_8940;
wire net_4021;
wire net_8999;
wire net_7026;
wire net_10960;
wire net_5461;
wire net_946;
wire net_1176;
wire net_2676;
wire net_6372;
wire net_7032;
wire net_4989;
wire net_2194;
wire net_11609;
wire net_1751;
wire net_13593;
wire net_5010;
wire net_3559;
wire net_8370;
wire net_4682;
wire net_6733;
wire net_10114;
wire net_3508;
wire net_10402;
wire net_12499;
wire net_10732;
wire net_2434;
wire net_3564;
wire net_1448;
wire net_2032;
wire net_392;
wire net_118;
wire net_2467;
wire net_5683;
wire net_11524;
wire net_7003;
wire net_2452;
wire net_14415;
wire net_11463;
wire net_9916;
wire net_12008;
wire net_10336;
wire net_3523;
wire net_4162;
wire net_5549;
wire net_3712;
wire net_6680;
wire net_8865;
wire net_7223;
wire net_6613;
wire net_246;
wire net_1186;
wire net_4747;
wire net_11269;
wire net_13041;
wire net_7074;
wire net_10607;
wire net_10437;
wire net_13436;
wire net_10121;
wire net_2216;
wire net_10410;
wire net_8968;
wire net_6725;
wire net_1378;
wire net_7399;
wire net_1773;
wire net_3773;
wire net_9057;
wire net_1600;
wire net_2531;
wire net_12440;
wire net_11971;
wire net_8731;
wire net_676;
wire net_11254;
wire net_12492;
wire net_6626;
wire net_4263;
wire net_5073;
wire net_2538;
wire net_4452;
wire net_2447;
wire net_7433;
wire net_5133;
wire net_5542;
wire net_14116;
wire net_5417;
wire net_5370;
wire net_4260;
wire net_3492;
wire net_8137;
wire net_6010;
wire net_182;
wire net_2462;
wire net_4359;
wire net_12760;
wire net_9635;
wire net_9018;
wire net_11260;
wire net_8820;
wire net_3324;
wire net_13485;
wire net_9547;
wire net_5426;
wire net_6450;
wire net_6138;
wire net_14237;
wire net_8398;
wire net_6979;
wire net_11442;
wire net_7893;
wire net_1435;
wire net_1370;
wire net_9600;
wire net_10429;
wire net_8112;
wire net_11274;
wire net_9462;
wire net_7939;
wire net_3568;
wire net_3207;
wire net_13920;
wire net_7810;
wire net_4482;
wire net_6470;
wire net_2204;
wire net_9668;
wire net_5088;
wire net_8459;
wire net_2492;
wire net_11188;
wire net_9088;
wire net_1970;
wire net_1306;
wire net_4045;
wire net_3843;
wire net_1858;
wire net_10223;
wire net_7635;
wire net_6543;
wire net_11005;
wire net_3038;
wire net_13560;
wire net_2690;
wire net_11332;
wire net_7016;
wire net_3924;
wire net_9825;
wire net_11196;
wire net_5226;
wire net_12242;
wire net_791;
wire net_14207;
wire net_10230;
wire net_9422;
wire net_1419;
wire net_3239;
wire net_8554;
wire net_2188;
wire net_8811;
wire net_10546;
wire net_1051;
wire net_12064;
wire net_13882;
wire net_10386;
wire net_10048;
wire net_7644;
wire net_11034;
wire net_7858;
wire net_7410;
wire net_12471;
wire net_1515;
wire net_1573;
wire net_10356;
wire net_7669;
wire net_7219;
wire net_13272;
wire net_6869;
wire net_4983;
wire net_6824;
wire net_361;
wire net_13932;
wire net_2890;
wire net_11547;
wire net_9984;
wire net_7100;
wire net_305;
wire net_4208;
wire net_4515;
wire net_1905;
wire net_12433;
wire net_2540;
wire net_12016;
wire net_12452;
wire net_9166;
wire net_1125;
wire net_2230;
wire net_10195;
wire net_227;
wire net_144;
wire net_13758;
wire net_4183;
wire net_10667;
wire net_10237;
wire net_3592;
wire net_5961;
wire net_13728;
wire net_12405;
wire net_12543;
wire net_6687;
wire net_8818;
wire net_13592;
wire net_7156;
wire net_14413;
wire net_12636;
wire net_4969;
wire net_9175;
wire net_1415;
wire net_3485;
wire net_7052;
wire net_8859;
wire net_6379;
wire net_2886;
wire net_3317;
wire net_14408;
wire net_11746;
wire net_8140;
wire net_1921;
wire net_11638;
wire net_10945;
wire net_9161;
wire net_3853;
wire net_9962;
wire net_10120;
wire net_11910;
wire net_9091;
wire net_1230;
wire net_2135;
wire net_667;
wire net_853;
wire net_212;
wire net_12265;
wire net_9508;
wire net_6047;
wire net_914;
wire net_10254;
wire net_9923;
wire net_12835;
wire net_6862;
wire net_6320;
wire net_6064;
wire net_6448;
wire x149;
wire net_875;
wire net_5619;
wire net_1092;
wire net_12046;
wire net_7585;
wire net_627;
wire net_10597;
wire net_8759;
wire net_2039;
wire net_11579;
wire net_12067;
wire net_1456;
wire net_9198;
wire net_11042;
wire net_2227;
wire net_5636;
wire net_10280;
wire net_8876;
wire net_12231;
wire net_2473;
wire net_6968;
wire net_399;
wire net_8107;
wire net_11041;
wire net_5949;
wire net_5069;
wire net_13509;
wire net_13844;
wire net_10678;
wire net_8752;
wire net_1390;
wire net_11209;
wire net_7180;
wire net_5565;
wire net_218;
wire net_12338;
wire net_10517;
wire net_7110;
wire net_1112;
wire net_9335;
wire net_5173;
wire net_1273;
wire net_3283;
wire net_10747;
wire net_9025;
wire net_4433;
wire net_13907;
wire net_11995;
wire net_8146;
wire net_5449;
wire net_2114;
wire net_2506;
wire net_11200;
wire net_12085;
wire net_5012;
wire net_9644;
wire net_3230;
wire net_13295;
wire net_7124;
wire net_11235;
wire net_11990;
wire net_10187;
wire net_14073;
wire net_285;
wire net_8316;
wire net_13585;
wire net_11486;
wire net_5677;
wire net_5296;
wire net_14171;
wire net_1310;
wire net_9634;
wire net_2499;
wire net_6057;
wire net_11567;
wire net_1297;
wire net_7579;
wire net_1304;
wire net_9471;
wire net_8901;
wire net_4381;
wire net_2177;
wire net_11918;
wire net_11378;
wire net_6674;
wire net_13427;
wire net_7863;
wire net_11450;
wire net_11587;
wire net_6581;
wire net_6916;
wire net_10370;
wire net_6127;
wire net_5030;
wire net_13417;
wire net_6058;
wire net_10919;
wire net_2449;
wire net_6070;
wire net_1317;
wire net_6588;
wire net_215;
wire net_416;
wire net_2394;
wire net_1382;
wire net_5629;
wire net_11593;
wire net_13408;
wire net_6896;
wire net_6442;
wire net_4508;
wire net_6642;
wire net_10760;
wire net_3498;
wire net_8093;
wire net_1377;
wire net_1786;
wire net_12831;
wire net_5620;
wire net_13580;
wire net_12031;
wire net_10253;
wire net_4513;
wire net_14025;
wire net_10940;
wire net_9658;
wire net_5965;
wire net_13428;
wire net_11118;
wire net_5586;
wire net_5430;
wire net_5954;
wire net_1393;
wire net_13724;
wire net_14321;
wire net_2169;
wire net_6119;
wire net_8758;
wire net_1324;
wire net_14020;
wire net_9960;
wire net_7114;
wire net_12058;
wire net_10672;
wire net_10476;
wire net_8017;
wire net_2207;
wire net_263;
wire net_6997;
wire net_9336;
wire net_4323;
wire net_8805;
wire net_1138;
wire net_3527;
wire net_8509;
wire net_14139;
wire net_3483;
wire net_6838;
wire net_10167;
wire net_10548;
wire net_1439;
wire net_3292;
wire net_8714;
wire net_12528;
wire net_13489;
wire net_9700;
wire net_508;
wire net_1778;
wire net_4189;
wire net_9256;
wire net_1090;
wire net_5098;
wire net_6907;
wire net_7438;
wire net_3685;
wire net_5355;
wire net_7030;
wire net_8149;
wire net_7012;
wire net_14107;
wire net_11962;
wire net_11453;
wire net_9007;
wire net_4285;
wire net_8643;
wire net_4434;
wire net_5413;
wire net_12068;
wire net_4744;
wire net_10726;
wire net_201;
wire net_5077;
wire net_9496;
wire net_6636;
wire net_3280;
wire net_9666;
wire net_3085;
wire net_4043;
wire net_2896;
wire net_8371;
wire net_4258;
wire net_7443;
wire net_12838;
wire net_12631;
wire net_12207;
wire net_12454;
wire net_13833;
wire net_9985;
wire net_1852;
wire net_11236;
wire net_11912;
wire net_9515;
wire net_6129;
wire net_1555;
wire net_7301;
wire net_10594;
wire net_2780;
wire net_9349;
wire net_4480;
wire net_789;
wire net_10131;
wire net_10769;
wire net_3244;
wire net_12819;
wire net_9041;
wire net_2171;
wire net_12080;
wire net_10233;
wire net_3833;
wire net_6338;
wire net_9967;
wire net_8664;
wire net_7256;
wire net_4521;
wire net_11245;
wire net_2425;
wire net_6112;
wire net_13691;
wire net_8319;
wire net_10573;
wire net_2509;
wire net_8143;
wire net_5137;
wire net_11569;
wire net_1860;
wire net_2156;
wire net_8025;
wire net_1432;
wire net_1312;
wire net_9474;
wire net_9177;
wire net_5463;
wire net_14188;
wire net_8843;
wire net_8488;
wire net_8435;
wire net_4801;
wire net_13246;
wire net_6831;
wire net_5334;
wire net_4314;
wire net_5290;
wire net_11640;
wire net_10005;
wire net_3343;
wire net_3546;
wire net_3326;
wire net_8002;
wire net_11877;
wire net_1453;
wire net_14328;
wire net_13802;
wire net_2239;
wire net_13075;
wire net_9603;
wire net_3394;
wire net_3542;
wire net_634;
wire net_5374;
wire net_8516;
wire net_14177;
wire net_12846;
wire net_9630;
wire net_4680;
wire net_8055;
wire net_14066;
wire net_371;
wire net_13786;
wire net_3903;
wire net_7752;
wire net_2787;
wire net_8879;
wire net_4050;
wire net_1571;
wire net_11467;
wire net_9248;
wire net_2466;
wire net_4904;
wire net_8580;
wire net_4699;
wire net_7710;
wire net_5090;
wire net_7975;
wire net_8872;
wire net_10530;
wire net_7574;
wire net_13921;
wire net_850;
wire net_5217;
wire net_12511;
wire net_679;
wire net_1168;
wire net_2680;
wire net_8116;
wire net_8924;
wire net_308;
wire net_10118;
wire net_11008;
wire net_12218;
wire net_9631;
wire net_5545;
wire net_10744;
wire net_6327;
wire net_3090;
wire net_8747;
wire net_8387;
wire net_1009;
wire net_715;
wire net_11444;
wire net_890;
wire net_13857;
wire net_8454;
wire net_11181;
wire net_2546;
wire net_7228;
wire net_12042;
wire net_7056;
wire net_9019;
wire net_13401;
wire net_9162;
wire net_13646;
wire net_13595;
wire net_2471;
wire net_6702;
wire net_11130;
wire net_312;
wire net_2404;
wire net_2627;
wire net_5386;
wire net_147;
wire net_481;
wire net_12490;
wire net_7182;
wire net_5346;
wire net_8589;
wire net_12137;
wire net_12335;
wire net_7750;
wire net_2444;
wire net_6891;
wire net_11482;
wire net_13496;
wire net_1188;
wire net_13855;
wire net_12936;
wire net_5297;
wire net_8148;
wire net_9625;
wire net_1446;
wire net_10122;
wire net_541;
wire net_8551;
wire net_13380;
wire net_1251;
wire net_8157;
wire net_14148;
wire net_10759;
wire net_8830;
wire net_1697;
wire net_4222;
wire net_7431;
wire net_12238;
wire net_1753;
wire net_4163;
wire net_5398;
wire net_5548;
wire net_245;
wire net_2435;
wire net_6990;
wire net_2383;
wire net_4858;
wire net_14298;
wire net_12177;
wire net_4264;
wire net_11013;
wire net_9749;
wire net_3491;
wire net_10829;
wire net_8380;
wire net_9908;
wire net_277;
wire net_1965;
wire net_4251;
wire net_11418;
wire net_7525;
wire net_13886;
wire net_3071;
wire net_8611;
wire net_680;
wire net_14238;
wire net_10925;
wire net_9568;
wire net_13435;
wire net_13230;
wire net_338;
wire net_7149;
wire net_9994;
wire net_4494;
wire net_7619;
wire net_8397;
wire net_2998;
wire net_243;
wire net_9971;
wire net_8905;
wire net_10705;
wire net_4089;
wire net_6882;
wire net_13721;
wire net_2854;
wire net_2009;
wire net_10730;
wire net_8867;
wire net_4026;
wire net_4132;
wire net_8925;
wire net_6697;
wire net_4990;
wire net_1380;
wire net_7721;
wire net_9292;
wire net_11056;
wire net_13588;
wire net_8326;
wire net_9340;
wire net_1915;
wire net_5176;
wire net_13566;
wire net_10992;
wire net_8280;
wire net_4334;
wire net_5936;
wire net_11956;
wire net_8937;
wire net_6987;
wire net_1997;
wire net_13206;
wire net_12738;
wire net_13779;
wire net_138;
wire net_12497;
wire net_7718;
wire net_13607;
wire net_8553;
wire net_6728;
wire net_13698;
wire net_13364;
wire net_11139;
wire net_9195;
wire net_12714;
wire net_14151;
wire net_7164;
wire net_12313;
wire net_6579;
wire net_9670;
wire net_7633;
wire net_1418;
wire net_13955;
wire net_8686;
wire net_13393;
wire net_5938;
wire net_8994;
wire net_3202;
wire net_13422;
wire net_8343;
wire net_4059;
wire net_5931;
wire net_6980;
wire net_6376;
wire net_6736;
wire net_7461;
wire net_12913;
wire net_1713;
wire net_10380;
wire net_5612;
wire net_2668;
wire net_4684;
wire net_13480;
wire net_11383;
wire net_2677;
wire net_8988;
wire net_10415;
wire net_2775;
wire x1527;
wire net_7001;
wire net_11540;
wire net_12007;
wire net_11741;
wire net_3916;
wire net_7654;
wire net_163;
wire net_6852;
wire net_6022;
wire net_8312;
wire net_5802;
wire net_13937;
wire net_11037;
wire net_8037;
wire net_12590;
wire net_9830;
wire net_8444;
wire net_5900;
wire net_6206;
wire net_13863;
wire net_11580;
wire net_6135;
wire net_3990;
wire net_12595;
wire net_2193;
wire net_12293;
wire net_12002;
wire net_11159;
wire net_10221;
wire net_3856;
wire net_9210;
wire net_5345;
wire net_6304;
wire net_8363;
wire net_4885;
wire net_11704;
wire net_5574;
wire net_5258;
wire net_1886;
wire net_2604;
wire net_3501;
wire net_13689;
wire net_14115;
wire net_12191;
wire net_7862;
wire net_12775;
wire net_4678;
wire net_14307;
wire net_6678;
wire net_7916;
wire net_14256;
wire net_13600;
wire net_4866;
wire net_5652;
wire net_8081;
wire net_13982;
wire net_14013;
wire net_8835;
wire net_1272;
wire net_1770;
wire net_2109;
wire net_10273;
wire net_3505;
wire net_4001;
wire net_5059;
wire net_655;
wire net_9326;
wire net_3536;
wire net_6878;
wire net_4703;
wire net_8534;
wire net_10059;
wire net_4770;
wire net_12961;
wire net_14049;
wire net_378;
wire net_7770;
wire net_14262;
wire net_9110;
wire net_3309;
wire net_14403;
wire net_5767;
wire net_423;
wire net_3036;
wire net_10032;
wire net_11628;
wire net_328;
wire net_4202;
wire net_10103;
wire net_10565;
wire net_1958;
wire net_7934;
wire net_1931;
wire net_7977;
wire net_9060;
wire net_14041;
wire net_3294;
wire net_1549;
wire net_6244;
wire net_10039;
wire net_3016;
wire net_4477;
wire net_7736;
wire net_2929;
wire net_7192;
wire net_12933;
wire net_9117;
wire net_7213;
wire net_5666;
wire net_11717;
wire net_11227;
wire net_8527;
wire net_818;
wire net_3749;
wire net_11275;
wire net_2746;
wire net_12592;
wire net_9403;
wire net_1211;
wire net_5024;
wire net_1183;
wire net_5448;
wire net_11863;
wire net_2594;
wire net_4248;
wire net_12337;
wire net_5944;
wire net_811;
wire net_1684;
wire net_7241;
wire net_9753;
wire net_1462;
wire net_9551;
wire net_9203;
wire net_4674;
wire net_2017;
wire net_6791;
wire net_9150;
wire net_4993;
wire net_5154;
wire net_11508;
wire net_1926;
wire net_12145;
wire net_2735;
wire net_3115;
wire net_8780;
wire net_14158;
wire net_8377;
wire net_3518;
wire net_13069;
wire x1209;
wire net_10261;
wire net_8800;
wire net_1621;
wire net_3680;
wire net_6926;
wire net_14319;
wire net_3984;
wire net_13317;
wire net_3615;
wire net_1035;
wire net_12253;
wire net_11331;
wire net_9559;
wire net_14076;
wire net_13172;
wire net_3055;
wire net_9844;
wire net_13035;
wire net_5597;
wire net_6914;
wire net_4656;
wire net_10264;
wire net_3593;
wire net_2845;
wire net_3095;
wire net_6510;
wire net_12585;
wire net_11358;
wire net_4586;
wire net_6748;
wire net_2641;
wire net_7711;
wire net_6688;
wire net_13141;
wire net_9389;
wire net_1763;
wire net_6168;
wire net_7291;
wire net_12321;
wire net_11067;
wire net_4035;
wire net_9362;
wire net_7816;
wire net_12999;
wire net_9881;
wire net_8948;
wire net_13464;
wire net_9092;
wire net_7919;
wire net_2882;
wire net_8131;
wire net_3278;
wire net_12277;
wire net_4386;
wire net_8837;
wire net_1513;
wire net_14191;
wire net_14253;
wire net_10668;
wire net_3064;
wire net_5731;
wire net_12701;
wire net_2276;
wire net_12748;
wire net_4613;
wire net_6369;
wire net_9302;
wire net_11639;
wire net_7763;
wire net_7748;
wire net_11388;
wire net_9426;
wire net_6745;
wire net_10084;
wire net_13716;
wire net_14149;
wire net_798;
wire net_3135;
wire net_5266;
wire net_5165;
wire net_2059;
wire net_8473;
wire net_9740;
wire net_8520;
wire net_8860;
wire net_8209;
wire net_1899;
wire net_6018;
wire net_8890;
wire net_1336;
wire net_4746;
wire net_12198;
wire net_9915;
wire net_10033;
wire net_1843;
wire net_6031;
wire net_11739;
wire net_6946;
wire net_12211;
wire net_7019;
wire net_534;
wire net_14114;
wire net_11534;
wire net_3793;
wire net_9261;
wire net_13523;
wire net_11671;
wire net_8659;
wire net_6823;
wire net_3336;
wire net_9561;
wire net_903;
wire net_1551;
wire net_10025;
wire net_12069;
wire net_486;
wire net_13796;
wire net_12898;
wire net_406;
wire net_11395;
wire net_8407;
wire net_7354;
wire net_5986;
wire net_4190;
wire net_2378;
wire net_5391;
wire net_12448;
wire net_11758;
wire net_10461;
wire net_6261;
wire net_8967;
wire net_10319;
wire net_8046;
wire net_13746;
wire net_7125;
wire net_3640;
wire net_748;
wire net_9865;
wire net_8605;
wire net_10587;
wire net_10010;
wire net_5566;
wire net_6917;
wire net_13124;
wire net_10778;
wire net_3958;
wire net_5281;
wire net_12270;
wire net_8776;
wire net_5427;
wire net_11621;
wire net_11684;
wire net_10868;
wire net_8772;
wire net_1003;
wire net_2327;
wire net_514;
wire net_11255;
wire net_3645;
wire net_7376;
wire net_10310;
wire net_1604;
wire net_6499;
wire net_5755;
wire net_14093;
wire net_5669;
wire net_6122;
wire net_524;
wire net_6497;
wire net_13387;
wire net_11991;
wire net_6060;
wire net_13816;
wire net_13554;
wire net_11513;
wire net_3742;
wire net_445;
wire net_4368;
wire net_7109;
wire net_13398;
wire net_13002;
wire net_10773;
wire net_6673;
wire net_3748;
wire net_12319;
wire net_13637;
wire net_10786;
wire net_9355;
wire net_8307;
wire net_2213;
wire net_12083;
wire net_2575;
wire net_5067;
wire net_11986;
wire net_10935;
wire net_1097;
wire net_11756;
wire net_12227;
wire net_14172;
wire net_9219;
wire net_12142;
wire net_762;
wire net_6921;
wire net_3589;
wire net_8445;
wire net_13517;
wire net_4943;
wire net_10876;
wire net_3713;
wire net_8400;
wire net_556;
wire net_6173;
wire net_893;
wire net_3330;
wire net_11163;
wire net_4121;
wire net_255;
wire net_3826;
wire net_620;
wire net_9641;
wire net_619;
wire net_13618;
wire net_9085;
wire net_8702;
wire net_4659;
wire net_7321;
wire net_3932;
wire net_7233;
wire net_14392;
wire net_11177;
wire net_4779;
wire net_5997;
wire net_11150;
wire net_7689;
wire net_8156;
wire net_5129;
wire net_7104;
wire net_10444;
wire net_7883;
wire net_3444;
wire net_4922;
wire net_6414;
wire net_3800;
wire net_5393;
wire net_3285;
wire net_6937;
wire net_7278;
wire net_7825;
wire net_4425;
wire net_4933;
wire net_5834;
wire net_4044;
wire net_13613;
wire net_8855;
wire net_11300;
wire net_1493;
wire net_9167;
wire net_13285;
wire net_11699;
wire net_5875;
wire net_4630;
wire net_11143;
wire net_976;
wire net_6287;
wire net_8498;
wire net_2709;
wire net_5309;
wire net_10321;
wire net_11630;
wire net_8897;
wire net_611;
wire net_7879;
wire net_2579;
wire net_3514;
wire net_4179;
wire net_5441;
wire net_8235;
wire net_9581;
wire net_10296;
wire net_6013;
wire net_7307;
wire net_5873;
wire net_12990;
wire net_1866;
wire net_6077;
wire net_10849;
wire net_4907;
wire net_6567;
wire net_4107;
wire net_6934;
wire net_5761;
wire net_2160;
wire net_3211;
wire net_3692;
wire net_13060;
wire net_10820;
wire net_3477;
wire net_391;
wire net_6361;
wire net_9268;
wire net_9723;
wire net_5927;
wire net_7634;
wire net_5040;
wire net_13894;
wire net_11738;
wire net_12754;
wire net_8625;
wire net_5820;
wire net_6692;
wire net_4172;
wire net_11732;
wire net_8342;
wire net_2516;
wire net_13892;
wire net_8123;
wire net_2807;
wire net_7553;
wire net_12417;
wire net_10676;
wire net_4687;
wire net_1141;
wire net_6253;
wire net_10621;
wire net_3243;
wire net_4867;
wire net_6321;
wire net_7871;
wire net_7584;
wire net_2104;
wire net_5564;
wire net_1288;
wire net_6190;
wire net_4708;
wire net_12554;
wire net_10511;
wire net_2766;
wire net_10559;
wire net_3771;
wire net_12469;
wire net_2300;
wire net_2417;
wire net_8119;
wire net_6710;
wire net_14406;
wire net_8426;
wire net_741;
wire net_7091;
wire net_13915;
wire net_6383;
wire net_4816;
wire net_5509;
wire net_6434;
wire net_11428;
wire net_6472;
wire net_7853;
wire net_13765;
wire net_11604;
wire net_3789;
wire net_13288;
wire net_5524;
wire net_9598;
wire net_4937;
wire net_11947;
wire net_4199;
wire net_11897;
wire net_1043;
wire net_12977;
wire net_2850;
wire net_770;
wire net_13905;
wire net_12901;
wire net_1005;
wire net_9737;
wire net_11792;
wire net_11198;
wire net_6389;
wire net_7493;
wire net_1059;
wire net_1630;
wire net_3891;
wire net_4918;
wire net_2956;
wire net_1082;
wire net_1796;
wire net_10328;
wire net_11170;
wire net_10405;
wire net_5187;
wire net_7501;
wire net_11368;
wire net_11291;
wire net_11861;
wire net_1507;
wire net_2310;
wire net_257;
wire net_3296;
wire net_11407;
wire net_10096;
wire net_8543;
wire net_7466;
wire net_9978;
wire net_474;
wire net_5500;
wire net_5770;
wire net_12518;
wire net_6576;
wire net_11421;
wire net_958;
wire net_12646;
wire net_11934;
wire net_11940;
wire net_4556;
wire net_6400;
wire net_7947;
wire net_11855;
wire net_11447;
wire net_12244;
wire net_12407;
wire net_944;
wire net_6199;
wire net_1734;
wire net_10189;
wire net_10008;
wire net_11175;
wire net_4308;
wire net_5534;
wire net_13477;
wire net_12538;
wire net_10987;
wire net_11002;
wire net_7199;
wire net_13450;
wire net_7166;
wire net_12580;
wire net_1728;
wire net_3050;
wire net_12883;
wire net_5963;
wire x1595;
wire net_3956;
wire net_12426;
wire net_10218;
wire net_8761;
wire net_8467;
wire net_13669;
wire net_425;
wire net_12028;
wire net_287;
wire net_189;
wire net_5204;
wire net_10414;
wire net_9893;
wire net_9860;
wire net_2205;
wire net_3755;
wire net_6036;
wire net_13154;
wire net_433;
wire net_11709;
wire net_8108;
wire net_8296;
wire net_4443;
wire net_11344;
wire net_13667;
wire net_368;
wire net_8064;
wire net_224;
wire net_4833;
wire net_1898;
wire net_10670;
wire net_9073;
wire net_608;
wire net_1212;
wire net_3604;
wire net_2000;
wire net_13089;
wire net_4383;
wire net_5331;
wire net_6226;
wire net_12502;
wire net_13194;
wire net_3706;
wire net_10603;
wire net_1020;
wire net_2984;
wire net_7062;
wire net_12879;
wire net_3282;
wire net_11997;
wire net_8299;
wire net_3122;
wire net_13989;
wire net_8546;
wire net_12832;
wire net_10164;
wire net_10763;
wire net_12521;
wire net_8594;
wire net_11965;
wire net_2094;
wire net_6416;
wire net_2543;
wire net_7282;
wire net_8275;
wire net_13227;
wire net_760;
wire net_2083;
wire net_12050;
wire net_8318;
wire net_873;
wire net_3851;
wire net_1811;
wire net_2488;
wire net_13884;
wire net_4536;
wire net_12374;
wire net_11080;
wire net_5034;
wire net_2588;
wire net_7802;
wire net_8192;
wire net_1870;
wire net_5200;
wire net_9771;
wire net_704;
wire net_12772;
wire net_12906;
wire net_2063;
wire net_3997;
wire net_192;
wire net_1356;
wire net_1739;
wire net_2912;
wire net_8913;
wire net_4140;
wire net_4393;
wire net_6541;
wire net_3816;
wire net_6101;
wire x1467;
wire net_13254;
wire net_13457;
wire net_735;
wire net_14269;
wire net_5539;
wire net_9056;
wire net_1711;
wire net_3809;
wire net_2084;
wire net_8186;
wire net_11590;
wire net_9442;
wire net_9530;
wire net_1081;
wire net_5085;
wire net_7031;
wire net_2037;
wire net_8163;
wire net_7349;
wire net_1237;
wire net_12478;
wire net_1420;
wire net_4789;
wire net_12653;
wire net_9112;
wire net_8680;
wire net_4836;
wire net_9587;
wire net_4064;
wire net_9712;
wire net_4237;
wire net_9602;
wire net_9542;
wire net_4559;
wire net_11663;
wire net_699;
wire net_3144;
wire net_7782;
wire net_7270;
wire net_359;
wire net_9283;
wire net_12892;
wire net_5239;
wire net_2526;
wire net_9414;
wire net_9068;
wire net_12862;
wire net_7338;
wire net_11316;
wire net_1644;
wire net_2819;
wire net_5827;
wire net_12126;
wire net_882;
wire net_2800;
wire net_14225;
wire net_7940;
wire net_1827;
wire net_6433;
wire net_8255;
wire net_12606;
wire net_1190;
wire net_3225;
wire net_4109;
wire net_8903;
wire net_3858;
wire net_14182;
wire net_10813;
wire net_7838;
wire net_4093;
wire net_6449;
wire net_4799;
wire net_13812;
wire net_8721;
wire net_12021;
wire net_1207;
wire net_2283;
wire net_10436;
wire net_9829;
wire net_6066;
wire net_8228;
wire net_2121;
wire net_2191;
wire net_14326;
wire net_13318;
wire net_13304;
wire net_2252;
wire net_10690;
wire net_4755;
wire net_13168;
wire net_12617;
wire net_7951;
wire net_12416;
wire net_12352;
wire net_14249;
wire net_2126;
wire net_5022;
wire net_1577;
wire net_1054;
wire net_4595;
wire net_10449;
wire net_9931;
wire net_7342;
wire net_9524;
wire net_2727;
wire net_12461;
wire net_5605;
wire net_2257;
wire net_6952;
wire net_10640;
wire net_3418;
wire net_3655;
wire net_2304;
wire net_5491;
wire net_14098;
wire net_13217;
wire net_12044;
wire net_2968;
wire net_7314;
wire net_12942;
wire net_10649;
wire net_5989;
wire net_12339;
wire net_7418;
wire net_1593;
wire net_2643;
wire net_5845;
wire net_8918;
wire net_10397;
wire net_9591;
wire net_3380;
wire net_3722;
wire net_12794;
wire net_11117;
wire net_11762;
wire net_1517;
wire net_5115;
wire net_4502;
wire net_12275;
wire net_11218;
wire net_5980;
wire net_13131;
wire net_12567;
wire net_2076;
wire net_2218;
wire net_4378;
wire net_6505;
wire net_6705;
wire net_9192;
wire net_6807;
wire net_10147;
wire net_1690;
wire net_9811;
wire net_1078;
wire net_12340;
wire net_9853;
wire net_11924;
wire net_2093;
wire net_2997;
wire net_6813;
wire net_6382;
wire net_5681;
wire net_13126;
wire net_14186;
wire net_10635;
wire net_9076;
wire net_7239;
wire net_14341;
wire net_12269;
wire net_11787;
wire net_5197;
wire net_12703;
wire net_13059;
wire net_12856;
wire net_2355;
wire net_13825;
wire net_9549;
wire net_4357;
wire net_3262;
wire net_139;
wire net_2536;
wire net_5890;
wire net_7968;
wire net_2949;
wire net_3429;
wire net_10954;
wire net_9032;
wire net_4495;
wire net_12587;
wire net_1708;
wire net_12398;
wire net_5519;
wire net_12824;
wire net_7454;
wire net_4196;
wire net_13678;
wire net_3974;
wire net_13112;
wire net_4626;
wire net_12575;
wire net_13050;
wire net_8532;
wire net_8478;
wire net_722;
wire net_2976;
wire net_13138;
wire net_5420;
wire net_12094;
wire net_988;
wire net_8221;
wire net_13099;
wire net_3621;
wire net_5798;
wire net_11351;
wire net_14313;
wire net_5223;
wire net_12441;
wire net_9820;
wire net_8216;
wire net_435;
wire net_12077;
wire net_1830;
wire net_4091;
wire net_12110;
wire net_132;
wire x1564;
wire net_2838;
wire net_5156;
wire net_6481;
wire net_1649;
wire net_6603;
wire net_1837;
wire net_1841;
wire net_5219;
wire net_5614;
wire net_6973;
wire net_1249;
wire net_2427;
wire net_4601;
wire net_1071;
wire net_3378;
wire net_8075;
wire net_7973;
wire net_3163;
wire net_4928;
wire net_5004;
wire net_5817;
wire net_6221;
wire net_9776;
wire x699;
wire net_1701;
wire net_4417;
wire net_5675;
wire net_11156;
wire net_822;
wire net_7145;
wire net_14007;
wire net_8678;
wire net_12175;
wire net_1633;
wire net_7084;
wire net_11132;
wire net_12150;
wire net_6561;
wire net_13470;
wire net_5251;
wire net_6842;
wire net_8694;
wire net_1974;
wire net_7701;
wire net_319;
wire net_8010;
wire net_2670;
wire net_4963;
wire net_1743;
wire net_2597;
wire net_5913;
wire net_11480;
wire net_9996;
wire net_9021;
wire net_1544;
wire net_7640;
wire net_11887;
wire net_7366;
wire net_4400;
wire net_10044;
wire net_4139;
wire net_2923;
wire net_10340;
wire net_7545;
wire net_512;
wire net_7929;
wire net_1174;
wire net_1109;
wire net_6664;
wire net_6731;
wire net_12326;
wire net_3102;
wire net_4224;
wire net_7510;
wire net_13733;
wire net_13513;
wire net_9683;
wire net_3457;
wire net_5780;
wire net_5721;
wire net_10963;
wire net_7904;
wire net_13119;
wire net_11721;
wire net_5276;
wire net_1102;
wire net_4471;
wire net_13644;
wire net_5487;
wire net_4976;
wire net_5640;
wire net_5245;
wire net_11205;
wire net_3371;
wire net_5317;
wire net_14175;
wire net_13953;
wire net_2692;
wire net_6800;
wire net_9375;
wire net_3777;
wire net_12673;
wire net_11322;
wire net_1875;
wire net_14355;
wire net_5862;
wire net_3420;
wire net_13353;
wire net_10285;
wire net_14382;
wire net_3887;
wire net_6279;
wire net_7050;
wire net_7516;
wire net_1487;
wire net_7037;
wire x681;
wire net_4572;
wire net_10020;
wire net_2759;
wire net_7484;
wire net_13373;
wire net_5408;
wire net_8243;
wire net_14128;
wire net_12486;
wire net_3634;
wire net_12189;
wire net_8736;
wire net_13348;
wire net_12953;
wire net_5178;
wire net_7678;
wire net_2835;
wire net_4543;
wire net_13705;
wire net_4871;
wire net_6599;
wire net_14215;
wire net_1240;
wire net_9213;
wire net_3000;
wire net_12200;
wire net_10338;
wire net_10349;
wire net_2564;
wire net_2821;
wire net_12674;
wire net_1658;
wire net_13048;
wire net_5481;
wire net_5688;
wire net_858;
wire net_7318;
wire net_3007;
wire net_9505;
wire net_9338;
wire net_7554;
wire net_4487;
wire net_8986;
wire net_4766;
wire net_9122;
wire net_3174;
wire net_6004;
wire x172;
wire net_2876;
wire net_6966;
wire net_8504;
wire net_844;
wire net_13549;
wire net_1496;
wire net_9867;
wire net_325;
wire net_3735;
wire net_7995;
wire net_1820;
wire net_10870;
wire net_11422;
wire net_1427;
wire net_5123;
wire net_8175;
wire net_3921;
wire net_5690;
wire net_7075;
wire net_13274;
wire net_5899;
wire net_4098;
wire net_5478;
wire net_7251;
wire net_10287;
wire net_5956;
wire net_12106;
wire net_9827;
wire net_5014;
wire net_11029;
wire net_4036;
wire net_7517;
wire net_11266;
wire net_1521;
wire net_4182;
wire net_6274;
wire net_10308;
wire net_6020;
wire net_7172;
wire net_1677;
wire net_11813;
wire net_7908;
wire net_11727;
wire net_4734;
wire net_7179;
wire net_2991;
wire net_13260;
wire net_10077;
wire net_564;
wire net_4276;
wire net_6154;
wire net_10618;
wire net_2050;
wire net_4086;
wire net_13992;
wire net_9082;
wire net_7089;
wire net_2811;
wire net_6788;
wire net_813;
wire net_14105;
wire net_10661;
wire net_5609;
wire net_1027;
wire net_2612;
wire net_8791;
wire net_5230;
wire net_2042;
wire net_12403;
wire net_1408;
wire net_265;
wire net_7189;
wire net_13626;
wire net_11649;
wire net_6649;
wire net_8110;
wire net_11720;
wire net_10949;
wire net_3488;
wire net_8673;
wire net_3023;
wire net_13538;
wire net_11097;
wire net_6774;
wire net_5584;
wire net_10834;
wire net_1202;
wire net_14373;
wire net_9351;
wire net_10890;
wire net_9258;
wire net_1155;
wire net_925;
wire net_4932;
wire net_6776;
wire net_7452;
wire net_9787;
wire net_12827;
wire net_5384;
wire net_7374;
wire net_12764;
wire net_11317;
wire net_10974;
wire net_12074;
wire net_4661;
wire net_2695;
wire net_10331;
wire net_864;
wire net_10196;
wire net_11054;
wire net_14337;
wire net_13336;
wire net_7691;
wire net_13004;
wire net_12851;
wire net_12611;
wire net_7404;
wire net_12787;
wire net_8564;
wire net_12285;
wire net_7783;
wire net_4113;
wire x1550;
wire net_8850;
wire net_10365;
wire net_6284;
wire net_660;
wire net_2298;
wire net_14060;
wire net_9436;
wire net_7132;
wire net_9707;
wire net_2313;
wire net_11655;
wire net_6580;
wire net_9044;
wire net_1908;
wire net_6172;
wire net_7595;
wire net_7647;
wire net_230;
wire net_4214;
wire net_9309;
wire net_3383;
wire net_13020;
wire net_12958;
wire net_6985;
wire net_7265;
wire net_3349;
wire net_4782;
wire net_6751;
wire net_1222;
wire net_3404;
wire net_14080;
wire net_14291;
wire net_3810;
wire net_9172;
wire net_3914;
wire net_7607;
wire net_12018;
wire net_6531;
wire net_14104;
wire net_6463;
wire net_11973;
wire net_4739;
wire net_6455;
wire net_4156;
wire net_10610;
wire net_5777;
wire net_8823;
wire net_12685;
wire x1006;
wire net_13449;
wire net_7576;
wire net_13693;
wire net_12459;
wire net_3440;
wire net_6904;
wire net_3358;
wire net_1776;
wire net_2145;
wire net_6488;
wire net_11109;
wire net_3368;
wire net_5747;
wire net_3311;
wire net_4014;
wire net_8874;
wire net_11020;
wire net_14036;
wire net_12729;
wire net_10887;
wire net_7204;
wire net_10454;
wire net_2132;
wire net_2292;
wire net_9313;
wire net_12367;
wire net_1880;
wire net_10716;
wire net_3862;
wire net_184;
wire net_5103;
wire net_13943;
wire net_4853;
wire net_8699;
wire net_5855;
wire net_10757;
wire net_14087;
wire net_11247;
wire net_10427;
wire net_10474;
wire net_7203;
wire net_13080;
wire net_11507;
wire net_3538;
wire net_1867;
wire net_9498;
wire net_8205;
wire net_1949;
wire net_2650;
wire net_13568;
wire net_10455;
wire net_1583;
wire net_1804;
wire net_9454;
wire net_2331;
wire net_4408;
wire net_6667;
wire net_1563;
wire net_4291;
wire net_3898;
wire net_13969;
wire net_12389;
wire net_4948;
wire net_8637;
wire net_7600;
wire net_13073;
wire net_5599;
wire net_3361;
wire net_1135;
wire net_1365;
wire net_13019;
wire net_11674;
wire net_10553;
wire net_1346;
wire net_5047;
wire net_14285;
wire net_8578;
wire net_1942;
wire net_11484;
wire net_11478;
wire net_13865;
wire net_10070;
wire net_13835;
wire net_9220;
wire net_12119;
wire net_9277;
wire net_1801;
wire net_13755;
wire net_7891;
wire net_14150;
wire net_1267;
wire net_14364;
wire net_6093;
wire net_12570;
wire net_11846;
wire net_3661;
wire net_3944;
wire net_9188;
wire net_4350;
wire net_6029;
wire net_4893;
wire net_12982;
wire net_8955;
wire net_669;
wire net_6526;
wire net_937;
wire net_11252;
wire net_10179;
wire net_5888;
wire net_8452;
wire net_9575;
wire net_5131;
wire net_8030;
wire net_2349;
wire net_479;
wire net_11074;
wire net_8740;
wire net_12769;
wire net_1294;
wire net_10350;
wire net_6086;
wire net_2030;
wire net_1587;
wire net_3520;
wire net_5006;
wire net_13232;
wire net_1354;
wire net_11025;
wire net_1308;
wire net_796;
wire net_2904;
wire net_7631;
wire net_12081;
wire net_4332;
wire net_9992;
wire net_1389;
wire net_648;
wire net_11901;
wire net_12114;
wire net_6884;
wire net_12040;
wire net_8150;
wire net_13818;
wire net_4748;
wire net_14300;
wire net_3250;
wire net_7054;
wire net_11950;
wire net_7625;
wire net_5304;
wire net_3658;
wire net_10737;
wire net_548;
wire net_12560;
wire net_2402;
wire net_4985;
wire net_6529;
wire net_14146;
wire net_5902;
wire net_6964;
wire net_9148;
wire net_5082;
wire net_636;
wire net_10239;
wire net_4269;
wire net_8237;
wire net_8159;
wire net_8556;
wire net_7649;
wire net_12179;
wire net_10739;
wire net_10232;
wire net_8725;
wire net_8471;
wire net_8218;
wire net_4492;
wire net_6700;
wire net_1961;
wire net_10831;
wire net_1260;
wire net_12678;
wire net_10124;
wire net_4165;
wire net_4262;
wire net_9832;
wire net_10228;
wire net_1185;
wire net_4506;
wire net_13868;
wire net_5001;
wire net_239;
wire net_13396;
wire net_310;
wire net_11216;
wire net_10367;
wire net_2437;
wire net_7942;
wire net_10792;
wire net_9401;
wire net_8982;
wire net_9917;
wire net_4826;
wire net_1912;
wire net_13498;
wire net_9566;
wire net_11353;
wire net_11263;
wire net_5886;
wire net_11416;
wire net_9118;
wire net_11542;
wire net_13711;
wire net_9906;
wire net_682;
wire net_1963;
wire net_7122;
wire net_1538;
wire net_14228;
wire net_13558;
wire net_9501;
wire net_12049;
wire net_11499;
wire net_8989;
wire net_13965;
wire net_3560;
wire net_5804;
wire net_1007;
wire net_1579;
wire net_7000;
wire net_13440;
wire net_4772;
wire net_7007;
wire net_11415;
wire net_1292;
wire net_7197;
wire net_10703;
wire net_10520;
wire net_6484;
wire net_7861;
wire net_10771;
wire net_12262;
wire net_1999;
wire net_1014;
wire net_6669;
wire net_11039;
wire net_1444;
wire net_2796;
wire net_11400;
wire net_2679;
wire net_5016;
wire net_4024;
wire net_6255;
wire net_4082;
wire net_6699;
wire net_11577;
wire net_9544;
wire net_9083;
wire net_538;
wire net_12994;
wire net_12443;
wire net_4130;
wire net_6280;
wire net_1937;
wire net_8043;
wire net_13306;
wire net_9965;
wire net_7215;
wire net_366;
wire net_1854;
wire net_1956;
wire net_11339;
wire net_1917;
wire net_13433;
wire net_1614;
wire net_1755;
wire net_13491;
wire net_12911;
wire net_1359;
wire net_11958;
wire net_7119;
wire net_2460;
wire net_13228;
wire net_8929;
wire net_10255;
wire net_3209;
wire net_12791;
wire net_11238;
wire net_4891;
wire net_8688;
wire net_13424;
wire net_11348;
wire net_10874;
wire net_8412;
wire net_12618;
wire net_209;
wire net_9242;
wire net_1282;
wire net_7716;
wire net_294;
wire net_8211;
wire net_13291;
wire net_9837;
wire net_4041;
wire net_10797;
wire net_2429;
wire net_9217;
wire net_1265;
wire net_3204;
wire net_10822;
wire net_8996;
wire net_6224;
wire net_8697;
wire net_11203;
wire net_12315;
wire net_3471;
wire net_9677;
wire net_12984;
wire net_1619;
wire net_5468;
wire net_8039;
wire net_12727;
wire net_2124;
wire net_5934;
wire net_9692;
wire net_12354;
wire net_12966;
wire net_1161;
wire net_3512;
wire net_7070;
wire net_4671;
wire net_13606;
wire net_12695;
wire net_8907;
wire net_7663;
wire net_11531;
wire net_9394;
wire net_11385;
wire net_10382;
wire net_10177;
wire net_2430;
wire net_10721;
wire net_8433;
wire net_4461;
wire net_7687;
wire net_13598;
wire net_8500;
wire net_1395;
wire net_11942;
wire net_3481;
wire net_8877;
wire net_9360;
wire net_1589;
wire net_11875;
wire net_8114;
wire net_5353;
wire net_2396;
wire net_9098;
wire net_8756;
wire net_5270;
wire net_9921;
wire net_13298;
wire net_12456;
wire net_8354;
wire net_2445;
wire net_5815;
wire net_3396;
wire net_6640;
wire net_2856;
wire net_5324;
wire net_10592;
wire net_787;
wire net_10789;
wire net_7777;
wire net_8125;
wire net_3603;
wire net_4511;
wire net_7395;
wire net_13419;
wire net_9656;
wire net_2894;
wire net_4187;
wire net_8095;
wire net_13714;
wire net_6999;
wire net_1988;
wire net_7388;
wire net_12071;
wire net_14323;
wire net_3718;
wire net_11001;
wire net_8463;
wire net_4419;
wire net_6195;
wire net_10767;
wire net_3579;
wire net_5284;
wire net_11125;
wire net_3525;
wire net_10696;
wire net_11069;
wire net_6850;
wire net_13508;
wire net_8870;
wire net_1608;
wire net_2139;
wire net_506;
wire net_5332;
wire net_3769;
wire net_12802;
wire net_8019;
wire net_10250;
wire net_9330;
wire net_12836;
wire net_1910;
wire net_3775;
wire net_8278;
wire net_8103;
wire net_12689;
wire net_5432;
wire net_6586;
wire net_3544;
wire net_9517;
wire net_3034;
wire net_5229;
wire net_9488;
wire net_5096;
wire net_7895;
wire net_7938;
wire net_6285;
wire net_7610;
wire net_12817;
wire net_11030;
wire net_9664;
wire net_2493;
wire net_11914;
wire net_919;
wire net_9009;
wire net_7589;
wire net_12055;
wire net_11574;
wire net_6909;
wire net_290;
wire net_6476;
wire net_7044;
wire net_13676;
wire net_6315;
wire net_6836;
wire net_10913;
wire net_3313;
wire net_4008;
wire net_6444;
wire net_12669;
wire net_9987;
wire net_2209;
wire net_1372;
wire net_8803;
wire net_11935;
wire net_1757;
wire x38;
wire net_5769;
wire x1203;
wire net_3591;
wire net_5729;
wire net_13341;
wire net_8816;
wire net_5215;
wire net_13084;
wire net_13015;
wire net_11926;
wire net_12430;
wire net_4436;
wire net_2682;
wire net_7151;
wire net_8053;
wire net_140;
wire net_11949;
wire net_2329;
wire net_6612;
wire net_8911;
wire x145;
wire net_7077;
wire net_2150;
wire net_3790;
wire net_7129;
wire net_9141;
wire net_2065;
wire net_10003;
wire net_13244;
wire net_10030;
wire net_4267;
wire net_8373;
wire net_2927;
wire net_12482;
wire net_7397;
wire net_7328;
wire net_11831;
wire net_11838;
wire net_194;
wire net_4856;
wire net_2178;
wire net_13941;
wire net_11264;
wire net_9448;
wire net_5292;
wire net_1128;
wire net_10134;
wire net_3073;
wire net_2713;
wire net_13161;
wire net_11582;
wire net_12539;
wire net_11320;
wire net_8840;
wire net_13846;
wire net_7949;
wire net_804;
wire net_10541;
wire net_1119;
wire net_9637;
wire net_3548;
wire net_1314;
wire net_9400;
wire net_4312;
wire net_8845;
wire net_6325;
wire net_5376;
wire net_531;
wire net_5299;
wire net_8582;
wire net_499;
wire net_8852;
wire net_3345;
wire net_2752;
wire net_10125;
wire net_7855;
wire net_11642;
wire net_11006;
wire net_9126;
wire net_7127;
wire net_7448;
wire net_10701;
wire net_11900;
wire net_9699;
wire net_9476;
wire net_10742;
wire net_3328;
wire net_13413;
wire net_3534;
wire net_4390;
wire net_8027;
wire net_12155;
wire net_1765;
wire net_8965;
wire net_10174;
wire net_2107;
wire net_10424;
wire net_180;
wire net_11231;
wire net_6208;
wire net_13462;
wire net_6859;
wire net_2420;
wire net_2774;
wire net_6068;
wire net_12437;
wire net_5657;
wire net_13410;
wire net_4367;
wire net_1979;
wire net_5135;
wire net_13927;
wire net_3290;
wire net_3731;
wire net_1475;
wire net_1460;
wire net_10241;
wire net_1451;
wire net_14112;
wire net_13978;
wire net_12246;
wire net_10601;
wire net_5446;
wire net_5008;
wire net_5065;
wire net_8419;
wire net_6619;
wire net_12719;
wire net_4803;
wire net_203;
wire net_2173;
wire net_9053;
wire net_6865;
wire net_6597;
wire net_7539;
wire net_11071;
wire net_1602;
wire net_12213;
wire net_6263;
wire net_5590;
wire net_9919;
wire net_613;
wire net_237;
wire net_13239;
wire net_11673;
wire net_14334;
wire net_5476;
wire net_14236;
wire net_3744;
wire net_11851;
wire net_4635;
wire net_1095;
wire net_12193;
wire net_578;
wire net_4729;
wire net_12236;
wire net_6570;
wire net_8309;
wire net_11288;
wire net_8514;
wire net_6939;
wire net_12968;
wire net_4485;
wire net_1558;
wire net_2743;
wire net_8603;
wire net_4641;
wire net_10958;
wire net_388;
wire net_2159;
wire net_10806;
wire net_14360;
wire net_3647;
wire net_14138;
wire net_536;
wire net_455;
wire net_11515;
wire net_1332;
wire net_10294;
wire net_115;
wire net_7498;
wire net_10589;
wire net_3276;
wire net_3339;
wire net_6303;
wire net_11980;
wire net_9428;
wire net_13525;
wire net_7352;
wire net_7468;
wire net_9130;
wire net_1832;
wire net_408;
wire net_12474;
wire net_12622;
wire net_10904;
wire net_1026;
wire net_10582;
wire net_2215;
wire net_3246;
wire net_1845;
wire net_6453;
wire net_2573;
wire net_10633;
wire net_12225;
wire net_9369;
wire net_9939;
wire net_10312;
wire net_7378;
wire net_3390;
wire net_3993;
wire net_13673;
wire net_1401;
wire net_2372;
wire net_12579;
wire net_3909;
wire net_12870;
wire net_868;
wire net_11858;
wire net_11223;
wire net_10979;
wire net_7889;
wire net_14394;
wire net_7248;
wire net_6079;
wire net_13311;
wire net_6821;
wire net_13750;
wire net_443;
wire x1193;
wire net_5029;
wire net_13871;
wire net_6367;
wire net_6495;
wire net_8486;
wire net_922;
wire net_522;
wire net_270;
wire net_2638;
wire net_9747;
wire net_13355;
wire net_12364;
wire net_7956;
wire net_5429;
wire net_14034;
wire x124;
wire net_11346;
wire net_1990;
wire net_4992;
wire net_7456;
wire net_10442;
wire net_5757;
wire net_6140;
wire net_2264;
wire net_11632;
wire net_977;
wire net_643;
wire net_4780;
wire net_9951;
wire x765;
wire net_7880;
wire net_11278;
wire net_11988;
wire net_11601;
wire net_622;
wire net_6876;
wire net_13564;
wire net_11993;
wire net_11165;
wire net_6175;
wire net_3587;
wire net_3762;
wire net_10580;
wire net_3687;
wire net_11277;
wire net_5909;
wire net_10056;
wire net_11225;
wire net_12015;
wire net_10483;
wire net_5307;
wire net_1338;
wire net_4920;
wire net_7842;
wire net_2045;
wire net_3874;
wire net_2053;
wire net_9357;
wire net_11790;
wire net_6623;
wire net_11829;
wire net_2180;
wire net_2869;
wire net_3332;
wire net_4242;
wire net_1892;
wire net_3446;
wire net_1798;
wire net_2119;
wire net_3220;
wire net_4427;
wire net_4720;
wire net_7401;
wire net_13108;
wire net_13109;
wire net_13287;
wire net_8627;
wire net_837;
wire net_7474;
wire net_10723;
wire net_3469;
wire net_9449;
wire net_5920;
wire net_6124;
wire net_8384;
wire net_6992;
wire net_927;
wire net_13519;
wire net_11686;
wire net_2007;
wire net_5143;
wire net_5763;
wire net_7703;
wire net_713;
wire net_10653;
wire net_1519;
wire net_693;
wire net_12633;
wire net_5711;
wire net_6378;
wire net_13338;
wire net_8700;
wire net_11104;
wire net_729;
wire net_11390;
wire net_9222;
wire net_4197;
wire net_13777;
wire net_3964;
wire net_12660;
wire net_13156;
wire net_4219;
wire net_7093;
wire net_7324;
wire net_13948;
wire net_9169;
wire net_8447;
wire net_9311;
wire net_5366;
wire net_9898;
wire net_11865;
wire net_8711;
wire net_13571;
wire net_10847;
wire net_341;
wire net_13611;
wire net_13391;
wire net_11651;
wire net_10208;
wire net_12992;
wire net_970;
wire net_13362;
wire net_488;
wire net_13389;
wire net_8653;
wire net_12009;
wire net_10460;
wire net_4909;
wire net_6034;
wire net_5452;
wire net_8088;
wire net_8324;
wire net_2319;
wire net_13917;
wire net_13184;
wire net_3044;
wire net_5929;
wire net_11785;
wire net_5458;
wire net_7102;
wire net_11145;
wire net_8440;
wire net_1532;
wire net_8971;
wire net_13726;
wire net_12308;
wire net_6653;
wire net_14071;
wire net_8207;
wire net_4475;
wire net_14233;
wire net_12038;
wire net_11595;
wire net_10100;
wire net_2163;
wire net_3417;
wire net_3307;
wire net_7765;
wire net_13301;
wire net_12534;
wire net_553;
wire net_4958;
wire net_4212;
wire net_5057;
wire net_6133;
wire net_1093;
wire net_2592;
wire net_7797;
wire net_6230;
wire net_7680;
wire net_8300;
wire x1572;
wire net_9876;
wire net_3580;
wire net_3259;
wire net_6239;
wire net_9877;
wire net_5260;
wire net_4701;
wire net_10057;
wire net_10889;
wire net_8833;
wire net_8922;
wire net_710;
wire net_462;
wire net_418;
wire net_3097;
wire net_5836;
wire net_161;
wire net_6478;
wire net_7988;
wire net_14401;
wire net_8660;
wire net_3970;
wire net_12516;
wire net_1486;
wire net_173;
wire net_2606;
wire net_3018;
wire net_14317;
wire net_1839;
wire net_2320;
wire net_1665;
wire net_11076;
wire net_9237;
wire net_3006;
wire net_6203;
wire net_13744;
wire net_10970;
wire net_8525;
wire net_8349;
wire net_1681;
wire net_7936;
wire net_3550;
wire net_12377;
wire net_11172;
wire net_7998;
wire net_6893;
wire net_9466;
wire net_2224;
wire net_7066;
wire net_10037;
wire net_4272;
wire net_6512;
wire net_5733;
wire net_10532;
wire net_746;
wire net_13406;
wire net_5877;
wire net_6147;
wire net_1274;
wire net_1682;
wire net_2458;
wire net_11302;
wire net_9324;
wire net_10788;
wire net_5743;
wire net_7910;
wire net_3435;
wire net_10109;
wire net_3466;
wire net_2635;
wire net_3374;
wire net_5207;
wire net_13540;
wire net_4995;
wire net_5572;
wire net_7834;
wire net_1663;
wire net_629;
wire net_8283;
wire net_1037;
wire net_8666;
wire net_2019;
wire net_4209;
wire net_4676;
wire net_9382;
wire net_8395;
wire net_3019;
wire net_6675;
wire net_13784;
wire net_13033;
wire net_7549;
wire net_5579;
wire net_2351;
wire net_6793;
wire net_9628;
wire net_1350;
wire net_1648;
wire net_6242;
wire net_12594;
wire net_1623;
wire net_2982;
wire net_6219;
wire net_631;
wire net_6948;
wire net_14201;
wire net_12128;
wire net_4410;
wire net_7230;
wire net_10086;
wire net_5785;
wire net_14047;
wire net_13143;
wire net_4007;
wire net_8566;
wire net_4499;
wire net_12100;
wire net_14251;
wire net_13657;
wire net_8650;
wire net_7190;
wire net_10907;
wire net_9910;
wire net_8596;
wire net_6928;
wire net_670;
wire net_10984;
wire net_6250;
wire net_12147;
wire net_2687;
wire net_12166;
wire net_6651;
wire net_9889;
wire net_5485;
wire net_7023;
wire net_7243;
wire net_12004;
wire net_10750;
wire net_3554;
wire net_9842;
wire net_9721;
wire net_12853;
wire net_12323;
wire net_1920;
wire net_4101;
wire net_3928;
wire net_13369;
wire net_2010;
wire net_3854;
wire net_7038;
wire net_11665;
wire net_8782;
wire net_6717;
wire net_6941;
wire net_9793;
wire net_9857;
wire net_8321;
wire net_9139;
wire net_5493;
wire net_13759;
wire net_4672;
wire net_8862;
wire net_6743;
wire net_755;
wire x744;
wire net_9557;
wire net_1723;
wire net_8465;
wire net_9285;
wire net_2900;
wire net_7754;
wire net_11015;
wire net_5152;
wire net_12545;
wire net_5718;
wire net_8190;
wire net_4376;
wire net_5892;
wire net_14397;
wire net_13468;
wire net_3151;
wire net_6763;
wire net_12890;
wire net_2306;
wire net_3628;
wire net_6053;
wire net_12382;
wire net_12023;
wire net_2873;
wire net_3272;
wire net_12829;
wire net_2254;
wire net_2861;
wire net_11319;
wire net_1652;
wire net_1429;
wire net_11844;
wire net_11061;
wire net_14343;
wire net_14223;
wire net_9570;
wire net_4574;
wire net_7130;
wire net_1209;
wire net_2725;
wire net_13166;
wire net_3613;
wire net_8964;
wire x1062;
wire net_4615;
wire net_13076;
wire net_4038;
wire net_727;
wire net_847;
wire net_11242;
wire net_10157;
wire net_4787;
wire net_9804;
wire net_11740;
wire net_283;
wire net_12864;
wire net_13505;
wire net_12559;
wire net_5117;
wire net_3190;
wire net_4955;
wire net_4690;
wire net_12796;
wire net_3757;
wire net_11457;
wire net_5020;
wire x342;
wire net_14126;
wire net_7316;
wire net_12658;
wire net_9224;
wire net_4445;
wire net_5445;
wire net_7428;
wire net_10023;
wire net_11115;
wire net_10990;
wire net_14247;
wire net_7958;
wire net_344;
wire net_14102;
wire net_3951;
wire net_4757;
wire net_2269;
wire net_884;
wire net_14184;
wire net_712;
wire net_13010;
wire net_11635;
wire net_1422;
wire net_2281;
wire net_12940;
wire net_2259;
wire net_12124;
wire net_4497;
wire net_11527;
wire net_10651;
wire net_6670;
wire net_1106;
wire net_4095;
wire net_13629;
wire net_8483;
wire net_2739;
wire net_2972;
wire net_13330;
wire net_5611;
wire net_11715;
wire net_10113;
wire net_2110;
wire net_11311;
wire net_10836;
wire net_2919;
wire net_10642;
wire net_2893;
wire net_11435;
wire net_2241;
wire net_13006;
wire net_2358;
wire net_3227;
wire net_12651;
wire net_9522;
wire net_8615;
wire net_8682;
wire net_3057;
wire net_1547;
wire net_9039;
wire net_571;
wire net_13053;
wire net_10692;
wire net_8768;
wire net_10543;
wire net_7569;
wire net_5122;
wire net_12495;
wire net_10400;
wire net_4935;
wire net_12168;
wire net_3934;
wire net_10385;
wire x1557;
wire net_11146;
wire net_5423;
wire net_13972;
wire net_1877;
wire net_720;
wire net_7971;
wire net_6507;
wire net_9912;
wire net_7653;
wire net_9038;
wire net_12152;
wire net_10395;
wire net_14005;
wire net_5209;
wire net_7344;
wire net_2199;
wire net_5055;
wire net_10628;
wire net_7303;
wire net_4794;
wire net_684;
wire net_2625;
wire net_4149;
wire net_2648;
wire net_5687;
wire net_7299;
wire net_7542;
wire net_3720;
wire net_510;
wire net_12922;
wire net_10909;
wire net_6849;
wire net_10292;
wire net_1595;
wire net_5849;
wire net_114;
wire net_8885;
wire net_12919;
wire net_2653;
wire net_3432;
wire net_2960;
wire net_2974;
wire net_9078;
wire net_6519;
wire net_3895;
wire net_8339;
wire net_8257;
wire net_13660;
wire net_6703;
wire net_12577;
wire net_11736;
wire net_2734;
wire net_12888;
wire net_13133;
wire net_494;
wire net_2782;
wire net_7043;
wire net_10637;
wire net_12569;
wire net_6761;
wire net_3146;
wire net_6294;
wire net_7827;
wire net_12877;
wire net_10999;
wire net_6390;
wire net_9347;
wire net_10496;
wire net_5237;
wire net_4283;
wire net_6592;
wire net_13830;
wire net_11553;
wire net_8953;
wire net_3022;
wire net_6084;
wire net_8226;
wire net_3461;
wire net_12365;
wire net_10989;
wire net_10956;
wire net_10327;
wire net_11747;
wire net_7495;
wire net_14366;
wire net_4610;
wire net_9616;
wire net_5741;
wire net_6391;
wire net_8476;
wire net_457;
wire net_4459;
wire net_12096;
wire net_8821;
wire net_2246;
wire net_772;
wire net_6308;
wire net_10180;
wire net_14375;
wire net_4371;
wire net_5700;
wire net_10190;
wire net_12773;
wire net_7441;
wire net_9671;
wire net_7966;
wire net_11807;
wire net_9159;
wire net_1277;
wire net_11899;
wire net_2661;
wire net_3893;
wire net_6113;
wire net_14260;
wire net_13459;
wire net_4706;
wire net_12467;
wire net_594;
wire net_5532;
wire net_11336;
wire net_9818;
wire net_4075;
wire net_6421;
wire net_7385;
wire net_14310;
wire net_6051;
wire net_11892;
wire net_8512;
wire net_11690;
wire net_1721;
wire net_2852;
wire net_6188;
wire net_7851;
wire net_12975;
wire net_4633;
wire net_4402;
wire net_6328;
wire net_6605;
wire net_6249;
wire net_5843;
wire net_2074;
wire net_8428;
wire net_5256;
wire net_5274;
wire net_10626;
wire net_10183;
wire net_2577;
wire net_11091;
wire net_8286;
wire net_2954;
wire net_1073;
wire net_8073;
wire net_11932;
wire x187;
wire net_1947;
wire net_3274;
wire net_2953;
wire net_141;
wire net_6380;
wire net_467;
wire net_879;
wire net_2910;
wire net_7227;
wire net_2415;
wire net_8728;
wire net_4851;
wire net_2081;
wire net_9245;
wire net_8738;
wire net_10522;
wire net_5195;
wire net_7312;
wire net_11426;
wire net_13225;
wire net_3165;
wire net_12644;
wire net_10740;
wire net_1348;
wire net_3197;
wire net_9774;
wire net_7276;
wire net_4965;
wire net_7201;
wire net_12295;
wire net_8648;
wire net_2302;
wire net_3422;
wire net_10151;
wire net_199;
wire net_12523;
wire net_2789;
wire net_7844;
wire net_12903;
wire net_431;
wire net_3835;
wire net_8545;
wire net_5783;
wire net_13649;
wire net_8250;
wire net_5502;
wire net_6805;
wire net_10898;
wire net_9373;
wire net_6387;
wire net_6403;
wire net_7734;
wire net_13873;
wire net_12409;
wire net_2368;
wire net_5186;
wire net_222;
wire net_4362;
wire net_13215;
wire net_12908;
wire net_4520;
wire net_3966;
wire net_3999;
wire net_7060;
wire net_7804;
wire net_1788;
wire net_6330;
wire net_12476;
wire net_607;
wire net_4301;
wire net_12392;
wire net_8106;
wire net_9739;
wire net_2935;
wire net_4142;
wire net_1045;
wire net_6166;
wire net_3497;
wire net_3905;
wire net_13087;
wire net_4345;
wire net_10507;
wire net_9318;
wire net_13249;
wire net_3516;
wire net_4939;
wire net_11799;
wire net_6547;
wire net_3601;
wire net_9933;
wire net_4588;
wire net_1438;
wire net_10374;
wire net_4395;
wire net_4538;
wire net_8502;
wire net_13044;
wire net_12052;
wire net_1143;
wire net_11167;
wire net_12662;
wire net_1088;
wire net_4527;
wire net_9434;
wire net_6410;
wire net_6419;
wire net_8548;
wire net_13262;
wire net_4144;
wire net_4716;
wire net_7586;
wire net_2079;
wire net_3885;
wire net_1731;
wire net_706;
wire net_2052;
wire net_6373;
wire net_9298;
wire net_9089;
wire net_14376;
wire net_9648;
wire net_9463;
wire net_2768;
wire net_6912;
wire net_12813;
wire net_5125;
wire net_13276;
wire net_13479;
wire net_12536;
wire net_551;
wire net_5952;
wire net_5368;
wire net_7873;
wire net_11769;
wire net_3636;
wire net_4617;
wire net_7184;
wire net_14095;
wire net_13182;
wire net_4727;
wire net_5032;
wire net_11046;
wire net_1536;
wire net_5852;
wire net_6232;
wire net_11033;
wire net_12504;
wire net_12419;
wire net_3478;
wire net_4168;
wire net_12376;
wire net_1498;
wire net_8117;
wire net_11371;
wire net_1199;
wire net_7986;
wire net_10815;
wire net_8930;
wire net_3627;
wire net_5561;
wire net_5530;
wire net_5626;
wire net_949;
wire net_4869;
wire net_289;
wire net_450;
wire net_14000;
wire net_12401;
wire net_10936;
wire net_8041;
wire net_7813;
wire net_9046;
wire net_4111;
wire net_14204;
wire net_9392;
wire net_10972;
wire net_1642;
wire net_2614;
wire net_14267;
wire net_12158;
wire net_10616;
wire net_5322;
wire net_12947;
wire net_12287;
wire net_12722;
wire net_14283;
wire net_2524;
wire net_11490;
wire net_8262;
wire net_1224;
wire net_9028;
wire net_2296;
wire net_6786;
wire net_9438;
wire net_13804;
wire net_13994;
wire net_768;
wire x1155;
wire net_3385;
wire net_11084;
wire net_357;
wire net_14068;
wire net_6954;
wire net_908;
wire net_9179;
wire net_12934;
wire net_13189;
wire net_7849;
wire net_519;
wire net_3451;
wire net_9697;
wire net_7085;
wire net_11773;
wire net_8790;
wire net_2694;
wire net_12280;
wire net_11052;
wire net_5607;
wire net_2096;
wire net_3118;
wire net_5555;
wire net_2697;
wire x821;
wire net_9184;
wire net_11501;
wire net_10808;
wire net_1829;
wire net_14240;
wire net_13904;
wire net_14082;
wire net_9190;
wire net_1204;
wire net_6282;
wire net_14089;
wire net_9780;
wire net_2342;
wire net_8331;
wire net_7336;
wire net_6628;
wire net_9969;
wire net_6778;
wire net_662;
wire net_862;
wire net_1986;
wire net_3214;
wire net_2307;
wire net_11472;
wire net_7168;
wire net_8127;
wire net_4174;
wire net_5396;
wire net_10864;
wire net_738;
wire net_4080;
wire net_4325;
wire net_12881;
wire net_1150;
wire net_504;
wire net_10333;
wire net_9789;
wire net_6634;
wire net_8203;
wire net_6467;
wire net_7527;
wire net_12613;
wire net_11537;
wire net_7698;
wire net_9164;
wire net_9012;
wire net_3406;
wire net_11657;
wire net_13110;
wire net_4229;
wire net_2130;
wire net_6474;
wire net_10198;
wire net_1148;
wire net_3362;
wire net_3120;
wire net_14324;
wire net_2382;
wire net_13620;
wire net_4504;
wire net_1561;
wire net_10698;
wire net_3442;
wire net_3864;
wire net_5942;
wire net_9271;
wire net_12161;
wire net_3269;
wire net_11455;
wire net_10472;
wire net_5796;
wire net_9730;
wire net_4421;
wire net_6666;
wire net_9416;
wire x1451;
wire net_6975;
wire net_13329;
wire net_9855;
wire net_1940;
wire net_4389;
wire net_13323;
wire net_11449;
wire net_13935;
wire net_11798;
wire net_10452;
wire net_10728;
wire net_8635;
wire net_11516;
wire net_12781;
wire net_10425;
wire net_4561;
wire net_11528;
wire net_991;
wire net_3912;
wire net_6528;
wire net_13204;
wire net_11676;
wire net_6753;
wire net_3088;
wire net_1473;
wire net_11107;
wire net_4607;
wire net_12484;
wire net_2979;
wire net_10714;
wire net_2772;
wire net_9564;
wire net_8491;
wire net_5775;
wire net_1674;
wire net_4180;
wire net_5582;
wire net_1651;
wire net_2375;
wire net_13582;
wire net_5109;
wire net_13839;
wire net_12116;
wire net_1806;
wire net_6422;
wire net_3234;
wire net_12180;
wire net_2347;
wire net_8746;
wire net_1363;
wire net_11710;
wire net_1869;
wire net_2684;
wire net_3806;
wire net_4053;
wire net_10795;
wire net_10352;
wire net_10526;
wire net_521;
wire net_3972;
wire net_14275;
wire net_13029;
wire net_9003;
wire net_2754;
wire net_267;
wire net_1585;
wire net_13748;
wire net_11613;
wire net_9143;
wire net_11099;
wire net_4012;
wire net_6898;
wire net_7421;
wire net_6169;
wire net_3663;
wire x77;
wire net_10885;
wire net_3260;
wire net_5110;
wire net_6647;
wire net_13017;
wire net_9186;
wire net_6465;
wire net_6486;
wire net_3681;
wire net_6048;
wire net_13177;
wire net_6621;
wire net_2716;
wire net_7902;
wire net_13097;
wire net_7503;
wire net_12717;
wire net_7857;
wire net_11815;
wire net_10015;
wire net_5246;
wire net_351;
wire net_8558;
wire net_6551;
wire net_4750;
wire net_7761;
wire net_13346;
wire net_4558;
wire net_12858;
wire net_12601;
wire net_10856;
wire net_6006;
wire net_4240;
wire net_7964;
wire net_2842;
wire net_8394;
wire net_1257;
wire net_2828;
wire net_3158;
wire net_939;
wire net_12749;
wire net_8365;
wire net_824;
wire net_3458;
wire net_1822;
wire x420;
wire net_13781;
wire net_7984;
wire net_9755;
wire net_14411;
wire net_13038;
wire net_10479;
wire net_1972;
wire net_2791;
wire net_10111;
wire net_11023;
wire net_12267;
wire net_3126;
wire net_993;
wire net_10555;
wire net_8795;
wire net_4271;
wire x561;
wire net_11817;
wire net_9895;
wire net_317;
wire net_856;
wire net_5974;
wire net_11853;
wire net_9456;
wire net_1100;
wire net_7035;
wire net_9944;
wire net_7920;
wire net_3845;
wire net_2817;
wire net_6686;
wire net_2026;
wire net_10046;
wire net_11822;
wire net_5727;
wire net_12195;
wire net_5673;
wire net_5996;
wire net_6730;
wire net_13823;
wire net_1326;
wire net_3033;
wire net_7488;
wire net_134;
wire net_546;
wire net_14059;
wire net_4648;
wire net_3373;
wire net_5382;
wire net_11471;
wire net_2672;
wire net_4546;
wire net_5351;
wire net_588;
wire net_10065;
wire net_13735;
wire net_13320;
wire net_2200;
wire net_8641;
wire net_8062;
wire net_1157;
wire net_12424;
wire net_3701;
wire net_14296;
wire net_4736;
wire net_7486;
wire net_7592;
wire net_7785;
wire net_5592;
wire net_5642;
wire net_4974;
wire net_7906;
wire net_8012;
wire net_3883;
wire net_6001;
wire net_9378;
wire net_1542;
wire net_1172;
wire net_14198;
wire net_9124;
wire net_13703;
wire net_8431;
wire net_4230;
wire net_6350;
wire net_7993;
wire net_9840;
wire net_14270;
wire net_10560;
wire net_11800;
wire net_13604;
wire net_5603;
wire net_9503;
wire net_1065;
wire net_13117;
wire net_4860;
wire net_2237;
wire net_2566;
wire net_8352;
wire net_3795;
wire net_3953;
wire net_13046;
wire net_3100;
wire net_13375;
wire net_241;
wire net_917;
wire net_9353;
wire net_3730;
wire net_13196;
wire net_13640;
wire net_13515;
wire net_12010;
wire net_2874;
wire net_10965;
wire net_8942;
wire net_13350;
wire net_4597;
wire net_13814;
wire net_599;
wire net_9685;
wire net_4589;
wire net_2993;
wire net_10921;
wire net_3067;
wire net_13950;
wire net_10075;
wire net_4844;
wire net_4288;
wire net_5860;
wire net_3111;
wire net_323;
wire net_5402;
wire net_963;
wire net_10301;
wire net_10346;
wire net_11880;
wire net_13543;
wire net_9653;
wire net_13575;
wire net_9482;
wire net_8692;
wire net_8356;
wire net_7368;
wire net_3737;
wire net_4689;
wire net_10216;
wire net_153;
wire net_2389;
wire net_12328;
wire net_6276;
wire net_7556;
wire net_375;
wire net_562;
wire net_6103;
wire net_364;
wire net_8675;
wire net_12260;
wire net_14380;
wire net_12770;
wire net_11723;
wire net_3172;
wire net_10485;
wire net_9686;
wire net_13772;
wire net_11706;
wire net_4239;
wire net_2849;
wire net_14011;
wire net_12671;
wire net_5516;
wire net_7177;
wire net_10799;
wire net_6313;
wire net_12693;
wire net_6341;
wire net_5589;
wire net_8161;
wire net_6840;
wire net_12810;
wire net_4873;
wire net_10851;
wire net_3171;
wire net_4298;
wire net_7514;
wire net_11286;
wire net_14217;
wire net_12742;
wire net_11250;
wire net_7170;
wire net_8004;
wire net_10091;
wire net_1247;
wire net_8173;
wire net_3673;
wire net_4137;
wire net_11149;
wire net_8528;
wire net_2388;
wire net_5162;
wire net_9870;
wire net_14006;
wire net_7561;
wire net_5765;
wire net_3496;
wire net_1215;
wire net_5169;
wire net_5248;
wire net_13361;
wire net_4216;
wire net_129;
wire net_4889;
wire net_10371;
wire net_151;
wire net_13638;
wire net_1625;
wire net_8784;
wire net_284;
wire net_6655;
wire net_9930;
wire net_12743;
wire net_439;
wire net_2513;
wire net_259;
wire net_3582;
wire net_3351;
wire net_4094;
wire net_8662;
wire net_7360;
wire net_7142;
wire net_10291;
wire net_10153;
wire net_3119;
wire net_1231;
wire net_187;
wire net_5841;
wire net_14072;
wire net_3305;
wire net_14045;
wire net_160;
wire net_6205;
wire x1034;
wire net_832;
wire net_12304;
wire net_815;
wire net_7875;
wire net_11304;
wire net_6514;
wire net_6749;
wire net_7728;
wire net_5578;
wire net_13742;
wire net_7670;
wire net_7897;
wire net_5632;
wire net_6501;
wire net_10279;
wire net_586;
wire net_9580;
wire net_10845;
wire net_1347;
wire net_5272;
wire net_1091;
wire net_6240;
wire net_13145;
wire net_3838;
wire net_7812;
wire net_7768;
wire net_11518;
wire net_3745;
wire net_120;
wire net_6260;
wire net_12489;
wire net_292;
wire net_5529;
wire net_11713;
wire net_9879;
wire net_3708;
wire net_12141;
wire net_9384;
wire net_167;
wire net_12371;
wire net_5830;
wire net_5227;
wire net_7536;
wire net_14259;
wire net_7042;
wire net_6073;
wire net_6170;
wire net_7308;
wire net_8864;
wire net_7478;
wire net_9847;
wire net_2556;
wire net_8599;
wire net_3519;
wire net_5735;
wire net_2740;
wire net_2806;
wire net_7294;
wire net_9679;
wire net_672;
wire net_13163;
wire net_4924;
wire net_8834;
wire net_4483;
wire net_8391;
wire net_5212;
wire net_2027;
wire net_9367;
wire net_5045;
wire net_13761;
wire net_11680;
wire net_7021;
wire net_11335;
wire net_6237;
wire net_2456;
wire net_3610;
wire net_2753;
wire net_8963;
wire net_10036;
wire net_1232;
wire net_9585;
wire net_4540;
wire net_5662;
wire net_5784;
wire net_1953;
wire net_3059;
wire net_11625;
wire net_13506;
wire net_10684;
wire net_12540;
wire net_14295;
wire net_3925;
wire net_5444;
wire net_13039;
wire net_464;
wire net_12003;
wire net_3847;
wire net_4473;
wire net_8230;
wire net_4582;
wire net_5699;
wire net_5089;
wire net_4200;
wire net_4547;
wire net_14205;
wire net_5867;
wire net_6300;
wire net_5362;
wire net_7819;
wire net_8954;
wire net_10136;
wire net_4640;
wire net_10926;
wire net_11602;
wire net_4658;
wire net_14195;
wire net_12625;
wire net_1256;
wire net_7071;
wire net_7982;
wire net_13264;
wire net_1413;
wire net_802;
wire net_12194;
wire net_14252;
wire net_3556;
wire net_13872;
wire net_3041;
wire net_1840;
wire net_12930;
wire net_12602;
wire net_4997;
wire net_14359;
wire net_9230;
wire net_6620;
wire net_5637;
wire net_8015;
wire net_3427;
wire net_7167;
wire net_1031;
wire net_4824;
wire net_13170;
wire net_7049;
wire net_14189;
wire net_13404;
wire net_1636;
wire net_7568;
wire net_9714;
wire net_3257;
wire net_10265;
wire net_13394;
wire net_4458;
wire net_7245;
wire net_10899;
wire net_9744;
wire net_7458;
wire net_10467;
wire net_10344;
wire net_10270;
wire net_10991;
wire net_1334;
wire net_10782;
wire net_757;
wire net_206;
wire net_8523;
wire net_2020;
wire net_1688;
wire net_10087;
wire net_13522;
wire net_10794;
wire net_13383;
wire net_10894;
wire net_7665;
wire net_14134;
wire net_235;
wire net_6126;
wire net_14056;
wire net_13121;
wire net_11695;
wire net_12223;
wire net_2961;
wire x1486;
wire net_4159;
wire net_4324;
wire net_5108;
wire net_2374;
wire net_7322;
wire net_9911;
wire net_4203;
wire net_7652;
wire net_5631;
wire net_3644;
wire net_10571;
wire net_12273;
wire net_250;
wire net_3600;
wire net_8655;
wire net_7260;
wire net_3081;
wire net_5882;
wire net_12927;
wire net_11279;
wire x1501;
wire net_2055;
wire net_10283;
wire net_4879;
wire net_6144;
wire net_12929;
wire net_2630;
wire net_7420;
wire net_10027;
wire net_1985;
wire net_403;
wire net_3524;
wire net_2340;
wire net_6265;
wire net_13680;
wire net_12219;
wire net_2275;
wire net_14302;
wire net_10752;
wire net_3976;
wire net_9619;
wire net_9899;
wire net_10939;
wire net_12562;
wire net_12202;
wire net_8602;
wire net_13128;
wire net_841;
wire net_10803;
wire net_1750;
wire net_6411;
wire net_794;
wire net_2397;
wire net_3346;
wire net_13277;
wire net_8136;
wire net_8269;
wire net_528;
wire net_10537;
wire net_3433;
wire net_335;
wire net_4878;
wire net_3464;
wire net_1468;
wire net_9132;
wire net_181;
wire net_9661;
wire net_4774;
wire net_6784;
wire net_11767;
wire net_12214;
wire net_3333;
wire net_11556;
wire net_6011;
wire net_10631;
wire net_9014;
wire net_8494;
wire net_7350;
wire net_13530;
wire net_6177;
wire net_6796;
wire net_3649;
wire net_2539;
wire net_1130;
wire net_5921;
wire net_6216;
wire net_8111;
wire net_386;
wire net_12680;
wire net_9421;
wire net_8239;
wire net_6150;
wire net_10051;
wire net_1790;
wire net_6451;
wire net_7918;
wire net_4103;
wire net_6493;
wire net_8166;
wire net_9281;
wire net_11221;
wire net_6130;
wire net_6309;
wire net_7745;
wire net_2318;
wire net_8787;
wire net_9207;
wire net_5562;
wire net_3449;
wire net_10583;
wire net_9134;
wire net_9004;
wire net_12718;
wire net_1039;
wire net_7573;
wire net_1709;
wire net_11972;
wire net_7822;
wire net_10981;
wire net_8629;
wire net_400;
wire net_4651;
wire net_10080;
wire net_9698;
wire net_1935;
wire net_5707;
wire net_11608;
wire net_13622;
wire net_175;
wire net_13102;
wire net_12650;
wire net_2925;
wire net_1850;
wire net_11873;
wire net_9142;
wire net_4429;
wire net_1855;
wire net_4882;
wire net_6365;
wire net_1992;
wire net_1177;
wire net_1163;
wire net_12346;
wire net_897;
wire net_7384;
wire net_13890;
wire net_11362;
wire net_10206;
wire net_5466;
wire net_9521;
wire net_2853;
wire net_10578;
wire net_2705;
wire net_7840;
wire net_5164;
wire net_9215;
wire net_615;
wire net_6712;
wire net_11494;
wire net_3273;
wire net_1559;
wire net_441;
wire net_8706;
wire net_5665;
wire net_1620;
wire net_13966;
wire net_2608;
wire net_14266;
wire net_14224;
wire net_6032;
wire net_9763;
wire net_2813;
wire net_2663;
wire net_728;
wire net_1276;
wire net_5473;
wire net_719;
wire net_7774;
wire net_10878;
wire net_170;
wire net_6873;
wire net_8068;
wire net_14032;
wire net_2571;
wire net_9888;
wire x14;
wire net_5305;
wire net_10741;
wire net_5703;
wire net_12264;
wire net_9418;
wire net_14325;
wire net_3479;
wire net_8609;
wire net_13617;
wire net_3222;
wire net_3321;
wire net_6393;
wire net_13764;
wire net_8410;
wire net_708;
wire net_3552;
wire net_696;
wire net_7685;
wire net_14079;
wire net_10824;
wire net_10777;
wire net_3216;
wire net_5713;
wire net_7427;
wire net_13175;
wire net_13947;
wire net_10401;
wire net_12972;
wire net_12256;
wire net_171;
wire net_10448;
wire net_9953;
wire net_9796;
wire net_10013;
wire net_6563;
wire net_3821;
wire net_9228;
wire net_10528;
wire net_604;
wire net_14101;
wire net_8403;
wire net_4503;
wire net_10872;
wire net_12385;
wire net_6938;
wire net_3486;
wire net_483;
wire net_7359;
wire net_1149;
wire net_9937;
wire net_8097;
wire net_5839;
wire net_7955;
wire net_11199;
wire net_8590;
wire net_8919;
wire net_9981;
wire net_8302;
wire net_1298;
wire net_296;
wire net_2131;
wire net_6681;
wire net_9733;
wire x315;
wire net_5651;
wire net_13461;
wire net_12845;
wire net_12053;
wire net_7004;
wire net_7153;
wire net_13632;
wire net_8941;
wire net_5435;
wire net_11369;
wire net_11461;
wire net_2228;
wire net_12357;
wire net_3020;
wire net_13720;
wire net_786;
wire net_5141;
wire net_11801;
wire net_11564;
wire net_8998;
wire net_9470;
wire net_127;
wire net_10518;
wire net_1339;
wire net_10608;
wire net_3781;
wire net_5685;
wire net_906;
wire net_9892;
wire net_9080;
wire net_8461;
wire net_2422;
wire net_5205;
wire net_3577;
wire net_13951;
wire net_10185;
wire net_652;
wire net_12955;
wire net_13958;
wire net_10137;
wire net_13707;
wire net_3840;
wire net_1815;
wire net_4361;
wire net_10590;
wire net_10211;
wire net_6145;
wire net_3782;
wire net_13250;
wire net_2505;
wire net_11185;
wire net_877;
wire net_2799;
wire net_10748;
wire net_6139;
wire net_6868;
wire net_6834;
wire net_3734;
wire net_8092;
wire net_14135;
wire net_2683;
wire net_8021;
wire net_4812;
wire net_9654;
wire net_2165;
wire net_4253;
wire net_11943;
wire net_11570;
wire net_11232;
wire net_8315;
wire net_4066;
wire net_13296;
wire net_6257;
wire net_3284;
wire net_8026;
wire net_1474;
wire net_4297;
wire net_12088;
wire net_2784;
wire net_6861;
wire net_11049;
wire net_13843;
wire net_8753;
wire net_675;
wire net_2562;
wire net_8355;
wire net_2867;
wire net_5134;
wire net_9129;
wire net_5293;
wire net_7195;
wire net_13841;
wire net_3472;
wire x620;
wire net_9120;
wire net_10700;
wire net_7578;
wire net_8151;
wire net_5172;
wire net_10092;
wire net_2182;
wire net_1768;
wire net_8145;
wire net_9928;
wire net_4718;
wire net_8032;
wire net_9295;
wire net_150;
wire net_12950;
wire net_6589;
wire net_7677;
wire net_11915;
wire net_304;
wire net_4351;
wire net_6993;
wire net_10951;
wire net_12436;
wire net_9791;
wire net_7326;
wire net_4347;
wire net_7666;
wire net_12768;
wire net_10551;
wire net_1703;
wire net_11004;
wire net_7848;
wire net_9420;
wire net_7731;
wire net_9690;
wire net_3693;
wire net_12731;
wire net_9027;
wire net_5100;
wire net_1316;
wire net_6845;
wire net_6545;
wire net_4319;
wire net_792;
wire net_13848;
wire net_13695;
wire net_3070;
wire net_6223;
wire net_13782;
wire net_8842;
wire net_3409;
wire net_9481;
wire net_2203;
wire net_4430;
wire net_13415;
wire net_5373;
wire net_4525;
wire net_1904;
wire net_9446;
wire net_3907;
wire net_5678;
wire net_6332;
wire net_219;
wire net_3609;
wire net_10001;
wire net_6584;
wire net_8617;
wire net_9976;
wire net_2187;
wire net_2476;
wire net_13798;
wire net_913;
wire net_10764;
wire net_4518;
wire net_5378;
wire net_5338;
wire net_13242;
wire net_3387;
wire net_13591;
wire net_1479;
wire net_7157;
wire net_4330;
wire net_7756;
wire net_10268;
wire net_4019;
wire net_4152;
wire net_6895;
wire net_10066;
wire net_10832;
wire net_3094;
wire net_360;
wire net_13561;
wire net_1927;
wire net_7017;
wire net_10243;
wire net_213;
wire net_6910;
wire net_2324;
wire net_11688;
wire net_9244;
wire net_947;
wire net_4805;
wire net_5359;
wire net_7970;
wire net_1126;
wire net_11538;
wire net_2004;
wire net_13259;
wire net_1325;
wire net_6943;
wire net_3316;
wire net_10162;
wire net_3032;
wire net_9507;
wire net_5094;
wire net_6298;
wire net_1373;
wire net_1352;
wire net_2885;
wire net_2567;
wire net_10735;
wire net_10258;
wire net_4696;
wire net_8814;
wire net_14029;
wire net_10944;
wire net_1187;
wire net_7643;
wire net_7408;
wire net_7411;
wire net_4988;
wire net_3206;
wire net_1303;
wire net_8050;
wire net_2858;
wire net_6334;
wire net_2102;
wire net_4451;
wire net_5569;
wire net_12234;
wire net_12047;
wire net_1442;
wire net_11903;
wire net_1807;
wire net_10042;
wire net_1943;
wire net_1930;
wire net_11544;
wire net_12298;
wire net_1894;
wire net_12113;
wire net_9645;
wire net_10694;
wire net_2431;
wire net_11555;
wire net_4054;
wire net_5544;
wire net_8213;
wire net_633;
wire net_113;
wire net_5054;
wire net_5750;
wire net_10115;
wire net_9674;
wire net_4848;
wire net_1914;
wire net_7791;
wire net_2408;
wire net_3889;
wire net_9904;
wire net_6627;
wire net_5943;
wire net_14039;
wire net_6974;
wire net_3567;
wire net_13717;
wire net_7831;
wire net_1457;
wire net_11525;
wire net_2741;
wire net_7010;
wire net_5414;
wire net_6483;
wire net_4011;
wire net_6616;
wire net_2448;
wire net_1436;
wire net_5424;
wire net_5541;
wire net_9199;
wire net_4338;
wire net_13234;
wire net_10719;
wire net_10054;
wire net_3400;
wire net_10725;
wire net_3392;
wire net_9571;
wire net_2551;
wire net_11572;
wire net_646;
wire net_12547;
wire net_2731;
wire net_5823;
wire net_14348;
wire net_11016;
wire net_2601;
wire net_6323;
wire net_8902;
wire net_2891;
wire net_8499;
wire net_520;
wire net_14314;
wire net_13482;
wire net_10159;
wire net_11201;
wire net_8928;
wire net_7237;
wire net_11261;
wire net_4722;
wire net_14110;
wire net_3231;
wire net_981;
wire net_2401;
wire x234;
wire net_9636;
wire net_8895;
wire net_1566;
wire net_1305;
wire net_11584;
wire net_2354;
wire net_12156;
wire net_9393;
wire net_1387;
wire net_1581;
wire net_10709;
wire net_10378;
wire net_10440;
wire net_8858;
wire net_5018;
wire net_7369;
wire net_11808;
wire net_4468;
wire net_2413;
wire net_5013;
wire net_7786;
wire net_11413;
wire net_559;
wire net_3042;
wire net_2792;
wire net_345;
wire net_2965;
wire net_2128;
wire net_12804;
wire net_1717;
wire net_7476;
wire net_9990;
wire net_11891;
wire net_6553;
wire net_398;
wire net_5302;
wire net_3399;
wire net_6976;
wire net_11489;
wire net_9344;
wire net_5080;
wire net_6693;
wire net_11140;
wire net_13584;
wire net_12834;
wire net_2117;
wire net_2461;
wire net_4085;
wire net_1766;
wire net_13493;
wire net_7393;
wire net_2582;
wire net_10099;
wire net_8974;
wire net_12472;
wire net_7898;
wire net_5905;
wire net_9788;
wire net_6724;
wire net_10419;
wire net_3872;
wire net_4956;
wire net_6054;
wire net_11867;
wire net_1572;
wire net_9407;
wire net_4447;
wire net_10357;
wire net_11647;
wire net_10226;
wire net_9265;
wire net_13933;
wire net_9235;
wire net_8990;
wire net_2134;
wire net_5179;
wire net_14166;
wire net_8794;
wire net_9834;
wire net_316;
wire net_5011;
wire net_13439;
wire net_4250;
wire net_4961;
wire net_4184;
wire net_11462;
wire net_12667;
wire net_14398;
wire net_13536;
wire net_13443;
wire net_10387;
wire net_1759;
wire net_12996;
wire net_7033;
wire net_12752;
wire net_3764;
wire net_4647;
wire net_12964;
wire net_4022;
wire net_11636;
wire net_2541;
wire net_12310;
wire net_9618;
wire net_3689;
wire net_12635;
wire net_533;
wire net_7436;
wire net_13282;
wire net_8347;
wire net_10040;
wire net_1695;
wire net_5932;
wire net_911;
wire net_1617;
wire net_7775;
wire net_12017;
wire net_7005;
wire net_10047;
wire net_9608;
wire net_6637;
wire net_9015;
wire net_7053;
wire net_5969;
wire net_5570;
wire net_9332;
wire net_11745;
wire net_9457;
wire net_568;
wire net_4579;
wire net_13709;
wire net_13809;
wire net_7962;
wire net_4807;
wire net_1227;
wire net_6046;
wire net_6485;
wire net_1008;
wire net_5312;
wire net_5340;
wire net_5861;
wire net_1443;
wire net_12178;
wire net_11888;
wire net_3069;
wire net_4862;
wire net_8691;
wire net_3170;
wire net_12239;
wire net_2840;
wire net_3463;
wire net_4005;
wire net_6008;
wire net_4819;
wire net_11883;
wire net_3199;
wire net_3597;
wire net_5671;
wire net_8001;
wire net_269;
wire net_5043;
wire net_3193;
wire net_3131;
wire net_469;
wire net_10107;
wire net_12171;
wire net_3179;
wire net_1978;
wire net_1945;
wire net_10064;
wire net_7207;
wire net_10858;
wire net_3167;
wire net_4073;
wire net_5159;
wire net_1170;
wire net_1833;
wire net_5656;
wire net_10144;
wire net_8496;
wire net_13202;
wire net_2280;
wire net_2831;
wire net_9174;
wire net_3029;
wire net_9622;
wire net_2366;
wire net_778;
wire net_7818;
wire net_5725;
wire net_12779;
wire net_2930;
wire net_1455;
wire net_9816;
wire net_8252;
wire net_6523;
wire net_14277;
wire net_5064;
wire net_5323;
wire net_6024;
wire net_12167;
wire net_6225;
wire net_11780;
wire net_6832;
wire net_5261;
wire net_4730;
wire net_12154;
wire net_6643;
wire net_11123;
wire net_8172;
wire net_7912;
wire net_5380;
wire net_10173;
wire net_8519;
wire net_4119;
wire net_5648;
wire net_14246;
wire net_11152;
wire net_13445;
wire net_11251;
wire net_9450;
wire net_9216;
wire net_10644;
wire net_3980;
wire net_10566;
wire net_10335;
wire net_1481;
wire net_10392;
wire net_995;
wire net_5645;
wire net_7922;
wire net_8328;
wire net_7088;
wire net_700;
wire net_5000;
wire net_12232;
wire net_7334;
wire net_11433;
wire net_9947;
wire net_8957;
wire net_1246;
wire net_13325;
wire net_11043;
wire net_6043;
wire net_7705;
wire net_5216;
wire net_1774;
wire net_4228;
wire net_11402;
wire net_11819;
wire net_1673;
wire net_3060;
wire net_10712;
wire net_2568;
wire net_11103;
wire net_11941;
wire net_3480;
wire net_321;
wire net_6715;
wire net_9465;
wire net_8933;
wire net_5518;
wire net_4135;
wire net_2995;
wire net_6982;
wire net_3526;
wire net_2945;
wire net_934;
wire net_3103;
wire net_12855;
wire net_5941;
wire net_3665;
wire net_544;
wire net_717;
wire net_4896;
wire net_12305;
wire net_10505;
wire net_8201;
wire net_11952;
wire net_3630;
wire net_1824;
wire net_12037;
wire net_9659;
wire net_3402;
wire net_2223;
wire net_7603;
wire net_4763;
wire net_5074;
wire net_6957;
wire net_2673;
wire net_5694;
wire net_8008;
wire net_3500;
wire net_6164;
wire net_3166;
wire net_9104;
wire net_7065;
wire net_10861;
wire net_9831;
wire net_9358;
wire net_5903;
wire net_8079;
wire net_7513;
wire net_10665;
wire net_9652;
wire net_1245;
wire net_5552;
wire net_3660;
wire net_860;
wire net_5806;
wire net_870;
wire net_9254;
wire net_7135;
wire net_2046;
wire net_7176;
wire net_11708;
wire net_7521;
wire net_7926;
wire net_10819;
wire net_7941;
wire net_2878;
wire net_2871;
wire net_13642;
wire net_12012;
wire net_9850;
wire net_3267;
wire net_2321;
wire net_6286;
wire net_9108;
wire net_12874;
wire net_12668;
wire net_11645;
wire net_817;
wire net_11667;
wire net_5127;
wire net_3414;
wire x1345;
wire net_7058;
wire net_14155;
wire net_10922;
wire net_10967;
wire net_7362;
wire net_14084;
wire net_13502;
wire net_9766;
wire net_4576;
wire net_13655;
wire net_2920;
wire net_1591;
wire net_14123;
wire net_13344;
wire net_7695;
wire net_13278;
wire net_1747;
wire net_5483;
wire net_2012;
wire net_650;
wire net_7139;
wire net_9761;
wire net_5557;
wire net_597;
wire net_9890;
wire net_14065;
wire net_743;
wire net_14387;
wire net_3770;
wire net_9062;
wire net_1922;
wire net_5984;
wire net_10482;
wire net_8272;
wire net_14281;
wire net_6336;
wire net_12481;
wire net_8889;
wire net_10853;
wire net_12384;
wire net_603;
wire net_6639;
wire net_8264;
wire net_4913;
wire net_13499;
wire net_2451;
wire net_14332;
wire net_642;
wire net_9806;
wire net_2699;
wire net_1522;
wire net_4031;
wire net_1158;
wire net_6989;
wire net_11496;
wire net_2926;
wire net_8006;
wire net_11082;
wire net_10775;
wire net_12782;
wire net_11530;
wire net_13964;
wire net_12289;
wire net_8042;
wire net_470;
wire net_13751;
wire net_2702;
wire net_430;
wire net_6991;
wire net_2834;
wire net_11659;
wire net_4551;
wire net_5972;
wire net_13557;
wire net_12945;
wire net_3943;
wire net_9370;
wire net_3129;
wire net_4438;
wire net_7675;
wire net_8568;
wire net_12353;
wire net_10839;
wire net_14154;
wire net_8557;
wire net_11771;
wire net_1063;
wire net_4218;
wire net_968;
wire net_13876;
wire net_13572;
wire net_9669;
wire net_12692;
wire net_10421;
wire net_12571;
wire net_9127;
wire net_2534;
wire net_6827;
wire net_7297;
wire net_4133;
wire net_13577;
wire net_1504;
wire net_475;
wire net_6737;
wire net_9432;
wire net_7216;
wire net_14272;
wire net_11137;
wire net_3732;
wire net_14024;
wire net_13768;
wire net_6903;
wire net_2309;
wire net_502;
wire net_8647;
wire net_2470;
wire net_1564;
wire net_11474;
wire net_1568;
wire net_6632;
wire net_14288;
wire net_12282;
wire net_3804;
wire net_10883;
wire net_6756;
wire net_9398;
wire net_1526;
wire net_13271;
wire net_13860;
wire net_8290;
wire net_1884;
wire net_12341;
wire net_12209;
wire net_13858;
wire net_3919;
wire net_7990;
wire net_4112;
wire net_2646;
wire net_3868;
wire net_3936;
wire net_7121;
wire net_4364;
wire net_13198;
wire net_5887;
wire net_6645;
wire net_13233;
wire net_2628;
wire net_4512;
wire net_6535;
wire net_9305;
wire net_11692;
wire net_5145;
wire net_12757;
wire net_11439;
wire net_11160;
wire net_1360;
wire net_6344;
wire net_10494;
wire net_9047;
wire net_3364;
wire net_11078;
wire net_13837;
wire net_13800;
wire net_5316;
wire net_664;
wire net_1364;
wire net_6003;
wire net_5050;
wire net_6292;
wire net_4622;
wire net_549;
wire net_827;
wire net_4605;
wire net_10192;
wire net_11050;
wire net_10450;
wire net_4295;
wire net_10687;
wire net_4563;
wire net_2337;
wire net_12533;
wire net_6945;
wire net_1369;
wire net_10614;
wire net_5773;
wire net_6900;
wire net_6405;
wire net_11068;
wire net_4695;
wire net_13550;
wire net_7469;
wire net_8622;
wire x1231;
wire net_1013;
wire net_1530;
wire net_6210;
wire net_13869;
wire net_3075;
wire net_2952;
wire net_842;
wire net_11783;
wire net_2336;
wire net_1705;
wire net_2035;
wire net_6571;
wire net_9500;
wire net_11215;
wire net_8951;
wire net_5070;
wire net_2826;
wire net_6560;
wire net_10325;
wire net_8199;
wire net_3739;
wire net_10451;
wire net_8455;
wire net_492;
wire net_11392;
wire net_3678;
wire net_6847;
wire net_2141;
wire net_7234;
wire net_8797;
wire net_2639;
wire net_14211;
wire net_10830;
wire net_8071;
wire net_11803;
wire net_13370;
wire net_11213;
wire net_3695;
wire net_3453;
wire net_12648;
wire net_5450;
wire net_5702;
wire net_1327;
wire net_8632;
wire net_10598;
wire net_9822;
wire net_4968;
wire net_1403;
wire net_6097;
wire net_4532;
wire net_12734;
wire net_2248;
wire net_2270;
wire net_1667;
wire net_4971;
wire net_11532;
wire net_7208;
wire net_3866;
wire net_8882;
wire net_1606;
wire x397;
wire net_6772;
wire net_3710;
wire net_13473;
wire net_7787;
wire net_13223;
wire net_12024;
wire net_3054;
wire net_12920;
wire net_4300;
wire net_9578;
wire net_7683;
wire net_4776;
wire net_8765;
wire net_3978;
wire net_10477;
wire net_4752;
wire net_12708;
wire net_13820;
wire net_2868;
wire net_2029;
wire net_6083;
wire net_5328;
wire net_3698;
wire net_8295;
wire net_11560;
wire net_4629;
wire net_2946;
wire net_2587;
wire net_11373;
wire net_1284;
wire net_4397;
wire net_2959;
wire net_13977;
wire net_13732;
wire net_11836;
wire net_1888;
wire net_13095;
wire net_6671;
wire net_9974;
wire net_4311;
wire net_3929;
wire net_9942;
wire net_12583;
wire net_1792;
wire net_2496;
wire net_4125;
wire net_13888;
wire net_7567;
wire net_10656;
wire net_3109;
wire net_2066;
wire net_13925;
wire net_9310;
wire net_1598;
wire net_7415;
wire net_14192;
wire net_14369;
wire net_731;
wire net_8109;
wire net_1146;
wire net_13042;
wire net_11679;
wire net_4612;
wire net_9704;
wire net_7287;
wire net_1733;
wire net_4519;
wire net_10576;
wire net_8584;
wire net_5853;
wire net_5511;
wire net_13881;
wire net_7590;
wire net_13962;
wire net_9897;
wire net_11093;
wire net_6708;
wire net_5495;
wire net_10412;
wire net_13071;
wire net_9511;
wire net_8284;
wire net_2762;
wire net_4146;
wire net_11828;
wire net_1724;
wire net_6106;
wire net_6439;
wire net_3703;
wire net_12551;
wire net_6247;
wire net_6424;
wire x657;
wire net_4619;
wire net_6377;
wire net_12682;
wire net_10161;
wire net_2089;
wire net_12506;
wire net_6352;
wire net_10843;
wire net_12429;
wire net_965;
wire net_12378;
wire net_3797;
wire net_9718;
wire net_3535;
wire net_12248;
wire net_1195;
wire net_2916;
wire net_11976;
wire net_8314;
wire net_421;
wire net_5348;
wire net_8184;
wire net_2502;
wire net_1396;
wire net_1104;
wire net_9783;
wire net_4069;
wire net_764;
wire net_4060;
wire net_7225;
wire net_13009;
wire net_5181;
wire net_2737;
wire net_6397;
wire net_5126;
wire net_5038;
wire net_12108;
wire net_2481;
wire net_12465;
wire net_4539;
wire net_1117;
wire net_7289;
wire net_13534;
wire net_10624;
wire x101;
wire net_6866;
wire net_7162;
wire net_13770;
wire net_3955;
wire net_8104;
wire net_14210;
wire net_2617;
wire net_1060;
wire net_5950;
wire net_12699;
wire net_11893;
wire net_8246;
wire net_9157;
wire net_4846;
wire x494;
wire net_5503;
wire net_7252;
wire net_8303;
wire net_2235;
wire net_11007;
wire net_12101;
wire net_11329;
wire net_1715;
wire net_5846;
wire net_2080;
wire net_3675;
wire net_9913;
wire net_2711;
wire net_6714;
wire net_2097;
wire net_7583;
wire net_9234;
wire net_6194;
wire net_11120;
wire net_6577;
wire net_3619;
wire net_1216;
wire net_4599;
wire net_2815;
wire net_3785;
wire net_11240;
wire net_1271;
wire net_1086;
wire net_1782;
wire net_9593;
wire net_10978;
wire net_11191;
wire net_8450;
wire net_13453;
wire net_1197;
wire net_7613;
wire net_1278;
wire net_273;
wire net_4863;
wire net_5744;
wire net_5858;
wire net_11752;
wire net_4714;
wire net_6430;
wire net_3182;
wire net_576;
wire net_8932;
wire net_1654;
wire net_12643;
wire net_2098;
wire net_3355;
wire net_177;
wire net_4232;
wire net_8438;
wire net_3005;
wire net_4305;
wire net_11183;
wire net_7806;
wire net_12902;
wire net_8739;
wire net_10679;
wire net_2803;
wire net_3301;
wire net_11272;
wire net_725;
wire net_12133;
wire net_6370;
wire net_3931;
wire net_6090;
wire net_953;
wire net_6183;
wire net_11600;
wire net_11171;
wire net_894;
wire net_1074;
wire net_13914;
wire net_10545;
wire net_1058;
wire net_7186;
wire net_12728;
wire net_11295;
wire net_9535;
wire net_1423;
wire net_13012;
wire net_2902;
wire net_1871;
wire net_517;
wire net_628;
wire net_14004;
wire net_9064;
wire x1215;
wire net_6159;
wire net_3494;
wire net_2489;
wire net_6962;
wire net_6600;
wire net_12123;
wire net_10377;
wire net_14018;
wire net_10204;
wire net_9555;
wire net_9036;
wire net_13829;
wire net_3160;
wire net_2125;
wire net_7622;
wire net_6406;
wire net_10322;
wire net_8179;
wire net_1289;
wire net_9546;
wire net_13078;
wire net_3138;
wire net_11982;
wire net_2623;
wire net_13377;
wire net_8448;
wire net_261;
wire net_10654;
wire net_12867;
wire net_2362;
wire net_6922;
wire net_12837;
wire net_11162;
wire net_5895;
wire net_8869;
wire net_12446;
wire net_4456;
wire net_5876;
wire net_4354;
wire net_1955;
wire net_5111;
wire net_2723;
wire net_5157;
wire net_13504;
wire net_2552;
wire net_8507;
wire net_3229;
wire net_1001;
wire net_8196;
wire net_13778;
wire net_3765;
wire net_781;
wire net_12886;
wire net_8479;
wire net_9729;
wire net_13063;
wire net_5241;
wire net_7506;
wire net_3012;
wire net_5967;
wire net_13134;
wire net_6818;
wire net_13188;
wire net_6014;
wire net_5367;
wire net_3754;
wire net_10432;
wire net_185;
wire net_7357;
wire net_6075;
wire net_9935;
wire net_11356;
wire net_3989;
wire net_13902;
wire net_10515;
wire net_7304;
wire net_11312;
wire net_10875;
wire net_4321;
wire net_4631;
wire net_5285;
wire net_1994;
wire net_1015;
wire net_10499;
wire net_2980;
wire net_8574;
wire net_4668;
wire net_3897;
wire net_9863;
wire net_9288;
wire net_3960;
wire net_4374;
wire net_3992;
wire net_6152;
wire net_9772;
wire net_2287;
wire net_4211;
wire net_11964;
wire net_5794;
wire net_448;
wire net_8224;
wire net_886;
wire net_7766;
wire net_3189;
wire net_11759;
wire net_6856;
wire net_2988;
wire net_2146;
wire net_405;
wire net_11927;
wire net_6811;
wire net_1111;
wire net_4592;
wire net_11614;
wire net_2651;
wire net_4281;
wire net_8259;
wire net_5279;
wire net_3651;
wire net_3971;
wire net_12182;
wire net_3155;
wire net_14345;
wire net_9059;
wire net_11440;
wire net_1470;
wire net_7969;
wire net_14053;
wire net_13358;
wire net_4627;
wire net_4423;
wire net_831;
wire net_4728;
wire net_5442;
wire net_451;
wire net_13674;
wire net_4233;
wire net_1234;
wire net_750;
wire net_12558;
wire net_4796;
wire net_7650;
wire net_8289;
wire net_7835;
wire net_9746;
wire net_13662;
wire net_2778;
wire net_2756;
wire net_12896;
wire net_13027;
wire net_12797;
wire net_7274;
wire net_11459;
wire net_9605;
wire net_8571;
wire net_1085;
wire net_5915;
wire net_5184;
wire net_592;
wire net_9528;
wire net_8983;
wire net_5788;
wire net_11920;
wire net_8472;
wire net_773;
wire net_4759;
wire net_7531;
wire net_2266;
wire net_11770;
wire net_281;
wire net_9590;
wire net_12493;
wire net_8337;
wire net_5254;
wire net_5193;
wire net_11796;
wire net_11622;
wire net_5235;
wire net_8537;
wire net_12098;
wire net_3727;
wire net_13986;
wire net_5520;
wire net_6766;
wire net_13269;
wire net_6355;
wire net_5052;
wire net_14400;
wire net_9997;
wire net_10801;
wire net_13532;
wire net_10281;
wire net_8305;
wire net_14091;
wire net_4205;
wire net_526;
wire net_2718;
wire net_834;
wire net_10298;
wire net_694;
wire net_13123;
wire net_13615;
wire net_13556;
wire net_2747;
wire net_13794;
wire net_5925;
wire net_14365;
wire net_9950;
wire net_7609;
wire net_12271;
wire net_9232;
wire net_8778;
wire net_8946;
wire net_8409;
wire net_974;
wire net_1570;
wire net_12348;
wire net_13385;
wire net_4645;
wire net_11777;
wire net_11100;
wire net_13853;
wire net_923;
wire net_10947;
wire net_1707;
wire net_12204;
wire net_9499;
wire net_2190;
wire net_4566;
wire net_1881;
wire net_11228;
wire net_7014;
wire net_10487;
wire net_7320;
wire net_10900;
wire net_12925;
wire net_8779;
wire net_124;
wire net_252;
wire net_10497;
wire net_3323;
wire net_11697;
wire net_6347;
wire net_7693;
wire net_7867;
wire net_2399;
wire net_11073;
wire net_8961;
wire net_901;
wire net_6267;
wire net_7846;
wire net_3425;
wire net_12221;
wire net_410;
wire net_1492;
wire net_8134;
wire x138;
wire net_14312;
wire net_4243;
wire net_6179;
wire net_10585;
wire net_10539;
wire net_6363;
wire net_9275;
wire net_8267;
wire net_9136;
wire net_2537;
wire net_11088;
wire net_6798;
wire net_6607;
wire net_3767;
wire net_6919;
wire net_12470;
wire net_6408;
wire net_7886;
wire net_4105;
wire net_11984;
wire net_11397;
wire net_2603;
wire net_5910;
wire net_7824;
wire net_1132;
wire net_5594;
wire net_14144;
wire net_5880;
wire net_6132;
wire net_10351;
wire net_9553;
wire net_9193;
wire net_2442;
wire net_4569;
wire net_5754;
wire net_3026;
wire net_7743;
wire net_13749;
wire net_12317;
wire net_9410;
wire net_5760;
wire x538;
wire net_5923;
wire net_13000;
wire net_2356;
wire net_3288;
wire net_971;
wire net_6214;
wire net_9798;
wire net_11558;
wire net_2273;
wire net_2049;
wire net_8194;
wire net_617;
wire net_11734;
wire net_11026;
wire net_2184;
wire net_6030;
wire net_13456;
wire net_11824;
wire net_8656;
wire net_554;
wire net_13625;
wire net_4176;
wire net_4653;
wire net_14232;
wire net_11187;
wire net_8704;
wire net_3740;
wire net_14221;
wire net_8317;
wire net_4032;
wire net_4154;
wire net_9294;
wire net_6306;
wire net_9413;
wire net_584;
wire net_13753;
wire net_10446;
wire net_12656;
wire net_10420;
wire net_9794;
wire net_7877;
wire net_9000;
wire net_5917;
wire net_3870;
wire net_2411;
wire net_5709;
wire net_6254;
wire net_13104;
wire net_11511;
wire net_5456;
wire net_165;
wire net_9226;
wire net_7105;
wire net_8310;
wire net_3438;
wire net_5946;
wire net_3824;
wire net_11662;
wire net_8789;
wire net_8742;
wire net_4440;
wire net_6854;
wire net_14132;
wire net_12216;
wire net_8576;
wire net_13766;
wire net_10082;
wire net_13612;
wire net_10170;
wire net_384;
wire net_12970;
wire net_3823;
wire net_9886;
wire net_4191;
wire net_8600;
wire net_3503;
wire net_5792;
wire net_9365;
wire net_13573;
wire net_13366;
wire net_3859;
wire net_2599;
wire net_8044;
wire net_2665;
wire net_9200;
wire net_3642;
wire net_7885;
wire net_3803;
wire net_2707;
wire net_8607;
wire net_7426;
wire net_11284;
wire net_485;
wire net_14338;
wire net_11179;
wire net_8880;
wire net_8592;
wire net_7707;
wire net_3334;
wire net_6789;
wire net_3224;
wire net_7772;
wire net_1719;
wire net_7348;
wire net_11364;
wire net_5715;
wire net_11562;
wire net_11589;
wire net_11081;
wire net_125;
wire net_11464;
wire net_9329;
wire net_13402;
wire net_8786;
wire net_8034;
wire net_11598;
wire net_2440;
wire net_1685;
wire net_9386;
wire net_6809;
wire net_14043;
wire net_12800;
wire net_4768;
wire net_1379;
wire net_1322;
wire net_12019;
wire net_14239;
wire net_13147;
wire net_2644;
wire net_6102;
wire net_12815;
wire net_9538;
wire net_13093;
wire net_8526;
wire net_12143;
wire net_10373;
wire net_1301;
wire net_12066;
wire net_14258;
wire net_12686;
wire net_286;
wire net_11668;
wire net_12487;
wire net_8749;
wire net_7596;
wire net_3584;
wire net_12756;
wire net_7051;
wire net_7247;
wire net_11591;
wire net_5588;
wire net_6932;
wire net_4999;
wire net_7116;
wire net_426;
wire net_5203;
wire net_10275;
wire net_4340;
wire net_4954;
wire net_6095;
wire net_414;
wire net_5878;
wire net_10277;
wire net_7793;
wire net_1048;
wire net_3048;
wire net_799;
wire net_5102;
wire net_3475;
wire net_8423;
wire net_5576;
wire net_14142;
wire net_5832;
wire net_5737;
wire net_12588;
wire net_2014;
wire net_9070;
wire net_8232;
wire net_12608;
wire net_1951;
wire net_7292;
wire net_12724;
wire net_9759;
wire net_8976;
wire x379;
wire net_6747;
wire net_13487;
wire net_5999;
wire net_7661;
wire net_12000;
wire net_11869;
wire net_9845;
wire net_5567;
wire net_2558;
wire net_4742;
wire net_2454;
wire net_8917;
wire net_8716;
wire net_2040;
wire net_1508;
wire net_3379;
wire net_4761;
wire net_931;
wire net_4466;
wire net_5983;
wire net_2242;
wire net_8505;
wire net_7672;
wire net_759;
wire net_6802;
wire net_7616;
wire net_6016;
wire net_7852;
wire net_11711;
wire net_11155;
wire net_8832;
wire net_10140;
wire net_12621;
wire net_247;
wire net_8083;
wire net_6428;
wire net_6742;
wire net_5242;
wire net_12573;
wire net_3413;
wire net_6516;
wire net_6924;
wire net_9742;
wire net_8619;
wire net_1341;
wire net_12627;
wire net_4541;
wire net_1934;
wire net_5210;
wire net_14180;
wire net_3242;
wire net_8138;
wire net_1835;
wire net_13740;
wire net_12513;
wire net_6235;
wire net_11327;
wire net_1848;
wire net_333;
wire net_639;
wire net_4724;
wire net_9583;
wire net_9322;
wire net_9114;
wire net_12309;
wire net_5697;
wire net_1238;
wire net_13697;
wire net_4664;
wire net_14074;
wire net_13547;
wire net_5976;
wire net_7599;
wire net_9483;
wire net_1033;
wire net_10155;
wire net_3923;
wire net_10604;
wire net_8839;
wire net_5560;
wire net_12458;
wire net_11333;
wire net_8333;
wire net_7210;
wire net_13149;
wire net_2554;
wire net_12196;
wire net_4479;
wire net_12005;
wire net_7931;
wire net_12302;
wire net_3107;
wire net_7069;
wire net_14100;
wire net_9716;
wire net_1686;
wire net_11860;
wire net_11481;
wire net_10686;
wire net_10263;
wire net_367;
wire net_3303;
wire net_6354;
wire net_13630;
wire net_9381;
wire net_10928;
wire net_6296;
wire net_10316;
wire net_10061;
wire net_1842;
wire net_7980;
wire net_204;
wire net_9849;
wire net_13037;
wire net_8774;
wire net_3957;
wire net_1180;
wire net_8561;
wire net_1627;
wire net_4596;
wire net_13065;
wire net_12932;
wire net_10235;
wire net_5869;
wire net_2002;
wire net_1069;
wire net_2022;
wire net_9932;
wire net_12014;
wire net_5406;
wire net_2385;
wire net_7626;
wire net_3431;
wire net_7382;
wire net_5829;
wire net_3565;
wire net_7009;
wire net_1416;
wire net_7656;
wire net_13484;
wire net_12045;
wire net_5416;
wire net_6065;
wire net_2433;
wire net_8142;
wire net_6726;
wire net_10784;
wire net_4029;
wire net_1601;
wire net_1916;
wire net_11419;
wire net_2468;
wire net_6614;
wire net_4087;
wire net_4255;
wire net_9854;
wire net_13437;
wire net_8866;
wire net_348;
wire net_7073;
wire net_7398;
wire net_14416;
wire net_9667;
wire net_626;
wire net_10796;
wire net_10953;
wire net_5068;
wire net_11257;
wire net_1809;
wire net_2195;
wire net_686;
wire net_1615;
wire net_11546;
wire net_11246;
wire net_3421;
wire net_1691;
wire net_10089;
wire net_14037;
wire net_7859;
wire net_9197;
wire net_4578;
wire net_2112;
wire net_5072;
wire net_595;
wire net_12312;
wire net_1320;
wire net_1828;
wire net_9461;
wire net_1466;
wire net_5320;
wire net_10438;
wire net_9573;
wire net_7434;
wire net_11268;
wire net_8960;
wire net_157;
wire net_6960;
wire net_1710;
wire net_10994;
wire net_14274;
wire net_11456;
wire net_9017;
wire net_11922;
wire net_6695;
wire net_9006;
wire net_7759;
wire net_11443;
wire net_1205;
wire net_11627;
wire net_10524;
wire net_8154;
wire net_5988;
wire net_6978;
wire net_466;
wire net_6969;
wire net_9612;
wire net_1179;
wire net_4336;
wire net_9601;
wire net_13030;
wire net_4161;
wire net_3039;
wire net_7833;
wire net_13057;
wire net_6207;
wire net_11021;
wire net_2217;
wire net_938;
wire net_1610;
wire net_1761;
wire net_12163;
wire net_3569;
wire net_5682;
wire net_4683;
wire net_183;
wire net_6814;
wire net_13236;
wire net_4246;
wire net_1440;
wire net_7330;
wire net_8893;
wire net_4020;
wire net_6539;
wire net_8389;
wire net_4453;
wire net_11018;
wire net_1011;
wire net_8792;
wire net_7118;
wire net_9902;
wire net_1355;
wire net_7040;
wire net_8420;
wire net_800;
wire net_9221;
wire net_644;
wire net_13495;
wire net_12111;
wire net_8847;
wire net_13586;
wire net_12063;
wire net_12750;
wire net_852;
wire net_5992;
wire net_11917;
wire net_11035;
wire net_11648;
wire net_9405;
wire net_4046;
wire net_2580;
wire net_13834;
wire net_7391;
wire net_13997;
wire net_9696;
wire net_8904;
wire net_13302;
wire net_9961;
wire net_8416;
wire net_8382;
wire net_1385;
wire net_1643;
wire x63;
wire net_1534;
wire net_1919;
wire net_11404;
wire net_9836;
wire net_14284;
wire net_12843;
wire net_10128;
wire net_8992;
wire net_14162;
wire net_8685;
wire net_11492;
wire net_9491;
wire net_8555;
wire net_4876;
wire net_11410;
wire net_9087;
wire net_659;
wire net_8993;
wire net_5871;
wire net_14061;
wire net_899;
wire net_1010;
wire net_1693;
wire net_10224;
wire net_13883;
wire net_10707;
wire net_3654;
wire net_8853;
wire net_10139;
wire net_3779;
wire net_4252;
wire net_2908;
wire net_2068;
wire net_4981;
wire net_3705;
wire net_5907;
wire net_11821;
wire net_5930;
wire net_6371;
wire net_13780;
wire net_13594;
wire net_13813;
wire net_4449;
wire net_11929;
wire net_8939;
wire x638;
wire net_6458;
wire net_7339;
wire net_2675;
wire net_13528;
wire net_2794;
wire net_13567;
wire net_6986;
wire net_314;
wire net_1752;
wire net_5395;
wire net_2527;
wire net_11906;
wire net_11381;
wire net_9765;
wire x1351;
wire net_2091;
wire net_2406;
wire net_6289;
wire net_8722;
wire net_12033;
wire net_8442;
wire net_4669;
wire net_807;
wire net_3405;
wire net_13791;
wire net_12422;
wire net_3270;
wire net_12665;
wire net_5460;
wire net_12479;
wire net_4286;
wire net_6880;
wire net_10238;
wire net_9872;
wire net_3484;
wire net_2474;
wire net_13931;
wire net_945;
wire net_6532;
wire net_2530;
wire net_4380;
wire net_6971;
wire net_12266;
wire net_11578;
wire net_2101;
wire net_7738;
wire net_9472;
wire net_6192;
wire net_6863;
wire net_11451;
wire net_8875;
wire net_8376;
wire net_217;
wire net_7679;
wire net_6582;
wire net_5800;
wire net_5601;
wire net_5336;
wire net_12086;
wire net_13426;
wire net_8844;
wire net_915;
wire net_2226;
wire net_5634;
wire net_3849;
wire net_8099;
wire net_12251;
wire net_8909;
wire net_8808;
wire net_6340;
wire net_8028;
wire net_13256;
wire net_10516;
wire net_9099;
wire net_5174;
wire net_11343;
wire net_8943;
wire net_1784;
wire net_1296;
wire net_8369;
wire net_13081;
wire net_4326;
wire net_2863;
wire net_3507;
wire net_1165;
wire net_5167;
wire net_10245;
wire net_677;
wire net_7159;
wire net_10762;
wire net_1472;
wire net_9735;
wire net_2939;
wire net_13294;
wire net_2424;
wire net_1113;
wire net_1968;
wire net_9945;
wire net_10746;
wire net_10407;
wire net_12291;
wire net_11208;
wire net_4488;
wire net_11619;
wire net_5092;
wire net_5295;
wire net_7464;
wire net_8362;
wire net_11040;
wire net_7713;
wire net_2507;
wire net_5120;
wire net_9633;
wire net_5948;
wire net_13908;
wire net_2685;
wire net_5676;
wire net_8357;
wire net_8340;
wire net_14264;
wire net_2898;
wire net_2658;
wire net_6197;
wire net_2174;
wire net_1391;
wire net_9334;
wire net_9926;
wire net_5132;
wire net_10304;
wire net_784;
wire net_1772;
wire net_3529;
wire net_6128;
wire net_5437;
wire net_8481;
wire net_8751;
wire net_2498;
wire net_381;
wire net_6021;
wire net_9144;
wire net_6574;
wire net_6889;
wire net_2326;
wire net_11566;
wire net_10710;
wire net_3540;
wire net_8094;
wire net_3783;
wire net_11234;
wire net_1857;
wire net_7445;
wire net_5375;
wire net_11586;
wire net_11010;
wire net_9489;
wire net_12078;
wire net_12059;
wire net_6109;
wire net_14414;
wire net_9883;
wire net_3238;
wire net_1318;
wire net_10677;
wire net_1557;
wire net_6843;
wire net_3852;
wire net_1514;
wire net_7668;
wire net_13072;
wire net_6825;
wire net_13874;
wire net_7155;
wire net_3092;
wire net_14407;
wire net_3575;
wire net_4349;
wire net_9209;
wire net_11195;
wire net_8802;
wire net_6995;
wire net_8023;
wire net_6440;
wire net_306;
wire net_4984;
wire net_4516;
wire net_13240;
wire net_9026;
wire net_5371;
wire net_12241;
wire net_500;
wire net_5061;
wire net_5357;
wire net_1906;
wire net_6471;
wire net_9094;
wire net_2610;
wire net_5660;
wire net_8056;
wire net_4432;
wire net_14391;
wire net_1329;
wire net_4584;
wire net_362;
wire net_11967;
wire net_3127;
wire net_9959;
wire net_1052;
wire net_14197;
wire net_10911;
wire net_3831;
wire net_14120;
wire net_13974;
wire net_11180;
wire net_10130;
wire net_11974;
wire net_9477;
wire net_4401;
wire net_3632;
wire net_2189;
wire net_2057;
wire net_4859;
wire net_226;
wire net_1124;
wire net_6413;
wire net_13945;
wire net_7645;
wire net_13737;
wire net_5960;
wire net_5615;
wire net_143;
wire net_12434;
wire net_9160;
wire net_190;
wire net_4964;
wire net_7015;
wire net_2887;
wire net_1447;
wire net_4207;
wire net_1929;
wire net_7741;
wire net_1983;
wire net_10129;
wire net_8735;
wire net_10248;
wire net_9423;
wire net_3493;
wire net_3030;
wire net_2061;
wire net_13466;
wire net_5288;
wire net_13956;
wire net_10251;
wire net_14030;
wire net_13910;
wire net_13727;
wire net_3842;
wire net_13710;
wire net_4266;
wire net_1553;
wire net_1895;
wire net_5360;
wire net_509;
wire net_4975;
wire net_13421;
wire net_10563;
wire net_9983;
wire net_8819;
wire net_2491;
wire net_211;
wire net_3208;
wire net_2704;
wire net_13430;
wire net_10079;
wire net_6752;
wire net_10933;
wire net_5771;
wire net_5819;
wire net_13541;
wire net_3910;
wire net_1851;
wire net_3941;
wire net_6630;
wire net_13684;
wire net_12604;
wire net_8645;
wire net_10976;
wire net_3445;
wire net_2233;
wire net_8709;
wire net_2941;
wire net_2033;
wire net_12726;
wire net_12091;
wire net_8487;
wire net_3348;
wire net_477;
wire net_2123;
wire net_10811;
wire net_12784;
wire net_2943;
wire net_12360;
wire net_9377;
wire net_9049;
wire net_3861;
wire net_5970;
wire net_10892;
wire net_2532;
wire net_6758;
wire net_6905;
wire net_2315;
wire net_8325;
wire net_12785;
wire net_13851;
wire net_2231;
wire net_11112;
wire net_1864;
wire net_11725;
wire net_3812;
wire net_1200;
wire net_6156;
wire net_12840;
wire net_9595;
wire net_2518;
wire net_9509;
wire net_6950;
wire net_10663;
wire net_12329;
wire net_4062;
wire net_7558;
wire net_12284;
wire net_14353;
wire net_7953;
wire net_1646;
wire net_4115;
wire net_11437;
wire net_11135;
wire net_2776;
wire net_13980;
wire net_11487;
wire net_3389;
wire net_3437;
wire net_12938;
wire net_1562;
wire net_2522;
wire net_472;
wire net_14286;
wire net_1510;
wire net_4178;
wire net_14022;
wire net_3077;
wire net_7267;
wire net_8671;
wire net_8639;
wire net_13608;
wire net_4829;
wire net_13878;
wire net_136;
wire net_12987;
wire net_9430;
wire net_1524;
wire net_4171;
wire net_1528;
wire net_10022;
wire net_13579;
wire net_12676;
wire net_9396;
wire net_1749;
wire net_3367;
wire net_4915;
wire net_8386;
wire net_4784;
wire net_12355;
wire net_601;
wire net_12531;
wire net_9785;
wire net_1362;
wire net_11670;
wire net_2346;
wire net_4385;
wire net_6461;
wire net_9315;
wire net_2511;
wire net_829;
wire net_13025;
wire net_2626;
wire net_12396;
wire net_11856;
wire net_2294;
wire net_2115;
wire net_4110;
wire net_4317;
wire net_13867;
wire net_2299;
wire net_14174;
wire net_4978;
wire net_9307;
wire net_10612;
wire net_2393;
wire net_7123;
wire net_3917;
wire net_8812;
wire net_8539;
wire net_13671;
wire net_3376;
wire net_7979;
wire net_1405;
wire net_13845;
wire net_7726;
wire net_10072;
wire net_13518;
wire net_7218;
wire net_10881;
wire net_6555;
wire net_5319;
wire net_716;
wire net_5147;
wire net_13273;
wire net_13200;
wire net_10489;
wire net_11445;
wire net_11045;
wire x1417;
wire net_1269;
wire net_6357;
wire net_13757;
wire net_8630;
wire net_3750;
wire net_12637;
wire net_5314;
wire net_3715;
wire net_3533;
wire net_5400;
wire net_5749;
wire net_12736;
wire net_11805;
wire net_10464;
wire net_9687;
wire net_2696;
wire net_14168;
wire net_6026;
wire net_8457;
wire net_10457;
wire net_12406;
wire net_1449;
wire net_4293;
wire net_9176;
wire net_6984;
wire net_5618;
wire net_666;
wire net_5310;
wire net_9725;
wire net_8620;
wire net_13114;
wire net_13776;
wire net_4809;
wire net_11308;
wire net_12989;
wire net_12706;
wire net_12184;
wire net_1220;
wire net_6212;
wire net_12343;
wire net_11394;
wire net_9702;
wire net_4017;
wire net_4693;
wire net_3946;
wire net_10596;
wire net_10194;
wire net_6346;
wire net_5522;
wire net_6319;
wire net_7636;
wire net_12716;
wire net_9024;
wire net_9824;
wire net_1657;
wire net_6063;
wire net_11781;
wire net_3084;
wire x106;
wire net_4945;
wire net_10689;
wire net_10863;
wire net_14208;
wire net_9859;
wire net_2334;
wire net_1367;
wire net_3994;
wire net_11764;
wire net_7943;
wire net_14213;
wire net_13645;
wire net_1976;
wire net_7960;
wire net_8510;
wire net_3169;
wire net_5647;
wire net_4079;
wire net_3792;
wire net_12104;
wire net_1371;
wire net_13511;
wire net_12542;
wire net_2758;
wire net_9972;
wire net_117;
wire net_1826;
wire net_5002;
wire net_8054;
wire net_6609;
wire net_7837;
wire net_4609;
wire net_10337;
wire net_6517;
wire net_2142;
wire net_4704;
wire net_5782;
wire net_11841;
wire net_9843;
wire net_7864;
wire net_11885;
wire net_7332;
wire net_920;
wire net_10359;
wire net_11826;
wire net_1461;
wire net_3009;
wire net_12980;
wire net_12799;
wire net_5596;
wire net_7512;
wire net_4226;
wire net_3177;
wire net_820;
wire net_7137;
wire net_11249;
wire net_11325;
wire net_8270;
wire net_12556;
wire net_10011;
wire net_9459;
wire net_7222;
wire net_13447;
wire net_8891;
wire net_10360;
wire net_6137;
wire net_13465;
wire net_10475;
wire net_10568;
wire net_437;
wire net_3573;
wire net_13208;
wire net_5959;
wire net_9681;
wire net_566;
wire net_10390;
wire net_9861;
wire net_11477;
wire net_5063;
wire net_7519;
wire net_9071;
wire net_7371;
wire net_12498;
wire net_10855;
wire net_7140;
wire net_9768;
wire net_624;
wire net_2148;
wire net_13173;
wire net_13811;
wire net_11616;
wire net_4735;
wire net_8517;
wire net_2108;
wire net_14063;
wire net_2529;
wire net_688;
wire net_6005;
wire net_6044;
wire net_4685;
wire net_4732;
wire net_9751;
wire net_8732;
wire net_5808;
wire net_8390;
wire net_5979;
wire net_7551;
wire net_11810;
wire net_8170;
wire net_3027;
wire net_12777;
wire net_5343;
wire net_14279;
wire net_6625;
wire net_4235;
wire net_14117;
wire net_11871;
wire net_9940;
wire net_13379;
wire net_4096;
wire net_5497;
wire net_7924;
wire net_9452;
wire net_4117;
wire net_1357;
wire net_5214;
wire net_13990;
wire net_3986;
wire net_4822;
wire net_3637;
wire net_11754;
wire net_5554;
wire net_1243;
wire net_7482;
wire net_12035;
wire net_1660;
wire net_6839;
wire net_1484;
wire net_5864;
wire net_8668;
wire net_4604;
wire net_7489;
wire net_6558;
wire net_12598;
wire net_3667;
wire net_419;
wire net_9949;
wire net_6566;
wire net_6041;
wire net_1635;
wire net_12463;
wire net_5027;
wire net_6779;
wire net_4840;
wire net_5658;
wire net_936;
wire net_12697;
wire net_9259;
wire net_7808;
wire net_8066;
wire net_819;
wire net_7133;
wire net_10969;
wire net_11954;
wire net_8241;
wire net_14121;
wire net_9106;
wire net_8828;
wire net_7523;
wire net_13653;
wire net_10306;
wire net_6871;
wire net_7174;
wire net_7020;
wire net_4070;
wire net_9327;
wire net_3002;
wire net_854;
wire net_11173;
wire net_8713;
wire net_2619;
wire net_6272;
wire net_3141;
wire net_5559;
wire net_1670;
wire net_2221;
wire net_11424;
wire net_4274;
wire net_3265;
wire net_2801;
wire net_10369;
wire net_5264;
wire net_6959;
wire net_2932;
wire net_4951;
wire net_6447;
wire net_7789;
wire net_13342;
wire net_12420;
wire net_7928;
wire net_8277;
wire net_9181;
wire net_5812;
wire net_1264;
wire net_5746;
wire net_8077;
wire net_4643;
wire net_13601;
wire net_9852;
wire net_332;
wire net_1745;
wire net_1679;
wire net_7364;
wire net_9058;
wire net_4883;
wire net_9300;
wire net_3148;
wire net_1229;
wire net_6316;
wire net_13739;
wire net_12746;
wire net_656;
wire net_5723;
wire net_14385;
wire net_4800;
wire net_6277;
wire net_8489;
wire net_766;
wire net_1153;
wire net_8935;
wire net_3014;
wire net_8469;
wire net_10961;
wire net_9102;
wire net_4284;
wire net_9252;
wire net_6734;
wire net_5692;
wire net_14241;
wire net_7027;
wire net_3113;
wire net_14157;
wire net_10924;
wire net_3454;
wire net_8826;
wire net_6816;
wire net_8614;
wire net_5113;
wire net_3969;
wire net_9533;
wire net_13682;
wire net_12333;
wire net_13266;
wire net_7232;
wire net_3729;
wire net_6602;
wire net_9873;
wire net_11164;
wire net_12615;
wire net_7688;
wire net_10465;
wire net_6162;
wire net_14347;
wire net_9589;
wire net_2251;
wire net_12914;
wire net_8898;
wire net_1698;
wire net_9623;
wire net_5897;
wire net_7439;
wire net_10418;
wire net_9727;
wire net_12391;
wire net_955;
wire net_1017;
wire net_2585;
wire net_14379;
wire net_14309;
wire net_1996;
wire net_7046;
wire net_13635;
wire net_1029;
wire net_14293;
wire net_13664;
wire net_13334;
wire net_9812;
wire net_9066;
wire net_412;
wire net_12566;
wire net_8887;
wire net_4798;
wire net_12762;
wire net_9869;
wire net_2986;
wire net_3162;
wire net_4034;
wire net_4791;
wire net_1873;
wire net_3801;
wire x1580;
wire net_13082;
wire net_453;
wire net_7547;
wire net_11937;
wire net_10209;
wire net_3510;
wire net_11848;
wire net_10492;
wire net_5835;
wire net_3180;
wire net_3249;
wire net_14002;
wire net_10439;
wire net_2263;
wire net_6157;
wire net_6181;
wire net_3624;
wire net_734;
wire net_14152;
wire net_12564;
wire net_2544;
wire net_7967;
wire net_9391;
wire net_11596;
wire net_2086;
wire net_951;
wire net_4930;
wire net_3186;
wire net_11314;
wire net_12869;
wire net_12278;
wire net_7272;
wire net_7096;
wire net_12654;
wire net_8977;
wire net_8177;
wire x1382;
wire net_13895;
wire net_14389;
wire net_10222;
wire net_10648;
wire net_12350;
wire net_12121;
wire net_5277;
wire net_7269;
wire net_2966;
wire net_4372;
wire net_13186;
wire net_1253;
wire net_2500;
wire net_10508;
wire net_9808;
wire net_13971;
wire net_1076;
wire net_3900;
wire net_14051;
wire net_10168;
wire net_8234;
wire net_13315;
wire net_10399;
wire net_9711;
wire net_4352;
wire net_3153;
wire net_681;
wire net_6721;
wire net_5155;
wire net_5471;
wire net_7346;
wire net_13136;
wire net_6533;
wire net_3598;
wire net_5252;
wire net_146;
wire net_9562;
wire net_8676;
wire net_3938;
wire net_7534;
wire net_11289;
wire net_5752;
wire net_4594;
wire net_9592;
wire net_1502;
wire net_4454;
wire net_6290;
wire net_4624;
wire net_11522;
wire net_11282;
wire net_6596;
wire net_7621;
wire net_428;
wire net_9675;
wire net_11065;
wire net_10557;
wire net_11306;
wire net_10329;
wire net_12138;
wire net_10117;
wire net_640;
wire net_7780;
wire net_4666;
wire net_2888;
wire net_7508;
wire net_12884;
wire net_775;
wire net_10903;
wire net_752;
wire net_14362;
wire net_3716;
wire net_888;
wire net_535;
wire net_498;
wire net_13066;
wire net_10772;
wire net_13212;
wire net_11298;
wire net_11095;
wire net_9526;
wire net_5191;
wire net_2721;
wire net_8480;
wire net_8900;
wire net_10513;
wire net_2637;
wire net_1023;
wire net_4814;
wire net_5233;
wire net_7499;
wire net_3623;
wire net_301;
wire net_4902;
wire net_6768;
wire net_2360;
wire net_5419;
wire net_3617;
wire net_12228;
wire net_299;
wire net_7432;
wire net_1343;
wire net_7147;
wire net_2285;
wire net_12894;
wire net_12690;
wire net_7355;
wire net_7413;
wire net_12387;
wire net_590;
wire net_3879;
wire net_11755;
wire net_2024;
wire net_3240;
wire net_8229;
wire net_11549;
wire net_3254;
wire net_9569;
wire net_9779;
wire net_9342;
wire net_9040;
wire net_3725;
wire net_12135;
wire net_10094;
wire net_4194;
wire net_12361;
wire net_5464;
wire net_9111;
wire net_8335;
wire net_6088;
wire net_8530;
wire net_5041;
wire net_5857;
wire net_407;
wire net_10145;
wire net_1736;
wire net_12807;
wire net_4405;
wire net_12258;
wire net_11793;
wire net_9814;
wire net_11660;
wire net_6947;
wire net_8723;
wire net_9801;
wire net_10314;
wire net_2312;
wire net_10574;
wire net_4148;
wire net_9155;
wire net_5048;
wire net_8586;
wire net_1669;
wire net_7869;
wire net_11505;
wire net_12408;
wire net_14096;
wire net_2073;
wire net_1041;
wire net_8189;
wire net_7628;
wire net_9146;
wire net_6385;
wire net_14027;
wire net_2950;
wire net_6056;
wire net_4057;
wire net_6108;
wire net_5851;
wire net_14350;
wire net_5105;
wire net_4778;
wire net_14244;
wire net_11211;
wire net_6081;
wire net_13159;
wire net_2364;
wire net_5507;
wire net_12173;
wire net_12526;
wire net_942;
wire net_12822;
wire net_8763;
wire net_7565;
wire net_1981;
wire x906;
wire net_4302;
wire net_1218;
wire net_6245;
wire net_10606;
wire net_13658;
wire net_10917;
wire net_6436;
wire net_1494;
wire net_3286;
wire net_4415;
wire x589;
wire net_2154;
wire net_1726;
wire net_5527;
wire net_4123;
wire net_7082;
wire net_11430;
wire net_5705;
wire net_12165;
wire net_3298;
wire net_3099;
wire net_1398;
wire net_12432;
wire net_10658;
wire net_13219;
wire net_10503;
wire net_6339;
wire net_4399;
wire net_7380;
wire net_8197;
wire net_1144;
wire net_6117;
wire net_1794;
wire net_9363;
wire net_8297;
wire net_12508;
wire net_6503;
wire net_10646;
wire net_5536;
wire net_1022;
wire net_4638;
wire net_11129;
wire net_2865;
wire net_2260;
wire net_6110;
wire net_8182;
wire net_9770;
wire net_3606;
wire net_702;
wire net_4328;
wire net_3195;
wire net_1477;
wire net_3210;
wire net_13960;
wire net_13221;
wire net_3318;
wire net_9270;
wire net_7800;
wire net_8188;
wire net_8122;
wire net_7571;
wire net_11682;
wire net_13152;
wire net_12948;
wire net_12904;
wire net_12439;
wire net_12979;
wire net_1193;
wire net_9412;
wire net_1425;
wire net_1122;
wire net_4911;
wire net_8436;
wire net_10790;
wire net_6228;
wire net_5505;
wire net_10622;
wire net_1813;
wire net_8540;
wire net_4534;
wire net_6252;
wire net_10673;
wire net_7945;
wire net_12411;
wire net_6491;
wire net_983;
wire net_355;
wire net_13898;
wire net_13702;
wire net_4713;
wire net_7258;
wire net_9709;
wire net_9513;
wire net_8102;
wire net_12427;
wire net_9002;
wire net_723;
wire net_4307;
wire net_7311;
wire net_11341;
wire net_8292;
wire net_7614;
wire net_2483;
wire net_5513;
wire net_8248;
wire net_3962;
wire net_12026;
wire net_11834;
wire net_4553;
wire net_275;
wire net_10501;
wire net_10202;
wire net_12641;
wire net_9486;
wire net_4831;
wire net_2914;
wire net_10547;
wire net_11366;
wire net_2590;
wire net_10841;
wire net_7280;
wire net_13293;
wire net_13351;
wire net_1137;
wire net_7424;
wire net_3948;
wire net_4830;
wire net_6142;
wire net_13475;
wire net_13455;
wire net_5036;
wire net_12414;
wire net_12872;
wire net_12860;
wire net_13909;
wire net_9493;
wire net_4865;
wire net_11765;
wire net_8254;
wire net_11945;
wire net_9955;
wire net_14370;
wire net_3819;
wire net_11978;
wire net_254;
wire net_11193;
wire net_12581;
wire net_11895;
wire net_1501;
wire net_3003;
wire net_5622;
wire net_12103;
wire net_574;
wire x868;
wire net_3357;
wire net_11375;
wire net_9467;
wire net_14054;
wire net_9694;
wire net_8425;

// Start cells
CLKBUF_X2 inst_12147 ( .A(net_10852), .Z(net_12109) );
OAI21_X2 inst_1783 ( .B1(net_5446), .ZN(net_5408), .A(net_4682), .B2(net_3988) );
CLKBUF_X2 inst_10910 ( .A(net_10871), .Z(net_10872) );
CLKBUF_X2 inst_13999 ( .A(net_11240), .Z(net_13961) );
DFF_X1 inst_6916 ( .D(net_2397), .Q(net_249), .CK(net_8025) );
NAND3_X2 inst_2685 ( .ZN(net_3178), .A3(net_2984), .A2(net_1962), .A1(net_1106) );
CLKBUF_X2 inst_9876 ( .A(net_9837), .Z(net_9838) );
NAND2_X2 inst_4123 ( .A2(net_1222), .ZN(net_1168), .A1(net_339) );
AOI21_X2 inst_7766 ( .B1(net_7132), .ZN(net_4445), .B2(net_2582), .A(net_2358) );
DFF_X1 inst_6919 ( .D(net_2388), .Q(net_254), .CK(net_10416) );
OAI21_X2 inst_1751 ( .ZN(net_5514), .A(net_4815), .B2(net_4153), .B1(net_1190) );
CLKBUF_X2 inst_8140 ( .A(net_7912), .Z(net_8102) );
INV_X4 inst_5359 ( .A(net_7408), .ZN(net_2107) );
NOR2_X4 inst_2235 ( .ZN(net_5663), .A1(net_5520), .A2(net_4491) );
SDFF_X2 inst_779 ( .D(net_7807), .SI(net_6907), .Q(net_6907), .SE(net_3781), .CK(net_11459) );
CLKBUF_X2 inst_13828 ( .A(net_13568), .Z(net_13790) );
CLKBUF_X2 inst_11465 ( .A(net_11426), .Z(net_11427) );
DFF_X1 inst_6439 ( .QN(net_6082), .D(net_5731), .CK(net_11680) );
INV_X4 inst_5306 ( .A(net_6004), .ZN(net_2600) );
NOR3_X2 inst_2205 ( .A3(net_5924), .ZN(net_3065), .A2(net_2807), .A1(net_2806) );
NAND2_X4 inst_2858 ( .A1(net_5878), .ZN(net_5074), .A2(net_4144) );
CLKBUF_X2 inst_10503 ( .A(net_10464), .Z(net_10465) );
CLKBUF_X2 inst_8981 ( .A(net_8618), .Z(net_8943) );
INV_X4 inst_5488 ( .A(net_6065), .ZN(net_3536) );
NAND2_X2 inst_4131 ( .A2(net_1225), .ZN(net_1063), .A1(net_362) );
CLKBUF_X2 inst_13591 ( .A(net_13552), .Z(net_13553) );
CLKBUF_X2 inst_9805 ( .A(net_9766), .Z(net_9767) );
CLKBUF_X2 inst_13926 ( .A(net_13094), .Z(net_13888) );
SDFF_X2 inst_214 ( .SI(net_6339), .Q(net_6300), .D(net_3703), .SE(net_392), .CK(net_13542) );
CLKBUF_X2 inst_13990 ( .A(net_13951), .Z(net_13952) );
CLKBUF_X2 inst_9115 ( .A(net_8416), .Z(net_9077) );
NAND2_X1 inst_4228 ( .ZN(net_4699), .A2(net_3989), .A1(net_2084) );
SDFF_X2 inst_548 ( .Q(net_6453), .D(net_6453), .SI(net_3821), .SE(net_3820), .CK(net_8427) );
CLKBUF_X2 inst_10808 ( .A(net_10769), .Z(net_10770) );
CLKBUF_X2 inst_12017 ( .A(net_11978), .Z(net_11979) );
INV_X4 inst_4647 ( .ZN(net_4175), .A(net_4010) );
NAND2_X1 inst_4372 ( .ZN(net_4355), .A2(net_3856), .A1(net_1799) );
AOI22_X2 inst_7408 ( .A2(net_3105), .B1(net_2970), .ZN(net_2827), .A1(net_730), .B2(net_258) );
CLKBUF_X2 inst_12796 ( .A(net_12757), .Z(net_12758) );
INV_X4 inst_4709 ( .ZN(net_2987), .A(net_2986) );
CLKBUF_X2 inst_10461 ( .A(net_10422), .Z(net_10423) );
CLKBUF_X2 inst_8488 ( .A(net_8449), .Z(net_8450) );
CLKBUF_X2 inst_14178 ( .A(net_14139), .Z(net_14140) );
CLKBUF_X2 inst_10820 ( .A(net_10781), .Z(net_10782) );
DFFR_X2 inst_7060 ( .QN(net_6032), .D(net_3059), .CK(net_10014), .RN(x1822) );
CLKBUF_X2 inst_14148 ( .A(net_14109), .Z(net_14110) );
CLKBUF_X2 inst_13127 ( .A(net_13088), .Z(net_13089) );
NAND2_X2 inst_3347 ( .ZN(net_3553), .A1(net_3552), .A2(net_3225) );
NAND2_X2 inst_3130 ( .ZN(net_4833), .A2(net_4153), .A1(net_2186) );
CLKBUF_X2 inst_11446 ( .A(net_11407), .Z(net_11408) );
CLKBUF_X2 inst_9568 ( .A(net_7943), .Z(net_9530) );
DFF_X1 inst_6406 ( .QN(net_6133), .D(net_5764), .CK(net_10964) );
INV_X4 inst_5341 ( .A(net_6155), .ZN(net_3611) );
NAND2_X2 inst_4136 ( .A2(net_1222), .ZN(net_1141), .A1(net_334) );
CLKBUF_X2 inst_12400 ( .A(net_12361), .Z(net_12362) );
CLKBUF_X2 inst_12585 ( .A(net_12546), .Z(net_12547) );
CLKBUF_X2 inst_9372 ( .A(net_9333), .Z(net_9334) );
SDFF_X2 inst_1228 ( .SI(net_7222), .Q(net_7222), .D(net_3794), .SE(net_3751), .CK(net_10611) );
CLKBUF_X2 inst_8913 ( .A(net_8874), .Z(net_8875) );
CLKBUF_X2 inst_13185 ( .A(net_7859), .Z(net_13147) );
CLKBUF_X2 inst_9653 ( .A(net_9614), .Z(net_9615) );
INV_X4 inst_4985 ( .A(net_3167), .ZN(net_744) );
NAND2_X1 inst_4221 ( .ZN(net_4739), .A2(net_3988), .A1(net_2109) );
SDFF_X2 inst_521 ( .Q(net_6704), .D(net_6704), .SI(net_3894), .SE(net_3871), .CK(net_11124) );
INV_X4 inst_5164 ( .ZN(net_641), .A(net_546) );
CLKBUF_X2 inst_9461 ( .A(net_9422), .Z(net_9423) );
DFF_X1 inst_6534 ( .QN(net_7481), .D(net_5417), .CK(net_12109) );
CLKBUF_X2 inst_9736 ( .A(net_9697), .Z(net_9698) );
INV_X2 inst_5947 ( .A(net_7688), .ZN(net_408) );
INV_X8 inst_4473 ( .ZN(net_5139), .A(net_4273) );
OAI21_X2 inst_1685 ( .ZN(net_5780), .B1(net_5778), .A(net_5715), .B2(net_5714) );
NOR2_X2 inst_2511 ( .A2(net_3232), .ZN(net_1171), .A1(net_1170) );
OAI221_X2 inst_1655 ( .ZN(net_4799), .A(net_4594), .C2(net_3977), .B2(net_3966), .C1(net_3770), .B1(net_1970) );
CLKBUF_X2 inst_12320 ( .A(net_11937), .Z(net_12282) );
CLKBUF_X2 inst_10720 ( .A(net_10505), .Z(net_10682) );
CLKBUF_X2 inst_9038 ( .A(net_8999), .Z(net_9000) );
DFF_X1 inst_6910 ( .D(net_2514), .QN(net_175), .CK(net_9853) );
NAND2_X2 inst_3578 ( .ZN(net_2436), .A2(net_2435), .A1(net_744) );
CLKBUF_X2 inst_9257 ( .A(net_9218), .Z(net_9219) );
CLKBUF_X2 inst_9938 ( .A(net_9899), .Z(net_9900) );
CLKBUF_X2 inst_14165 ( .A(net_14126), .Z(net_14127) );
AOI22_X2 inst_7415 ( .B1(net_5939), .ZN(net_2779), .A1(net_2777), .B2(net_218), .A2(net_181) );
CLKBUF_X2 inst_8731 ( .A(net_8692), .Z(net_8693) );
CLKBUF_X2 inst_12238 ( .A(net_12199), .Z(net_12200) );
INV_X4 inst_4847 ( .ZN(net_5100), .A(net_1063) );
INV_X2 inst_6010 ( .A(net_6164), .ZN(net_2700) );
INV_X2 inst_5940 ( .A(net_7314), .ZN(net_1785) );
CLKBUF_X2 inst_14010 ( .A(net_13971), .Z(net_13972) );
CLKBUF_X2 inst_13236 ( .A(net_11274), .Z(net_13198) );
SDFF_X2 inst_1066 ( .D(net_7802), .SI(net_7204), .Q(net_7204), .SE(net_3750), .CK(net_13319) );
CLKBUF_X2 inst_10825 ( .A(net_10786), .Z(net_10787) );
CLKBUF_X2 inst_9978 ( .A(net_9939), .Z(net_9940) );
CLKBUF_X2 inst_7977 ( .A(net_7938), .Z(net_7939) );
NAND2_X2 inst_3392 ( .ZN(net_3763), .A2(net_3365), .A1(net_2889) );
CLKBUF_X2 inst_12122 ( .A(net_12083), .Z(net_12084) );
CLKBUF_X2 inst_10377 ( .A(net_9000), .Z(net_10339) );
INV_X4 inst_5063 ( .ZN(net_728), .A(net_634) );
DFF_X2 inst_6232 ( .QN(net_6062), .D(net_3457), .CK(net_12382) );
NOR2_X2 inst_2342 ( .A2(net_6047), .A1(net_5778), .ZN(net_5683) );
INV_X4 inst_4608 ( .ZN(net_4236), .A(net_4090) );
NOR2_X4 inst_2294 ( .ZN(net_2712), .A1(net_2711), .A2(net_736) );
CLKBUF_X2 inst_9143 ( .A(net_9104), .Z(net_9105) );
CLKBUF_X2 inst_14321 ( .A(net_14282), .Z(net_14283) );
CLKBUF_X2 inst_12495 ( .A(net_12456), .Z(net_12457) );
OAI22_X2 inst_1617 ( .B1(net_5942), .ZN(net_2789), .A1(net_2784), .B2(net_211), .A2(net_174) );
CLKBUF_X2 inst_12553 ( .A(net_12514), .Z(net_12515) );
SDFF_X2 inst_151 ( .Q(net_6227), .SI(net_6226), .SE(net_392), .D(net_133), .CK(net_14095) );
NOR2_X4 inst_2256 ( .ZN(net_5630), .A1(net_5475), .A2(net_4433) );
INV_X4 inst_4821 ( .ZN(net_3055), .A(net_1092) );
CLKBUF_X2 inst_8696 ( .A(net_8657), .Z(net_8658) );
AOI222_X2 inst_7519 ( .B1(net_7377), .C1(net_7313), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2012), .A1(net_2011) );
NAND2_X2 inst_3931 ( .A1(net_6710), .A2(net_1497), .ZN(net_1367) );
INV_X4 inst_4880 ( .A(net_3048), .ZN(net_2965) );
CLKBUF_X2 inst_12409 ( .A(net_12370), .Z(net_12371) );
CLKBUF_X2 inst_11637 ( .A(net_11598), .Z(net_11599) );
CLKBUF_X2 inst_12682 ( .A(net_11834), .Z(net_12644) );
CLKBUF_X2 inst_10370 ( .A(net_9100), .Z(net_10332) );
NAND2_X2 inst_3867 ( .A1(net_6565), .A2(net_1705), .ZN(net_1462) );
OAI21_X2 inst_2072 ( .B1(net_5910), .B2(net_4436), .ZN(net_4421), .A(net_3624) );
OAI22_X2 inst_1603 ( .B2(net_3200), .A2(net_3187), .ZN(net_3132), .A1(net_3131), .B1(net_731) );
CLKBUF_X2 inst_13237 ( .A(net_13198), .Z(net_13199) );
CLKBUF_X2 inst_9634 ( .A(net_9595), .Z(net_9596) );
SDFF_X2 inst_340 ( .Q(net_6364), .SI(net_6363), .D(net_3560), .SE(net_392), .CK(net_13605) );
CLKBUF_X2 inst_11590 ( .A(net_11551), .Z(net_11552) );
CLKBUF_X2 inst_10785 ( .A(net_9093), .Z(net_10747) );
CLKBUF_X2 inst_13098 ( .A(net_13059), .Z(net_13060) );
CLKBUF_X2 inst_8109 ( .A(net_7872), .Z(net_8071) );
CLKBUF_X2 inst_8864 ( .A(net_8825), .Z(net_8826) );
CLKBUF_X2 inst_11075 ( .A(net_11009), .Z(net_11037) );
NAND2_X1 inst_4280 ( .ZN(net_4587), .A2(net_3867), .A1(net_1852) );
SDFF_X2 inst_158 ( .Q(net_6256), .SI(net_6255), .D(net_3546), .SE(net_392), .CK(net_13990) );
CLKBUF_X2 inst_8171 ( .A(net_8132), .Z(net_8133) );
AOI222_X2 inst_7493 ( .C1(net_7527), .B1(net_7495), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2094), .A1(net_2093) );
INV_X4 inst_5411 ( .A(net_7680), .ZN(net_797) );
CLKBUF_X2 inst_14279 ( .A(net_14240), .Z(net_14241) );
CLKBUF_X2 inst_13529 ( .A(net_11044), .Z(net_13491) );
NAND2_X1 inst_4244 ( .ZN(net_4683), .A2(net_3988), .A1(net_2172) );
OAI22_X2 inst_1490 ( .B1(net_4666), .A1(net_4132), .B2(net_4124), .ZN(net_4121), .A2(net_4120) );
SDFF_X2 inst_507 ( .Q(net_6474), .D(net_6474), .SE(net_3904), .SI(net_3897), .CK(net_8793) );
INV_X8 inst_4559 ( .ZN(net_1651), .A(net_476) );
NAND2_X1 inst_4289 ( .ZN(net_4578), .A2(net_3867), .A1(net_1191) );
NAND2_X2 inst_3709 ( .A1(net_6897), .ZN(net_1640), .A2(net_1639) );
CLKBUF_X2 inst_14365 ( .A(net_11181), .Z(net_14327) );
CLKBUF_X2 inst_10566 ( .A(net_10527), .Z(net_10528) );
CLKBUF_X2 inst_10934 ( .A(net_10895), .Z(net_10896) );
DFF_X2 inst_6319 ( .QN(net_7800), .CK(net_8160), .D(x1542) );
CLKBUF_X2 inst_12311 ( .A(net_12272), .Z(net_12273) );
SDFF_X2 inst_884 ( .Q(net_7114), .D(net_7114), .SE(net_3888), .SI(net_3787), .CK(net_7870) );
SDFF_X2 inst_711 ( .SI(net_6784), .Q(net_6784), .SE(net_3816), .D(net_3790), .CK(net_8359) );
SDFF_X2 inst_827 ( .Q(net_6996), .D(net_6996), .SE(net_3899), .SI(net_3797), .CK(net_9097) );
DFF_X1 inst_6542 ( .QN(net_7474), .D(net_5574), .CK(net_9260) );
CLKBUF_X2 inst_11477 ( .A(net_11438), .Z(net_11439) );
CLKBUF_X2 inst_14452 ( .A(net_14413), .Z(net_14414) );
CLKBUF_X2 inst_9573 ( .A(net_8074), .Z(net_9535) );
CLKBUF_X2 inst_10730 ( .A(net_10691), .Z(net_10692) );
CLKBUF_X2 inst_10574 ( .A(net_10535), .Z(net_10536) );
CLKBUF_X2 inst_11213 ( .A(net_11174), .Z(net_11175) );
CLKBUF_X2 inst_8465 ( .A(net_8426), .Z(net_8427) );
NAND2_X2 inst_3040 ( .A1(net_6992), .A2(net_4977), .ZN(net_4967) );
CLKBUF_X2 inst_12937 ( .A(net_12898), .Z(net_12899) );
NAND2_X2 inst_4191 ( .A2(net_6021), .ZN(net_1739), .A1(net_472) );
NAND2_X2 inst_3870 ( .A1(net_6572), .A2(net_1705), .ZN(net_1458) );
CLKBUF_X2 inst_14171 ( .A(net_11005), .Z(net_14133) );
INV_X4 inst_5675 ( .A(net_7529), .ZN(net_705) );
NAND2_X1 inst_4269 ( .ZN(net_4648), .A2(net_3993), .A1(net_1507) );
CLKBUF_X2 inst_8559 ( .A(net_8520), .Z(net_8521) );
INV_X4 inst_4640 ( .ZN(net_4182), .A(net_4023) );
XNOR2_X2 inst_18 ( .ZN(net_2633), .B(net_2632), .A(net_2475) );
INV_X2 inst_6047 ( .ZN(net_398), .A(x837) );
NAND2_X2 inst_4128 ( .ZN(net_1235), .A2(net_1225), .A1(net_365) );
CLKBUF_X2 inst_9040 ( .A(net_9001), .Z(net_9002) );
CLKBUF_X2 inst_10154 ( .A(net_10115), .Z(net_10116) );
NOR2_X4 inst_2263 ( .ZN(net_5623), .A1(net_5468), .A2(net_4420) );
INV_X4 inst_5608 ( .A(net_7736), .ZN(net_2673) );
INV_X4 inst_4861 ( .A(net_7802), .ZN(net_3291) );
INV_X4 inst_4796 ( .A(net_2855), .ZN(net_2805) );
INV_X4 inst_5183 ( .A(net_530), .ZN(net_520) );
NAND2_X2 inst_3549 ( .ZN(net_2518), .A2(net_2064), .A1(net_1758) );
CLKBUF_X2 inst_12602 ( .A(net_12563), .Z(net_12564) );
NAND2_X2 inst_3501 ( .A1(net_6401), .ZN(net_2718), .A2(net_2564) );
CLKBUF_X2 inst_10035 ( .A(net_9996), .Z(net_9997) );
NAND2_X2 inst_3936 ( .A1(net_7464), .A2(net_1696), .ZN(net_1357) );
CLKBUF_X2 inst_13029 ( .A(net_12877), .Z(net_12991) );
CLKBUF_X2 inst_13738 ( .A(net_13699), .Z(net_13700) );
NAND2_X2 inst_4175 ( .A1(net_6553), .ZN(net_780), .A2(net_666) );
INV_X2 inst_6069 ( .A(net_7285), .ZN(net_2007) );
DFF_X1 inst_6675 ( .QN(net_7252), .D(net_5151), .CK(net_12726) );
CLKBUF_X2 inst_9783 ( .A(net_8009), .Z(net_9745) );
CLKBUF_X2 inst_8535 ( .A(net_8496), .Z(net_8497) );
DFFR_X2 inst_7076 ( .D(net_2811), .QN(net_298), .CK(net_11420), .RN(x1822) );
INV_X2 inst_6020 ( .A(net_6038), .ZN(net_2609) );
CLKBUF_X2 inst_14217 ( .A(net_12732), .Z(net_14179) );
CLKBUF_X2 inst_12739 ( .A(net_12700), .Z(net_12701) );
DFFS_X2 inst_6954 ( .QN(net_6404), .D(net_2653), .CK(net_14397), .SN(x1822) );
CLKBUF_X2 inst_9416 ( .A(net_9377), .Z(net_9378) );
AOI22_X2 inst_7378 ( .B1(net_7741), .A1(net_7712), .A2(net_5916), .B2(net_2957), .ZN(net_2943) );
CLKBUF_X2 inst_9217 ( .A(net_9074), .Z(net_9179) );
DFF_X1 inst_6475 ( .QN(net_6088), .D(net_5584), .CK(net_12956) );
NAND2_X1 inst_4397 ( .A2(net_5891), .ZN(net_3237), .A1(net_3236) );
CLKBUF_X2 inst_10818 ( .A(net_10779), .Z(net_10780) );
AOI22_X2 inst_7392 ( .ZN(net_2926), .A2(net_2925), .B2(net_2924), .A1(net_1200), .B1(net_1199) );
NAND2_X2 inst_3102 ( .A1(net_6581), .ZN(net_4901), .A2(net_4897) );
CLKBUF_X2 inst_12847 ( .A(net_10412), .Z(net_12809) );
AOI22_X2 inst_7364 ( .A2(net_5916), .ZN(net_2961), .B2(net_2957), .B1(net_2658), .A1(net_853) );
INV_X2 inst_5816 ( .A(net_1639), .ZN(net_1097) );
NAND3_X2 inst_2695 ( .ZN(net_2980), .A3(net_2895), .A2(net_2754), .A1(net_1713) );
CLKBUF_X2 inst_13801 ( .A(net_13762), .Z(net_13763) );
CLKBUF_X2 inst_12748 ( .A(net_12709), .Z(net_12710) );
NAND2_X2 inst_3860 ( .A1(net_7102), .A2(net_1675), .ZN(net_1473) );
CLKBUF_X2 inst_12515 ( .A(net_12379), .Z(net_12477) );
OAI21_X2 inst_2063 ( .B2(net_4436), .ZN(net_4432), .B1(net_4056), .A(net_3549) );
CLKBUF_X2 inst_13635 ( .A(net_10114), .Z(net_13597) );
CLKBUF_X2 inst_10692 ( .A(net_10653), .Z(net_10654) );
INV_X4 inst_4801 ( .ZN(net_5099), .A(net_1235) );
CLKBUF_X2 inst_14150 ( .A(net_14111), .Z(net_14112) );
NAND2_X2 inst_3723 ( .A1(net_6896), .A2(net_1639), .ZN(net_1622) );
CLKBUF_X2 inst_13228 ( .A(net_13189), .Z(net_13190) );
NAND2_X2 inst_3521 ( .ZN(net_2546), .A2(net_2116), .A1(net_1412) );
CLKBUF_X2 inst_9346 ( .A(net_9307), .Z(net_9308) );
CLKBUF_X2 inst_8969 ( .A(net_8242), .Z(net_8931) );
NAND2_X2 inst_3440 ( .ZN(net_3207), .A2(net_3169), .A1(net_3109) );
CLKBUF_X2 inst_12286 ( .A(net_12247), .Z(net_12248) );
CLKBUF_X2 inst_14350 ( .A(net_14311), .Z(net_14312) );
INV_X4 inst_5386 ( .A(net_7684), .ZN(net_886) );
NAND2_X2 inst_3985 ( .ZN(net_1285), .A1(net_885), .A2(net_323) );
OAI21_X2 inst_2036 ( .B1(net_4600), .B2(net_4476), .ZN(net_4467), .A(net_3588) );
INV_X2 inst_5802 ( .ZN(net_1836), .A(net_1835) );
NAND2_X2 inst_4001 ( .ZN(net_1155), .A1(net_919), .A2(net_690) );
CLKBUF_X2 inst_12249 ( .A(net_12210), .Z(net_12211) );
CLKBUF_X2 inst_11107 ( .A(net_11068), .Z(net_11069) );
CLKBUF_X2 inst_9853 ( .A(net_8232), .Z(net_9815) );
CLKBUF_X2 inst_7897 ( .A(net_7838), .Z(net_7859) );
OAI21_X2 inst_2049 ( .B2(net_4457), .ZN(net_4451), .B1(net_4074), .A(net_3708) );
SDFF_X2 inst_868 ( .SI(net_7055), .Q(net_7055), .SE(net_3818), .D(net_3789), .CK(net_10984) );
CLKBUF_X2 inst_10747 ( .A(net_8043), .Z(net_10709) );
CLKBUF_X2 inst_8187 ( .A(net_8110), .Z(net_8149) );
CLKBUF_X2 inst_9188 ( .A(net_8249), .Z(net_9150) );
DFF_X1 inst_6625 ( .QN(net_7595), .D(net_5262), .CK(net_10578) );
CLKBUF_X2 inst_11240 ( .A(net_11201), .Z(net_11202) );
DFF_X2 inst_6184 ( .Q(net_6396), .D(net_6395), .CK(net_14186) );
SDFF_X2 inst_201 ( .Q(net_6313), .SI(net_6312), .D(net_3695), .SE(net_392), .CK(net_13577) );
CLKBUF_X2 inst_10958 ( .A(net_10919), .Z(net_10920) );
NAND2_X2 inst_3627 ( .ZN(net_1956), .A1(net_1292), .A2(net_1126) );
SDFF_X2 inst_1084 ( .SI(net_7062), .Q(net_7062), .D(net_3802), .SE(net_3747), .CK(net_9087) );
SDFF_X2 inst_304 ( .SI(net_7525), .Q(net_7525), .D(net_5100), .SE(net_3988), .CK(net_12455) );
CLKBUF_X2 inst_14388 ( .A(net_10118), .Z(net_14350) );
CLKBUF_X2 inst_10106 ( .A(net_10067), .Z(net_10068) );
NAND2_X2 inst_4157 ( .A1(net_7228), .ZN(net_881), .A2(net_611) );
SDFF_X2 inst_1027 ( .SI(net_6514), .Q(net_6514), .SE(net_3889), .D(net_3790), .CK(net_11229) );
CLKBUF_X2 inst_8432 ( .A(net_8393), .Z(net_8394) );
INV_X2 inst_5793 ( .A(net_5969), .ZN(net_2235) );
SDFF_X2 inst_1143 ( .SI(net_6803), .Q(net_6803), .D(net_3811), .SE(net_3729), .CK(net_11136) );
CLKBUF_X2 inst_12823 ( .A(net_11001), .Z(net_12785) );
CLKBUF_X2 inst_11336 ( .A(net_11297), .Z(net_11298) );
CLKBUF_X2 inst_10670 ( .A(net_10631), .Z(net_10632) );
SDFFR_X2 inst_1345 ( .Q(net_7713), .D(net_7713), .SI(net_3804), .SE(net_3405), .CK(net_10708), .RN(x1822) );
NAND2_X2 inst_2947 ( .ZN(net_5499), .A1(net_4958), .A2(net_4957) );
CLKBUF_X2 inst_12024 ( .A(net_9670), .Z(net_11986) );
CLKBUF_X2 inst_10457 ( .A(net_7886), .Z(net_10419) );
INV_X4 inst_5122 ( .A(net_597), .ZN(net_595) );
CLKBUF_X2 inst_14225 ( .A(net_13616), .Z(net_14187) );
CLKBUF_X2 inst_12951 ( .A(net_12912), .Z(net_12913) );
CLKBUF_X2 inst_12679 ( .A(net_12640), .Z(net_12641) );
CLKBUF_X2 inst_11824 ( .A(net_11785), .Z(net_11786) );
INV_X4 inst_5638 ( .A(net_7730), .ZN(net_2685) );
CLKBUF_X2 inst_8503 ( .A(net_8464), .Z(net_8465) );
NAND2_X2 inst_3608 ( .ZN(net_2388), .A2(net_1890), .A1(net_1337) );
CLKBUF_X2 inst_10724 ( .A(net_10685), .Z(net_10686) );
AOI22_X2 inst_7306 ( .B1(net_6679), .A1(net_6647), .A2(net_5139), .B2(net_5138), .ZN(net_5137) );
SDFF_X2 inst_1016 ( .SI(net_6510), .Q(net_6510), .SE(net_3889), .D(net_3775), .CK(net_8401) );
NAND2_X2 inst_4147 ( .ZN(net_1689), .A2(net_894), .A1(net_715) );
OAI22_X2 inst_1538 ( .B1(net_4637), .A1(net_4030), .B2(net_4022), .ZN(net_4019), .A2(net_4018) );
SDFF_X2 inst_848 ( .Q(net_7000), .D(net_7000), .SE(net_3899), .SI(net_3799), .CK(net_11949) );
CLKBUF_X2 inst_13394 ( .A(net_13355), .Z(net_13356) );
CLKBUF_X2 inst_10349 ( .A(net_10310), .Z(net_10311) );
CLKBUF_X2 inst_12525 ( .A(net_12486), .Z(net_12487) );
NOR2_X2 inst_2479 ( .A2(net_5778), .ZN(net_2666), .A1(net_505) );
CLKBUF_X2 inst_14333 ( .A(net_14294), .Z(net_14295) );
DFF_X1 inst_6465 ( .QN(net_6150), .D(net_5594), .CK(net_11980) );
DFF_X2 inst_6312 ( .Q(net_7802), .CK(net_8163), .D(x1527) );
NOR4_X2 inst_2179 ( .A2(net_7756), .ZN(net_3313), .A3(net_3208), .A1(net_2921), .A4(net_617) );
NAND3_X2 inst_2578 ( .ZN(net_5761), .A1(net_5656), .A2(net_5278), .A3(net_4315) );
AOI222_X2 inst_7514 ( .B1(net_7374), .C1(net_7310), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2026), .A1(net_2025) );
OAI21_X2 inst_1996 ( .B2(net_4518), .ZN(net_4517), .B1(net_4134), .A(net_3698) );
OAI22_X2 inst_1554 ( .B2(net_3405), .A2(net_3360), .ZN(net_3351), .A1(net_3201), .B1(net_544) );
OAI22_X2 inst_1542 ( .B1(net_4637), .B2(net_4418), .A2(net_4032), .A1(net_4030), .ZN(net_4011) );
INV_X8 inst_4511 ( .ZN(net_3893), .A(net_3165) );
CLKBUF_X2 inst_8849 ( .A(net_8810), .Z(net_8811) );
AND2_X4 inst_7830 ( .ZN(net_3014), .A2(net_2815), .A1(net_2251) );
CLKBUF_X2 inst_11580 ( .A(net_11541), .Z(net_11542) );
CLKBUF_X2 inst_12838 ( .A(net_12799), .Z(net_12800) );
NAND2_X2 inst_3340 ( .ZN(net_3567), .A1(net_3566), .A2(net_3225) );
SDFF_X2 inst_644 ( .SI(net_6628), .Q(net_6628), .SE(net_3850), .D(net_3798), .CK(net_12900) );
INV_X4 inst_4683 ( .ZN(net_3740), .A(net_3368) );
INV_X4 inst_5015 ( .A(net_7806), .ZN(net_3811) );
OR2_X4 inst_1380 ( .ZN(net_4155), .A2(net_3402), .A1(net_3222) );
NAND3_X2 inst_2806 ( .ZN(net_2292), .A3(net_1540), .A1(net_1331), .A2(net_973) );
NAND2_X2 inst_3891 ( .A1(net_6695), .A2(net_1497), .ZN(net_1425) );
CLKBUF_X2 inst_11298 ( .A(net_11259), .Z(net_11260) );
CLKBUF_X2 inst_12484 ( .A(net_12445), .Z(net_12446) );
DFF_X1 inst_6736 ( .QN(net_7355), .D(net_5319), .CK(net_12975) );
NAND2_X2 inst_4008 ( .ZN(net_1685), .A2(net_886), .A1(net_862) );
CLKBUF_X2 inst_8318 ( .A(net_8165), .Z(net_8280) );
DFF_X1 inst_6449 ( .QN(net_6100), .D(net_5721), .CK(net_9220) );
CLKBUF_X2 inst_10652 ( .A(net_10613), .Z(net_10614) );
INV_X4 inst_4834 ( .A(net_3849), .ZN(net_3052) );
NAND2_X2 inst_3472 ( .ZN(net_2742), .A1(net_2708), .A2(net_266) );
CLKBUF_X2 inst_12229 ( .A(net_12190), .Z(net_12191) );
INV_X4 inst_4896 ( .ZN(net_909), .A(net_872) );
CLKBUF_X2 inst_8736 ( .A(net_8697), .Z(net_8698) );
CLKBUF_X2 inst_9933 ( .A(net_9566), .Z(net_9895) );
SDFF_X2 inst_432 ( .Q(net_7388), .D(net_7388), .SE(net_3994), .SI(net_353), .CK(net_12433) );
SDFF_X2 inst_282 ( .D(net_6397), .SE(net_5800), .SI(net_362), .Q(net_362), .CK(net_13675) );
CLKBUF_X2 inst_8906 ( .A(net_8867), .Z(net_8868) );
CLKBUF_X2 inst_11584 ( .A(net_11545), .Z(net_11546) );
CLKBUF_X2 inst_8428 ( .A(net_8389), .Z(net_8390) );
CLKBUF_X2 inst_12533 ( .A(net_12494), .Z(net_12495) );
CLKBUF_X2 inst_9605 ( .A(net_8852), .Z(net_9567) );
NOR2_X2 inst_2322 ( .A2(net_6296), .A1(net_5843), .ZN(net_5819) );
SDFF_X2 inst_513 ( .SI(net_6783), .Q(net_6783), .D(net_3898), .SE(net_3872), .CK(net_8381) );
NAND2_X2 inst_3266 ( .ZN(net_4137), .A1(net_3849), .A2(net_3461) );
NAND2_X2 inst_3171 ( .ZN(net_4762), .A2(net_3941), .A1(net_2059) );
CLKBUF_X2 inst_14340 ( .A(net_14301), .Z(net_14302) );
CLKBUF_X2 inst_8725 ( .A(net_8410), .Z(net_8687) );
AOI21_X2 inst_7694 ( .B1(net_6737), .ZN(net_4131), .B2(net_2581), .A(net_2369) );
CLKBUF_X2 inst_14060 ( .A(net_10265), .Z(net_14022) );
OAI22_X1 inst_1630 ( .B2(net_4157), .ZN(net_3832), .A2(net_3402), .A1(net_1710), .B1(net_1271) );
CLKBUF_X2 inst_12479 ( .A(net_12440), .Z(net_12441) );
OAI22_X2 inst_1586 ( .B2(net_3200), .ZN(net_3189), .A1(net_3188), .A2(net_3187), .B1(net_545) );
CLKBUF_X2 inst_9318 ( .A(net_9279), .Z(net_9280) );
CLKBUF_X2 inst_7887 ( .A(net_7844), .Z(net_7849) );
CLKBUF_X2 inst_10296 ( .A(net_8913), .Z(net_10258) );
SDFF_X2 inst_774 ( .SI(net_7802), .Q(net_6870), .D(net_6870), .SE(net_3901), .CK(net_11800) );
NOR2_X4 inst_2292 ( .A2(net_7791), .ZN(net_2864), .A1(net_803) );
CLKBUF_X2 inst_13954 ( .A(net_7940), .Z(net_13916) );
INV_X2 inst_6083 ( .A(net_7596), .ZN(net_1428) );
NAND2_X1 inst_4256 ( .ZN(net_4670), .A2(net_3993), .A1(net_1488) );
CLKBUF_X2 inst_10773 ( .A(net_10734), .Z(net_10735) );
INV_X4 inst_5300 ( .A(net_7734), .ZN(net_2949) );
CLKBUF_X2 inst_12340 ( .A(net_12301), .Z(net_12302) );
NAND3_X2 inst_2766 ( .ZN(net_2334), .A3(net_1579), .A1(net_1511), .A2(net_984) );
NAND2_X1 inst_4326 ( .ZN(net_4538), .A2(net_3870), .A1(net_2099) );
OAI22_X2 inst_1508 ( .B1(net_4650), .ZN(net_4084), .A2(net_4083), .B2(net_4082), .A1(net_4080) );
SDFF_X2 inst_1222 ( .SI(net_7196), .Q(net_7196), .D(net_3806), .SE(net_3751), .CK(net_13309) );
CLKBUF_X2 inst_9151 ( .A(net_8696), .Z(net_9113) );
CLKBUF_X2 inst_7938 ( .A(net_7846), .Z(net_7900) );
CLKBUF_X2 inst_13985 ( .A(net_13946), .Z(net_13947) );
CLKBUF_X2 inst_11366 ( .A(net_10816), .Z(net_11328) );
NAND2_X2 inst_3407 ( .ZN(net_3746), .A2(net_3339), .A1(net_872) );
SDFF_X2 inst_1073 ( .SI(net_7224), .Q(net_7224), .D(net_3821), .SE(net_3751), .CK(net_10621) );
NOR2_X2 inst_2323 ( .A2(net_6295), .A1(net_5843), .ZN(net_5818) );
NAND2_X2 inst_3741 ( .A1(net_6625), .A2(net_1624), .ZN(net_1604) );
OAI22_X2 inst_1449 ( .B1(net_4855), .ZN(net_4625), .B2(net_4624), .A2(net_4622), .A1(net_4220) );
SDFF_X2 inst_127 ( .QN(net_6194), .SI(net_6193), .D(net_3920), .SE(net_392), .CK(net_13749) );
CLKBUF_X2 inst_11279 ( .A(net_11240), .Z(net_11241) );
CLKBUF_X2 inst_10657 ( .A(net_8137), .Z(net_10619) );
INV_X4 inst_5657 ( .A(net_7417), .ZN(net_2166) );
CLKBUF_X2 inst_11614 ( .A(net_11575), .Z(net_11576) );
CLKBUF_X2 inst_7872 ( .A(net_7827), .Z(net_7834) );
SDFF_X2 inst_187 ( .Q(net_6267), .SI(net_6266), .D(net_3519), .SE(net_392), .CK(net_13477) );
SDFF_X2 inst_206 ( .Q(net_6308), .SI(net_6307), .D(net_3671), .SE(net_392), .CK(net_13564) );
CLKBUF_X2 inst_14270 ( .A(net_14231), .Z(net_14232) );
NAND2_X2 inst_3739 ( .A1(net_6626), .A2(net_1624), .ZN(net_1606) );
NAND2_X2 inst_3029 ( .A1(net_7019), .ZN(net_4980), .A2(net_4979) );
SDFF_X2 inst_1268 ( .Q(net_6691), .D(net_3435), .SI(net_3434), .SE(net_2241), .CK(net_9689) );
XNOR2_X2 inst_122 ( .ZN(net_5868), .B(net_1645), .A(net_831) );
CLKBUF_X2 inst_8944 ( .A(net_7898), .Z(net_8906) );
SDFF_X2 inst_405 ( .SI(net_7369), .Q(net_7369), .D(net_4781), .SE(net_3853), .CK(net_9902) );
CLKBUF_X2 inst_9740 ( .A(net_9701), .Z(net_9702) );
DFF_X1 inst_6436 ( .QN(net_6079), .D(net_5734), .CK(net_11286) );
INV_X4 inst_4788 ( .A(net_3044), .ZN(net_1717) );
CLKBUF_X2 inst_10505 ( .A(net_10466), .Z(net_10467) );
HA_X1 inst_6166 ( .S(net_1708), .CO(net_1707), .B(net_1228), .A(net_1043) );
DFF_X2 inst_6281 ( .QN(net_7689), .D(net_2563), .CK(net_9498) );
AOI222_X2 inst_7540 ( .C1(net_7675), .A1(net_7643), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1882), .B1(net_1881) );
CLKBUF_X2 inst_10077 ( .A(net_10038), .Z(net_10039) );
NAND2_X2 inst_3912 ( .A1(net_6969), .A2(net_1833), .ZN(net_1394) );
CLKBUF_X2 inst_12833 ( .A(net_12794), .Z(net_12795) );
CLKBUF_X2 inst_8499 ( .A(net_8286), .Z(net_8461) );
NOR2_X2 inst_2306 ( .A2(net_6208), .A1(net_5840), .ZN(net_5835) );
DFF_X1 inst_6776 ( .QN(net_6104), .D(net_4326), .CK(net_11170) );
CLKBUF_X2 inst_13087 ( .A(net_13048), .Z(net_13049) );
CLKBUF_X2 inst_9191 ( .A(net_9152), .Z(net_9153) );
INV_X4 inst_5645 ( .A(net_7413), .ZN(net_2194) );
CLKBUF_X2 inst_13046 ( .A(net_13007), .Z(net_13008) );
CLKBUF_X2 inst_14008 ( .A(net_13969), .Z(net_13970) );
OAI221_X2 inst_1646 ( .ZN(net_5384), .C2(net_5383), .B2(net_5089), .A(net_4528), .B1(net_2425), .C1(net_1083) );
NOR4_X2 inst_2176 ( .A2(net_7750), .ZN(net_3319), .A3(net_3208), .A1(net_2923), .A4(net_687) );
DFF_X1 inst_6748 ( .QN(net_7603), .D(net_4852), .CK(net_10825) );
INV_X2 inst_5773 ( .ZN(net_2972), .A(net_2875) );
NAND2_X4 inst_2892 ( .ZN(net_3869), .A2(net_3437), .A1(net_3259) );
AOI222_X2 inst_7547 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1863), .A1(net_1862), .B1(net_1861), .C1(net_1860) );
CLKBUF_X2 inst_13664 ( .A(net_10103), .Z(net_13626) );
DFF_X1 inst_6741 ( .QN(net_7316), .D(net_4862), .CK(net_12685) );
DFF_X2 inst_6294 ( .QN(net_5965), .D(net_1660), .CK(net_12529) );
DFF_X1 inst_6339 ( .D(net_5847), .CK(net_14388), .Q(x14) );
INV_X4 inst_5550 ( .A(net_6172), .ZN(net_3552) );
SDFF_X2 inst_1102 ( .SI(net_6791), .Q(net_6791), .D(net_3806), .SE(net_3729), .CK(net_8269) );
CLKBUF_X2 inst_13024 ( .A(net_12985), .Z(net_12986) );
DFF_X1 inst_6368 ( .QN(net_6294), .D(net_5816), .CK(net_13789) );
CLKBUF_X2 inst_11663 ( .A(net_10290), .Z(net_11625) );
AND3_X2 inst_7804 ( .ZN(net_1667), .A1(net_1666), .A3(net_1665), .A2(net_684) );
CLKBUF_X2 inst_13329 ( .A(net_13290), .Z(net_13291) );
CLKBUF_X2 inst_9795 ( .A(net_9756), .Z(net_9757) );
INV_X4 inst_5365 ( .A(net_7725), .ZN(net_2931) );
SDFF_X2 inst_702 ( .SI(net_6773), .Q(net_6773), .SE(net_3872), .D(net_3787), .CK(net_8517) );
NOR2_X2 inst_2482 ( .A2(net_5778), .ZN(net_2675), .A1(net_2597) );
INV_X2 inst_5860 ( .ZN(net_920), .A(net_612) );
NAND2_X2 inst_2957 ( .ZN(net_5483), .A1(net_4936), .A2(net_4935) );
CLKBUF_X2 inst_12448 ( .A(net_12409), .Z(net_12410) );
CLKBUF_X2 inst_10880 ( .A(net_10841), .Z(net_10842) );
CLKBUF_X2 inst_9297 ( .A(net_9258), .Z(net_9259) );
NAND3_X2 inst_2711 ( .ZN(net_2466), .A2(net_1818), .A3(net_1597), .A1(net_1379) );
CLKBUF_X2 inst_12808 ( .A(net_12769), .Z(net_12770) );
CLKBUF_X2 inst_9980 ( .A(net_9941), .Z(net_9942) );
NAND2_X2 inst_3531 ( .ZN(net_2536), .A2(net_2072), .A1(net_1453) );
NAND3_X2 inst_2753 ( .ZN(net_2348), .A3(net_1566), .A1(net_1371), .A2(net_1002) );
NAND2_X2 inst_3672 ( .A2(net_1798), .ZN(net_1786), .A1(net_1785) );
CLKBUF_X2 inst_14329 ( .A(net_13944), .Z(net_14291) );
SDFF_X2 inst_132 ( .Q(net_6218), .SI(net_6217), .SE(net_392), .D(net_152), .CK(net_14239) );
CLKBUF_X2 inst_10353 ( .A(net_10314), .Z(net_10315) );
CLKBUF_X2 inst_13900 ( .A(net_13861), .Z(net_13862) );
CLKBUF_X2 inst_11502 ( .A(net_11463), .Z(net_11464) );
CLKBUF_X2 inst_12233 ( .A(net_12194), .Z(net_12195) );
CLKBUF_X2 inst_12619 ( .A(net_12580), .Z(net_12581) );
CLKBUF_X2 inst_13912 ( .A(net_13831), .Z(net_13874) );
CLKBUF_X2 inst_9049 ( .A(net_9010), .Z(net_9011) );
CLKBUF_X2 inst_10369 ( .A(net_9660), .Z(net_10331) );
CLKBUF_X2 inst_7935 ( .A(net_7896), .Z(net_7897) );
INV_X1 inst_6149 ( .A(net_3401), .ZN(net_3328) );
NAND2_X2 inst_3545 ( .ZN(net_2522), .A2(net_2080), .A1(net_1752) );
CLKBUF_X2 inst_12365 ( .A(net_12326), .Z(net_12327) );
CLKBUF_X2 inst_13335 ( .A(net_13296), .Z(net_13297) );
NAND2_X2 inst_3611 ( .ZN(net_2336), .A2(net_1834), .A1(net_1644) );
NAND2_X2 inst_2928 ( .ZN(net_5525), .A1(net_4999), .A2(net_4998) );
NAND2_X2 inst_3813 ( .A1(net_6907), .A2(net_1639), .ZN(net_1532) );
SDFF_X2 inst_400 ( .SI(net_7342), .Q(net_7342), .D(net_4784), .SE(net_3856), .CK(net_12355) );
NAND2_X2 inst_2991 ( .A1(net_6755), .A2(net_5033), .ZN(net_5020) );
CLKBUF_X2 inst_8895 ( .A(net_8055), .Z(net_8857) );
CLKBUF_X2 inst_12612 ( .A(net_12068), .Z(net_12574) );
DFF_X2 inst_6309 ( .QN(net_7794), .CK(net_11827), .D(x1587) );
NAND2_X2 inst_3513 ( .ZN(net_2554), .A2(net_2153), .A1(net_1519) );
SDFF_X2 inst_261 ( .Q(net_6373), .SI(net_6372), .D(net_3491), .SE(net_392), .CK(net_14086) );
CLKBUF_X2 inst_12418 ( .A(net_12379), .Z(net_12380) );
SDFF_X2 inst_268 ( .D(net_6400), .SE(net_5800), .SI(net_365), .Q(net_365), .CK(net_14161) );
OAI22_X2 inst_1518 ( .B1(net_4650), .B2(net_4460), .A2(net_4082), .A1(net_4080), .ZN(net_4060) );
CLKBUF_X2 inst_10985 ( .A(net_10946), .Z(net_10947) );
CLKBUF_X2 inst_8198 ( .A(net_8115), .Z(net_8160) );
CLKBUF_X2 inst_8586 ( .A(net_8262), .Z(net_8548) );
NAND2_X2 inst_3975 ( .ZN(net_1295), .A1(net_885), .A2(net_322) );
CLKBUF_X2 inst_11025 ( .A(net_10986), .Z(net_10987) );
CLKBUF_X2 inst_10976 ( .A(net_10701), .Z(net_10938) );
SDFF_X2 inst_327 ( .SI(net_7492), .Q(net_7492), .D(net_5101), .SE(net_3989), .CK(net_9773) );
CLKBUF_X2 inst_9199 ( .A(net_9160), .Z(net_9161) );
CLKBUF_X2 inst_12264 ( .A(net_10329), .Z(net_12226) );
CLKBUF_X2 inst_8874 ( .A(net_8835), .Z(net_8836) );
AND3_X2 inst_7801 ( .ZN(net_2592), .A1(net_2591), .A2(net_2590), .A3(net_2584) );
AOI22_X2 inst_7245 ( .B1(net_6813), .A1(net_6781), .ZN(net_5317), .A2(net_5316), .B2(net_5315) );
CLKBUF_X2 inst_14118 ( .A(net_14079), .Z(net_14080) );
NAND2_X2 inst_3509 ( .ZN(net_2558), .A2(net_2187), .A1(net_1396) );
CLKBUF_X2 inst_13936 ( .A(net_13897), .Z(net_13898) );
CLKBUF_X2 inst_9431 ( .A(net_9392), .Z(net_9393) );
CLKBUF_X2 inst_10746 ( .A(net_10707), .Z(net_10708) );
CLKBUF_X2 inst_7971 ( .A(net_7932), .Z(net_7933) );
NAND2_X2 inst_3853 ( .A1(net_6698), .A2(net_1497), .ZN(net_1482) );
CLKBUF_X2 inst_8044 ( .A(net_7895), .Z(net_8006) );
DFF_X1 inst_6702 ( .QN(net_7285), .D(net_5373), .CK(net_9446) );
CLKBUF_X2 inst_11511 ( .A(net_11472), .Z(net_11473) );
CLKBUF_X2 inst_14304 ( .A(net_14265), .Z(net_14266) );
CLKBUF_X2 inst_12421 ( .A(net_9511), .Z(net_12383) );
CLKBUF_X2 inst_7905 ( .A(net_7866), .Z(net_7867) );
DFF_X1 inst_6348 ( .QN(net_6210), .D(net_5836), .CK(net_13936) );
CLKBUF_X2 inst_9229 ( .A(net_9190), .Z(net_9191) );
CLKBUF_X2 inst_8357 ( .A(net_8318), .Z(net_8319) );
NAND2_X2 inst_3097 ( .A1(net_6444), .A2(net_4925), .ZN(net_4906) );
CLKBUF_X2 inst_10739 ( .A(net_9743), .Z(net_10701) );
CLKBUF_X2 inst_9625 ( .A(net_8747), .Z(net_9587) );
NAND2_X2 inst_3661 ( .A1(net_7068), .ZN(net_1802), .A2(net_791) );
CLKBUF_X2 inst_13678 ( .A(net_13639), .Z(net_13640) );
SDFF_X2 inst_502 ( .SI(net_6900), .Q(net_6900), .D(net_3883), .SE(net_3781), .CK(net_8894) );
CLKBUF_X2 inst_14244 ( .A(net_9097), .Z(net_14206) );
CLKBUF_X2 inst_13976 ( .A(net_13937), .Z(net_13938) );
CLKBUF_X2 inst_9001 ( .A(net_8408), .Z(net_8963) );
CLKBUF_X2 inst_11836 ( .A(net_11797), .Z(net_11798) );
CLKBUF_X2 inst_8745 ( .A(net_8706), .Z(net_8707) );
NAND2_X2 inst_3221 ( .ZN(net_4705), .A2(net_3986), .A1(net_1841) );
NAND2_X2 inst_3645 ( .A1(net_7073), .ZN(net_1818), .A2(net_791) );
OAI22_X2 inst_1598 ( .A1(net_3287), .B2(net_3200), .A2(net_3144), .ZN(net_3138), .B1(net_697) );
CLKBUF_X2 inst_12335 ( .A(net_12296), .Z(net_12297) );
SDFF_X2 inst_357 ( .SI(net_7604), .Q(net_7604), .D(net_4792), .SE(net_3870), .CK(net_13258) );
CLKBUF_X2 inst_11083 ( .A(net_11044), .Z(net_11045) );
DFFR_X2 inst_6969 ( .QN(net_6004), .D(net_4005), .CK(net_12568), .RN(x1822) );
CLKBUF_X2 inst_10028 ( .A(net_9103), .Z(net_9990) );
CLKBUF_X2 inst_10167 ( .A(net_9061), .Z(net_10129) );
HA_X1 inst_6173 ( .B(net_6413), .A(net_6412), .S(net_693), .CO(net_692) );
NAND2_X2 inst_4092 ( .A1(net_7206), .A2(net_1648), .ZN(net_960) );
CLKBUF_X2 inst_13865 ( .A(net_8652), .Z(net_13827) );
CLKBUF_X2 inst_10098 ( .A(net_9499), .Z(net_10060) );
CLKBUF_X2 inst_7880 ( .A(net_7841), .Z(net_7842) );
NAND2_X2 inst_3980 ( .ZN(net_1290), .A1(net_885), .A2(net_314) );
NAND2_X2 inst_3152 ( .ZN(net_4811), .A2(net_4153), .A1(net_2115) );
CLKBUF_X2 inst_11438 ( .A(net_11399), .Z(net_11400) );
NAND2_X2 inst_4161 ( .ZN(net_1048), .A2(net_609), .A1(net_563) );
NAND2_X2 inst_3758 ( .A1(net_6639), .A2(net_1624), .ZN(net_1587) );
SDFF_X2 inst_912 ( .Q(net_7246), .D(net_7246), .SE(net_3822), .SI(net_342), .CK(net_12671) );
CLKBUF_X2 inst_10065 ( .A(net_10026), .Z(net_10027) );
CLKBUF_X2 inst_11678 ( .A(net_8333), .Z(net_11640) );
CLKBUF_X2 inst_10117 ( .A(net_10078), .Z(net_10079) );
INV_X2 inst_5869 ( .A(net_816), .ZN(net_507) );
NAND2_X2 inst_3196 ( .ZN(net_4730), .A2(net_3986), .A1(net_1851) );
CLKBUF_X2 inst_12724 ( .A(net_10823), .Z(net_12686) );
INV_X2 inst_5872 ( .A(net_820), .ZN(net_430) );
DFF_X1 inst_6525 ( .QN(net_7441), .D(net_5426), .CK(net_12110) );
NAND2_X2 inst_4025 ( .A1(net_6797), .A2(net_1651), .ZN(net_1027) );
SDFF_X2 inst_322 ( .SI(net_7487), .Q(net_7487), .D(net_5105), .SE(net_3989), .CK(net_9781) );
CLKBUF_X2 inst_10070 ( .A(net_10031), .Z(net_10032) );
NAND2_X2 inst_3516 ( .ZN(net_2551), .A2(net_2155), .A1(net_1357) );
DFFR_X2 inst_6988 ( .QN(net_7694), .D(net_3348), .CK(net_10371), .RN(x1822) );
NAND2_X2 inst_4200 ( .ZN(net_1826), .A1(net_629), .A2(net_308) );
NAND2_X2 inst_4188 ( .ZN(net_1747), .A1(net_565), .A2(net_271) );
CLKBUF_X2 inst_14405 ( .A(net_13511), .Z(net_14367) );
NAND2_X2 inst_4169 ( .ZN(net_923), .A1(net_601), .A2(net_498) );
NAND2_X2 inst_3902 ( .A1(net_6971), .A2(net_1833), .ZN(net_1408) );
CLKBUF_X2 inst_10858 ( .A(net_10694), .Z(net_10820) );
CLKBUF_X2 inst_9894 ( .A(net_9855), .Z(net_9856) );
DFF_X2 inst_6191 ( .QN(net_7094), .D(net_5058), .CK(net_12205) );
DFF_X1 inst_6863 ( .D(net_2535), .QN(net_212), .CK(net_12613) );
CLKBUF_X2 inst_10647 ( .A(net_10608), .Z(net_10609) );
DFF_X2 inst_6243 ( .QN(net_7753), .D(net_3025), .CK(net_10403) );
CLKBUF_X2 inst_8302 ( .A(net_8263), .Z(net_8264) );
DFF_X1 inst_6908 ( .D(net_2501), .Q(net_160), .CK(net_12218) );
INV_X4 inst_5346 ( .A(net_6112), .ZN(net_3671) );
DFF_X2 inst_6289 ( .Q(net_6384), .D(net_6383), .CK(net_14168) );
NAND2_X2 inst_4181 ( .ZN(net_706), .A1(net_705), .A2(net_473) );
CLKBUF_X2 inst_12662 ( .A(net_12623), .Z(net_12624) );
NOR2_X2 inst_2315 ( .A2(net_6239), .A1(net_5840), .ZN(net_5826) );
SDFF_X2 inst_962 ( .Q(net_6440), .D(net_6440), .SE(net_3820), .SI(net_3809), .CK(net_8494) );
CLKBUF_X2 inst_10865 ( .A(net_10826), .Z(net_10827) );
DFF_X1 inst_6350 ( .QN(net_6208), .D(net_5834), .CK(net_13716) );
OAI21_X2 inst_2008 ( .B1(net_5904), .B2(net_4518), .ZN(net_4503), .A(net_3672) );
SDFF_X2 inst_641 ( .SI(net_6653), .Q(net_6653), .SE(net_3850), .D(net_3801), .CK(net_9103) );
SDFF_X2 inst_498 ( .SI(net_6491), .Q(net_6491), .D(net_3892), .SE(net_3886), .CK(net_8796) );
OAI21_X2 inst_1988 ( .B1(net_4851), .ZN(net_4841), .A(net_4561), .B2(net_3866) );
CLKBUF_X2 inst_11489 ( .A(net_11450), .Z(net_11451) );
CLKBUF_X2 inst_9673 ( .A(net_9634), .Z(net_9635) );
CLKBUF_X2 inst_8374 ( .A(net_8335), .Z(net_8336) );
CLKBUF_X2 inst_12346 ( .A(net_8981), .Z(net_12308) );
CLKBUF_X2 inst_8287 ( .A(net_8248), .Z(net_8249) );
CLKBUF_X2 inst_11971 ( .A(net_8376), .Z(net_11933) );
CLKBUF_X2 inst_7955 ( .A(net_7916), .Z(net_7917) );
INV_X4 inst_5517 ( .A(net_6170), .ZN(net_3556) );
OAI21_X2 inst_1912 ( .ZN(net_5156), .B1(net_4870), .A(net_4758), .B2(net_3941) );
CLKBUF_X2 inst_14044 ( .A(net_14005), .Z(net_14006) );
OAI21_X2 inst_1831 ( .ZN(net_5348), .B1(net_5347), .A(net_4358), .B2(net_3856) );
CLKBUF_X2 inst_13438 ( .A(net_12580), .Z(net_13400) );
CLKBUF_X2 inst_9308 ( .A(net_9269), .Z(net_9270) );
DFF_X1 inst_6714 ( .QN(net_7330), .D(net_5352), .CK(net_9878) );
DFF_X1 inst_6683 ( .QN(net_7271), .D(net_5121), .CK(net_9887) );
CLKBUF_X2 inst_14339 ( .A(net_14300), .Z(net_14301) );
CLKBUF_X2 inst_13671 ( .A(net_13632), .Z(net_13633) );
NAND2_X2 inst_3468 ( .A1(net_7743), .A2(net_2957), .ZN(net_2756) );
CLKBUF_X2 inst_11876 ( .A(net_11837), .Z(net_11838) );
SDFF_X2 inst_350 ( .SI(net_7645), .Q(net_7645), .D(net_4802), .SE(net_3867), .CK(net_10280) );
CLKBUF_X2 inst_11322 ( .A(net_11283), .Z(net_11284) );
NOR2_X2 inst_2395 ( .A2(net_3996), .ZN(net_3990), .A1(net_890) );
SDFF_X2 inst_231 ( .Q(net_6323), .SI(net_6322), .D(net_3639), .SE(net_392), .CK(net_14016) );
CLKBUF_X2 inst_9024 ( .A(net_8098), .Z(net_8986) );
CLKBUF_X2 inst_10403 ( .A(net_10364), .Z(net_10365) );
NAND2_X2 inst_3309 ( .ZN(net_3628), .A1(net_3627), .A2(net_3229) );
CLKBUF_X2 inst_14437 ( .A(net_14398), .Z(net_14399) );
INV_X4 inst_5104 ( .A(net_7795), .ZN(net_3802) );
CLKBUF_X2 inst_9952 ( .A(net_9606), .Z(net_9914) );
INV_X4 inst_5676 ( .A(net_7278), .ZN(net_2025) );
CLKBUF_X2 inst_12851 ( .A(net_12812), .Z(net_12813) );
NOR2_X2 inst_2317 ( .A2(net_6221), .A1(net_5840), .ZN(net_5824) );
CLKBUF_X2 inst_11901 ( .A(net_11862), .Z(net_11863) );
CLKBUF_X2 inst_11365 ( .A(net_10882), .Z(net_11327) );
CLKBUF_X2 inst_8518 ( .A(net_8093), .Z(net_8480) );
AOI222_X2 inst_7506 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2048), .A1(net_2047), .B1(net_2046), .C1(net_2045) );
OAI22_X2 inst_1452 ( .B1(net_4855), .A2(net_4622), .ZN(net_4618), .B2(net_4617), .A1(net_4214) );
CLKBUF_X2 inst_13740 ( .A(net_10385), .Z(net_13702) );
CLKBUF_X2 inst_11867 ( .A(net_11816), .Z(net_11829) );
DFF_X1 inst_6756 ( .QN(net_7300), .D(net_4873), .CK(net_12683) );
DFF_X1 inst_6549 ( .Q(net_7774), .D(net_5608), .CK(net_13291) );
INV_X4 inst_5000 ( .A(net_1730), .ZN(net_869) );
CLKBUF_X2 inst_12967 ( .A(net_10152), .Z(net_12929) );
NAND2_X2 inst_4077 ( .A1(net_6930), .A2(net_1654), .ZN(net_975) );
NAND2_X2 inst_3139 ( .ZN(net_4824), .A2(net_4153), .A1(net_2156) );
CLKBUF_X2 inst_12801 ( .A(net_12762), .Z(net_12763) );
NAND4_X2 inst_2558 ( .A4(net_7690), .ZN(net_2616), .A3(net_1218), .A2(net_836), .A1(x1155) );
OR2_X4 inst_1396 ( .A2(net_6689), .A1(net_6688), .ZN(net_528) );
SDFF_X2 inst_352 ( .SI(net_7637), .Q(net_7637), .D(net_4801), .SE(net_3867), .CK(net_8007) );
SDFF_X2 inst_286 ( .D(net_6396), .SE(net_5800), .SI(net_361), .Q(net_361), .CK(net_13673) );
CLKBUF_X2 inst_13354 ( .A(net_11479), .Z(net_13316) );
CLKBUF_X2 inst_10112 ( .A(net_10073), .Z(net_10074) );
DFF_X1 inst_6880 ( .D(net_2523), .Q(net_236), .CK(net_13055) );
CLKBUF_X2 inst_8901 ( .A(net_8311), .Z(net_8863) );
CLKBUF_X2 inst_10447 ( .A(net_10408), .Z(net_10409) );
CLKBUF_X2 inst_12984 ( .A(net_12945), .Z(net_12946) );
CLKBUF_X2 inst_13006 ( .A(net_12967), .Z(net_12968) );
CLKBUF_X2 inst_7961 ( .A(net_7922), .Z(net_7923) );
NAND2_X2 inst_3003 ( .A1(net_6851), .ZN(net_5008), .A2(net_5004) );
DFF_X1 inst_6792 ( .D(net_3947), .CK(net_12470), .Q(x561) );
CLKBUF_X2 inst_12169 ( .A(net_12130), .Z(net_12131) );
INV_X4 inst_5579 ( .A(net_6141), .ZN(net_3651) );
NAND2_X2 inst_3841 ( .A1(net_6700), .ZN(net_1498), .A2(net_1497) );
CLKBUF_X2 inst_13134 ( .A(net_13095), .Z(net_13096) );
CLKBUF_X2 inst_9555 ( .A(net_9516), .Z(net_9517) );
CLKBUF_X2 inst_9165 ( .A(net_9126), .Z(net_9127) );
CLKBUF_X2 inst_8550 ( .A(net_8511), .Z(net_8512) );
NOR3_X4 inst_2185 ( .ZN(net_1672), .A2(net_624), .A3(net_615), .A1(net_483) );
NAND2_X2 inst_4050 ( .A1(net_6942), .A2(net_1654), .ZN(net_1002) );
AOI21_X2 inst_7737 ( .B1(net_7141), .ZN(net_4083), .B2(net_2582), .A(net_2325) );
DFFR_X2 inst_6972 ( .QN(net_6037), .D(net_4000), .CK(net_10531), .RN(x1822) );
CLKBUF_X2 inst_12203 ( .A(net_12164), .Z(net_12165) );
CLKBUF_X2 inst_9427 ( .A(net_7953), .Z(net_9389) );
NOR2_X2 inst_2370 ( .ZN(net_5215), .A2(net_4616), .A1(net_4448) );
CLKBUF_X2 inst_14069 ( .A(net_14030), .Z(net_14031) );
INV_X2 inst_5887 ( .A(net_7499), .ZN(net_2069) );
NAND2_X2 inst_3882 ( .A1(net_6560), .A2(net_1705), .ZN(net_1437) );
CLKBUF_X2 inst_11598 ( .A(net_11559), .Z(net_11560) );
CLKBUF_X2 inst_13452 ( .A(net_8634), .Z(net_13414) );
NAND3_X2 inst_2811 ( .ZN(net_2287), .A3(net_1529), .A1(net_1312), .A2(net_944) );
CLKBUF_X2 inst_12001 ( .A(net_8769), .Z(net_11963) );
INV_X16 inst_6120 ( .ZN(net_5031), .A(net_4270) );
INV_X4 inst_4615 ( .ZN(net_4207), .A(net_4075) );
SDFF_X2 inst_137 ( .Q(net_6213), .SI(net_6212), .SE(net_392), .D(net_147), .CK(net_14227) );
DFF_X1 inst_6889 ( .D(net_2495), .Q(net_235), .CK(net_13049) );
SDFF_X2 inst_425 ( .SI(net_7758), .Q(net_7758), .SE(net_5925), .D(net_3907), .CK(net_12518) );
NAND3_X4 inst_2567 ( .A2(net_5934), .ZN(net_3297), .A1(net_2907), .A3(net_689) );
CLKBUF_X2 inst_11384 ( .A(net_11345), .Z(net_11346) );
NAND2_X2 inst_3206 ( .ZN(net_4720), .A2(net_3986), .A1(net_1891) );
CLKBUF_X2 inst_11742 ( .A(net_11703), .Z(net_11704) );
CLKBUF_X2 inst_8416 ( .A(net_8305), .Z(net_8378) );
CLKBUF_X2 inst_8591 ( .A(net_8552), .Z(net_8553) );
NAND3_X2 inst_2572 ( .ZN(net_5767), .A1(net_5662), .A2(net_5290), .A3(net_4236) );
CLKBUF_X2 inst_13764 ( .A(net_13725), .Z(net_13726) );
CLKBUF_X2 inst_9380 ( .A(net_9341), .Z(net_9342) );
DFF_X1 inst_6755 ( .QN(net_6147), .D(net_4856), .CK(net_11972) );
CLKBUF_X2 inst_13111 ( .A(net_13072), .Z(net_13073) );
CLKBUF_X2 inst_10245 ( .A(net_10206), .Z(net_10207) );
NAND2_X2 inst_4046 ( .A1(net_6938), .A2(net_1654), .ZN(net_1006) );
NAND2_X2 inst_3365 ( .ZN(net_3516), .A1(net_3515), .A2(net_3223) );
NAND2_X2 inst_3254 ( .ZN(net_5043), .A1(net_3849), .A2(net_3462) );
CLKBUF_X2 inst_11752 ( .A(net_10324), .Z(net_11714) );
SDFF_X2 inst_983 ( .Q(net_6468), .D(net_6468), .SE(net_3904), .SI(net_3812), .CK(net_11256) );
INV_X4 inst_4980 ( .A(net_6823), .ZN(net_686) );
CLKBUF_X2 inst_8026 ( .A(net_7987), .Z(net_7988) );
CLKBUF_X2 inst_8112 ( .A(net_8073), .Z(net_8074) );
CLKBUF_X2 inst_8511 ( .A(net_8472), .Z(net_8473) );
OAI21_X2 inst_1897 ( .B1(net_5204), .ZN(net_5179), .A(net_4556), .B2(net_3866) );
CLKBUF_X2 inst_10615 ( .A(net_10576), .Z(net_10577) );
AOI21_X2 inst_7773 ( .B1(net_6599), .ZN(net_4032), .B2(net_2583), .A(net_2293) );
CLKBUF_X2 inst_11810 ( .A(net_11771), .Z(net_11772) );
NAND2_X2 inst_3159 ( .ZN(net_4774), .A2(net_3941), .A1(net_2117) );
CLKBUF_X2 inst_11291 ( .A(net_11072), .Z(net_11253) );
CLKBUF_X2 inst_11196 ( .A(net_10546), .Z(net_11158) );
INV_X4 inst_4776 ( .ZN(net_1716), .A(net_1715) );
DFF_X2 inst_6237 ( .D(net_3069), .QN(net_113), .CK(net_10217) );
OAI22_X2 inst_1569 ( .A2(net_3297), .B2(net_3286), .ZN(net_3281), .A1(net_3280), .B1(net_753) );
CLKBUF_X2 inst_11722 ( .A(net_11683), .Z(net_11684) );
CLKBUF_X2 inst_12990 ( .A(net_12951), .Z(net_12952) );
NAND3_X2 inst_2633 ( .ZN(net_5696), .A1(net_5673), .A2(net_5307), .A3(net_4247) );
CLKBUF_X2 inst_13565 ( .A(net_13526), .Z(net_13527) );
AOI22_X2 inst_7314 ( .B1(net_6675), .A1(net_6643), .A2(net_5139), .B2(net_5138), .ZN(net_5125) );
DFFR_X2 inst_7080 ( .QN(net_7732), .D(net_2802), .CK(net_10743), .RN(x1822) );
OAI21_X2 inst_1772 ( .B1(net_5444), .ZN(net_5422), .A(net_4701), .B2(net_3989) );
DFF_X1 inst_6947 ( .Q(net_6380), .CK(net_13836), .D(x806) );
DFF_X2 inst_6274 ( .Q(net_6386), .D(net_6385), .CK(net_14175) );
CLKBUF_X2 inst_13725 ( .A(net_13686), .Z(net_13687) );
OAI21_X2 inst_2143 ( .B1(net_5778), .ZN(net_2801), .A(net_2680), .B2(net_2678) );
CLKBUF_X2 inst_14233 ( .A(net_13519), .Z(net_14195) );
SDFF_X2 inst_1291 ( .D(net_7802), .SE(net_3256), .SI(net_139), .Q(net_139), .CK(net_8460) );
AOI21_X2 inst_7671 ( .B1(net_7006), .ZN(net_4231), .A(net_2457), .B2(net_1100) );
DFFR_X2 inst_7029 ( .QN(net_6012), .D(net_3143), .CK(net_10448), .RN(x1822) );
OAI21_X2 inst_2130 ( .ZN(net_2906), .A(net_2905), .B2(net_2895), .B1(net_903) );
SDFF_X2 inst_359 ( .SI(net_7607), .Q(net_7607), .D(net_4790), .SE(net_3870), .CK(net_8000) );
CLKBUF_X2 inst_8239 ( .A(net_8200), .Z(net_8201) );
NAND2_X1 inst_4388 ( .ZN(net_4339), .A2(net_3859), .A1(net_2214) );
SDFF_X2 inst_1055 ( .Q(net_7134), .D(net_7134), .SE(net_3903), .SI(net_3892), .CK(net_13323) );
CLKBUF_X2 inst_12382 ( .A(net_11351), .Z(net_12344) );
CLKBUF_X2 inst_13114 ( .A(net_10960), .Z(net_13076) );
OAI21_X2 inst_2100 ( .B2(net_7770), .ZN(net_4803), .A(net_4304), .B1(net_407) );
NOR2_X4 inst_2284 ( .ZN(net_5917), .A2(net_5870), .A1(net_3024) );
OAI21_X2 inst_1962 ( .B1(net_5399), .ZN(net_5048), .A(net_4656), .B2(net_3993) );
INV_X4 inst_4829 ( .ZN(net_4792), .A(net_1081) );
INV_X4 inst_4757 ( .A(net_3252), .ZN(net_2578) );
SDFF_X2 inst_923 ( .Q(net_7133), .D(net_7133), .SE(net_3903), .SI(net_3802), .CK(net_13352) );
CLKBUF_X2 inst_13037 ( .A(net_12998), .Z(net_12999) );
CLKBUF_X2 inst_12153 ( .A(net_9460), .Z(net_12115) );
CLKBUF_X2 inst_13582 ( .A(net_13543), .Z(net_13544) );
CLKBUF_X2 inst_10492 ( .A(net_10453), .Z(net_10454) );
CLKBUF_X2 inst_8671 ( .A(net_7885), .Z(net_8633) );
CLKBUF_X2 inst_11551 ( .A(net_11232), .Z(net_11513) );
CLKBUF_X2 inst_8599 ( .A(net_8560), .Z(net_8561) );
CLKBUF_X2 inst_11604 ( .A(net_11565), .Z(net_11566) );
CLKBUF_X2 inst_12925 ( .A(net_12702), .Z(net_12887) );
INV_X4 inst_5283 ( .A(net_7266), .ZN(net_2075) );
CLKBUF_X2 inst_13470 ( .A(net_13431), .Z(net_13432) );
DFFR_X2 inst_6975 ( .QN(net_7786), .D(net_3998), .CK(net_13031), .RN(x1822) );
CLKBUF_X2 inst_8168 ( .A(net_8015), .Z(net_8130) );
DFF_X2 inst_6174 ( .Q(net_6400), .D(net_6399), .CK(net_14199) );
CLKBUF_X2 inst_11819 ( .A(net_9299), .Z(net_11781) );
AOI222_X2 inst_7564 ( .A1(net_7243), .ZN(net_5335), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_337), .C2(net_335) );
SDFF_X2 inst_194 ( .SI(net_6299), .Q(net_6260), .D(net_3517), .SE(net_392), .CK(net_13775) );
CLKBUF_X2 inst_8421 ( .A(net_8322), .Z(net_8383) );
DFFR_X2 inst_7109 ( .D(net_1950), .QN(net_121), .CK(net_12312), .RN(x1822) );
INV_X2 inst_5890 ( .A(net_7474), .ZN(net_2189) );
NAND2_X2 inst_3453 ( .A2(net_5925), .ZN(net_2919), .A1(net_1211) );
CLKBUF_X2 inst_8793 ( .A(net_8754), .Z(net_8755) );
AOI21_X2 inst_7686 ( .B1(net_6605), .ZN(net_4022), .B2(net_2583), .A(net_2289) );
CLKBUF_X2 inst_12946 ( .A(net_12907), .Z(net_12908) );
NAND2_X2 inst_3766 ( .A1(net_7178), .A2(net_1637), .ZN(net_1579) );
CLKBUF_X2 inst_12480 ( .A(net_8941), .Z(net_12442) );
CLKBUF_X2 inst_14181 ( .A(net_14142), .Z(net_14143) );
INV_X2 inst_5935 ( .A(net_7284), .ZN(net_2019) );
CLKBUF_X2 inst_8714 ( .A(net_8675), .Z(net_8676) );
INV_X16 inst_6136 ( .ZN(net_1675), .A(net_881) );
AOI21_X2 inst_7704 ( .B1(net_6734), .ZN(net_4134), .B2(net_2581), .A(net_2374) );
CLKBUF_X2 inst_11317 ( .A(net_11278), .Z(net_11279) );
NOR2_X2 inst_2536 ( .A2(net_6827), .ZN(net_1251), .A1(net_571) );
CLKBUF_X2 inst_11730 ( .A(net_11691), .Z(net_11692) );
CLKBUF_X2 inst_13103 ( .A(net_13064), .Z(net_13065) );
CLKBUF_X2 inst_9389 ( .A(net_9350), .Z(net_9351) );
DFFR_X2 inst_7100 ( .D(net_1946), .QN(net_120), .CK(net_9591), .RN(x1822) );
SDFF_X2 inst_442 ( .Q(net_7396), .D(net_7396), .SE(net_3994), .SI(net_361), .CK(net_9631) );
CLKBUF_X2 inst_9618 ( .A(net_9579), .Z(net_9580) );
NOR2_X2 inst_2507 ( .ZN(net_1237), .A2(net_669), .A1(net_666) );
CLKBUF_X2 inst_9337 ( .A(net_9298), .Z(net_9299) );
CLKBUF_X2 inst_8338 ( .A(net_8299), .Z(net_8300) );
NOR2_X4 inst_2245 ( .ZN(net_5641), .A1(net_5487), .A2(net_4453) );
CLKBUF_X2 inst_14036 ( .A(net_12302), .Z(net_13998) );
CLKBUF_X2 inst_12620 ( .A(net_12581), .Z(net_12582) );
DFF_X1 inst_6870 ( .D(net_2545), .Q(net_220), .CK(net_9529) );
INV_X4 inst_5237 ( .A(net_845), .ZN(net_454) );
CLKBUF_X2 inst_13300 ( .A(net_13261), .Z(net_13262) );
INV_X2 inst_5915 ( .A(net_7359), .ZN(net_2062) );
INV_X2 inst_6097 ( .A(net_7349), .ZN(net_2008) );
CLKBUF_X2 inst_10998 ( .A(net_9158), .Z(net_10960) );
OAI21_X2 inst_1925 ( .ZN(net_5120), .A(net_4771), .B2(net_3941), .B1(net_1267) );
NAND2_X1 inst_4298 ( .ZN(net_4568), .A2(net_3866), .A1(net_1893) );
CLKBUF_X2 inst_11242 ( .A(net_11203), .Z(net_11204) );
XNOR2_X2 inst_40 ( .ZN(net_2422), .B(net_2421), .A(net_1272) );
NAND2_X1 inst_4437 ( .A2(net_2131), .ZN(net_1373), .A1(net_1372) );
SDFF_X2 inst_1249 ( .SI(net_6545), .Q(net_6545), .D(net_3902), .SE(net_3756), .CK(net_8392) );
NAND2_X2 inst_4099 ( .A1(net_6670), .A2(net_1655), .ZN(net_953) );
CLKBUF_X2 inst_8765 ( .A(net_8404), .Z(net_8727) );
INV_X4 inst_5403 ( .A(net_7254), .ZN(net_2216) );
INV_X4 inst_4740 ( .ZN(net_2751), .A(net_2750) );
OR2_X2 inst_1416 ( .ZN(net_3770), .A2(net_788), .A1(net_596) );
INV_X2 inst_5967 ( .ZN(net_406), .A(x889) );
CLKBUF_X2 inst_12066 ( .A(net_8767), .Z(net_12028) );
SDFF_X2 inst_1318 ( .D(net_6381), .SE(net_5801), .SI(net_326), .Q(net_326), .CK(net_13860) );
DFF_X1 inst_6894 ( .D(net_2494), .Q(net_171), .CK(net_12225) );
AOI22_X2 inst_7280 ( .B1(net_7217), .A1(net_7185), .ZN(net_5250), .A2(net_5244), .B2(net_5243) );
SDFF_X2 inst_439 ( .Q(net_7390), .D(net_7390), .SE(net_3994), .SI(net_355), .CK(net_9636) );
CLKBUF_X2 inst_11567 ( .A(net_9555), .Z(net_11529) );
INV_X8 inst_4529 ( .A(net_3297), .ZN(net_3286) );
INV_X4 inst_4584 ( .A(net_5049), .ZN(net_4328) );
SDFF_X2 inst_1070 ( .SI(net_6521), .Q(net_6521), .D(net_3806), .SE(net_3755), .CK(net_11547) );
CLKBUF_X2 inst_12037 ( .A(net_8190), .Z(net_11999) );
NOR2_X2 inst_2454 ( .ZN(net_2816), .A2(net_2692), .A1(net_1171) );
CLKBUF_X2 inst_12255 ( .A(net_12216), .Z(net_12217) );
CLKBUF_X2 inst_8280 ( .A(net_7907), .Z(net_8242) );
NAND2_X2 inst_3601 ( .ZN(net_2399), .A2(net_1870), .A1(net_1316) );
CLKBUF_X2 inst_9693 ( .A(net_9654), .Z(net_9655) );
INV_X8 inst_4536 ( .A(net_6053), .ZN(net_5801) );
CLKBUF_X2 inst_13309 ( .A(net_9253), .Z(net_13271) );
CLKBUF_X2 inst_13475 ( .A(net_13436), .Z(net_13437) );
CLKBUF_X2 inst_9478 ( .A(net_9439), .Z(net_9440) );
CLKBUF_X2 inst_11854 ( .A(net_10309), .Z(net_11816) );
INV_X4 inst_5601 ( .A(net_6556), .ZN(net_491) );
DFF_X1 inst_6763 ( .QN(net_6086), .D(net_4641), .CK(net_12949) );
SDFF_X2 inst_654 ( .Q(net_6711), .D(net_6711), .SE(net_3871), .SI(net_3808), .CK(net_8522) );
OAI221_X2 inst_1673 ( .C2(net_4300), .ZN(net_4169), .B2(net_4168), .C1(net_4152), .A(net_3984), .B1(net_1927) );
INV_X2 inst_5745 ( .ZN(net_3719), .A(net_3416) );
CLKBUF_X2 inst_13616 ( .A(net_8327), .Z(net_13578) );
CLKBUF_X2 inst_14373 ( .A(net_14334), .Z(net_14335) );
CLKBUF_X2 inst_13656 ( .A(net_12017), .Z(net_13618) );
OAI21_X2 inst_1708 ( .ZN(net_5586), .A(net_5153), .B2(net_4439), .B1(net_4057) );
SDFF_X2 inst_1153 ( .SI(net_6815), .Q(net_6815), .D(net_3898), .SE(net_3722), .CK(net_8340) );
CLKBUF_X2 inst_7959 ( .A(net_7911), .Z(net_7921) );
AOI21_X2 inst_7632 ( .ZN(net_4296), .B2(net_3450), .B1(net_3178), .A(x868) );
NAND2_X2 inst_3823 ( .A1(net_6840), .ZN(net_1522), .A2(net_1521) );
CLKBUF_X2 inst_10905 ( .A(net_10866), .Z(net_10867) );
AOI22_X2 inst_7325 ( .ZN(net_3427), .A2(net_3426), .B2(net_3425), .A1(net_1335), .B1(net_901) );
SDFF_X2 inst_391 ( .SI(net_7312), .Q(net_7312), .D(net_4777), .SE(net_3859), .CK(net_12211) );
CLKBUF_X2 inst_11997 ( .A(net_11958), .Z(net_11959) );
NAND2_X2 inst_4107 ( .A1(net_6535), .A2(net_1645), .ZN(net_945) );
CLKBUF_X2 inst_10440 ( .A(net_9207), .Z(net_10402) );
CLKBUF_X2 inst_11004 ( .A(net_10965), .Z(net_10966) );
NAND3_X2 inst_2738 ( .ZN(net_2363), .A3(net_1564), .A1(net_1433), .A2(net_1019) );
SDFF_X2 inst_634 ( .SI(net_6646), .Q(net_6646), .SE(net_3850), .D(net_3803), .CK(net_10657) );
NAND2_X2 inst_3122 ( .A1(net_6579), .A2(net_4897), .ZN(net_4879) );
CLKBUF_X2 inst_14092 ( .A(net_14053), .Z(net_14054) );
CLKBUF_X2 inst_9090 ( .A(net_9051), .Z(net_9052) );
CLKBUF_X2 inst_10896 ( .A(net_10625), .Z(net_10858) );
CLKBUF_X2 inst_8035 ( .A(net_7996), .Z(net_7997) );
CLKBUF_X2 inst_9232 ( .A(net_8768), .Z(net_9194) );
CLKBUF_X2 inst_10420 ( .A(net_7945), .Z(net_10382) );
INV_X2 inst_6074 ( .A(net_7466), .ZN(net_2181) );
OAI22_X2 inst_1477 ( .B1(net_4855), .A1(net_4228), .B2(net_4218), .ZN(net_4215), .A2(net_4214) );
CLKBUF_X2 inst_13774 ( .A(net_13735), .Z(net_13736) );
CLKBUF_X2 inst_9263 ( .A(net_9078), .Z(net_9225) );
CLKBUF_X2 inst_8403 ( .A(net_8343), .Z(net_8365) );
DFFR_X2 inst_7043 ( .QN(net_6008), .D(net_3175), .CK(net_11424), .RN(x1822) );
OAI21_X2 inst_1799 ( .ZN(net_5391), .A(net_4718), .B2(net_3986), .B1(net_1163) );
CLKBUF_X2 inst_9813 ( .A(net_8256), .Z(net_9775) );
SDFF_X2 inst_529 ( .Q(net_6616), .D(net_6616), .SI(net_3902), .SE(net_3830), .CK(net_12042) );
NAND2_X1 inst_4442 ( .A1(net_7608), .A2(net_2131), .ZN(net_1337) );
AOI22_X2 inst_7385 ( .A2(net_5916), .B2(net_2957), .ZN(net_2935), .B1(net_2934), .A1(net_710) );
OAI22_X2 inst_1528 ( .B1(net_4644), .A1(net_4057), .B2(net_4043), .ZN(net_4040), .A2(net_4039) );
CLKBUF_X2 inst_11192 ( .A(net_8881), .Z(net_11154) );
CLKBUF_X2 inst_9326 ( .A(net_8637), .Z(net_9288) );
NAND2_X2 inst_3458 ( .ZN(net_2978), .A2(net_2740), .A1(net_263) );
INV_X2 inst_5788 ( .A(net_5965), .ZN(net_2240) );
CLKBUF_X2 inst_11788 ( .A(net_11749), .Z(net_11750) );
INV_X4 inst_4694 ( .ZN(net_4138), .A(net_3323) );
SDFF_X2 inst_1313 ( .D(net_6382), .SE(net_5800), .SI(net_347), .Q(net_347), .CK(net_14140) );
CLKBUF_X2 inst_14267 ( .A(net_9772), .Z(net_14229) );
CLKBUF_X2 inst_11030 ( .A(net_10991), .Z(net_10992) );
CLKBUF_X2 inst_11104 ( .A(net_11065), .Z(net_11066) );
CLKBUF_X2 inst_8098 ( .A(net_8059), .Z(net_8060) );
SDFF_X2 inst_675 ( .Q(net_6739), .D(net_6739), .SE(net_3815), .SI(net_3811), .CK(net_11157) );
CLKBUF_X2 inst_8632 ( .A(net_8593), .Z(net_8594) );
NAND2_X2 inst_4068 ( .A1(net_7210), .A2(net_1648), .ZN(net_984) );
CLKBUF_X2 inst_11953 ( .A(net_11914), .Z(net_11915) );
CLKBUF_X2 inst_13706 ( .A(net_13667), .Z(net_13668) );
INV_X2 inst_5729 ( .ZN(net_3966), .A(net_3965) );
NAND2_X2 inst_4116 ( .A2(net_1222), .ZN(net_1177), .A1(net_337) );
NAND2_X4 inst_2886 ( .ZN(net_3992), .A2(net_3743), .A1(net_3340) );
NAND3_X2 inst_2705 ( .ZN(net_2472), .A2(net_1808), .A3(net_1581), .A1(net_1388) );
DFF_X1 inst_6523 ( .QN(net_7439), .D(net_5428), .CK(net_9278) );
INV_X4 inst_5150 ( .ZN(net_639), .A(net_566) );
CLKBUF_X2 inst_13291 ( .A(net_13252), .Z(net_13253) );
CLKBUF_X2 inst_13747 ( .A(net_13708), .Z(net_13709) );
CLKBUF_X2 inst_12902 ( .A(net_12863), .Z(net_12864) );
CLKBUF_X2 inst_9613 ( .A(net_9574), .Z(net_9575) );
CLKBUF_X2 inst_12924 ( .A(net_12885), .Z(net_12886) );
CLKBUF_X2 inst_10978 ( .A(net_10939), .Z(net_10940) );
INV_X2 inst_5737 ( .ZN(net_3728), .A(net_3436) );
CLKBUF_X2 inst_13199 ( .A(net_8636), .Z(net_13161) );
INV_X4 inst_5332 ( .A(net_6072), .ZN(net_3623) );
NAND3_X2 inst_2773 ( .ZN(net_2327), .A3(net_1577), .A1(net_1383), .A2(net_954) );
OAI21_X2 inst_2081 ( .B2(net_4415), .ZN(net_4409), .B1(net_4024), .A(net_3502) );
NAND2_X2 inst_3261 ( .ZN(net_4148), .A2(net_3468), .A1(net_1216) );
CLKBUF_X2 inst_8717 ( .A(net_8678), .Z(net_8679) );
CLKBUF_X2 inst_13606 ( .A(net_11633), .Z(net_13568) );
CLKBUF_X2 inst_11144 ( .A(net_9504), .Z(net_11106) );
SDFF_X2 inst_1211 ( .SI(net_7067), .Q(net_7067), .D(net_3883), .SE(net_3747), .CK(net_11835) );
CLKBUF_X2 inst_9078 ( .A(net_9039), .Z(net_9040) );
NAND2_X2 inst_3751 ( .A1(net_7038), .A2(net_1975), .ZN(net_1594) );
SDFF_X2 inst_1192 ( .SI(net_7073), .Q(net_7073), .D(net_3811), .SE(net_3742), .CK(net_8993) );
SDFF_X2 inst_682 ( .Q(net_6746), .D(net_6746), .SE(net_3815), .SI(net_3805), .CK(net_10923) );
SDFF_X2 inst_238 ( .Q(net_6356), .SI(net_6355), .D(net_3523), .SE(net_392), .CK(net_13956) );
CLKBUF_X2 inst_12463 ( .A(net_11352), .Z(net_12425) );
CLKBUF_X2 inst_12394 ( .A(net_10378), .Z(net_12356) );
DFF_X1 inst_6735 ( .QN(net_7354), .D(net_5320), .CK(net_12699) );
DFF_X1 inst_6643 ( .QN(net_7632), .D(net_5223), .CK(net_13427) );
CLKBUF_X2 inst_9123 ( .A(net_9084), .Z(net_9085) );
NOR2_X4 inst_2222 ( .ZN(net_5676), .A1(net_5550), .A2(net_4513) );
INV_X4 inst_4578 ( .ZN(net_5496), .A(net_5495) );
NAND2_X2 inst_3333 ( .ZN(net_3580), .A1(net_3579), .A2(net_3228) );
CLKBUF_X2 inst_10021 ( .A(net_9432), .Z(net_9983) );
CLKBUF_X2 inst_12102 ( .A(net_11193), .Z(net_12064) );
NAND2_X2 inst_4059 ( .A1(net_7205), .A2(net_1648), .ZN(net_993) );
NAND2_X2 inst_3109 ( .A1(net_6617), .A2(net_4899), .ZN(net_4892) );
CLKBUF_X2 inst_10046 ( .A(net_10007), .Z(net_10008) );
OAI21_X2 inst_1755 ( .ZN(net_5447), .B1(net_5446), .A(net_4670), .B2(net_3993) );
NOR2_X4 inst_2240 ( .ZN(net_5646), .A1(net_5492), .A2(net_4461) );
CLKBUF_X2 inst_11680 ( .A(net_11641), .Z(net_11642) );
SDFF_X2 inst_1210 ( .D(net_7799), .SI(net_7066), .Q(net_7066), .SE(net_3742), .CK(net_11920) );
INV_X2 inst_6090 ( .A(net_7660), .ZN(net_1893) );
CLKBUF_X2 inst_12759 ( .A(net_12720), .Z(net_12721) );
NOR2_X2 inst_2437 ( .ZN(net_3425), .A1(net_3046), .A2(net_3045) );
CLKBUF_X2 inst_12715 ( .A(net_12676), .Z(net_12677) );
SDFF_X2 inst_806 ( .Q(net_6979), .D(net_6979), .SE(net_3891), .SI(net_3787), .CK(net_8088) );
INV_X8 inst_4521 ( .ZN(net_3741), .A(net_3116) );
CLKBUF_X2 inst_8324 ( .A(net_8285), .Z(net_8286) );
DFFR_X1 inst_7119 ( .QN(net_5851), .D(net_5685), .CK(net_12352), .RN(x1822) );
OAI21_X2 inst_1981 ( .ZN(net_4850), .B1(net_4849), .A(net_4538), .B2(net_3870) );
DFF_X2 inst_6324 ( .QN(net_7809), .CK(net_8680), .D(x1467) );
SDFF_X2 inst_491 ( .Q(net_6989), .D(net_6989), .SI(net_3902), .SE(net_3891), .CK(net_10874) );
INV_X2 inst_5960 ( .A(net_7357), .ZN(net_2014) );
CLKBUF_X2 inst_10485 ( .A(net_10446), .Z(net_10447) );
INV_X2 inst_6027 ( .A(net_7588), .ZN(net_1977) );
INV_X4 inst_4943 ( .ZN(net_3940), .A(net_745) );
CLKBUF_X2 inst_13219 ( .A(net_9039), .Z(net_13181) );
CLKBUF_X2 inst_13515 ( .A(net_13476), .Z(net_13477) );
CLKBUF_X2 inst_8309 ( .A(net_8270), .Z(net_8271) );
CLKBUF_X2 inst_10987 ( .A(net_10948), .Z(net_10949) );
NAND2_X2 inst_3775 ( .A1(net_6504), .A2(net_1642), .ZN(net_1570) );
CLKBUF_X2 inst_13762 ( .A(net_10457), .Z(net_13724) );
CLKBUF_X2 inst_12097 ( .A(net_9463), .Z(net_12059) );
NOR2_X2 inst_2472 ( .A2(net_5778), .ZN(net_2678), .A1(net_2610) );
CLKBUF_X2 inst_9441 ( .A(net_9402), .Z(net_9403) );
NAND2_X2 inst_3086 ( .A1(net_6483), .A2(net_4927), .ZN(net_4917) );
NAND3_X2 inst_2791 ( .ZN(net_2309), .A3(net_1536), .A1(net_1501), .A2(net_994) );
CLKBUF_X2 inst_12090 ( .A(net_12051), .Z(net_12052) );
CLKBUF_X2 inst_11239 ( .A(net_11200), .Z(net_11201) );
INV_X4 inst_5583 ( .A(net_6411), .ZN(net_429) );
CLKBUF_X2 inst_10243 ( .A(net_10204), .Z(net_10205) );
CLKBUF_X2 inst_8293 ( .A(net_8254), .Z(net_8255) );
SDFF_X2 inst_872 ( .SI(net_7058), .Q(net_7058), .SE(net_3818), .D(net_3801), .CK(net_8206) );
DFF_X1 inst_6641 ( .QN(net_7629), .D(net_5231), .CK(net_13070) );
CLKBUF_X2 inst_11479 ( .A(net_8000), .Z(net_11441) );
CLKBUF_X2 inst_9210 ( .A(net_9171), .Z(net_9172) );
NAND2_X1 inst_4419 ( .ZN(net_2277), .A1(net_1725), .A2(net_915) );
INV_X4 inst_5234 ( .ZN(net_3922), .A(net_801) );
CLKBUF_X2 inst_12579 ( .A(net_9315), .Z(net_12541) );
DFF_X1 inst_6850 ( .D(net_2560), .Q(net_204), .CK(net_9744) );
OAI221_X2 inst_1667 ( .C2(net_5901), .ZN(net_4645), .B1(net_4644), .B2(net_4424), .C1(net_4057), .A(net_3578) );
DFF_X1 inst_6698 ( .QN(net_7296), .D(net_5377), .CK(net_12992) );
SDFFR_X2 inst_1349 ( .D(net_3805), .SE(net_3256), .SI(net_150), .Q(net_150), .CK(net_8549), .RN(x1822) );
SDFF_X2 inst_462 ( .Q(net_6999), .D(net_6999), .SE(net_3899), .SI(net_3892), .CK(net_11971) );
DFFR_X2 inst_7012 ( .D(net_3290), .QN(net_282), .CK(net_12871), .RN(x1822) );
CLKBUF_X2 inst_12744 ( .A(net_12705), .Z(net_12706) );
CLKBUF_X2 inst_10261 ( .A(net_9169), .Z(net_10223) );
NAND2_X2 inst_3745 ( .A1(net_6493), .A2(net_1642), .ZN(net_1600) );
CLKBUF_X2 inst_9398 ( .A(net_9359), .Z(net_9360) );
INV_X4 inst_5572 ( .A(net_6039), .ZN(net_538) );
NAND2_X1 inst_4347 ( .ZN(net_4380), .A2(net_3856), .A1(net_1751) );
CLKBUF_X2 inst_10579 ( .A(net_10540), .Z(net_10541) );
INV_X2 inst_5962 ( .A(net_7348), .ZN(net_2020) );
NOR2_X4 inst_2224 ( .ZN(net_5674), .A1(net_5544), .A2(net_4511) );
CLKBUF_X2 inst_13381 ( .A(net_13342), .Z(net_13343) );
CLKBUF_X2 inst_10002 ( .A(net_8261), .Z(net_9964) );
CLKBUF_X2 inst_10185 ( .A(net_10146), .Z(net_10147) );
DFF_X1 inst_6661 ( .QN(net_7653), .D(net_5179), .CK(net_13142) );
INV_X4 inst_5226 ( .A(net_1223), .ZN(net_463) );
CLKBUF_X2 inst_13012 ( .A(net_12973), .Z(net_12974) );
CLKBUF_X2 inst_10389 ( .A(net_10350), .Z(net_10351) );
INV_X4 inst_4909 ( .A(net_3797), .ZN(net_3128) );
DFFR_X1 inst_7114 ( .QN(net_5856), .D(net_5796), .CK(net_13303), .RN(x1822) );
INV_X4 inst_5310 ( .A(net_6552), .ZN(net_447) );
DFF_X1 inst_6836 ( .Q(net_391), .D(net_388), .CK(net_10543) );
CLKBUF_X2 inst_8412 ( .A(net_8373), .Z(net_8374) );
AOI221_X2 inst_7611 ( .C2(net_3105), .ZN(net_2971), .B1(net_2970), .A(net_2783), .C1(net_766), .B2(net_250) );
OAI21_X2 inst_1914 ( .ZN(net_5151), .B1(net_4866), .A(net_4769), .B2(net_3941) );
DFF_X2 inst_6219 ( .Q(net_6392), .D(net_6391), .CK(net_13846) );
INV_X4 inst_4996 ( .A(net_3003), .ZN(net_866) );
OAI21_X2 inst_1975 ( .B1(net_4872), .ZN(net_4861), .A(net_4366), .B2(net_3853) );
OAI21_X2 inst_1890 ( .B1(net_5230), .ZN(net_5191), .A(net_4567), .B2(net_3866) );
NOR2_X2 inst_2308 ( .A2(net_6206), .A1(net_5840), .ZN(net_5833) );
DFF_X1 inst_6647 ( .QN(net_7621), .D(net_5205), .CK(net_13153) );
NAND2_X2 inst_4093 ( .A1(net_7202), .A2(net_1648), .ZN(net_959) );
CLKBUF_X2 inst_9728 ( .A(net_9501), .Z(net_9690) );
INV_X4 inst_4806 ( .ZN(net_5098), .A(net_1176) );
CLKBUF_X2 inst_9585 ( .A(net_9546), .Z(net_9547) );
NAND2_X4 inst_2879 ( .A1(net_4272), .ZN(net_4260), .A2(net_1705) );
CLKBUF_X2 inst_8117 ( .A(net_8070), .Z(net_8079) );
CLKBUF_X2 inst_12362 ( .A(net_12323), .Z(net_12324) );
AOI222_X2 inst_7482 ( .ZN(net_2137), .A1(net_2136), .A2(net_2135), .B1(net_2134), .B2(net_2133), .C1(net_2132), .C2(net_2131) );
NOR2_X2 inst_2338 ( .A2(net_6280), .A1(net_5840), .ZN(net_5803) );
CLKBUF_X2 inst_11893 ( .A(net_11854), .Z(net_11855) );
NAND2_X2 inst_3475 ( .ZN(net_2857), .A2(net_2708), .A1(net_2629) );
NAND2_X2 inst_3017 ( .A1(net_6858), .A2(net_5004), .ZN(net_4992) );
DFF_X1 inst_6389 ( .QN(net_6120), .D(net_5699), .CK(net_11194) );
CLKBUF_X2 inst_13170 ( .A(net_13131), .Z(net_13132) );
AND2_X4 inst_7818 ( .ZN(net_3262), .A2(net_3166), .A1(net_558) );
CLKBUF_X2 inst_11431 ( .A(net_8180), .Z(net_11393) );
SDFF_X2 inst_845 ( .Q(net_6998), .D(net_6998), .SE(net_3899), .SI(net_3802), .CK(net_9092) );
NAND2_X2 inst_3554 ( .ZN(net_2513), .A2(net_2040), .A1(net_1765) );
OR2_X4 inst_1367 ( .ZN(net_3979), .A2(net_3740), .A1(net_687) );
DFF_X1 inst_6516 ( .QN(net_7447), .D(net_5439), .CK(net_9287) );
CLKBUF_X2 inst_8649 ( .A(net_8610), .Z(net_8611) );
INV_X4 inst_5198 ( .ZN(net_1140), .A(net_502) );
INV_X2 inst_5909 ( .A(net_7360), .ZN(net_2058) );
CLKBUF_X2 inst_10980 ( .A(net_10941), .Z(net_10942) );
CLKBUF_X2 inst_9175 ( .A(net_9136), .Z(net_9137) );
CLKBUF_X2 inst_10898 ( .A(net_9793), .Z(net_10860) );
OAI21_X2 inst_2016 ( .B2(net_4497), .ZN(net_4492), .B1(net_4101), .A(net_3654) );
NAND2_X2 inst_3687 ( .A2(net_1798), .ZN(net_1760), .A1(net_1759) );
CLKBUF_X2 inst_10837 ( .A(net_8127), .Z(net_10799) );
CLKBUF_X2 inst_12723 ( .A(net_12684), .Z(net_12685) );
CLKBUF_X2 inst_8434 ( .A(net_8395), .Z(net_8396) );
NAND2_X2 inst_4012 ( .ZN(net_1265), .A2(net_1228), .A1(net_375) );
CLKBUF_X2 inst_10103 ( .A(net_10064), .Z(net_10065) );
NAND2_X2 inst_3053 ( .A1(net_7121), .ZN(net_4953), .A2(net_4950) );
CLKBUF_X2 inst_8385 ( .A(net_8299), .Z(net_8347) );
CLKBUF_X2 inst_9289 ( .A(net_8643), .Z(net_9251) );
AOI21_X2 inst_7630 ( .ZN(net_4170), .B2(net_4145), .A(net_2847), .B1(net_155) );
CLKBUF_X2 inst_9920 ( .A(net_9595), .Z(net_9882) );
AND2_X4 inst_7829 ( .ZN(net_3016), .A2(net_2818), .A1(net_2261) );
SDFF_X2 inst_393 ( .SI(net_7334), .Q(net_7334), .D(net_4783), .SE(net_3856), .CK(net_12756) );
CLKBUF_X2 inst_10409 ( .A(net_10370), .Z(net_10371) );
INV_X4 inst_4810 ( .ZN(net_4875), .A(net_1168) );
CLKBUF_X2 inst_9962 ( .A(net_8130), .Z(net_9924) );
INV_X2 inst_5969 ( .ZN(net_1131), .A(net_118) );
OAI21_X2 inst_1813 ( .ZN(net_5375), .B1(net_5351), .A(net_4345), .B2(net_3859) );
XNOR2_X2 inst_92 ( .B(net_3001), .ZN(net_1662), .A(net_1153) );
CLKBUF_X2 inst_11168 ( .A(net_11129), .Z(net_11130) );
CLKBUF_X2 inst_10708 ( .A(net_9140), .Z(net_10670) );
SDFF_X2 inst_345 ( .SI(net_7311), .Q(net_7311), .D(net_4876), .SE(net_3859), .CK(net_9410) );
NAND2_X2 inst_3103 ( .A1(net_6614), .ZN(net_4900), .A2(net_4899) );
CLKBUF_X2 inst_9086 ( .A(net_9047), .Z(net_9048) );
CLKBUF_X2 inst_11985 ( .A(net_11946), .Z(net_11947) );
CLKBUF_X2 inst_11856 ( .A(net_8235), .Z(net_11818) );
AOI222_X2 inst_7520 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2010), .A1(net_2009), .B1(net_2008), .C1(net_2007) );
NAND2_X2 inst_3304 ( .ZN(net_3638), .A1(net_3637), .A2(net_3229) );
CLKBUF_X2 inst_10233 ( .A(net_9219), .Z(net_10195) );
AOI21_X2 inst_7762 ( .B1(net_6463), .ZN(net_4437), .B2(net_2580), .A(net_2304) );
CLKBUF_X2 inst_10087 ( .A(net_10048), .Z(net_10049) );
DFF_X1 inst_6362 ( .QN(net_6220), .D(net_5822), .CK(net_14119) );
INV_X4 inst_5384 ( .A(net_6169), .ZN(net_3571) );
CLKBUF_X2 inst_8076 ( .A(net_7830), .Z(net_8038) );
CLKBUF_X2 inst_13806 ( .A(net_8603), .Z(net_13768) );
CLKBUF_X2 inst_11009 ( .A(net_10970), .Z(net_10971) );
CLKBUF_X2 inst_10585 ( .A(net_8336), .Z(net_10547) );
XNOR2_X2 inst_57 ( .ZN(net_1931), .B(net_1699), .A(net_1698) );
INV_X4 inst_4723 ( .A(net_5967), .ZN(net_3049) );
NAND2_X2 inst_3655 ( .A1(net_7060), .ZN(net_1808), .A2(net_791) );
AOI222_X2 inst_7532 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1908), .A1(net_1907), .B1(net_1906), .C1(net_1905) );
CLKBUF_X2 inst_12145 ( .A(net_12106), .Z(net_12107) );
DFF_X1 inst_6692 ( .QN(net_7281), .D(net_5112), .CK(net_12798) );
CLKBUF_X2 inst_9312 ( .A(net_9273), .Z(net_9274) );
DFF_X1 inst_6617 ( .QN(net_7578), .D(net_5390), .CK(net_13446) );
NAND2_X4 inst_2843 ( .ZN(net_5535), .A1(net_5012), .A2(net_5011) );
OAI21_X2 inst_1888 ( .B1(net_5235), .ZN(net_5193), .A(net_4569), .B2(net_3866) );
NAND2_X2 inst_3379 ( .ZN(net_3488), .A1(net_3487), .A2(net_3223) );
OAI21_X2 inst_1763 ( .B1(net_5554), .ZN(net_5431), .A(net_4649), .B2(net_3993) );
SDFF_X2 inst_1307 ( .D(net_6386), .SE(net_5800), .SI(net_351), .Q(net_351), .CK(net_13658) );
CLKBUF_X2 inst_13071 ( .A(net_13032), .Z(net_13033) );
AOI21_X2 inst_7759 ( .B1(net_6457), .ZN(net_4424), .B2(net_2580), .A(net_2308) );
CLKBUF_X2 inst_10878 ( .A(net_10839), .Z(net_10840) );
CLKBUF_X2 inst_8565 ( .A(net_8494), .Z(net_8527) );
DFF_X1 inst_6789 ( .D(net_3932), .CK(net_12843), .Q(x657) );
CLKBUF_X2 inst_13685 ( .A(net_11561), .Z(net_13647) );
CLKBUF_X2 inst_14309 ( .A(net_14270), .Z(net_14271) );
SDFF_X2 inst_1094 ( .SI(net_6944), .Q(net_6944), .D(net_3784), .SE(net_3741), .CK(net_11702) );
CLKBUF_X2 inst_12960 ( .A(net_12921), .Z(net_12922) );
NAND2_X2 inst_4145 ( .A1(net_1152), .ZN(net_910), .A2(net_879) );
INV_X4 inst_4590 ( .ZN(net_4308), .A(net_4213) );
DFFR_X1 inst_7124 ( .Q(net_5992), .D(net_4800), .CK(net_10381), .RN(x1822) );
DFF_X1 inst_6376 ( .QN(net_6286), .D(net_5808), .CK(net_14259) );
NAND2_X2 inst_3680 ( .A2(net_1798), .ZN(net_1773), .A1(net_1772) );
INV_X4 inst_4878 ( .ZN(net_2853), .A(net_903) );
OAI21_X2 inst_1699 ( .ZN(net_5595), .A(net_5269), .B2(net_4617), .B1(net_4228) );
CLKBUF_X2 inst_8616 ( .A(net_8577), .Z(net_8578) );
SDFF_X2 inst_851 ( .Q(net_7004), .D(net_7004), .SE(net_3899), .SI(net_3814), .CK(net_9029) );
CLKBUF_X2 inst_12685 ( .A(net_12646), .Z(net_12647) );
SDFF_X2 inst_831 ( .SI(net_7807), .Q(net_7010), .D(net_7010), .SE(net_3899), .CK(net_10865) );
XNOR2_X2 inst_50 ( .ZN(net_2255), .A(net_1917), .B(net_895) );
CLKBUF_X2 inst_11762 ( .A(net_8653), .Z(net_11724) );
INV_X2 inst_5824 ( .ZN(net_932), .A(net_931) );
NAND2_X1 inst_4264 ( .ZN(net_4656), .A2(net_3993), .A1(net_1431) );
NAND3_X2 inst_2589 ( .ZN(net_5750), .A1(net_5645), .A2(net_5245), .A3(net_4209) );
CLKBUF_X2 inst_10626 ( .A(net_10587), .Z(net_10588) );
CLKBUF_X2 inst_11448 ( .A(net_10754), .Z(net_11410) );
NAND2_X1 inst_4430 ( .A1(net_7614), .A2(net_2131), .ZN(net_1439) );
CLKBUF_X2 inst_8699 ( .A(net_8660), .Z(net_8661) );
OAI221_X2 inst_1650 ( .ZN(net_5053), .C2(net_5052), .B2(net_5049), .A(net_4524), .B1(net_2427), .C1(net_1056) );
CLKBUF_X2 inst_11174 ( .A(net_11135), .Z(net_11136) );
OAI22_X2 inst_1497 ( .B1(net_4660), .ZN(net_4106), .A1(net_4105), .A2(net_4104), .B2(net_4103) );
CLKBUF_X2 inst_8250 ( .A(net_7895), .Z(net_8212) );
AOI222_X2 inst_7469 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2175), .A1(net_2174), .B1(net_2173), .C1(net_2172) );
NAND2_X1 inst_4439 ( .A2(net_2131), .ZN(net_1353), .A1(net_1352) );
INV_X2 inst_5706 ( .ZN(net_4312), .A(net_4221) );
NAND2_X4 inst_2872 ( .A1(net_4280), .ZN(net_4267), .A2(net_1521) );
CLKBUF_X2 inst_8683 ( .A(net_8644), .Z(net_8645) );
SDFF_X2 inst_1002 ( .Q(net_6461), .D(net_6461), .SE(net_3904), .SI(net_3798), .CK(net_11654) );
CLKBUF_X2 inst_12076 ( .A(net_9573), .Z(net_12038) );
CLKBUF_X2 inst_8057 ( .A(net_8018), .Z(net_8019) );
CLKBUF_X2 inst_13179 ( .A(net_11420), .Z(net_13141) );
SDFF_X2 inst_478 ( .Q(net_6832), .D(net_6832), .SE(net_3893), .SI(net_3892), .CK(net_8976) );
CLKBUF_X2 inst_8630 ( .A(net_8163), .Z(net_8592) );
NAND2_X2 inst_3380 ( .ZN(net_3486), .A1(net_3485), .A2(net_3223) );
INV_X4 inst_5666 ( .A(net_6414), .ZN(net_1700) );
SDFF_X2 inst_804 ( .Q(net_6977), .D(net_6977), .SE(net_3891), .SI(net_3811), .CK(net_11911) );
NAND2_X2 inst_3290 ( .ZN(net_3666), .A1(net_3665), .A2(net_3229) );
CLKBUF_X2 inst_13953 ( .A(net_12636), .Z(net_13915) );
CLKBUF_X2 inst_8824 ( .A(net_8750), .Z(net_8786) );
XNOR2_X2 inst_13 ( .ZN(net_2643), .B(net_2642), .A(net_2483) );
CLKBUF_X2 inst_12173 ( .A(net_12134), .Z(net_12135) );
CLKBUF_X2 inst_14126 ( .A(net_14087), .Z(net_14088) );
INV_X4 inst_5378 ( .A(net_6146), .ZN(net_3591) );
NAND3_X2 inst_2584 ( .ZN(net_5755), .A1(net_5650), .A2(net_5272), .A3(net_4310) );
INV_X4 inst_5665 ( .A(net_6176), .ZN(net_3566) );
INV_X4 inst_4931 ( .ZN(net_767), .A(net_766) );
CLKBUF_X2 inst_11540 ( .A(net_8642), .Z(net_11502) );
AOI22_X2 inst_7334 ( .B2(net_3439), .ZN(net_3308), .A2(net_2712), .B1(net_763), .A1(net_150) );
SDFF_X2 inst_799 ( .SI(net_6901), .Q(net_6901), .D(net_3814), .SE(net_3781), .CK(net_11789) );
CLKBUF_X2 inst_12906 ( .A(net_12867), .Z(net_12868) );
NAND2_X2 inst_3481 ( .ZN(net_2677), .A1(net_2676), .A2(net_2675) );
SDFF_X2 inst_738 ( .Q(net_6856), .D(net_6856), .SE(net_3893), .SI(net_3789), .CK(net_11502) );
CLKBUF_X2 inst_13666 ( .A(net_8183), .Z(net_13628) );
DFF_X1 inst_6481 ( .QN(net_7412), .D(net_5571), .CK(net_10101) );
NAND3_X2 inst_2755 ( .ZN(net_2346), .A3(net_1613), .A1(net_1443), .A2(net_1010) );
CLKBUF_X2 inst_9393 ( .A(net_9354), .Z(net_9355) );
CLKBUF_X2 inst_9101 ( .A(net_9062), .Z(net_9063) );
OAI21_X2 inst_1819 ( .ZN(net_5369), .B1(net_5339), .A(net_4336), .B2(net_3859) );
CLKBUF_X2 inst_14284 ( .A(net_14245), .Z(net_14246) );
SDFF_X2 inst_255 ( .Q(net_6379), .SI(net_6378), .D(net_3532), .SE(net_392), .CK(net_13513) );
NAND3_X2 inst_2726 ( .ZN(net_2375), .A3(net_1634), .A1(net_1498), .A2(net_1009) );
SDFF_X2 inst_453 ( .Q(net_6060), .SI(net_3921), .SE(net_3318), .D(net_3317), .CK(net_10326) );
SDFF_X2 inst_493 ( .Q(net_6847), .D(net_6847), .SI(net_3897), .SE(net_3893), .CK(net_8897) );
CLKBUF_X2 inst_10555 ( .A(net_8553), .Z(net_10517) );
NAND3_X2 inst_2674 ( .ZN(net_3749), .A3(net_3308), .A1(net_2971), .A2(net_2944) );
XNOR2_X2 inst_23 ( .ZN(net_2576), .B(net_2575), .A(net_2449) );
CLKBUF_X2 inst_10390 ( .A(net_10351), .Z(net_10352) );
CLKBUF_X2 inst_10279 ( .A(net_8609), .Z(net_10241) );
DFF_X1 inst_6686 ( .QN(net_7274), .D(net_5118), .CK(net_9456) );
CLKBUF_X2 inst_8784 ( .A(net_8341), .Z(net_8746) );
SDFF_X2 inst_1113 ( .SI(net_6671), .Q(net_6671), .D(net_3785), .SE(net_3465), .CK(net_7845) );
OAI21_X2 inst_1822 ( .ZN(net_5366), .B1(net_5365), .A(net_4385), .B2(net_3856) );
NAND2_X2 inst_3790 ( .A1(net_6772), .A2(net_1635), .ZN(net_1555) );
CLKBUF_X2 inst_12438 ( .A(net_10376), .Z(net_12400) );
NAND2_X2 inst_4206 ( .A2(net_6020), .A1(net_6019), .ZN(net_3238) );
CLKBUF_X2 inst_12551 ( .A(net_11369), .Z(net_12513) );
INV_X4 inst_5415 ( .A(net_6181), .ZN(net_3707) );
DFF_X1 inst_6701 ( .QN(net_7299), .D(net_5374), .CK(net_9881) );
CLKBUF_X2 inst_10340 ( .A(net_10301), .Z(net_10302) );
CLKBUF_X2 inst_10347 ( .A(net_10308), .Z(net_10309) );
SDFF_X2 inst_812 ( .Q(net_6986), .D(net_6986), .SE(net_3891), .SI(net_3804), .CK(net_11027) );
SDFF_X2 inst_179 ( .Q(net_6275), .SI(net_6274), .D(net_3505), .SE(net_392), .CK(net_13481) );
INV_X4 inst_5698 ( .ZN(net_5927), .A(net_5925) );
OAI21_X2 inst_1730 ( .ZN(net_5564), .B1(net_5399), .A(net_4829), .B2(net_4153) );
NAND2_X2 inst_3799 ( .A1(net_7174), .A2(net_1637), .ZN(net_1546) );
CLKBUF_X2 inst_8101 ( .A(net_8062), .Z(net_8063) );
NAND2_X2 inst_3734 ( .A1(net_7182), .A2(net_1637), .ZN(net_1611) );
NOR3_X2 inst_2191 ( .ZN(net_5954), .A2(net_3951), .A3(net_3879), .A1(net_3759) );
XNOR2_X2 inst_76 ( .ZN(net_1936), .B(net_668), .A(net_611) );
INV_X4 inst_5296 ( .A(net_5861), .ZN(net_549) );
SDFF_X2 inst_1127 ( .SI(net_6677), .Q(net_6677), .D(net_3775), .SE(net_3471), .CK(net_9076) );
DFF_X1 inst_6769 ( .QN(net_6167), .D(net_4651), .CK(net_7949) );
SDFF_X2 inst_172 ( .Q(net_6242), .SI(net_6241), .D(net_3534), .SE(net_392), .CK(net_13527) );
CLKBUF_X2 inst_12184 ( .A(net_7862), .Z(net_12146) );
CLKBUF_X2 inst_11228 ( .A(net_11189), .Z(net_11190) );
SDFF_X2 inst_362 ( .SI(net_7611), .Q(net_7611), .D(net_4787), .SE(net_3870), .CK(net_8312) );
NAND2_X1 inst_4366 ( .ZN(net_4361), .A2(net_3853), .A1(net_1996) );
SDFF_X2 inst_277 ( .D(net_6398), .SE(net_5800), .SI(net_363), .Q(net_363), .CK(net_13680) );
AOI21_X2 inst_7787 ( .ZN(net_2233), .A(net_2232), .B1(net_1154), .B2(net_1069) );
XNOR2_X2 inst_83 ( .B(net_2241), .ZN(net_1309), .A(net_1308) );
SDFF_X2 inst_306 ( .SI(net_7523), .Q(net_7523), .D(net_5102), .SE(net_3988), .CK(net_9797) );
NAND2_X2 inst_4186 ( .A2(net_5999), .ZN(net_1741), .A1(net_541) );
INV_X4 inst_5566 ( .A(net_7745), .ZN(net_2670) );
CLKBUF_X2 inst_8662 ( .A(net_8623), .Z(net_8624) );
CLKBUF_X2 inst_13499 ( .A(net_13460), .Z(net_13461) );
CLKBUF_X2 inst_9460 ( .A(net_9421), .Z(net_9422) );
CLKBUF_X2 inst_7946 ( .A(net_7907), .Z(net_7908) );
NAND2_X2 inst_3386 ( .ZN(net_3474), .A1(net_3473), .A2(net_3231) );
NAND2_X2 inst_3095 ( .A1(net_6455), .A2(net_4925), .ZN(net_4908) );
CLKBUF_X2 inst_9884 ( .A(net_9845), .Z(net_9846) );
OAI21_X2 inst_1715 ( .ZN(net_5579), .B1(net_5551), .A(net_4689), .B2(net_3989) );
CLKBUF_X2 inst_13673 ( .A(net_13634), .Z(net_13635) );
DFF_X1 inst_6396 ( .QN(net_6135), .D(net_5692), .CK(net_11767) );
AOI22_X2 inst_7355 ( .B2(net_3105), .ZN(net_3095), .A2(net_2712), .A1(net_1125), .B1(net_440) );
SDFF_X2 inst_140 ( .Q(net_6238), .SI(net_6237), .SE(net_392), .D(net_144), .CK(net_13625) );
SDFF_X2 inst_267 ( .D(net_6400), .SE(net_5801), .SI(net_345), .Q(net_345), .CK(net_14341) );
CLKBUF_X2 inst_7990 ( .A(net_7951), .Z(net_7952) );
NAND3_X2 inst_2824 ( .A1(net_6415), .ZN(net_1929), .A2(net_1700), .A3(net_692) );
INV_X2 inst_5945 ( .A(net_7451), .ZN(net_1431) );
SDFF_X2 inst_716 ( .SI(net_6788), .Q(net_6788), .SE(net_3872), .D(net_3801), .CK(net_8358) );
NAND2_X2 inst_3594 ( .ZN(net_2406), .A2(net_1880), .A1(net_1454) );
OAI21_X2 inst_1906 ( .B1(net_5357), .ZN(net_5163), .A(net_4763), .B2(net_3941) );
SDFF_X2 inst_792 ( .SI(net_6922), .Q(net_6922), .D(net_3821), .SE(net_3781), .CK(net_11713) );
CLKBUF_X2 inst_8155 ( .A(net_8116), .Z(net_8117) );
OAI21_X2 inst_2024 ( .B1(net_5906), .B2(net_4497), .ZN(net_4482), .A(net_3630) );
NAND2_X2 inst_3124 ( .A1(net_6580), .A2(net_4897), .ZN(net_4877) );
CLKBUF_X2 inst_9984 ( .A(net_9945), .Z(net_9946) );
CLKBUF_X2 inst_7993 ( .A(net_7954), .Z(net_7955) );
NAND2_X2 inst_2952 ( .ZN(net_5488), .A1(net_4945), .A2(net_4944) );
CLKBUF_X2 inst_11896 ( .A(net_11857), .Z(net_11858) );
CLKBUF_X2 inst_9061 ( .A(net_9022), .Z(net_9023) );
CLKBUF_X2 inst_10476 ( .A(net_10437), .Z(net_10438) );
CLKBUF_X2 inst_8933 ( .A(net_8499), .Z(net_8895) );
NOR2_X4 inst_2216 ( .ZN(net_5682), .A1(net_5563), .A2(net_4522) );
CLKBUF_X2 inst_11558 ( .A(net_11519), .Z(net_11520) );
SDFF_X2 inst_174 ( .SI(net_6279), .Q(net_6240), .D(net_3585), .SE(net_392), .CK(net_13968) );
NAND2_X2 inst_2988 ( .A1(net_6721), .A2(net_5031), .ZN(net_5023) );
CLKBUF_X2 inst_8658 ( .A(net_8449), .Z(net_8620) );
INV_X8 inst_4494 ( .ZN(net_3830), .A(net_3153) );
CLKBUF_X2 inst_12293 ( .A(net_11687), .Z(net_12255) );
CLKBUF_X2 inst_8942 ( .A(net_8903), .Z(net_8904) );
CLKBUF_X2 inst_11186 ( .A(net_11147), .Z(net_11148) );
OAI21_X2 inst_2105 ( .ZN(net_3974), .A(net_3973), .B2(net_3875), .B1(net_1059) );
SDFF_X2 inst_1199 ( .SI(net_7081), .Q(net_7081), .D(net_3836), .SE(net_3747), .CK(net_8987) );
XOR2_X2 inst_5 ( .A(net_2571), .Z(net_1244), .B(net_1243) );
SDFF_X2 inst_729 ( .Q(net_6845), .D(net_6845), .SE(net_3893), .SI(net_3809), .CK(net_8504) );
DFF_X1 inst_6567 ( .QN(net_7503), .D(net_5106), .CK(net_9255) );
CLKBUF_X2 inst_11520 ( .A(net_10896), .Z(net_11482) );
DFF_X1 inst_6506 ( .QN(net_7428), .D(net_5519), .CK(net_9680) );
OAI21_X2 inst_2157 ( .ZN(net_2491), .A(net_2225), .B2(net_1916), .B1(net_1667) );
OAI221_X2 inst_1662 ( .C2(net_5896), .ZN(net_4663), .B1(net_4660), .B2(net_4487), .C1(net_4105), .A(net_3642) );
CLKBUF_X2 inst_10891 ( .A(net_10852), .Z(net_10853) );
INV_X8 inst_4553 ( .ZN(net_1910), .A(net_812) );
NAND3_X2 inst_2783 ( .ZN(net_2317), .A3(net_1618), .A1(net_1341), .A2(net_1011) );
AOI222_X2 inst_7508 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2040), .A1(net_2039), .B1(net_2038), .C1(net_2037) );
INV_X2 inst_5804 ( .ZN(net_1713), .A(net_191) );
SDFF_X2 inst_604 ( .Q(net_6608), .D(net_6608), .SE(net_3830), .SI(net_3808), .CK(net_12170) );
CLKBUF_X2 inst_9004 ( .A(net_7908), .Z(net_8966) );
CLKBUF_X2 inst_13240 ( .A(net_10391), .Z(net_13202) );
CLKBUF_X2 inst_11251 ( .A(net_11212), .Z(net_11213) );
CLKBUF_X2 inst_13872 ( .A(net_13833), .Z(net_13834) );
AOI222_X2 inst_7539 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1886), .A1(net_1885), .B1(net_1884), .C1(net_1883) );
DFFR_X2 inst_7085 ( .QN(net_7730), .D(net_2803), .CK(net_10431), .RN(x1822) );
SDFF_X2 inst_1285 ( .D(net_3802), .SE(net_3256), .SI(net_132), .Q(net_132), .CK(net_8477) );
SDFF_X2 inst_380 ( .SI(net_7675), .Q(net_7675), .D(net_4787), .SE(net_3866), .CK(net_8309) );
NAND2_X2 inst_4057 ( .A1(net_6674), .A2(net_1655), .ZN(net_995) );
SDFF_X2 inst_1179 ( .SI(net_6952), .Q(net_6952), .D(net_3789), .SE(net_3741), .CK(net_8119) );
SDFF_X2 inst_292 ( .D(net_6395), .SE(net_5800), .SI(net_360), .Q(net_360), .CK(net_14156) );
NAND2_X2 inst_3650 ( .A1(net_7072), .ZN(net_1813), .A2(net_791) );
CLKBUF_X2 inst_11661 ( .A(net_11622), .Z(net_11623) );
CLKBUF_X2 inst_13508 ( .A(net_13469), .Z(net_13470) );
OAI21_X2 inst_2012 ( .B2(net_4497), .ZN(net_4496), .B1(net_4109), .A(net_3662) );
CLKBUF_X2 inst_11350 ( .A(net_11311), .Z(net_11312) );
CLKBUF_X2 inst_10900 ( .A(net_10861), .Z(net_10862) );
AOI22_X2 inst_7423 ( .A1(net_2970), .B1(net_2772), .ZN(net_2769), .A2(net_230), .B2(net_156) );
INV_X4 inst_4970 ( .ZN(net_697), .A(net_696) );
CLKBUF_X2 inst_12583 ( .A(net_8504), .Z(net_12545) );
SDFF_X2 inst_706 ( .SI(net_6759), .Q(net_6759), .SE(net_3872), .D(net_3806), .CK(net_8274) );
CLKBUF_X2 inst_10874 ( .A(net_9929), .Z(net_10836) );
DFF_X1 inst_6605 ( .QN(net_7512), .D(net_5403), .CK(net_12474) );
CLKBUF_X2 inst_9834 ( .A(net_9795), .Z(net_9796) );
SDFF_X2 inst_839 ( .Q(net_7019), .D(net_7019), .SE(net_3899), .SI(net_3803), .CK(net_8080) );
CLKBUF_X2 inst_13366 ( .A(net_13327), .Z(net_13328) );
CLKBUF_X2 inst_7985 ( .A(net_7946), .Z(net_7947) );
INV_X4 inst_4734 ( .A(net_5982), .ZN(net_3873) );
SDFF_X2 inst_240 ( .Q(net_6354), .SI(net_6353), .D(net_3603), .SE(net_392), .CK(net_13949) );
CLKBUF_X2 inst_13055 ( .A(net_11825), .Z(net_13017) );
INV_X4 inst_5455 ( .A(net_7531), .ZN(net_1204) );
AOI222_X2 inst_7501 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2068), .A1(net_2067), .B1(net_2066), .C1(net_2065) );
NAND2_X2 inst_3966 ( .A1(net_6562), .A2(net_1705), .ZN(net_1314) );
XNOR2_X2 inst_110 ( .A(net_2571), .ZN(net_832), .B(net_831) );
CLKBUF_X2 inst_13681 ( .A(net_8565), .Z(net_13643) );
OAI21_X2 inst_2047 ( .B2(net_4457), .ZN(net_4453), .B1(net_4079), .A(net_3706) );
INV_X8 inst_4545 ( .ZN(net_1798), .A(net_1107) );
NAND2_X2 inst_3825 ( .A1(net_7456), .A2(net_1696), .ZN(net_1519) );
DFF_X1 inst_6634 ( .QN(net_7590), .D(net_5248), .CK(net_10573) );
XNOR2_X2 inst_99 ( .ZN(net_2242), .A(net_1151), .B(net_1145) );
CLKBUF_X2 inst_9997 ( .A(net_9958), .Z(net_9959) );
CLKBUF_X2 inst_13210 ( .A(net_8690), .Z(net_13172) );
CLKBUF_X2 inst_7876 ( .A(net_7837), .Z(net_7838) );
CLKBUF_X2 inst_13152 ( .A(net_13113), .Z(net_13114) );
CLKBUF_X2 inst_10842 ( .A(net_10803), .Z(net_10804) );
CLKBUF_X2 inst_11927 ( .A(net_11888), .Z(net_11889) );
CLKBUF_X2 inst_11050 ( .A(net_11011), .Z(net_11012) );
NAND2_X1 inst_4384 ( .ZN(net_4343), .A2(net_3859), .A1(net_2045) );
AND2_X4 inst_7846 ( .ZN(net_1962), .A2(net_707), .A1(net_620) );
OAI21_X2 inst_2059 ( .ZN(net_4438), .B1(net_4437), .B2(net_4436), .A(net_3559) );
CLKBUF_X2 inst_13851 ( .A(net_13812), .Z(net_13813) );
DFFR_X2 inst_7023 ( .D(net_3294), .QN(net_273), .CK(net_12335), .RN(x1822) );
CLKBUF_X2 inst_9473 ( .A(net_9434), .Z(net_9435) );
CLKBUF_X2 inst_9445 ( .A(net_9406), .Z(net_9407) );
NAND2_X2 inst_2949 ( .ZN(net_5491), .A1(net_4952), .A2(net_4951) );
NOR2_X2 inst_2414 ( .A1(net_5986), .ZN(net_3409), .A2(net_3401) );
CLKBUF_X2 inst_9656 ( .A(net_9617), .Z(net_9618) );
SDFF_X2 inst_311 ( .SI(net_7453), .Q(net_7453), .D(net_5098), .SE(net_3993), .CK(net_9792) );
CLKBUF_X2 inst_12461 ( .A(net_11141), .Z(net_12423) );
CLKBUF_X2 inst_9914 ( .A(net_9875), .Z(net_9876) );
CLKBUF_X2 inst_13205 ( .A(net_13166), .Z(net_13167) );
CLKBUF_X2 inst_10429 ( .A(net_8441), .Z(net_10391) );
CLKBUF_X2 inst_13180 ( .A(net_13141), .Z(net_13142) );
CLKBUF_X2 inst_8139 ( .A(net_8100), .Z(net_8101) );
NOR3_X2 inst_2203 ( .ZN(net_3149), .A1(net_2987), .A3(net_1745), .A2(net_1105) );
CLKBUF_X2 inst_11132 ( .A(net_10530), .Z(net_11094) );
CLKBUF_X2 inst_7901 ( .A(net_7862), .Z(net_7863) );
CLKBUF_X2 inst_10495 ( .A(net_10456), .Z(net_10457) );
DFFR_X2 inst_6981 ( .D(net_3438), .QN(net_299), .CK(net_10829), .RN(x1822) );
CLKBUF_X2 inst_14413 ( .A(net_14374), .Z(net_14375) );
CLKBUF_X2 inst_11695 ( .A(net_11656), .Z(net_11657) );
AOI22_X2 inst_7316 ( .ZN(net_4595), .B2(net_3980), .A2(net_3453), .A1(net_1738), .B1(net_1047) );
OAI21_X2 inst_1930 ( .ZN(net_5115), .A(net_4770), .B2(net_3941), .B1(net_1169) );
CLKBUF_X2 inst_14440 ( .A(net_14401), .Z(net_14402) );
SDFF_X2 inst_889 ( .Q(net_7119), .D(net_7119), .SE(net_3888), .SI(net_3805), .CK(net_8785) );
SDFF_X2 inst_577 ( .Q(net_6574), .D(net_6574), .SE(net_3823), .SI(net_3810), .CK(net_12191) );
INV_X4 inst_5536 ( .A(net_6060), .ZN(net_800) );
CLKBUF_X2 inst_12305 ( .A(net_12266), .Z(net_12267) );
CLKBUF_X2 inst_8935 ( .A(net_8896), .Z(net_8897) );
CLKBUF_X2 inst_13497 ( .A(net_8147), .Z(net_13459) );
CLKBUF_X2 inst_8533 ( .A(net_8253), .Z(net_8495) );
INV_X4 inst_4975 ( .A(net_2891), .ZN(net_809) );
DFF_X1 inst_6760 ( .QN(net_7315), .D(net_4863), .CK(net_12795) );
CLKBUF_X2 inst_12457 ( .A(net_11309), .Z(net_12419) );
INV_X4 inst_5188 ( .A(net_896), .ZN(net_515) );
NOR2_X2 inst_2379 ( .ZN(net_5128), .A2(net_4606), .A1(net_4404) );
NAND2_X2 inst_3938 ( .A1(net_6976), .A2(net_1833), .ZN(net_1355) );
CLKBUF_X2 inst_10358 ( .A(net_7830), .Z(net_10320) );
CLKBUF_X2 inst_8774 ( .A(net_8246), .Z(net_8736) );
CLKBUF_X2 inst_11754 ( .A(net_11715), .Z(net_11716) );
CLKBUF_X2 inst_11244 ( .A(net_11205), .Z(net_11206) );
NAND2_X4 inst_2865 ( .ZN(net_4286), .A1(net_4276), .A2(net_1648) );
CLKBUF_X2 inst_10382 ( .A(net_10343), .Z(net_10344) );
INV_X2 inst_5986 ( .A(net_7299), .ZN(net_2049) );
INV_X4 inst_4916 ( .A(net_3821), .ZN(net_827) );
CLKBUF_X2 inst_8149 ( .A(net_8110), .Z(net_8111) );
INV_X4 inst_4891 ( .ZN(net_1181), .A(net_875) );
NAND2_X2 inst_3571 ( .ZN(net_2496), .A2(net_2213), .A1(net_1762) );
INV_X16 inst_6132 ( .ZN(net_3405), .A(net_3360) );
SDFF_X2 inst_1190 ( .SI(net_7070), .Q(net_7070), .D(net_3894), .SE(net_3742), .CK(net_8189) );
SDFF_X2 inst_444 ( .Q(net_7395), .D(net_7395), .SE(net_3994), .SI(net_360), .CK(net_9623) );
CLKBUF_X2 inst_8865 ( .A(net_8826), .Z(net_8827) );
AOI222_X2 inst_7460 ( .ZN(net_2217), .A1(net_2216), .B1(net_2215), .C1(net_2214), .A2(net_2211), .B2(net_2209), .C2(net_2207) );
CLKBUF_X2 inst_11092 ( .A(net_11053), .Z(net_11054) );
CLKBUF_X2 inst_11016 ( .A(net_10540), .Z(net_10978) );
AOI222_X2 inst_7489 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2108), .A1(net_2107), .B1(net_2106), .C1(net_2105) );
CLKBUF_X2 inst_8246 ( .A(net_8207), .Z(net_8208) );
DFF_X2 inst_6264 ( .QN(net_5966), .D(net_2643), .CK(net_12533) );
CLKBUF_X2 inst_12816 ( .A(net_12777), .Z(net_12778) );
CLKBUF_X2 inst_9064 ( .A(net_8169), .Z(net_9026) );
CLKBUF_X2 inst_10033 ( .A(net_9994), .Z(net_9995) );
CLKBUF_X2 inst_14196 ( .A(net_14157), .Z(net_14158) );
CLKBUF_X2 inst_8705 ( .A(net_8666), .Z(net_8667) );
CLKBUF_X2 inst_11720 ( .A(net_11681), .Z(net_11682) );
DFFR_X2 inst_7040 ( .QN(net_6000), .D(net_3138), .CK(net_10017), .RN(x1822) );
INV_X4 inst_4905 ( .A(net_3854), .ZN(net_3046) );
XNOR2_X2 inst_63 ( .ZN(net_1729), .B(net_1728), .A(net_1090) );
INV_X2 inst_5833 ( .A(net_1334), .ZN(net_901) );
CLKBUF_X2 inst_12047 ( .A(net_8226), .Z(net_12009) );
XNOR2_X2 inst_119 ( .ZN(net_5865), .B(net_1654), .A(net_829) );
NAND2_X2 inst_3181 ( .ZN(net_4752), .A2(net_3941), .A1(net_2027) );
SDFF_X2 inst_939 ( .SI(net_7182), .Q(net_7182), .SE(net_3819), .D(net_3784), .CK(net_13339) );
CLKBUF_X2 inst_7968 ( .A(net_7923), .Z(net_7930) );
CLKBUF_X2 inst_9722 ( .A(net_8083), .Z(net_9684) );
CLKBUF_X2 inst_10770 ( .A(net_10731), .Z(net_10732) );
INV_X4 inst_5469 ( .A(net_6134), .ZN(net_3665) );
SDFF_X2 inst_1233 ( .SI(net_7200), .Q(net_7200), .D(net_3798), .SE(net_3750), .CK(net_13308) );
CLKBUF_X2 inst_10445 ( .A(net_10406), .Z(net_10407) );
CLKBUF_X2 inst_8205 ( .A(net_8166), .Z(net_8167) );
NAND2_X2 inst_2924 ( .ZN(net_5533), .A1(net_5009), .A2(net_5008) );
CLKBUF_X2 inst_11117 ( .A(net_11078), .Z(net_11079) );
SDFF_X2 inst_1019 ( .SI(net_6515), .Q(net_6515), .SE(net_3886), .D(net_3789), .CK(net_11244) );
CLKBUF_X2 inst_13490 ( .A(net_11978), .Z(net_13452) );
OAI21_X2 inst_2006 ( .B1(net_5894), .B2(net_4518), .ZN(net_4505), .A(net_3676) );
CLKBUF_X2 inst_10337 ( .A(net_7850), .Z(net_10299) );
OAI21_X2 inst_1827 ( .ZN(net_5356), .B1(net_5355), .A(net_4379), .B2(net_3856) );
CLKBUF_X2 inst_10830 ( .A(net_10791), .Z(net_10792) );
SDFF_X2 inst_742 ( .Q(net_6859), .D(net_6859), .SE(net_3893), .SI(net_3801), .CK(net_11495) );
CLKBUF_X2 inst_13372 ( .A(net_11339), .Z(net_13334) );
NAND3_X2 inst_2619 ( .ZN(net_5720), .A1(net_5615), .A2(net_5132), .A3(net_4179) );
DFFR_X2 inst_7057 ( .QN(net_5991), .D(net_3112), .CK(net_12856), .RN(x1822) );
NAND2_X2 inst_3465 ( .A2(net_3439), .ZN(net_2856), .A1(net_2855) );
OAI21_X2 inst_2033 ( .B2(net_4476), .ZN(net_4470), .B1(net_4222), .A(net_3600) );
CLKBUF_X2 inst_14131 ( .A(net_14092), .Z(net_14093) );
AND2_X4 inst_7850 ( .A2(net_6406), .A1(net_6405), .ZN(net_825) );
INV_X8 inst_4481 ( .ZN(net_4276), .A(net_3927) );
AOI21_X2 inst_7675 ( .B1(net_7011), .ZN(net_4223), .A(net_2455), .B2(net_1100) );
NAND4_X2 inst_2559 ( .A1(net_6422), .A3(net_2453), .ZN(net_2263), .A2(net_897), .A4(net_503) );
CLKBUF_X2 inst_13898 ( .A(net_13859), .Z(net_13860) );
CLKBUF_X2 inst_13545 ( .A(net_13506), .Z(net_13507) );
CLKBUF_X2 inst_13336 ( .A(net_13297), .Z(net_13298) );
AOI22_X2 inst_7345 ( .ZN(net_3107), .B1(net_3106), .B2(net_3105), .A2(net_2712), .A1(net_1135) );
CLKBUF_X2 inst_12039 ( .A(net_12000), .Z(net_12001) );
INV_X4 inst_5289 ( .A(net_6827), .ZN(net_558) );
CLKBUF_X2 inst_10201 ( .A(net_7827), .Z(net_10163) );
CLKBUF_X2 inst_9121 ( .A(net_8466), .Z(net_9083) );
CLKBUF_X2 inst_8386 ( .A(net_8347), .Z(net_8348) );
DFFR_X2 inst_6997 ( .QN(net_7707), .D(net_3355), .CK(net_10751), .RN(x1822) );
OAI21_X2 inst_1955 ( .B1(net_5208), .ZN(net_5065), .A(net_4710), .B2(net_3986) );
CLKBUF_X2 inst_8837 ( .A(net_8798), .Z(net_8799) );
INV_X16 inst_6125 ( .ZN(net_4897), .A(net_4260) );
CLKBUF_X2 inst_12657 ( .A(net_12618), .Z(net_12619) );
NAND2_X2 inst_3618 ( .ZN(net_1972), .A2(net_1971), .A1(net_1715) );
SDFF_X2 inst_1269 ( .Q(net_6961), .D(net_3429), .SI(net_3428), .SE(net_2259), .CK(net_8539) );
CLKBUF_X2 inst_13575 ( .A(net_13333), .Z(net_13537) );
CLKBUF_X2 inst_14430 ( .A(net_14391), .Z(net_14392) );
CLKBUF_X2 inst_9181 ( .A(net_7835), .Z(net_9143) );
CLKBUF_X2 inst_9781 ( .A(net_9742), .Z(net_9743) );
NAND2_X2 inst_3241 ( .ZN(net_4159), .A2(net_3868), .A1(net_1731) );
NAND3_X2 inst_2704 ( .ZN(net_2473), .A2(net_1811), .A3(net_1558), .A1(net_1338) );
CLKBUF_X2 inst_11842 ( .A(net_11803), .Z(net_11804) );
OAI22_X2 inst_1620 ( .B1(net_5942), .ZN(net_2785), .A1(net_2784), .B2(net_212), .A2(net_175) );
INV_X4 inst_4958 ( .ZN(net_4152), .A(net_724) );
CLKBUF_X2 inst_13344 ( .A(net_13305), .Z(net_13306) );
CLKBUF_X2 inst_8349 ( .A(net_8310), .Z(net_8311) );
CLKBUF_X2 inst_11461 ( .A(net_11422), .Z(net_11423) );
CLKBUF_X2 inst_10572 ( .A(net_9329), .Z(net_10534) );
INV_X2 inst_5924 ( .A(net_7443), .ZN(net_1488) );
SDFF_X2 inst_347 ( .SI(net_7303), .Q(net_7303), .D(net_4874), .SE(net_3859), .CK(net_9848) );
INV_X4 inst_5438 ( .A(net_7723), .ZN(net_2661) );
CLKBUF_X2 inst_11600 ( .A(net_11561), .Z(net_11562) );
CLKBUF_X2 inst_13327 ( .A(net_13288), .Z(net_13289) );
SDFF_X2 inst_755 ( .Q(net_6877), .D(net_6877), .SE(net_3901), .SI(net_3786), .CK(net_8500) );
CLKBUF_X2 inst_9508 ( .A(net_9469), .Z(net_9470) );
OAI21_X2 inst_1724 ( .ZN(net_5570), .B1(net_5442), .A(net_4835), .B2(net_4153) );
CLKBUF_X2 inst_7918 ( .A(net_7864), .Z(net_7880) );
CLKBUF_X2 inst_9701 ( .A(net_9662), .Z(net_9663) );
INV_X2 inst_5855 ( .ZN(net_668), .A(net_667) );
CLKBUF_X2 inst_13149 ( .A(net_13110), .Z(net_13111) );
INV_X8 inst_4505 ( .ZN(net_3781), .A(net_3261) );
NAND3_X2 inst_2610 ( .ZN(net_5729), .A1(net_5624), .A2(net_5149), .A3(net_4189) );
CLKBUF_X2 inst_8819 ( .A(net_8780), .Z(net_8781) );
INV_X4 inst_5473 ( .A(net_6111), .ZN(net_3673) );
SDFF_X2 inst_1043 ( .Q(net_7234), .D(net_7234), .SE(net_3822), .SI(net_330), .CK(net_12670) );
CLKBUF_X2 inst_12327 ( .A(net_12288), .Z(net_12289) );
NAND2_X2 inst_4030 ( .A1(net_7209), .A2(net_1648), .ZN(net_1022) );
CLKBUF_X2 inst_9234 ( .A(net_7868), .Z(net_9196) );
INV_X4 inst_4817 ( .ZN(net_4876), .A(net_1137) );
NAND2_X1 inst_4456 ( .A2(net_1256), .ZN(net_1118), .A1(net_1117) );
INV_X4 inst_4926 ( .A(net_3811), .ZN(net_3287) );
CLKBUF_X2 inst_9769 ( .A(net_8355), .Z(net_9731) );
DFF_X1 inst_6846 ( .D(net_2533), .QN(net_213), .CK(net_9545) );
OAI21_X2 inst_1792 ( .B1(net_5414), .ZN(net_5398), .A(net_4673), .B2(net_3988) );
NAND2_X1 inst_4426 ( .A1(net_7612), .A2(net_2131), .ZN(net_1454) );
CLKBUF_X2 inst_13840 ( .A(net_13801), .Z(net_13802) );
INV_X2 inst_6017 ( .A(net_7590), .ZN(net_2089) );
INV_X4 inst_4571 ( .ZN(net_5792), .A(net_5791) );
CLKBUF_X2 inst_10231 ( .A(net_10192), .Z(net_10193) );
INV_X4 inst_5111 ( .ZN(net_609), .A(net_608) );
NAND2_X2 inst_3928 ( .A1(net_7108), .A2(net_1675), .ZN(net_1370) );
NAND2_X2 inst_3353 ( .ZN(net_3539), .A1(net_3538), .A2(net_3226) );
NAND2_X2 inst_3634 ( .ZN(net_1949), .A1(net_1285), .A2(net_1122) );
CLKBUF_X2 inst_12877 ( .A(net_12838), .Z(net_12839) );
CLKBUF_X2 inst_12212 ( .A(net_12173), .Z(net_12174) );
CLKBUF_X2 inst_11849 ( .A(net_11810), .Z(net_11811) );
NAND2_X2 inst_4017 ( .A1(net_7198), .A2(net_1648), .ZN(net_1035) );
DFFR_X1 inst_7121 ( .Q(net_6025), .D(net_4796), .CK(net_10765), .RN(x1822) );
INV_X4 inst_4598 ( .ZN(net_5055), .A(net_4291) );
INV_X4 inst_4681 ( .ZN(net_3381), .A(net_3380) );
INV_X4 inst_5135 ( .ZN(net_666), .A(net_581) );
CLKBUF_X2 inst_12879 ( .A(net_10122), .Z(net_12841) );
CLKBUF_X2 inst_13050 ( .A(net_13011), .Z(net_13012) );
CLKBUF_X2 inst_9772 ( .A(net_9733), .Z(net_9734) );
CLKBUF_X2 inst_11204 ( .A(net_11165), .Z(net_11166) );
INV_X2 inst_5760 ( .ZN(net_3035), .A(net_2992) );
AOI222_X2 inst_7556 ( .A1(net_7550), .ZN(net_5227), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_382), .C2(net_380) );
CLKBUF_X2 inst_11513 ( .A(net_9835), .Z(net_11475) );
DFFR_X2 inst_7037 ( .QN(net_5997), .D(net_3161), .CK(net_10348), .RN(x1822) );
AOI22_X2 inst_7294 ( .B1(net_6544), .A1(net_6512), .A2(net_5184), .B2(net_5183), .ZN(net_5181) );
INV_X4 inst_5095 ( .A(net_7797), .ZN(net_3799) );
SDFF_X2 inst_426 ( .SI(net_7750), .Q(net_7750), .SE(net_5925), .D(net_3915), .CK(net_10329) );
NAND2_X2 inst_3145 ( .ZN(net_4818), .A2(net_4153), .A1(net_2103) );
INV_X4 inst_5144 ( .ZN(net_640), .A(net_572) );
SDFF_X2 inst_648 ( .Q(net_6694), .D(net_6694), .SE(net_3871), .SI(net_3792), .CK(net_11113) );
CLKBUF_X2 inst_10600 ( .A(net_10561), .Z(net_10562) );
INV_X2 inst_6035 ( .ZN(net_3075), .A(net_273) );
AND2_X2 inst_7857 ( .ZN(net_2701), .A1(net_2700), .A2(net_2699) );
CLKBUF_X2 inst_13718 ( .A(net_13679), .Z(net_13680) );
SDFF_X2 inst_270 ( .D(net_6400), .SE(net_6052), .SI(net_325), .Q(net_325), .CK(net_14222) );
OAI21_X2 inst_1901 ( .B1(net_5196), .ZN(net_5174), .A(net_4552), .B2(net_3866) );
CLKBUF_X2 inst_13856 ( .A(net_13817), .Z(net_13818) );
NAND2_X1 inst_4302 ( .ZN(net_4564), .A2(net_3866), .A1(net_1854) );
CLKBUF_X2 inst_11654 ( .A(net_11615), .Z(net_11616) );
CLKBUF_X2 inst_11068 ( .A(net_11029), .Z(net_11030) );
CLKBUF_X2 inst_8092 ( .A(net_7902), .Z(net_8054) );
DFF_X1 inst_6560 ( .QN(net_7658), .D(net_5194), .CK(net_10601) );
AOI21_X2 inst_7725 ( .B1(net_6459), .ZN(net_5901), .B2(net_2580), .A(net_2347) );
NAND2_X2 inst_4104 ( .A1(net_6666), .A2(net_1655), .ZN(net_948) );
DFF_X1 inst_6341 ( .Q(net_6190), .D(net_5845), .CK(net_13770) );
CLKBUF_X2 inst_11826 ( .A(net_11474), .Z(net_11788) );
CLKBUF_X2 inst_8608 ( .A(net_7900), .Z(net_8570) );
NOR2_X2 inst_2552 ( .A2(net_6012), .A1(net_6006), .ZN(net_2883) );
CLKBUF_X2 inst_11809 ( .A(net_11770), .Z(net_11771) );
SDFF_X2 inst_631 ( .SI(net_6624), .Q(net_6624), .SE(net_3850), .D(net_3806), .CK(net_9332) );
CLKBUF_X2 inst_11163 ( .A(net_9413), .Z(net_11125) );
CLKBUF_X2 inst_8544 ( .A(net_8505), .Z(net_8506) );
CLKBUF_X2 inst_9247 ( .A(net_9208), .Z(net_9209) );
DFF_X1 inst_6427 ( .QN(net_6182), .D(net_5743), .CK(net_10676) );
NAND2_X2 inst_3674 ( .A1(net_7336), .A2(net_1798), .ZN(net_1783) );
CLKBUF_X2 inst_9904 ( .A(net_7975), .Z(net_9866) );
CLKBUF_X2 inst_12835 ( .A(net_12796), .Z(net_12797) );
CLKBUF_X2 inst_11346 ( .A(net_11307), .Z(net_11308) );
CLKBUF_X2 inst_13505 ( .A(net_13466), .Z(net_13467) );
CLKBUF_X2 inst_13789 ( .A(net_13750), .Z(net_13751) );
CLKBUF_X2 inst_12558 ( .A(net_12519), .Z(net_12520) );
CLKBUF_X2 inst_8136 ( .A(net_8097), .Z(net_8098) );
NAND2_X2 inst_3995 ( .A2(net_1910), .ZN(net_1194), .A1(net_1193) );
NAND2_X2 inst_4211 ( .A2(net_5998), .A1(net_5997), .ZN(net_3243) );
INV_X4 inst_5074 ( .A(net_6688), .ZN(net_1151) );
OAI21_X2 inst_1745 ( .ZN(net_5526), .A(net_4822), .B2(net_4153), .B1(net_1260) );
NAND2_X2 inst_3831 ( .A1(net_6833), .A2(net_1521), .ZN(net_1509) );
OAI21_X2 inst_2079 ( .B2(net_4415), .ZN(net_4411), .B1(net_4029), .A(net_3506) );
XNOR2_X2 inst_102 ( .ZN(net_1918), .A(net_745), .B(net_417) );
CLKBUF_X2 inst_10534 ( .A(net_10495), .Z(net_10496) );
NOR2_X2 inst_2527 ( .ZN(net_3834), .A1(net_1726), .A2(net_568) );
DFF_X1 inst_6819 ( .QN(net_5960), .D(net_3013), .CK(net_10736) );
NAND2_X2 inst_3277 ( .ZN(net_3692), .A1(net_3691), .A2(net_3231) );
CLKBUF_X2 inst_12042 ( .A(net_12003), .Z(net_12004) );
CLKBUF_X2 inst_9299 ( .A(net_8759), .Z(net_9261) );
CLKBUF_X2 inst_14053 ( .A(net_14014), .Z(net_14015) );
INV_X4 inst_5352 ( .A(net_6555), .ZN(net_831) );
NAND3_X2 inst_2786 ( .ZN(net_2314), .A3(net_1626), .A1(net_1486), .A2(net_980) );
CLKBUF_X2 inst_11045 ( .A(net_11006), .Z(net_11007) );
CLKBUF_X2 inst_10043 ( .A(net_10004), .Z(net_10005) );
SDFF_X2 inst_1224 ( .SI(net_7217), .Q(net_7217), .D(net_3775), .SE(net_3750), .CK(net_11536) );
NAND2_X2 inst_3905 ( .A1(net_6966), .A2(net_1833), .ZN(net_1405) );
AOI21_X2 inst_7666 ( .ZN(net_3011), .B1(net_2867), .B2(net_2745), .A(net_1048) );
DFF_X1 inst_6554 ( .QN(net_7253), .D(net_5150), .CK(net_9465) );
INV_X4 inst_5615 ( .A(net_7256), .ZN(net_2001) );
CLKBUF_X2 inst_11797 ( .A(net_10858), .Z(net_11759) );
CLKBUF_X2 inst_8929 ( .A(net_8867), .Z(net_8891) );
SDFF_X2 inst_1170 ( .SI(net_6941), .Q(net_6941), .D(net_3785), .SE(net_3734), .CK(net_8488) );
CLKBUF_X2 inst_14246 ( .A(net_9848), .Z(net_14208) );
CLKBUF_X2 inst_12081 ( .A(net_11624), .Z(net_12043) );
NAND3_X2 inst_2596 ( .ZN(net_5743), .A1(net_5638), .A2(net_5217), .A3(net_4187) );
CLKBUF_X2 inst_11659 ( .A(net_11620), .Z(net_11621) );
DFF_X1 inst_6599 ( .QN(net_7497), .D(net_5409), .CK(net_9656) );
DFF_X2 inst_6242 ( .QN(net_7768), .D(net_3008), .CK(net_10407) );
CLKBUF_X2 inst_8752 ( .A(net_8713), .Z(net_8714) );
CLKBUF_X2 inst_8579 ( .A(net_8540), .Z(net_8541) );
NAND2_X2 inst_3022 ( .A1(net_6881), .A2(net_5006), .ZN(net_4987) );
CLKBUF_X2 inst_12133 ( .A(net_12094), .Z(net_12095) );
SDFF_X2 inst_680 ( .Q(net_6745), .D(net_6745), .SE(net_3815), .SI(net_3807), .CK(net_11338) );
DFF_X1 inst_6575 ( .QN(net_7565), .D(net_5079), .CK(net_13096) );
SDFF_X2 inst_785 ( .SI(net_6913), .Q(net_6913), .D(net_3805), .SE(net_3781), .CK(net_8147) );
NOR2_X2 inst_2362 ( .ZN(net_5288), .A2(net_4631), .A1(net_4488) );
CLKBUF_X2 inst_10323 ( .A(net_10284), .Z(net_10285) );
NAND2_X2 inst_3299 ( .ZN(net_3648), .A1(net_3647), .A2(net_3226) );
NAND2_X4 inst_2856 ( .A1(net_5877), .ZN(net_5089), .A2(net_4151) );
CLKBUF_X2 inst_9280 ( .A(net_9241), .Z(net_9242) );
CLKBUF_X2 inst_10417 ( .A(net_7873), .Z(net_10379) );
AND2_X4 inst_7820 ( .ZN(net_3260), .A2(net_3169), .A1(net_598) );
DFFR_X2 inst_7065 ( .QN(net_6044), .D(net_3058), .CK(net_10008), .RN(x1822) );
AOI21_X2 inst_7643 ( .B1(net_5890), .ZN(net_3910), .B2(net_3909), .A(net_2611) );
CLKBUF_X2 inst_7945 ( .A(net_7906), .Z(net_7907) );
AOI222_X2 inst_7551 ( .C1(net_7674), .A1(net_7642), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1849), .B1(net_1848) );
SDFF_X2 inst_527 ( .SI(net_6633), .Q(net_6633), .D(net_3894), .SE(net_3851), .CK(net_9199) );
CLKBUF_X2 inst_12697 ( .A(net_12658), .Z(net_12659) );
NAND2_X2 inst_3567 ( .ZN(net_2500), .A2(net_2006), .A1(net_1777) );
SDFF_X2 inst_226 ( .Q(net_6328), .SI(net_6327), .D(net_3629), .SE(net_392), .CK(net_14028) );
SDFF_X2 inst_1180 ( .SI(net_6953), .Q(net_6953), .D(net_3788), .SE(net_3741), .CK(net_11446) );
INV_X4 inst_5509 ( .A(net_7424), .ZN(net_2152) );
SDFF_X2 inst_414 ( .D(net_6392), .SE(net_5800), .SI(net_357), .Q(net_357), .CK(net_13666) );
CLKBUF_X2 inst_13861 ( .A(net_13822), .Z(net_13823) );
CLKBUF_X2 inst_8223 ( .A(net_8184), .Z(net_8185) );
CLKBUF_X2 inst_11232 ( .A(net_8549), .Z(net_11194) );
SDFF_X2 inst_531 ( .Q(net_6612), .D(net_6612), .SI(net_3900), .SE(net_3830), .CK(net_12200) );
CLKBUF_X2 inst_11688 ( .A(net_11649), .Z(net_11650) );
SDFF_X2 inst_212 ( .Q(net_6302), .SI(net_6301), .D(net_3625), .SE(net_392), .CK(net_13547) );
NAND3_X2 inst_2732 ( .ZN(net_2369), .A3(net_1630), .A1(net_1492), .A2(net_996) );
CLKBUF_X2 inst_9315 ( .A(net_9276), .Z(net_9277) );
DFF_X2 inst_6321 ( .QN(net_7815), .CK(net_10886), .D(x1417) );
OAI21_X2 inst_1952 ( .ZN(net_5068), .B1(net_4851), .A(net_4725), .B2(net_3986) );
CLKBUF_X2 inst_9323 ( .A(net_9284), .Z(net_9285) );
CLKBUF_X2 inst_10013 ( .A(net_9697), .Z(net_9975) );
CLKBUF_X2 inst_8827 ( .A(net_8375), .Z(net_8789) );
INV_X2 inst_6060 ( .A(net_7598), .ZN(net_1389) );
INV_X4 inst_5431 ( .A(net_7685), .ZN(net_449) );
INV_X4 inst_5023 ( .A(net_6408), .ZN(net_1683) );
CLKBUF_X2 inst_8330 ( .A(net_8291), .Z(net_8292) );
INV_X4 inst_5617 ( .A(net_6073), .ZN(net_3528) );
NAND2_X2 inst_3698 ( .ZN(net_1732), .A1(net_1280), .A2(net_1099) );
NAND2_X2 inst_4155 ( .ZN(net_929), .A1(net_572), .A2(net_468) );
DFFR_X2 inst_6962 ( .QN(net_7746), .D(net_4602), .CK(net_13232), .RN(x1822) );
INV_X4 inst_5118 ( .ZN(net_635), .A(net_600) );
NAND2_X2 inst_2966 ( .ZN(net_5461), .A1(net_4888), .A2(net_4887) );
CLKBUF_X2 inst_14223 ( .A(net_14184), .Z(net_14185) );
NAND2_X2 inst_3246 ( .A2(net_3992), .ZN(net_3988), .A1(net_1652) );
CLKBUF_X2 inst_9686 ( .A(net_9647), .Z(net_9648) );
CLKBUF_X2 inst_10208 ( .A(net_10169), .Z(net_10170) );
INV_X4 inst_4904 ( .A(net_3854), .ZN(net_865) );
CLKBUF_X2 inst_10699 ( .A(net_10560), .Z(net_10661) );
INV_X4 inst_4887 ( .ZN(net_1300), .A(net_880) );
CLKBUF_X2 inst_11272 ( .A(net_11233), .Z(net_11234) );
INV_X2 inst_5823 ( .ZN(net_934), .A(net_933) );
NOR2_X2 inst_2381 ( .ZN(net_5126), .A2(net_4603), .A1(net_4401) );
CLKBUF_X2 inst_11538 ( .A(net_8861), .Z(net_11500) );
INV_X4 inst_5338 ( .A(net_7700), .ZN(net_844) );
SDFF_X2 inst_570 ( .SI(net_6768), .Q(net_6768), .D(net_3894), .SE(net_3816), .CK(net_11122) );
OAI22_X2 inst_1570 ( .A2(net_3297), .B2(net_3286), .ZN(net_3279), .A1(net_3128), .B1(net_1716) );
CLKBUF_X2 inst_11284 ( .A(net_11245), .Z(net_11246) );
CLKBUF_X2 inst_12055 ( .A(net_9047), .Z(net_12017) );
OAI22_X2 inst_1612 ( .A1(net_3280), .A2(net_3087), .B2(net_3084), .ZN(net_3060), .B1(net_727) );
INV_X4 inst_4645 ( .ZN(net_4177), .A(net_4013) );
SDFF_X2 inst_454 ( .Q(net_6059), .SI(net_3920), .SE(net_3316), .D(net_3315), .CK(net_10386) );
CLKBUF_X2 inst_13947 ( .A(net_11179), .Z(net_13909) );
CLKBUF_X2 inst_13753 ( .A(net_13714), .Z(net_13715) );
CLKBUF_X2 inst_14299 ( .A(net_14260), .Z(net_14261) );
CLKBUF_X2 inst_12545 ( .A(net_9931), .Z(net_12507) );
CLKBUF_X2 inst_8251 ( .A(net_8107), .Z(net_8213) );
CLKBUF_X2 inst_7899 ( .A(net_7860), .Z(net_7861) );
CLKBUF_X2 inst_11419 ( .A(net_11380), .Z(net_11381) );
NAND2_X2 inst_3718 ( .A1(net_6770), .A2(net_1635), .ZN(net_1628) );
CLKBUF_X2 inst_12592 ( .A(net_12553), .Z(net_12554) );
CLKBUF_X2 inst_11130 ( .A(net_10776), .Z(net_11092) );
NAND2_X2 inst_3077 ( .A1(net_6479), .ZN(net_4928), .A2(net_4927) );
CLKBUF_X2 inst_11067 ( .A(net_11028), .Z(net_11029) );
DFFR_X2 inst_6990 ( .QN(net_7698), .D(net_3344), .CK(net_12879), .RN(x1822) );
CLKBUF_X2 inst_13622 ( .A(net_13583), .Z(net_13584) );
CLKBUF_X2 inst_12974 ( .A(net_11672), .Z(net_12936) );
CLKBUF_X2 inst_12599 ( .A(net_12560), .Z(net_12561) );
INV_X4 inst_5224 ( .ZN(net_466), .A(net_465) );
CLKBUF_X2 inst_8099 ( .A(net_7984), .Z(net_8061) );
CLKBUF_X2 inst_9566 ( .A(net_8233), .Z(net_9528) );
OR2_X2 inst_1423 ( .A2(net_7228), .A1(net_7227), .ZN(net_667) );
NOR2_X2 inst_2419 ( .A2(net_7768), .ZN(net_4146), .A1(net_153) );
SDFF_X2 inst_1034 ( .Q(net_7550), .D(net_7550), .SE(net_3896), .SI(net_384), .CK(net_13109) );
CLKBUF_X2 inst_11612 ( .A(net_11573), .Z(net_11574) );
CLKBUF_X2 inst_9484 ( .A(net_9445), .Z(net_9446) );
CLKBUF_X2 inst_9855 ( .A(net_9816), .Z(net_9817) );
SDFF_X2 inst_1207 ( .SI(net_7091), .Q(net_7091), .D(net_3800), .SE(net_3742), .CK(net_11838) );
SDFF_X2 inst_613 ( .Q(net_6619), .D(net_6619), .SE(net_3830), .SI(net_3793), .CK(net_12023) );
CLKBUF_X2 inst_9945 ( .A(net_9906), .Z(net_9907) );
NAND2_X1 inst_4275 ( .ZN(net_4593), .A2(net_3867), .A1(net_1193) );
CLKBUF_X2 inst_8694 ( .A(net_8655), .Z(net_8656) );
INV_X4 inst_5041 ( .A(net_2275), .ZN(net_2232) );
DFF_X1 inst_6444 ( .QN(net_6095), .D(net_5726), .CK(net_9224) );
OR2_X2 inst_1428 ( .A2(net_6553), .A1(net_6552), .ZN(net_669) );
CLKBUF_X2 inst_11089 ( .A(net_10312), .Z(net_11051) );
SDFF_X2 inst_483 ( .Q(net_7106), .D(net_7106), .SI(net_3890), .SE(net_3888), .CK(net_11594) );
INV_X4 inst_5005 ( .A(net_7815), .ZN(net_3804) );
CLKBUF_X2 inst_9907 ( .A(net_9428), .Z(net_9869) );
CLKBUF_X2 inst_9456 ( .A(net_9417), .Z(net_9418) );
NAND3_X2 inst_2739 ( .ZN(net_2362), .A3(net_1525), .A1(net_1313), .A2(net_1014) );
SDFF_X2 inst_259 ( .Q(net_6375), .SI(net_6374), .D(net_3705), .SE(net_392), .CK(net_13960) );
CLKBUF_X2 inst_12691 ( .A(net_12652), .Z(net_12653) );
DFF_X1 inst_6845 ( .D(net_2562), .Q(net_203), .CK(net_10068) );
SDFF_X2 inst_1046 ( .Q(net_7247), .D(net_7247), .SE(net_3822), .SI(net_343), .CK(net_9831) );
DFF_X1 inst_6812 ( .D(net_3301), .CK(net_13212), .Q(x287) );
INV_X2 inst_5955 ( .A(net_7622), .ZN(net_1195) );
CLKBUF_X2 inst_10152 ( .A(net_10113), .Z(net_10114) );
NAND2_X1 inst_4355 ( .ZN(net_4372), .A2(net_3853), .A1(net_2014) );
INV_X4 inst_5426 ( .A(net_7732), .ZN(net_2682) );
INV_X4 inst_4707 ( .ZN(net_3031), .A(net_2953) );
DFF_X2 inst_6206 ( .QN(net_7534), .D(net_4169), .CK(net_12600) );
INV_X4 inst_4846 ( .ZN(net_4778), .A(net_1064) );
CLKBUF_X2 inst_9515 ( .A(net_8253), .Z(net_9477) );
CLKBUF_X2 inst_8621 ( .A(net_8582), .Z(net_8583) );
AOI222_X2 inst_7592 ( .A1(net_7390), .ZN(net_5548), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_353), .C2(net_351) );
CLKBUF_X2 inst_13197 ( .A(net_12567), .Z(net_13159) );
CLKBUF_X2 inst_10517 ( .A(net_10478), .Z(net_10479) );
SDFF_X2 inst_909 ( .Q(net_7146), .D(net_7146), .SE(net_3903), .SI(net_3787), .CK(net_7854) );
NOR2_X2 inst_2484 ( .A2(net_5778), .ZN(net_2657), .A1(net_2595) );
CLKBUF_X2 inst_9927 ( .A(net_8003), .Z(net_9889) );
INV_X2 inst_5758 ( .ZN(net_3089), .A(net_2712) );
DFF_X1 inst_6494 ( .QN(net_7406), .D(net_5549), .CK(net_12123) );
CLKBUF_X2 inst_10686 ( .A(net_8843), .Z(net_10648) );
NAND2_X2 inst_2919 ( .A2(net_7773), .ZN(net_5773), .A1(net_5609) );
SDFF_X2 inst_894 ( .Q(net_7126), .D(net_7126), .SE(net_3888), .SI(net_3794), .CK(net_8715) );
INV_X4 inst_5039 ( .A(net_7805), .ZN(net_3812) );
NOR2_X2 inst_2425 ( .A2(net_5893), .ZN(net_3223), .A1(net_682) );
OAI21_X2 inst_1872 ( .ZN(net_5236), .B1(net_5235), .A(net_4591), .B2(net_3867) );
CLKBUF_X2 inst_10795 ( .A(net_10756), .Z(net_10757) );
CLKBUF_X2 inst_10827 ( .A(net_10788), .Z(net_10789) );
SDFF_X2 inst_994 ( .Q(net_6482), .D(net_6482), .SE(net_3904), .SI(net_3790), .CK(net_8412) );
CLKBUF_X2 inst_9803 ( .A(net_9764), .Z(net_9765) );
CLKBUF_X2 inst_12003 ( .A(net_11964), .Z(net_11965) );
NAND2_X2 inst_4028 ( .A1(net_6803), .A2(net_1651), .ZN(net_1024) );
CLKBUF_X2 inst_8478 ( .A(net_8439), .Z(net_8440) );
OAI21_X2 inst_1879 ( .ZN(net_5209), .B1(net_5208), .A(net_4579), .B2(net_3867) );
OAI21_X2 inst_1863 ( .ZN(net_5252), .B1(net_5208), .A(net_4536), .B2(net_3870) );
OAI21_X2 inst_2135 ( .ZN(net_2849), .B2(net_2820), .A(net_2710), .B1(net_898) );
CLKBUF_X2 inst_13556 ( .A(net_13517), .Z(net_13518) );
CLKBUF_X2 inst_14082 ( .A(net_14043), .Z(net_14044) );
NAND2_X2 inst_3119 ( .A1(net_6622), .A2(net_4899), .ZN(net_4882) );
INV_X4 inst_5138 ( .A(net_710), .ZN(net_577) );
NAND2_X2 inst_3777 ( .A1(net_6774), .A2(net_1635), .ZN(net_1568) );
SDFF_X2 inst_764 ( .Q(net_6888), .D(net_6888), .SE(net_3901), .SI(net_3794), .CK(net_11479) );
CLKBUF_X2 inst_10961 ( .A(net_10922), .Z(net_10923) );
CLKBUF_X2 inst_12015 ( .A(net_11976), .Z(net_11977) );
OAI22_X2 inst_1547 ( .B2(net_3405), .A2(net_3360), .ZN(net_3358), .A1(net_3287), .B1(net_461) );
XNOR2_X2 inst_29 ( .ZN(net_2485), .A(net_2484), .B(net_911) );
CLKBUF_X2 inst_9900 ( .A(net_9861), .Z(net_9862) );
CLKBUF_X2 inst_8469 ( .A(net_8430), .Z(net_8431) );
DFF_X1 inst_6937 ( .D(net_2406), .Q(net_258), .CK(net_13267) );
CLKBUF_X2 inst_9713 ( .A(net_9674), .Z(net_9675) );
AOI21_X2 inst_7782 ( .B1(net_6609), .ZN(net_4014), .B2(net_2583), .A(net_2284) );
CLKBUF_X2 inst_11745 ( .A(net_11339), .Z(net_11707) );
NOR2_X2 inst_2369 ( .ZN(net_5267), .A2(net_4618), .A1(net_4464) );
OAI21_X2 inst_2152 ( .B1(net_5778), .ZN(net_2792), .A(net_2656), .B2(net_2654) );
INV_X2 inst_6105 ( .A(net_7634), .ZN(net_1862) );
CLKBUF_X2 inst_10540 ( .A(net_9926), .Z(net_10502) );
NAND2_X2 inst_3947 ( .A1(net_7101), .A2(net_1675), .ZN(net_1341) );
SDFF_X2 inst_1274 ( .D(net_6388), .SE(net_5800), .SI(net_353), .Q(net_353), .CK(net_13664) );
CLKBUF_X2 inst_13270 ( .A(net_13231), .Z(net_13232) );
AOI21_X2 inst_7740 ( .B1(net_7143), .ZN(net_4076), .B2(net_2582), .A(net_2313) );
NAND2_X2 inst_3838 ( .A1(net_6443), .A2(net_1677), .ZN(net_1501) );
CLKBUF_X2 inst_11152 ( .A(net_8287), .Z(net_11114) );
CLKBUF_X2 inst_10590 ( .A(net_10551), .Z(net_10552) );
CLKBUF_X2 inst_12775 ( .A(net_12736), .Z(net_12737) );
INV_X4 inst_5495 ( .A(net_7564), .ZN(net_1894) );
INV_X4 inst_5326 ( .A(net_7707), .ZN(net_847) );
DFF_X2 inst_6207 ( .QN(net_7535), .D(net_4302), .CK(net_9527) );
CLKBUF_X2 inst_11396 ( .A(net_11265), .Z(net_11358) );
SDFF_X2 inst_538 ( .Q(net_6584), .D(net_6584), .SI(net_3898), .SE(net_3823), .CK(net_12037) );
NAND3_X2 inst_2831 ( .A1(net_7782), .A3(net_7781), .ZN(net_936), .A2(net_510) );
CLKBUF_X2 inst_12785 ( .A(net_7954), .Z(net_12747) );
CLKBUF_X2 inst_8344 ( .A(net_8305), .Z(net_8306) );
SDFF_X2 inst_1300 ( .D(net_6387), .SE(net_5800), .SI(net_352), .Q(net_352), .CK(net_13663) );
INV_X4 inst_5280 ( .A(net_7262), .ZN(net_2079) );
INV_X8 inst_4537 ( .ZN(net_2644), .A(net_2488) );
CLKBUF_X2 inst_12022 ( .A(net_11983), .Z(net_11984) );
XNOR2_X2 inst_35 ( .ZN(net_2454), .B(net_2453), .A(net_1939) );
INV_X4 inst_5317 ( .A(net_6108), .ZN(net_3679) );
CLKBUF_X2 inst_13698 ( .A(net_13659), .Z(net_13660) );
CLKBUF_X2 inst_8890 ( .A(net_8851), .Z(net_8852) );
INV_X4 inst_4765 ( .ZN(net_2427), .A(net_1936) );
CLKBUF_X2 inst_13693 ( .A(net_13654), .Z(net_13655) );
CLKBUF_X2 inst_10599 ( .A(net_10041), .Z(net_10561) );
CLKBUF_X2 inst_11146 ( .A(net_11107), .Z(net_11108) );
AOI22_X2 inst_7309 ( .B1(net_6682), .A1(net_6650), .A2(net_5139), .B2(net_5138), .ZN(net_5134) );
NOR2_X4 inst_2279 ( .ZN(net_3839), .A1(net_3401), .A2(net_3232) );
CLKBUF_X2 inst_12572 ( .A(net_10390), .Z(net_12534) );
NAND3_X2 inst_2600 ( .ZN(net_5739), .A1(net_5634), .A2(net_5186), .A3(net_4201) );
CLKBUF_X2 inst_14158 ( .A(net_11010), .Z(net_14120) );
OAI21_X2 inst_2038 ( .B1(net_4624), .B2(net_4476), .ZN(net_4465), .A(net_3584) );
OAI21_X2 inst_2044 ( .B2(net_4457), .ZN(net_4456), .B1(net_4082), .A(net_3567) );
AND2_X4 inst_7833 ( .ZN(net_2993), .A1(net_2855), .A2(net_227) );
INV_X4 inst_5178 ( .ZN(net_772), .A(net_527) );
NOR2_X4 inst_2274 ( .ZN(net_5612), .A1(net_5457), .A2(net_4400) );
CLKBUF_X2 inst_10055 ( .A(net_10016), .Z(net_10017) );
SDFF_X2 inst_695 ( .SI(net_7799), .Q(net_6732), .D(net_6732), .SE(net_3815), .CK(net_11097) );
CLKBUF_X2 inst_13630 ( .A(net_8170), .Z(net_13592) );
DFF_X2 inst_6249 ( .QN(net_7759), .D(net_3019), .CK(net_10516) );
NAND2_X2 inst_4038 ( .A1(net_6659), .A2(net_1655), .ZN(net_1014) );
CLKBUF_X2 inst_13711 ( .A(net_13672), .Z(net_13673) );
CLKBUF_X2 inst_10606 ( .A(net_10567), .Z(net_10568) );
INV_X4 inst_5492 ( .A(net_5993), .ZN(net_2594) );
CLKBUF_X2 inst_10663 ( .A(net_10624), .Z(net_10625) );
CLKBUF_X2 inst_14001 ( .A(net_13962), .Z(net_13963) );
CLKBUF_X2 inst_10782 ( .A(net_9894), .Z(net_10744) );
DFF_X1 inst_6877 ( .D(net_2496), .Q(net_165), .CK(net_10229) );
DFF_X1 inst_6610 ( .QN(net_7498), .D(net_5397), .CK(net_12549) );
NOR2_X2 inst_2493 ( .ZN(net_2584), .A2(net_1832), .A1(net_624) );
CLKBUF_X2 inst_14376 ( .A(net_14337), .Z(net_14338) );
INV_X1 inst_6154 ( .A(net_5859), .ZN(x131) );
SDFF_X2 inst_511 ( .SI(net_6914), .Q(net_6914), .D(net_3900), .SE(net_3887), .CK(net_8157) );
CLKBUF_X2 inst_9593 ( .A(net_9554), .Z(net_9555) );
CLKBUF_X2 inst_8665 ( .A(net_8626), .Z(net_8627) );
NAND2_X2 inst_3559 ( .ZN(net_2508), .A2(net_2032), .A1(net_1801) );
INV_X2 inst_5720 ( .ZN(net_4246), .A(net_4113) );
CLKBUF_X2 inst_12277 ( .A(net_10823), .Z(net_12239) );
NAND3_X2 inst_2645 ( .ZN(net_5949), .A3(net_3963), .A2(net_1386), .A1(net_806) );
SDFF_X2 inst_1164 ( .SI(net_7198), .Q(net_7198), .D(net_3892), .SE(net_3750), .CK(net_10481) );
CLKBUF_X2 inst_9449 ( .A(net_8311), .Z(net_9411) );
NAND2_X2 inst_3112 ( .A1(net_6586), .A2(net_4897), .ZN(net_4889) );
CLKBUF_X2 inst_14025 ( .A(net_13986), .Z(net_13987) );
CLKBUF_X2 inst_11772 ( .A(net_11733), .Z(net_11734) );
CLKBUF_X2 inst_8328 ( .A(net_8289), .Z(net_8290) );
CLKBUF_X2 inst_12790 ( .A(net_12751), .Z(net_12752) );
CLKBUF_X2 inst_11410 ( .A(net_11371), .Z(net_11372) );
AOI22_X2 inst_7276 ( .B1(net_7090), .A1(net_7058), .A2(net_5280), .B2(net_5279), .ZN(net_5272) );
DFFR_X2 inst_7004 ( .QN(net_7696), .D(net_3346), .CK(net_12876), .RN(x1822) );
INV_X2 inst_6001 ( .A(net_7282), .ZN(net_2160) );
CLKBUF_X2 inst_12506 ( .A(net_12467), .Z(net_12468) );
CLKBUF_X2 inst_11416 ( .A(net_11377), .Z(net_11378) );
CLKBUF_X2 inst_8193 ( .A(net_8024), .Z(net_8155) );
SDFF_X2 inst_1242 ( .SI(net_6537), .Q(net_6537), .D(net_3776), .SE(net_3755), .CK(net_8483) );
CLKBUF_X2 inst_14086 ( .A(net_14047), .Z(net_14048) );
CLKBUF_X2 inst_11646 ( .A(net_8953), .Z(net_11608) );
CLKBUF_X2 inst_11525 ( .A(net_11486), .Z(net_11487) );
CLKBUF_X2 inst_10751 ( .A(net_10712), .Z(net_10713) );
CLKBUF_X2 inst_10666 ( .A(net_8010), .Z(net_10628) );
DFF_X1 inst_6592 ( .QN(net_7570), .D(net_5069), .CK(net_8043) );
CLKBUF_X2 inst_13363 ( .A(net_13324), .Z(net_13325) );
INV_X4 inst_5217 ( .A(net_578), .ZN(net_477) );
CLKBUF_X2 inst_8362 ( .A(net_8323), .Z(net_8324) );
CLKBUF_X2 inst_8069 ( .A(net_8029), .Z(net_8031) );
SDFF_X2 inst_388 ( .SI(net_7308), .Q(net_7308), .D(net_4779), .SE(net_3859), .CK(net_9923) );
INV_X4 inst_4600 ( .ZN(net_4244), .A(net_4111) );
CLKBUF_X2 inst_11574 ( .A(net_11535), .Z(net_11536) );
CLKBUF_X2 inst_9273 ( .A(net_9234), .Z(net_9235) );
DFF_X1 inst_6923 ( .D(net_2404), .Q(net_260), .CK(net_12391) );
NAND2_X2 inst_3872 ( .A2(net_1696), .ZN(net_1453), .A1(net_1452) );
CLKBUF_X2 inst_12374 ( .A(net_11832), .Z(net_12336) );
SDFF_X2 inst_489 ( .Q(net_7124), .D(net_7124), .SI(net_3902), .SE(net_3888), .CK(net_8732) );
CLKBUF_X2 inst_9278 ( .A(net_9239), .Z(net_9240) );
CLKBUF_X2 inst_10227 ( .A(net_8022), .Z(net_10189) );
INV_X4 inst_5502 ( .A(net_6020), .ZN(net_2843) );
NAND2_X2 inst_3622 ( .ZN(net_1963), .A2(net_1962), .A1(net_1719) );
CLKBUF_X2 inst_11625 ( .A(net_11586), .Z(net_11587) );
OR2_X2 inst_1411 ( .ZN(net_1231), .A1(net_861), .A2(net_825) );
SDFF_X2 inst_149 ( .Q(net_6229), .SI(net_6228), .SE(net_392), .D(net_135), .CK(net_14102) );
XNOR2_X2 inst_39 ( .ZN(net_2437), .A(net_1688), .B(net_425) );
CLKBUF_X2 inst_11028 ( .A(net_10432), .Z(net_10990) );
CLKBUF_X2 inst_12527 ( .A(net_10434), .Z(net_12489) );
CLKBUF_X2 inst_8854 ( .A(net_8389), .Z(net_8816) );
DFF_X1 inst_6924 ( .D(net_2412), .Q(net_245), .CK(net_13134) );
NAND3_X2 inst_2627 ( .ZN(net_5702), .A1(net_5679), .A2(net_5313), .A3(net_4253) );
CLKBUF_X2 inst_8987 ( .A(net_8948), .Z(net_8949) );
CLKBUF_X2 inst_9542 ( .A(net_8197), .Z(net_9504) );
AOI21_X2 inst_7771 ( .B1(net_6740), .ZN(net_4124), .B2(net_2581), .A(net_2367) );
NOR2_X2 inst_2320 ( .A2(net_6298), .A1(net_5843), .ZN(net_5821) );
NAND2_X2 inst_3173 ( .ZN(net_4760), .A2(net_3941), .A1(net_2075) );
SDFF_X2 inst_125 ( .Q(net_6197), .SI(net_6196), .D(net_3922), .SE(net_392), .CK(net_13758) );
NOR2_X2 inst_2534 ( .A2(net_7754), .A1(net_3208), .ZN(net_680) );
INV_X4 inst_4770 ( .ZN(net_1930), .A(net_1929) );
CLKBUF_X2 inst_10775 ( .A(net_9241), .Z(net_10737) );
INV_X4 inst_5377 ( .A(net_6107), .ZN(net_3683) );
AOI21_X2 inst_7696 ( .B1(net_6739), .ZN(net_4126), .B2(net_2581), .A(net_2368) );
NAND2_X2 inst_3737 ( .A1(net_6893), .A2(net_1639), .ZN(net_1608) );
CLKBUF_X2 inst_11919 ( .A(net_11880), .Z(net_11881) );
OAI222_X2 inst_1636 ( .A1(net_5868), .C2(net_5043), .ZN(net_5042), .A2(net_5041), .B2(net_5040), .B1(net_2443), .C1(net_580) );
SDFF_X2 inst_430 ( .SI(net_7760), .Q(net_7760), .SE(net_5925), .D(net_3905), .CK(net_12512) );
SDFF_X2 inst_515 ( .Q(net_6723), .D(net_6723), .SE(net_3871), .SI(net_3821), .CK(net_11398) );
CLKBUF_X2 inst_8501 ( .A(net_8056), .Z(net_8463) );
CLKBUF_X2 inst_12242 ( .A(net_9002), .Z(net_12204) );
AOI22_X2 inst_7278 ( .B1(net_7080), .A1(net_7048), .A2(net_5280), .B2(net_5279), .ZN(net_5266) );
OAI22_X2 inst_1501 ( .B1(net_4660), .A1(net_4105), .B2(net_4099), .ZN(net_4096), .A2(net_4095) );
CLKBUF_X2 inst_11800 ( .A(net_11761), .Z(net_11762) );
NAND2_X2 inst_3212 ( .ZN(net_4714), .A2(net_3986), .A1(net_1877) );
NAND4_X2 inst_2565 ( .ZN(net_1234), .A3(net_660), .A1(net_659), .A2(net_658), .A4(net_628) );
DFFR_X2 inst_7061 ( .QN(net_6042), .D(net_3064), .CK(net_10526), .RN(x1822) );
NAND2_X2 inst_2945 ( .ZN(net_5501), .A1(net_4962), .A2(net_4961) );
OAI22_X2 inst_1584 ( .A1(net_3270), .B2(net_3200), .ZN(net_3192), .A2(net_3187), .B1(net_441) );
SDFF_X2 inst_642 ( .SI(net_6654), .Q(net_6654), .SE(net_3851), .D(net_3800), .CK(net_12008) );
CLKBUF_X2 inst_14183 ( .A(net_14144), .Z(net_14145) );
CLKBUF_X2 inst_13035 ( .A(net_12996), .Z(net_12997) );
NAND2_X2 inst_2993 ( .A1(net_6756), .A2(net_5033), .ZN(net_5018) );
CLKBUF_X2 inst_9361 ( .A(net_9322), .Z(net_9323) );
CLKBUF_X2 inst_13168 ( .A(net_9007), .Z(net_13130) );
CLKBUF_X2 inst_11023 ( .A(net_9121), .Z(net_10985) );
CLKBUF_X2 inst_7933 ( .A(net_7864), .Z(net_7895) );
SDFF_X2 inst_1018 ( .SI(net_6512), .Q(net_6512), .SE(net_3889), .D(net_3779), .CK(net_11645) );
CLKBUF_X2 inst_10726 ( .A(net_10687), .Z(net_10688) );
CLKBUF_X2 inst_10655 ( .A(net_9527), .Z(net_10617) );
CLKBUF_X2 inst_8129 ( .A(net_8090), .Z(net_8091) );
CLKBUF_X2 inst_14160 ( .A(net_14121), .Z(net_14122) );
NAND2_X2 inst_2933 ( .ZN(net_5516), .A1(net_4989), .A2(net_4988) );
SDFF_X2 inst_700 ( .SI(net_6770), .Q(net_6770), .SE(net_3816), .D(net_3812), .CK(net_8279) );
CLKBUF_X2 inst_13507 ( .A(net_8319), .Z(net_13469) );
CLKBUF_X2 inst_12295 ( .A(net_12256), .Z(net_12257) );
CLKBUF_X2 inst_8706 ( .A(net_8667), .Z(net_8668) );
DFF_X1 inst_6467 ( .QN(net_6168), .D(net_5592), .CK(net_7972) );
CLKBUF_X2 inst_13323 ( .A(net_13284), .Z(net_13285) );
CLKBUF_X2 inst_8107 ( .A(net_8068), .Z(net_8069) );
CLKBUF_X2 inst_9152 ( .A(net_9113), .Z(net_9114) );
CLKBUF_X2 inst_8555 ( .A(net_8516), .Z(net_8517) );
SDFF_X2 inst_979 ( .Q(net_6432), .D(net_6432), .SE(net_3820), .SI(net_3814), .CK(net_11263) );
NAND3_X2 inst_2713 ( .ZN(net_2463), .A2(net_1810), .A3(net_1562), .A1(net_1368) );
SDFF_X2 inst_1008 ( .SI(net_6500), .Q(net_6500), .SE(net_3889), .D(net_3812), .CK(net_8635) );
CLKBUF_X2 inst_7877 ( .A(net_7838), .Z(net_7839) );
INV_X8 inst_4568 ( .ZN(net_5926), .A(net_5925) );
SDFF_X2 inst_559 ( .SI(net_7170), .Q(net_7170), .D(net_3890), .SE(net_3819), .CK(net_8729) );
CLKBUF_X2 inst_8872 ( .A(net_8833), .Z(net_8834) );
INV_X2 inst_5989 ( .A(net_7483), .ZN(net_2169) );
CLKBUF_X2 inst_9785 ( .A(net_9746), .Z(net_9747) );
CLKBUF_X2 inst_9476 ( .A(net_9437), .Z(net_9438) );
AOI21_X2 inst_7706 ( .B1(net_6458), .ZN(net_5900), .B2(net_2580), .A(net_2307) );
DFF_X1 inst_6725 ( .QN(net_7358), .D(net_5331), .CK(net_12979) );
NOR2_X4 inst_2296 ( .A1(net_7093), .ZN(net_791), .A2(net_570) );
CLKBUF_X2 inst_11596 ( .A(net_11557), .Z(net_11558) );
CLKBUF_X2 inst_9250 ( .A(net_8592), .Z(net_9212) );
CLKBUF_X2 inst_13092 ( .A(net_13053), .Z(net_13054) );
CLKBUF_X2 inst_12477 ( .A(net_9203), .Z(net_12439) );
CLKBUF_X2 inst_12012 ( .A(net_11973), .Z(net_11974) );
INV_X4 inst_4964 ( .ZN(net_2259), .A(net_716) );
CLKBUF_X2 inst_9587 ( .A(net_8799), .Z(net_9549) );
NAND2_X2 inst_3405 ( .A2(net_5972), .ZN(net_3382), .A1(net_2879) );
CLKBUF_X2 inst_14133 ( .A(net_14094), .Z(net_14095) );
CLKBUF_X2 inst_8979 ( .A(net_8940), .Z(net_8941) );
NAND2_X2 inst_3888 ( .A1(net_6832), .A2(net_1521), .ZN(net_1430) );
CLKBUF_X2 inst_12831 ( .A(net_12792), .Z(net_12793) );
NAND2_X1 inst_4258 ( .ZN(net_4665), .A2(net_3993), .A1(net_1381) );
CLKBUF_X2 inst_7889 ( .A(net_7850), .Z(net_7851) );
CLKBUF_X2 inst_9797 ( .A(net_9758), .Z(net_9759) );
CLKBUF_X2 inst_9607 ( .A(net_9568), .Z(net_9569) );
CLKBUF_X2 inst_9764 ( .A(net_9725), .Z(net_9726) );
CLKBUF_X2 inst_9018 ( .A(net_8979), .Z(net_8980) );
NAND2_X2 inst_4040 ( .A1(net_6795), .A2(net_1651), .ZN(net_1012) );
CLKBUF_X2 inst_12221 ( .A(net_12182), .Z(net_12183) );
AOI22_X2 inst_7366 ( .A2(net_5916), .B2(net_2957), .ZN(net_2956), .B1(net_2685), .A1(net_845) );
NAND2_X1 inst_4334 ( .ZN(net_4530), .A2(net_3870), .A1(net_1315) );
SDFF_X2 inst_1059 ( .SI(net_6903), .Q(net_6903), .D(net_3894), .SE(net_3781), .CK(net_11784) );
CLKBUF_X2 inst_8017 ( .A(net_7978), .Z(net_7979) );
SDFF_X2 inst_1075 ( .SI(net_7220), .Q(net_7220), .D(net_3902), .SE(net_3751), .CK(net_8696) );
CLKBUF_X2 inst_13987 ( .A(net_13948), .Z(net_13949) );
CLKBUF_X2 inst_14227 ( .A(net_14188), .Z(net_14189) );
CLKBUF_X2 inst_10215 ( .A(net_8779), .Z(net_10177) );
CLKBUF_X2 inst_12701 ( .A(net_12662), .Z(net_12663) );
CLKBUF_X2 inst_9230 ( .A(net_9191), .Z(net_9192) );
NAND2_X1 inst_4328 ( .ZN(net_4536), .A2(net_3870), .A1(net_2132) );
CLKBUF_X2 inst_11504 ( .A(net_8143), .Z(net_11466) );
NOR2_X4 inst_2257 ( .ZN(net_5629), .A1(net_5474), .A2(net_4432) );
CLKBUF_X2 inst_11781 ( .A(net_11742), .Z(net_11743) );
NAND2_X2 inst_4173 ( .A1(net_6958), .ZN(net_789), .A2(net_639) );
INV_X2 inst_6039 ( .A(net_7600), .ZN(net_1352) );
CLKBUF_X2 inst_12454 ( .A(net_11500), .Z(net_12416) );
DFF_X1 inst_6425 ( .QN(net_6180), .D(net_5745), .CK(net_10681) );
SDFF_X2 inst_1104 ( .SI(net_6806), .Q(net_6806), .D(net_3786), .SE(net_3729), .CK(net_11305) );
NOR2_X2 inst_2355 ( .ZN(net_5649), .A1(net_5501), .A2(net_4468) );
CLKBUF_X2 inst_14306 ( .A(net_12783), .Z(net_14268) );
CLKBUF_X2 inst_13641 ( .A(net_13602), .Z(net_13603) );
CLKBUF_X2 inst_10886 ( .A(net_8873), .Z(net_10848) );
DFF_X1 inst_6536 ( .QN(net_7468), .D(net_5580), .CK(net_9668) );
INV_X2 inst_5753 ( .ZN(net_3907), .A(net_3736) );
DFFR_X2 inst_7058 ( .QN(net_5996), .D(net_3206), .CK(net_9605), .RN(x1822) );
CLKBUF_X2 inst_12535 ( .A(net_12496), .Z(net_12497) );
CLKBUF_X2 inst_9742 ( .A(net_9703), .Z(net_9704) );
DFF_X1 inst_6434 ( .QN(net_6077), .D(net_5736), .CK(net_8442) );
INV_X2 inst_6110 ( .ZN(net_5918), .A(net_5862) );
SDFF_X2 inst_329 ( .SI(net_7495), .Q(net_7495), .D(net_5097), .SE(net_3989), .CK(net_12441) );
SDFF_X2 inst_494 ( .SI(net_6896), .Q(net_6896), .D(net_3892), .SE(net_3887), .CK(net_8973) );
AOI22_X2 inst_7287 ( .B1(net_7224), .A1(net_7192), .A2(net_5244), .B2(net_5243), .ZN(net_5218) );
SDFF_X2 inst_574 ( .Q(net_6570), .D(net_6570), .SE(net_3823), .SI(net_3813), .CK(net_9360) );
CLKBUF_X2 inst_12446 ( .A(net_12407), .Z(net_12408) );
INV_X4 inst_5552 ( .A(net_6012), .ZN(net_474) );
INV_X2 inst_5942 ( .A(net_7503), .ZN(net_2109) );
CLKBUF_X2 inst_13845 ( .A(net_13806), .Z(net_13807) );
NOR2_X2 inst_2347 ( .ZN(net_5657), .A1(net_5509), .A2(net_4478) );
CLKBUF_X2 inst_14349 ( .A(net_14310), .Z(net_14311) );
CLKBUF_X2 inst_13085 ( .A(net_13046), .Z(net_13047) );
CLKBUF_X2 inst_8087 ( .A(net_8048), .Z(net_8049) );
NAND2_X2 inst_4102 ( .A1(net_6655), .A2(net_1655), .ZN(net_950) );
SDFF_X2 inst_1229 ( .SI(net_7223), .Q(net_7223), .D(net_3793), .SE(net_3751), .CK(net_10606) );
CLKBUF_X2 inst_10512 ( .A(net_9217), .Z(net_10474) );
CLKBUF_X2 inst_14167 ( .A(net_14128), .Z(net_14129) );
AOI222_X2 inst_7545 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1870), .A1(net_1869), .B1(net_1868), .C1(net_1867) );
CLKBUF_X2 inst_13780 ( .A(net_9411), .Z(net_13742) );
CLKBUF_X2 inst_13604 ( .A(net_13565), .Z(net_13566) );
INV_X4 inst_5219 ( .A(net_600), .ZN(net_473) );
NAND2_X4 inst_2894 ( .ZN(net_3743), .A1(net_3339), .A2(net_3338) );
NOR2_X2 inst_2358 ( .ZN(net_5306), .A2(net_4636), .A1(net_4509) );
CLKBUF_X2 inst_13139 ( .A(net_13100), .Z(net_13101) );
DFFR_X2 inst_7045 ( .QN(net_5985), .D(net_3186), .CK(net_9610), .RN(x1822) );
INV_X2 inst_5949 ( .ZN(net_1121), .A(net_127) );
OAI21_X2 inst_2125 ( .B1(net_3293), .B2(net_3087), .ZN(net_3062), .A(net_2910) );
INV_X2 inst_6085 ( .A(net_7512), .ZN(net_2176) );
CLKBUF_X2 inst_10192 ( .A(net_8790), .Z(net_10154) );
CLKBUF_X2 inst_11572 ( .A(net_10357), .Z(net_11534) );
CLKBUF_X2 inst_10549 ( .A(net_10502), .Z(net_10511) );
NAND2_X2 inst_2959 ( .ZN(net_5481), .A1(net_4932), .A2(net_4931) );
SDFF_X2 inst_599 ( .Q(net_6602), .D(net_6602), .SE(net_3830), .SI(net_3813), .CK(net_12175) );
CLKBUF_X2 inst_13906 ( .A(net_13867), .Z(net_13868) );
OAI221_X2 inst_1683 ( .A(net_2724), .ZN(net_2689), .B2(net_2417), .C2(net_2234), .C1(net_1821), .B1(net_1232) );
CLKBUF_X2 inst_10714 ( .A(net_10675), .Z(net_10676) );
NAND2_X2 inst_3865 ( .A1(net_6701), .A2(net_1497), .ZN(net_1467) );
CLKBUF_X2 inst_13382 ( .A(net_12459), .Z(net_13344) );
SDFF_X2 inst_541 ( .Q(net_7551), .D(net_7551), .SE(net_3896), .SI(net_385), .CK(net_13118) );
NAND2_X2 inst_4047 ( .A1(net_6939), .A2(net_1654), .ZN(net_1005) );
CLKBUF_X2 inst_10459 ( .A(net_10420), .Z(net_10421) );
CLKBUF_X2 inst_13910 ( .A(net_13871), .Z(net_13872) );
CLKBUF_X2 inst_13109 ( .A(net_12237), .Z(net_13071) );
SDFF_X2 inst_505 ( .SI(net_7035), .Q(net_7035), .D(net_3890), .SE(net_3777), .CK(net_8093) );
DFF_X1 inst_6366 ( .QN(net_6296), .D(net_5818), .CK(net_13792) );
SDFFR_X2 inst_1365 ( .SI(net_7742), .Q(net_7742), .D(net_4596), .SE(net_2603), .CK(net_13171), .RN(x1822) );
AOI22_X2 inst_7247 ( .B1(net_6815), .A1(net_6783), .A2(net_5316), .B2(net_5315), .ZN(net_5313) );
CLKBUF_X2 inst_9896 ( .A(net_7988), .Z(net_9858) );
CLKBUF_X2 inst_7936 ( .A(net_7897), .Z(net_7898) );
SDFF_X2 inst_198 ( .Q(net_6316), .SI(net_6315), .D(net_3691), .SE(net_392), .CK(net_13590) );
CLKBUF_X2 inst_13624 ( .A(net_13585), .Z(net_13586) );
NAND2_X2 inst_4125 ( .A2(net_1225), .ZN(net_1166), .A1(net_355) );
OR2_X4 inst_1371 ( .ZN(net_3971), .A2(net_3736), .A1(net_3227) );
CLKBUF_X2 inst_10809 ( .A(net_10770), .Z(net_10771) );
INV_X4 inst_5622 ( .A(net_7788), .ZN(net_2272) );
NAND2_X1 inst_4321 ( .ZN(net_4543), .A2(net_3870), .A1(net_1455) );
OAI221_X2 inst_1644 ( .ZN(net_5451), .B2(net_5052), .C2(net_5050), .A(net_4922), .C1(net_1149), .B1(net_874) );
DFF_X1 inst_6346 ( .QN(net_6185), .D(net_5838), .CK(net_13768) );
NAND2_X2 inst_3543 ( .ZN(net_2524), .A2(net_1980), .A1(net_1192) );
CLKBUF_X2 inst_12645 ( .A(net_12606), .Z(net_12607) );
DFF_X1 inst_6712 ( .QN(net_7328), .D(net_5356), .CK(net_10150) );
CLKBUF_X2 inst_10737 ( .A(net_10698), .Z(net_10699) );
CLKBUF_X2 inst_8946 ( .A(net_8907), .Z(net_8908) );
AOI222_X2 inst_7529 ( .A2(net_2135), .B2(net_2133), .C2(net_2131), .ZN(net_1980), .A1(net_1979), .B1(net_1978), .C1(net_1977) );
CLKBUF_X2 inst_13867 ( .A(net_10096), .Z(net_13829) );
CLKBUF_X2 inst_13333 ( .A(net_13294), .Z(net_13295) );
CLKBUF_X2 inst_11361 ( .A(net_11322), .Z(net_11323) );
CLKBUF_X2 inst_9351 ( .A(net_7952), .Z(net_9313) );
CLKBUF_X2 inst_8158 ( .A(net_7894), .Z(net_8120) );
CLKBUF_X2 inst_12423 ( .A(net_12384), .Z(net_12385) );
CLKBUF_X2 inst_10974 ( .A(net_10935), .Z(net_10936) );
NAND2_X2 inst_3461 ( .A2(net_5974), .ZN(net_2890), .A1(net_2889) );
CLKBUF_X2 inst_9754 ( .A(net_9715), .Z(net_9716) );
INV_X4 inst_4969 ( .ZN(net_1334), .A(net_699) );
NAND2_X2 inst_3511 ( .ZN(net_2556), .A2(net_2175), .A1(net_1460) );
CLKBUF_X2 inst_8546 ( .A(net_8086), .Z(net_8508) );
CLKBUF_X2 inst_8244 ( .A(net_8205), .Z(net_8206) );
INV_X4 inst_4692 ( .ZN(net_4140), .A(net_3325) );
DFF_X1 inst_6726 ( .QN(net_7359), .D(net_5330), .CK(net_10128) );
INV_X4 inst_4883 ( .A(net_3852), .ZN(net_884) );
CLKBUF_X2 inst_10487 ( .A(net_7949), .Z(net_10449) );
CLKBUF_X2 inst_10363 ( .A(net_10324), .Z(net_10325) );
CLKBUF_X2 inst_8580 ( .A(net_8541), .Z(net_8542) );
INV_X4 inst_5693 ( .A(net_6080), .ZN(net_3546) );
CLKBUF_X2 inst_9992 ( .A(net_9953), .Z(net_9954) );
AOI222_X2 inst_7538 ( .C1(net_7673), .A1(net_7641), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1888), .B1(net_1887) );
NOR4_X2 inst_2178 ( .A2(net_7754), .ZN(net_3315), .A4(net_3230), .A3(net_3208), .A1(net_2922) );
SDFF_X2 inst_263 ( .Q(net_6371), .SI(net_6370), .D(net_3711), .SE(net_392), .CK(net_14080) );
CLKBUF_X2 inst_10889 ( .A(net_10850), .Z(net_10851) );
SDFF_X2 inst_185 ( .Q(net_6269), .SI(net_6268), .D(net_3475), .SE(net_392), .CK(net_13915) );
CLKBUF_X2 inst_9498 ( .A(net_9459), .Z(net_9460) );
AOI22_X2 inst_7399 ( .A1(net_6035), .B1(net_5939), .ZN(net_2841), .A2(net_2838), .B2(net_200) );
INV_X2 inst_5953 ( .A(net_7352), .ZN(net_2000) );
SDFF_X2 inst_166 ( .Q(net_6248), .SI(net_6247), .D(net_3623), .SE(net_392), .CK(net_13973) );
DFF_X1 inst_6742 ( .QN(net_7650), .D(net_4839), .CK(net_13060) );
NAND2_X2 inst_3815 ( .A1(net_6503), .A2(net_1642), .ZN(net_1530) );
INV_X4 inst_4786 ( .A(net_2703), .ZN(net_1965) );
CLKBUF_X2 inst_13822 ( .A(net_13783), .Z(net_13784) );
CLKBUF_X2 inst_12617 ( .A(net_10932), .Z(net_12579) );
DFF_X2 inst_6307 ( .QN(net_7813), .CK(net_8438), .D(x1432) );
AOI22_X2 inst_7371 ( .A2(net_5916), .B2(net_2957), .ZN(net_2951), .B1(net_2679), .A1(net_841) );
OAI21_X2 inst_1757 ( .ZN(net_5443), .B1(net_5442), .A(net_4665), .B2(net_3993) );
NAND2_X2 inst_3851 ( .ZN(net_1485), .A2(net_1484), .A1(net_1092) );
CLKBUF_X2 inst_10650 ( .A(net_10189), .Z(net_10612) );
CLKBUF_X2 inst_10121 ( .A(net_10082), .Z(net_10083) );
DFF_X1 inst_6772 ( .QN(net_6087), .D(net_4638), .CK(net_12947) );
DFF_X1 inst_6370 ( .QN(net_6292), .D(net_5814), .CK(net_13781) );
CLKBUF_X2 inst_12358 ( .A(net_12319), .Z(net_12320) );
CLKBUF_X2 inst_11923 ( .A(net_11884), .Z(net_11885) );
DFF_X1 inst_6359 ( .Q(net_6223), .D(net_5825), .CK(net_14125) );
NAND2_X2 inst_4118 ( .A2(net_1222), .ZN(net_1073), .A1(net_335) );
CLKBUF_X2 inst_12026 ( .A(net_11987), .Z(net_11988) );
CLKBUF_X2 inst_13410 ( .A(net_13371), .Z(net_13372) );
OAI22_X2 inst_1605 ( .B2(net_3200), .A2(net_3144), .ZN(net_3129), .A1(net_3128), .B1(net_1722) );
INV_X4 inst_5440 ( .A(net_7415), .ZN(net_2186) );
INV_X4 inst_4849 ( .A(net_3855), .ZN(net_1059) );
CLKBUF_X2 inst_10206 ( .A(net_10167), .Z(net_10168) );
CLKBUF_X2 inst_11635 ( .A(net_11596), .Z(net_11597) );
CLKBUF_X2 inst_13593 ( .A(net_11093), .Z(net_13555) );
INV_X4 inst_4649 ( .ZN(net_4634), .A(net_4282) );
CLKBUF_X2 inst_12904 ( .A(net_12865), .Z(net_12866) );
CLKBUF_X2 inst_10558 ( .A(net_10112), .Z(net_10520) );
CLKBUF_X2 inst_8185 ( .A(net_8146), .Z(net_8147) );
CLKBUF_X2 inst_11223 ( .A(net_11184), .Z(net_11185) );
CLKBUF_X2 inst_12922 ( .A(net_12883), .Z(net_12884) );
INV_X4 inst_5308 ( .A(net_6957), .ZN(net_567) );
AOI22_X2 inst_7413 ( .A1(net_3855), .A2(net_3105), .B1(net_2970), .ZN(net_2822), .B2(net_254) );
CLKBUF_X2 inst_14263 ( .A(net_9533), .Z(net_14225) );
INV_X8 inst_4475 ( .ZN(net_4954), .A(net_4269) );
AOI222_X2 inst_7590 ( .A1(net_7386), .ZN(net_5412), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_349), .C2(net_347) );
CLKBUF_X2 inst_8698 ( .A(net_8659), .Z(net_8660) );
INV_X4 inst_5034 ( .A(net_7798), .ZN(net_3798) );
INV_X4 inst_4853 ( .ZN(net_1053), .A(net_1052) );
DFF_X2 inst_6322 ( .QN(net_7819), .CK(net_11036), .D(x1382) );
AOI21_X2 inst_7757 ( .B1(net_6474), .ZN(net_4041), .B2(net_2580), .A(net_2310) );
CLKBUF_X2 inst_11077 ( .A(net_11038), .Z(net_11039) );
NAND2_X2 inst_3898 ( .A1(net_6970), .A2(net_1833), .ZN(net_1416) );
INV_X4 inst_5254 ( .A(net_709), .ZN(net_436) );
INV_X4 inst_5201 ( .ZN(net_685), .A(net_499) );
NOR2_X2 inst_2373 ( .ZN(net_5212), .A2(net_4612), .A1(net_4443) );
CLKBUF_X2 inst_9370 ( .A(net_9331), .Z(net_9332) );
CLKBUF_X2 inst_11949 ( .A(net_11910), .Z(net_11911) );
CLKBUF_X2 inst_11436 ( .A(net_11397), .Z(net_11398) );
NAND2_X2 inst_3503 ( .A1(net_6401), .ZN(net_2820), .A2(net_2263) );
CLKBUF_X2 inst_13974 ( .A(net_13935), .Z(net_13936) );
CLKBUF_X2 inst_9215 ( .A(net_9176), .Z(net_9177) );
CLKBUF_X2 inst_7973 ( .A(net_7934), .Z(net_7935) );
SDFFR_X2 inst_1331 ( .SI(net_7767), .Q(net_7767), .SE(net_4259), .D(net_4258), .CK(net_12367), .RN(x1822) );
CLKBUF_X2 inst_12322 ( .A(net_10817), .Z(net_12284) );
AOI222_X2 inst_7604 ( .A1(net_7236), .ZN(net_4866), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_330), .C2(net_328) );
NAND2_X2 inst_4138 ( .A2(net_1222), .ZN(net_1175), .A1(net_338) );
XNOR2_X2 inst_52 ( .ZN(net_2251), .A(net_2250), .B(net_2249) );
AOI22_X2 inst_7404 ( .A1(net_6046), .B1(net_5939), .A2(net_2838), .ZN(net_2833), .B2(net_208) );
CLKBUF_X2 inst_12600 ( .A(net_10003), .Z(net_12562) );
SDFF_X2 inst_668 ( .Q(net_6699), .D(net_6699), .SE(net_3871), .SI(net_3798), .CK(net_8288) );
NAND2_X2 inst_3223 ( .ZN(net_4679), .A2(net_3988), .A1(net_2083) );
NAND2_X2 inst_3049 ( .A1(net_7017), .A2(net_4979), .ZN(net_4958) );
CLKBUF_X2 inst_11987 ( .A(net_11948), .Z(net_11949) );
NAND2_X2 inst_3560 ( .ZN(net_2507), .A2(net_2030), .A1(net_1792) );
NAND2_X2 inst_4159 ( .A2(net_6408), .ZN(net_1052), .A1(net_529) );
NAND3_X2 inst_2683 ( .ZN(net_3203), .A2(net_3159), .A3(net_3051), .A1(net_3001) );
CLKBUF_X2 inst_13736 ( .A(net_13697), .Z(net_13698) );
CLKBUF_X2 inst_12567 ( .A(net_12528), .Z(net_12529) );
NAND2_X1 inst_4223 ( .ZN(net_4736), .A2(net_3988), .A1(net_2188) );
NAND2_X2 inst_3349 ( .ZN(net_3549), .A1(net_3548), .A2(net_3226) );
CLKBUF_X2 inst_11444 ( .A(net_11405), .Z(net_11406) );
CLKBUF_X2 inst_14277 ( .A(net_10158), .Z(net_14239) );
CLKBUF_X2 inst_14152 ( .A(net_14113), .Z(net_14114) );
CLKBUF_X2 inst_10057 ( .A(net_10018), .Z(net_10019) );
NOR2_X2 inst_2545 ( .A2(net_6557), .ZN(net_1243), .A1(net_491) );
CLKBUF_X2 inst_8220 ( .A(net_8099), .Z(net_8182) );
CLKBUF_X2 inst_12390 ( .A(net_12351), .Z(net_12352) );
CLKBUF_X2 inst_10722 ( .A(net_10446), .Z(net_10684) );
CLKBUF_X2 inst_7999 ( .A(net_7960), .Z(net_7961) );
CLKBUF_X2 inst_13283 ( .A(net_12945), .Z(net_13245) );
CLKBUF_X2 inst_13077 ( .A(net_13038), .Z(net_13039) );
NAND3_X2 inst_2768 ( .ZN(net_2332), .A3(net_1609), .A1(net_1436), .A2(net_1004) );
DFF_X1 inst_6677 ( .QN(net_7255), .D(net_5147), .CK(net_10178) );
CLKBUF_X2 inst_9878 ( .A(net_9839), .Z(net_9840) );
OAI21_X2 inst_1835 ( .ZN(net_5340), .B1(net_5339), .A(net_4355), .B2(net_3856) );
OAI21_X2 inst_1910 ( .B1(net_5349), .ZN(net_5158), .A(net_4773), .B2(net_3941) );
CLKBUF_X2 inst_13777 ( .A(net_13738), .Z(net_13739) );
CLKBUF_X2 inst_13420 ( .A(net_13381), .Z(net_13382) );
INV_X4 inst_4639 ( .ZN(net_4183), .A(net_4025) );
CLKBUF_X2 inst_12399 ( .A(net_10356), .Z(net_12361) );
CLKBUF_X2 inst_9670 ( .A(net_9185), .Z(net_9632) );
AND3_X4 inst_7797 ( .ZN(net_2588), .A1(net_2393), .A3(net_2231), .A2(net_1707) );
SDFF_X2 inst_621 ( .Q(net_6599), .D(net_6599), .SE(net_3830), .SI(net_3814), .CK(net_9338) );
CLKBUF_X2 inst_10272 ( .A(net_10233), .Z(net_10234) );
AOI21_X2 inst_7764 ( .B1(net_6610), .ZN(net_4012), .B2(net_2583), .A(net_2283) );
CLKBUF_X2 inst_9265 ( .A(net_8954), .Z(net_9227) );
INV_X2 inst_5814 ( .A(net_1624), .ZN(net_1099) );
NAND2_X2 inst_3115 ( .A1(net_6620), .A2(net_4899), .ZN(net_4886) );
NAND4_X2 inst_2560 ( .ZN(net_3452), .A1(net_2272), .A3(net_1928), .A2(net_889), .A4(net_651) );
CLKBUF_X2 inst_10867 ( .A(net_10828), .Z(net_10829) );
NAND2_X2 inst_3219 ( .ZN(net_4707), .A2(net_3986), .A1(net_2091) );
INV_X4 inst_5673 ( .A(net_7575), .ZN(net_1909) );
CLKBUF_X2 inst_10025 ( .A(net_9986), .Z(net_9987) );
CLKBUF_X2 inst_12236 ( .A(net_12197), .Z(net_12198) );
CLKBUF_X2 inst_9651 ( .A(net_9612), .Z(net_9613) );
CLKBUF_X2 inst_14435 ( .A(net_14396), .Z(net_14397) );
OR2_X4 inst_1387 ( .ZN(net_2997), .A2(net_2735), .A1(net_1657) );
OAI21_X2 inst_1991 ( .B1(net_5778), .ZN(net_4602), .A(net_4167), .B2(net_4166) );
CLKBUF_X2 inst_13687 ( .A(net_11572), .Z(net_13649) );
NOR2_X2 inst_2365 ( .ZN(net_5285), .A2(net_4627), .A1(net_4483) );
CLKBUF_X2 inst_13054 ( .A(net_13015), .Z(net_13016) );
NAND2_X2 inst_3066 ( .A1(net_7128), .A2(net_4950), .ZN(net_4939) );
CLKBUF_X2 inst_12094 ( .A(net_12055), .Z(net_12056) );
NOR2_X4 inst_2250 ( .ZN(net_5636), .A1(net_5482), .A2(net_4442) );
AND2_X2 inst_7861 ( .ZN(net_1233), .A1(net_1232), .A2(net_1231) );
CLKBUF_X2 inst_14129 ( .A(net_14090), .Z(net_14091) );
CLKBUF_X2 inst_11630 ( .A(net_10242), .Z(net_11592) );
DFF_X1 inst_6629 ( .QN(net_7600), .D(net_5256), .CK(net_13433) );
AOI22_X2 inst_7419 ( .A1(net_2970), .ZN(net_2774), .B1(net_2772), .A2(net_237), .B2(net_163) );
NOR3_X2 inst_2187 ( .ZN(net_5946), .A2(net_3955), .A3(net_3884), .A1(net_3771) );
CLKBUF_X2 inst_13221 ( .A(net_8141), .Z(net_13183) );
CLKBUF_X2 inst_11215 ( .A(net_11176), .Z(net_11177) );
DFF_X1 inst_6771 ( .QN(net_6067), .D(net_4645), .CK(net_11604) );
INV_X2 inst_5747 ( .ZN(net_3717), .A(net_3414) );
CLKBUF_X2 inst_14323 ( .A(net_10950), .Z(net_14285) );
CLKBUF_X2 inst_8173 ( .A(net_7844), .Z(net_8135) );
AOI22_X2 inst_7448 ( .A2(net_2676), .B2(net_2673), .ZN(net_849), .A1(net_848), .B1(net_847) );
DFF_X1 inst_6640 ( .QN(net_7628), .D(net_5233), .CK(net_13075) );
INV_X4 inst_4703 ( .ZN(net_3337), .A(net_3258) );
NAND3_X2 inst_2672 ( .ZN(net_3754), .A3(net_3302), .A1(net_2962), .A2(net_2942) );
XNOR2_X2 inst_25 ( .ZN(net_2572), .B(net_2571), .A(net_2442) );
CLKBUF_X2 inst_9043 ( .A(net_9004), .Z(net_9005) );
INV_X4 inst_5239 ( .ZN(net_3004), .A(net_451) );
NAND2_X2 inst_3527 ( .ZN(net_2540), .A2(net_2108), .A1(net_1449) );
INV_X4 inst_5032 ( .A(net_3000), .ZN(net_702) );
CLKBUF_X2 inst_13924 ( .A(net_13885), .Z(net_13886) );
INV_X4 inst_5166 ( .A(net_856), .ZN(net_544) );
CLKBUF_X2 inst_13637 ( .A(net_13598), .Z(net_13599) );
CLKBUF_X2 inst_9691 ( .A(net_9652), .Z(net_9653) );
CLKBUF_X2 inst_9558 ( .A(net_9519), .Z(net_9520) );
NOR2_X2 inst_2500 ( .A1(net_3052), .ZN(net_1738), .A2(net_1737) );
CLKBUF_X2 inst_12119 ( .A(net_12080), .Z(net_12081) );
CLKBUF_X2 inst_9734 ( .A(net_9695), .Z(net_9696) );
INV_X2 inst_6045 ( .A(net_7350), .ZN(net_2215) );
NAND2_X1 inst_4395 ( .A2(net_5893), .ZN(net_3244), .A1(net_3243) );
NAND2_X2 inst_3434 ( .ZN(net_3214), .A2(net_3098), .A1(net_2763) );
CLKBUF_X2 inst_9042 ( .A(net_8704), .Z(net_9004) );
DFF_X1 inst_6408 ( .QN(net_6155), .D(net_5762), .CK(net_11917) );
NAND2_X1 inst_4296 ( .ZN(net_4570), .A2(net_3866), .A1(net_1905) );
NAND2_X2 inst_3764 ( .A1(net_7028), .A2(net_1975), .ZN(net_1581) );
CLKBUF_X2 inst_8764 ( .A(net_8725), .Z(net_8726) );
CLKBUF_X2 inst_11912 ( .A(net_9808), .Z(net_11874) );
CLKBUF_X2 inst_13101 ( .A(net_13062), .Z(net_13063) );
AOI22_X2 inst_7330 ( .A2(net_3429), .B2(net_3428), .ZN(net_3416), .B1(net_2573), .A1(net_1250) );
AOI222_X2 inst_7581 ( .A1(net_7247), .ZN(net_5357), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_341), .C2(net_339) );
NOR2_X2 inst_2340 ( .A2(net_6025), .A1(net_5778), .ZN(net_5714) );
NAND2_X2 inst_3204 ( .ZN(net_4722), .A2(net_3986), .A1(net_1865) );
CLKBUF_X2 inst_14219 ( .A(net_14180), .Z(net_14181) );
NAND2_X2 inst_3421 ( .ZN(net_3402), .A2(net_3240), .A1(net_719) );
NAND2_X1 inst_4444 ( .A2(net_2131), .ZN(net_1316), .A1(net_1315) );
CLKBUF_X2 inst_12019 ( .A(net_8858), .Z(net_11981) );
NAND3_X2 inst_2679 ( .ZN(net_3336), .A3(net_3104), .A1(net_2856), .A2(net_2773) );
XNOR2_X2 inst_16 ( .ZN(net_2637), .B(net_2636), .A(net_2479) );
DFF_X1 inst_6935 ( .Q(net_6053), .D(net_2381), .CK(net_14368) );
CLKBUF_X2 inst_14173 ( .A(net_7994), .Z(net_14135) );
NAND2_X2 inst_3949 ( .A1(net_6708), .A2(net_1497), .ZN(net_1339) );
NAND3_X2 inst_2808 ( .ZN(net_2290), .A3(net_1538), .A1(net_1324), .A2(net_988) );
SDFF_X2 inst_156 ( .Q(net_6258), .SI(net_6257), .D(net_3542), .SE(net_392), .CK(net_13997) );
INV_X4 inst_4617 ( .ZN(net_4205), .A(net_4071) );
OAI21_X2 inst_1777 ( .B1(net_5434), .ZN(net_5417), .A(net_4696), .B2(net_3989) );
DFF_X2 inst_6239 ( .QN(net_7379), .D(net_3035), .CK(net_9513) );
SDFF_X2 inst_1068 ( .SI(net_6543), .Q(net_6543), .D(net_3780), .SE(net_3755), .CK(net_11629) );
SDFF_X2 inst_886 ( .Q(net_7116), .D(net_7116), .SE(net_3888), .SI(net_3808), .CK(net_7865) );
CLKBUF_X2 inst_12799 ( .A(net_12760), .Z(net_12761) );
CLKBUF_X2 inst_11799 ( .A(net_11760), .Z(net_11761) );
NAND2_X2 inst_3442 ( .ZN(net_3165), .A2(net_3164), .A1(net_3150) );
CLKBUF_X2 inst_12509 ( .A(net_8236), .Z(net_12471) );
NAND3_X2 inst_2693 ( .ZN(net_2984), .A3(net_2897), .A2(net_2753), .A1(net_1924) );
INV_X4 inst_5350 ( .A(net_6123), .ZN(net_3687) );
CLKBUF_X2 inst_10307 ( .A(net_10268), .Z(net_10269) );
INV_X4 inst_5380 ( .A(net_6825), .ZN(net_818) );
CLKBUF_X2 inst_10936 ( .A(net_10897), .Z(net_10898) );
CLKBUF_X2 inst_13319 ( .A(net_13280), .Z(net_13281) );
DFF_X1 inst_6473 ( .QN(net_6070), .D(net_5586), .CK(net_8103) );
INV_X8 inst_4468 ( .ZN(net_5316), .A(net_4283) );
CLKBUF_X2 inst_11740 ( .A(net_11701), .Z(net_11702) );
NAND2_X2 inst_3020 ( .A1(net_6892), .A2(net_5006), .ZN(net_4989) );
OAI22_X2 inst_1549 ( .B2(net_3405), .A2(net_3360), .ZN(net_3356), .A1(net_3198), .B1(net_610) );
CLKBUF_X2 inst_12894 ( .A(net_12855), .Z(net_12856) );
CLKBUF_X2 inst_11533 ( .A(net_11494), .Z(net_11495) );
CLKBUF_X2 inst_9239 ( .A(net_9200), .Z(net_9201) );
DFF_X2 inst_6186 ( .QN(net_6690), .D(net_5091), .CK(net_9724) );
CLKBUF_X2 inst_14450 ( .A(net_14411), .Z(net_14412) );
CLKBUF_X2 inst_11484 ( .A(net_9829), .Z(net_11446) );
CLKBUF_X2 inst_11270 ( .A(net_11231), .Z(net_11232) );
CLKBUF_X2 inst_12380 ( .A(net_12341), .Z(net_12342) );
CLKBUF_X2 inst_13477 ( .A(net_13438), .Z(net_13439) );
CLKBUF_X2 inst_10576 ( .A(net_10537), .Z(net_10538) );
CLKBUF_X2 inst_8844 ( .A(net_8058), .Z(net_8806) );
OAI21_X2 inst_1969 ( .ZN(net_4869), .B1(net_4868), .A(net_4341), .B2(net_3859) );
CLKBUF_X2 inst_9113 ( .A(net_9074), .Z(net_9075) );
AND2_X4 inst_7837 ( .A2(net_1823), .ZN(net_1069), .A1(net_1068) );
NAND2_X4 inst_2881 ( .ZN(net_3927), .A1(net_3841), .A2(net_433) );
SDFF_X2 inst_821 ( .Q(net_6995), .D(net_6995), .SE(net_3891), .SI(net_3800), .CK(net_10868) );
CLKBUF_X2 inst_11382 ( .A(net_10042), .Z(net_11344) );
CLKBUF_X2 inst_8879 ( .A(net_8840), .Z(net_8841) );
CLKBUF_X2 inst_9128 ( .A(net_9089), .Z(net_9090) );
CLKBUF_X2 inst_9348 ( .A(net_9309), .Z(net_9310) );
CLKBUF_X2 inst_8183 ( .A(net_8144), .Z(net_8145) );
DFF_X1 inst_6914 ( .D(net_2413), .Q(net_241), .CK(net_13138) );
SDFF_X2 inst_980 ( .SI(net_7802), .Q(net_6433), .D(net_6433), .SE(net_3820), .CK(net_11258) );
DFF_X1 inst_6540 ( .QN(net_7472), .D(net_5576), .CK(net_10079) );
CLKBUF_X2 inst_8486 ( .A(net_8447), .Z(net_8448) );
CLKBUF_X2 inst_13136 ( .A(net_13097), .Z(net_13098) );
OAI21_X2 inst_1785 ( .B1(net_5442), .ZN(net_5406), .A(net_4680), .B2(net_3988) );
CLKBUF_X2 inst_10104 ( .A(net_10065), .Z(net_10066) );
CLKBUF_X2 inst_12939 ( .A(net_12359), .Z(net_12901) );
NAND2_X2 inst_4213 ( .ZN(net_3338), .A2(net_281), .A1(net_280) );
NAND2_X2 inst_3150 ( .ZN(net_4813), .A2(net_4153), .A1(net_2125) );
CLKBUF_X2 inst_9341 ( .A(net_9302), .Z(net_9303) );
CLKBUF_X2 inst_10761 ( .A(net_10722), .Z(net_10723) );
CLKBUF_X2 inst_9575 ( .A(net_9536), .Z(net_9537) );
CLKBUF_X2 inst_12765 ( .A(net_8128), .Z(net_12727) );
CLKBUF_X2 inst_12118 ( .A(net_12079), .Z(net_12080) );
CLKBUF_X2 inst_10694 ( .A(net_10655), .Z(net_10656) );
CLKBUF_X2 inst_8522 ( .A(net_8215), .Z(net_8484) );
INV_X2 inst_6022 ( .A(net_7318), .ZN(net_1759) );
NOR2_X4 inst_2286 ( .ZN(net_5891), .A2(net_5873), .A1(net_3018) );
DFF_X2 inst_6216 ( .QN(net_7532), .D(net_3981), .CK(net_12598) );
INV_X2 inst_5791 ( .A(net_5977), .ZN(net_2237) );
SDFF_X2 inst_866 ( .SI(net_7052), .Q(net_7052), .D(net_3779), .SE(net_3777), .CK(net_9016) );
AOI222_X2 inst_7512 ( .B1(net_7371), .C1(net_7307), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2030), .A1(net_2029) );
OAI21_X2 inst_2137 ( .ZN(net_2813), .A(net_518), .B1(net_190), .B2(net_188) );
CLKBUF_X2 inst_11061 ( .A(net_9226), .Z(net_11023) );
CLKBUF_X2 inst_9406 ( .A(net_9367), .Z(net_9368) );
OAI22_X2 inst_1439 ( .B1(net_5850), .ZN(net_5684), .A2(net_5494), .B2(net_5493), .A1(net_5253) );
NAND2_X2 inst_3640 ( .ZN(net_1943), .A1(net_1294), .A2(net_1112) );
DFFR_X2 inst_7107 ( .D(net_1947), .QN(net_129), .CK(net_9584), .RN(x1822) );
CLKBUF_X2 inst_12367 ( .A(net_12328), .Z(net_12329) );
CLKBUF_X2 inst_8444 ( .A(net_8405), .Z(net_8406) );
INV_X4 inst_5604 ( .A(net_6405), .ZN(net_460) );
SDFF_X2 inst_248 ( .Q(net_6346), .SI(net_6345), .D(net_3583), .SE(net_392), .CK(net_13653) );
OAI22_X2 inst_1613 ( .A1(net_3282), .A2(net_3087), .B2(net_3084), .ZN(net_3059), .B1(net_743) );
NAND2_X2 inst_3107 ( .A1(net_6616), .A2(net_4899), .ZN(net_4894) );
DFF_X1 inst_6624 ( .QN(net_7594), .D(net_5263), .CK(net_10580) );
OAI21_X2 inst_1919 ( .B1(net_5337), .ZN(net_5144), .A(net_4768), .B2(net_3941) );
INV_X4 inst_5659 ( .A(net_6011), .ZN(net_592) );
INV_X2 inst_5965 ( .A(net_7441), .ZN(net_1327) );
CLKBUF_X2 inst_12222 ( .A(net_12183), .Z(net_12184) );
SDFF_X2 inst_1141 ( .SI(net_6800), .Q(net_6800), .D(net_3894), .SE(net_3729), .CK(net_11074) );
NAND2_X2 inst_3589 ( .ZN(net_2411), .A2(net_1908), .A1(net_1466) );
NOR2_X2 inst_2488 ( .ZN(net_2628), .A2(net_2616), .A1(net_624) );
CLKBUF_X2 inst_10528 ( .A(net_9677), .Z(net_10490) );
SDFF_X2 inst_932 ( .SI(net_7174), .Q(net_7174), .SE(net_3819), .D(net_3813), .CK(net_12154) );
CLKBUF_X2 inst_12891 ( .A(net_12852), .Z(net_12853) );
SDFF_X2 inst_180 ( .Q(net_6274), .SI(net_6273), .D(net_3507), .SE(net_392), .CK(net_13927) );
CLKBUF_X2 inst_13472 ( .A(net_12832), .Z(net_13434) );
OAI21_X2 inst_1960 ( .B1(net_5198), .ZN(net_5060), .A(net_4705), .B2(net_3986) );
CLKBUF_X2 inst_9057 ( .A(net_8439), .Z(net_9019) );
CLKBUF_X2 inst_8003 ( .A(net_7964), .Z(net_7965) );
CLKBUF_X2 inst_11995 ( .A(net_8415), .Z(net_11957) );
CLKBUF_X2 inst_8475 ( .A(net_8436), .Z(net_8437) );
CLKBUF_X2 inst_8712 ( .A(net_8673), .Z(net_8674) );
DFF_X1 inst_6455 ( .QN(net_6108), .D(net_5604), .CK(net_11182) );
CLKBUF_X2 inst_13273 ( .A(net_13234), .Z(net_13235) );
CLKBUF_X2 inst_12635 ( .A(net_12596), .Z(net_12597) );
CLKBUF_X2 inst_11886 ( .A(net_11847), .Z(net_11848) );
CLKBUF_X2 inst_10283 ( .A(net_10244), .Z(net_10245) );
CLKBUF_X2 inst_10659 ( .A(net_10620), .Z(net_10621) );
CLKBUF_X2 inst_12654 ( .A(net_12615), .Z(net_12616) );
CLKBUF_X2 inst_10744 ( .A(net_9005), .Z(net_10706) );
INV_X4 inst_4636 ( .ZN(net_4186), .A(net_4034) );
SDFF_X2 inst_302 ( .SI(net_7520), .Q(net_7520), .D(net_5104), .SE(net_3988), .CK(net_12073) );
CLKBUF_X2 inst_13527 ( .A(net_13488), .Z(net_13489) );
CLKBUF_X2 inst_10318 ( .A(net_8745), .Z(net_10280) );
SDFF_X2 inst_673 ( .Q(net_6737), .D(net_6737), .SE(net_3815), .SI(net_3813), .CK(net_8286) );
NAND2_X2 inst_3585 ( .ZN(net_2598), .A2(net_2417), .A1(net_1824) );
NAND2_X2 inst_3287 ( .ZN(net_3672), .A1(net_3671), .A2(net_3231) );
CLKBUF_X2 inst_11628 ( .A(net_11589), .Z(net_11590) );
INV_X2 inst_5892 ( .A(net_7292), .ZN(net_2065) );
SDFF_X2 inst_211 ( .Q(net_6303), .SI(net_6302), .D(net_3683), .SE(net_392), .CK(net_13551) );
SDFF_X2 inst_1151 ( .SI(net_6812), .Q(net_6812), .D(net_3804), .SE(net_3722), .CK(net_11132) );
CLKBUF_X2 inst_11399 ( .A(net_10579), .Z(net_11361) );
INV_X4 inst_4659 ( .ZN(net_5882), .A(net_3927) );
NAND2_X2 inst_3120 ( .A1(net_6590), .A2(net_4897), .ZN(net_4881) );
INV_X2 inst_5917 ( .A(net_7472), .ZN(net_2106) );
INV_X2 inst_5735 ( .ZN(net_5887), .A(net_4139) );
SDFF_X2 inst_561 ( .SI(net_7188), .Q(net_7188), .D(net_3902), .SE(net_3817), .CK(net_8726) );
CLKBUF_X2 inst_13417 ( .A(net_10653), .Z(net_13379) );
CLKBUF_X2 inst_11565 ( .A(net_11526), .Z(net_11527) );
CLKBUF_X2 inst_12999 ( .A(net_11747), .Z(net_12961) );
CLKBUF_X2 inst_10903 ( .A(net_10724), .Z(net_10865) );
NOR2_X2 inst_2505 ( .ZN(net_1239), .A2(net_673), .A1(net_632) );
DFF_X1 inst_6504 ( .QN(net_7426), .D(net_5523), .CK(net_9817) );
CLKBUF_X2 inst_12253 ( .A(net_8085), .Z(net_12215) );
OAI221_X2 inst_1641 ( .ZN(net_5454), .B2(net_5087), .C2(net_5085), .A(net_5010), .C1(net_1150), .B1(net_741) );
CLKBUF_X2 inst_12806 ( .A(net_9995), .Z(net_12768) );
DFF_X1 inst_6945 ( .Q(net_7790), .D(net_1681), .CK(net_14349) );
DFF_X1 inst_6765 ( .QN(net_6107), .D(net_4667), .CK(net_11128) );
NAND3_X2 inst_2736 ( .ZN(net_2365), .A3(net_1559), .A1(net_1276), .A2(net_998) );
CLKBUF_X2 inst_12524 ( .A(net_12485), .Z(net_12486) );
CLKBUF_X2 inst_11749 ( .A(net_11710), .Z(net_11711) );
AOI21_X2 inst_7636 ( .ZN(net_3954), .B2(net_3766), .B1(net_2884), .A(net_925) );
SDFF_X2 inst_196 ( .Q(net_6318), .SI(net_6317), .D(net_3689), .SE(net_392), .CK(net_13593) );
OAI22_X2 inst_1567 ( .A2(net_3297), .B2(net_3286), .ZN(net_3284), .A1(net_3139), .B1(net_738) );
NAND2_X2 inst_3451 ( .A2(net_5925), .ZN(net_2921), .A1(net_1830) );
INV_X8 inst_4489 ( .ZN(net_4855), .A(net_3410) );
NOR2_X2 inst_2417 ( .ZN(net_3470), .A2(net_3392), .A1(net_2804) );
INV_X4 inst_5523 ( .A(net_7577), .ZN(net_1887) );
CLKBUF_X2 inst_13481 ( .A(net_10845), .Z(net_13443) );
CLKBUF_X2 inst_12828 ( .A(net_12789), .Z(net_12790) );
CLKBUF_X2 inst_10637 ( .A(net_10598), .Z(net_10599) );
CLKBUF_X2 inst_8405 ( .A(net_7904), .Z(net_8367) );
OR2_X2 inst_1403 ( .ZN(net_3184), .A2(net_3183), .A1(net_2996) );
INV_X4 inst_5606 ( .A(net_7718), .ZN(net_856) );
CLKBUF_X2 inst_14371 ( .A(net_12780), .Z(net_14333) );
SDFF_X2 inst_298 ( .D(net_6394), .SE(net_6052), .SI(net_319), .Q(net_319), .CK(net_13743) );
NOR4_X2 inst_2180 ( .A2(net_7758), .ZN(net_3311), .A4(net_3227), .A3(net_3208), .A1(net_2920) );
OAI21_X2 inst_1856 ( .ZN(net_5262), .B1(net_5235), .A(net_4547), .B2(net_3870) );
CLKBUF_X2 inst_9379 ( .A(net_9340), .Z(net_9341) );
INV_X4 inst_5507 ( .A(net_6178), .ZN(net_3521) );
XNOR2_X2 inst_42 ( .B(net_6825), .ZN(net_2449), .A(net_1242) );
DFF_X1 inst_6594 ( .QN(net_7483), .D(net_5039), .CK(net_9659) );
CLKBUF_X2 inst_13535 ( .A(net_13496), .Z(net_13497) );
CLKBUF_X2 inst_10521 ( .A(net_10482), .Z(net_10483) );
NAND2_X2 inst_4084 ( .A1(net_6525), .A2(net_1645), .ZN(net_968) );
OAI22_X2 inst_1479 ( .B1(net_4855), .B2(net_4477), .A1(net_4228), .ZN(net_4212), .A2(net_4211) );
CLKBUF_X2 inst_11390 ( .A(net_11351), .Z(net_11352) );
CLKBUF_X2 inst_11124 ( .A(net_8941), .Z(net_11086) );
DFF_X2 inst_6180 ( .QN(net_7093), .D(net_5452), .CK(net_9383) );
NAND2_X2 inst_3529 ( .ZN(net_2538), .A2(net_2221), .A1(net_1366) );
OAI21_X2 inst_2040 ( .B1(net_4619), .B2(net_4476), .ZN(net_4463), .A(net_3620) );
SDFF_X2 inst_437 ( .Q(net_7391), .D(net_7391), .SE(net_3994), .SI(net_356), .CK(net_12066) );
CLKBUF_X2 inst_10834 ( .A(net_10795), .Z(net_10796) );
CLKBUF_X2 inst_11606 ( .A(net_8557), .Z(net_11568) );
CLKBUF_X2 inst_13307 ( .A(net_13268), .Z(net_13269) );
AOI22_X2 inst_7327 ( .ZN(net_3421), .A2(net_3420), .B2(net_3419), .A1(net_1301), .B1(net_907) );
INV_X4 inst_4742 ( .ZN(net_2747), .A(net_2746) );
CLKBUF_X2 inst_8316 ( .A(net_8277), .Z(net_8278) );
DFF_X1 inst_6527 ( .QN(net_7465), .D(net_5424), .CK(net_9813) );
CLKBUF_X2 inst_14391 ( .A(net_14352), .Z(net_14353) );
CLKBUF_X2 inst_12782 ( .A(net_12743), .Z(net_12744) );
CLKBUF_X2 inst_10451 ( .A(net_10412), .Z(net_10413) );
CLKBUF_X2 inst_9425 ( .A(net_8285), .Z(net_9387) );
INV_X2 inst_6099 ( .A(net_7508), .ZN(net_2201) );
OAI21_X2 inst_1706 ( .B2(net_5910), .ZN(net_5588), .A(net_5161), .B1(net_4057) );
CLKBUF_X2 inst_12687 ( .A(net_7947), .Z(net_12649) );
DFF_X1 inst_6733 ( .QN(net_7352), .D(net_5322), .CK(net_12978) );
INV_X8 inst_4561 ( .A(net_3338), .ZN(net_1225) );
CLKBUF_X2 inst_11315 ( .A(net_11276), .Z(net_11277) );
CLKBUF_X2 inst_9324 ( .A(net_9285), .Z(net_9286) );
DFF_X1 inst_6778 ( .QN(net_6125), .D(net_4323), .CK(net_11828) );
CLKBUF_X2 inst_9611 ( .A(net_9572), .Z(net_9573) );
DFF_X2 inst_6221 ( .QN(net_6827), .D(net_3727), .CK(net_10790) );
NOR2_X4 inst_2220 ( .ZN(net_5678), .A1(net_5556), .A2(net_4515) );
NAND3_X2 inst_2743 ( .ZN(net_2358), .A3(net_1557), .A1(net_1505), .A2(net_961) );
OAI21_X2 inst_2083 ( .B2(net_4415), .ZN(net_4407), .B1(net_4020), .A(net_3498) );
OAI22_X2 inst_1470 ( .B1(net_4855), .ZN(net_4232), .A2(net_4231), .B2(net_4230), .A1(net_4228) );
CLKBUF_X2 inst_9958 ( .A(net_7917), .Z(net_9920) );
CLKBUF_X2 inst_8019 ( .A(net_7980), .Z(net_7981) );
NOR2_X4 inst_2247 ( .ZN(net_5639), .A1(net_5485), .A2(net_4451) );
SDFF_X2 inst_1213 ( .D(net_7799), .SI(net_7201), .Q(net_7201), .SE(net_3750), .CK(net_8691) );
CLKBUF_X2 inst_13517 ( .A(net_13478), .Z(net_13479) );
CLKBUF_X2 inst_9706 ( .A(net_9667), .Z(net_9668) );
NAND2_X2 inst_3072 ( .A1(net_7119), .A2(net_4950), .ZN(net_4933) );
AOI222_X2 inst_7524 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_1994), .A1(net_1993), .B1(net_1992), .C1(net_1991) );
CLKBUF_X2 inst_12128 ( .A(net_12089), .Z(net_12090) );
CLKBUF_X2 inst_11852 ( .A(net_10949), .Z(net_11814) );
CLKBUF_X2 inst_14094 ( .A(net_14055), .Z(net_14056) );
NOR2_X2 inst_2452 ( .ZN(net_2818), .A2(net_2695), .A1(net_1139) );
CLKBUF_X2 inst_11370 ( .A(net_11331), .Z(net_11332) );
SDFF_X2 inst_428 ( .SI(net_7754), .Q(net_7754), .SE(net_5925), .D(net_3911), .CK(net_10391) );
CLKBUF_X2 inst_11821 ( .A(net_11782), .Z(net_11783) );
INV_X2 inst_5786 ( .ZN(net_2439), .A(net_2438) );
NAND2_X2 inst_3418 ( .A2(net_5890), .ZN(net_3331), .A1(net_619) );
NAND2_X2 inst_3334 ( .ZN(net_3578), .A1(net_3577), .A2(net_3226) );
SDFF_X2 inst_407 ( .SI(net_7371), .Q(net_7371), .D(net_4875), .SE(net_3853), .CK(net_9898) );
CLKBUF_X2 inst_9093 ( .A(net_8566), .Z(net_9055) );
NAND2_X2 inst_3558 ( .ZN(net_2509), .A2(net_2159), .A1(net_1784) );
SDFF_X2 inst_1208 ( .SI(net_7063), .Q(net_7063), .D(net_3892), .SE(net_3747), .CK(net_9059) );
XNOR2_X2 inst_97 ( .ZN(net_2260), .A(net_1148), .B(net_1147) );
INV_X2 inst_5843 ( .A(net_1152), .ZN(net_746) );
SDFF_X2 inst_775 ( .SI(net_6893), .Q(net_6893), .D(net_3792), .SE(net_3781), .CK(net_8930) );
CLKBUF_X2 inst_8120 ( .A(net_8052), .Z(net_8082) );
INV_X4 inst_4652 ( .ZN(net_4610), .A(net_4274) );
SDFF_X2 inst_652 ( .Q(net_6709), .D(net_6709), .SE(net_3871), .SI(net_3810), .CK(net_8526) );
AOI21_X2 inst_7642 ( .B1(net_5917), .ZN(net_3912), .B2(net_3911), .A(net_2596) );
CLKBUF_X2 inst_11102 ( .A(net_11063), .Z(net_11064) );
CLKBUF_X2 inst_9935 ( .A(net_9896), .Z(net_9897) );
CLKBUF_X2 inst_11812 ( .A(net_11773), .Z(net_11774) );
CLKBUF_X2 inst_14281 ( .A(net_11753), .Z(net_14243) );
SDFF_X2 inst_677 ( .Q(net_6741), .D(net_6741), .SE(net_3815), .SI(net_3787), .CK(net_11347) );
CLKBUF_X2 inst_12155 ( .A(net_12011), .Z(net_12117) );
SDFF_X2 inst_130 ( .Q(net_6191), .SI(net_6190), .D(net_3917), .SE(net_392), .CK(net_13631) );
OAI22_X2 inst_1566 ( .A2(net_3297), .B2(net_3286), .ZN(net_3285), .A1(net_3133), .B1(net_764) );
CLKBUF_X2 inst_12468 ( .A(net_12429), .Z(net_12430) );
CLKBUF_X2 inst_10829 ( .A(net_10192), .Z(net_10791) );
AOI21_X2 inst_7711 ( .B1(net_6875), .ZN(net_4097), .B2(net_2579), .A(net_2350) );
NOR2_X4 inst_2242 ( .ZN(net_5644), .A1(net_5490), .A2(net_4456) );
CLKBUF_X2 inst_10489 ( .A(net_10450), .Z(net_10451) );
SDFF_X2 inst_1054 ( .Q(net_7003), .D(net_7003), .SE(net_3899), .SI(net_3890), .CK(net_11861) );
CLKBUF_X2 inst_11420 ( .A(net_11381), .Z(net_11382) );
CLKBUF_X2 inst_12954 ( .A(net_10820), .Z(net_12916) );
SDFF_X2 inst_972 ( .Q(net_6452), .D(net_6452), .SE(net_3820), .SI(net_3788), .CK(net_10847) );
OAI221_X2 inst_1671 ( .ZN(net_4299), .B2(net_4157), .C2(net_4154), .A(net_3929), .B1(net_815), .C1(net_814) );
CLKBUF_X2 inst_13992 ( .A(net_8958), .Z(net_13954) );
OAI21_X2 inst_1843 ( .B1(net_5355), .ZN(net_5329), .A(net_4369), .B2(net_3853) );
INV_X4 inst_4581 ( .A(net_5084), .ZN(net_4331) );
CLKBUF_X2 inst_10044 ( .A(net_9132), .Z(net_10006) );
CLKBUF_X2 inst_13203 ( .A(net_13164), .Z(net_13165) );
CLKBUF_X2 inst_11113 ( .A(net_8314), .Z(net_11075) );
NAND2_X4 inst_2884 ( .ZN(net_3924), .A1(net_3843), .A2(net_502) );
SDFF_X2 inst_600 ( .Q(net_6603), .D(net_6603), .SE(net_3830), .SI(net_3812), .CK(net_9175) );
CLKBUF_X2 inst_13662 ( .A(net_13623), .Z(net_13624) );
CLKBUF_X2 inst_11951 ( .A(net_8983), .Z(net_11913) );
CLKBUF_X2 inst_10224 ( .A(net_10185), .Z(net_10186) );
INV_X4 inst_5319 ( .A(net_7568), .ZN(net_1855) );
INV_X8 inst_4498 ( .ZN(net_3850), .A(net_3264) );
SDFF_X2 inst_1194 ( .SI(net_7076), .Q(net_7076), .D(net_3785), .SE(net_3742), .CK(net_11855) );
CLKBUF_X2 inst_11480 ( .A(net_11441), .Z(net_11442) );
CLKBUF_X2 inst_12717 ( .A(net_12678), .Z(net_12679) );
CLKBUF_X2 inst_14292 ( .A(net_14253), .Z(net_14254) );
SDFF_X2 inst_204 ( .Q(net_6310), .SI(net_6309), .D(net_3701), .SE(net_392), .CK(net_13568) );
XNOR2_X2 inst_49 ( .ZN(net_2258), .A(net_2257), .B(net_2256) );
OAI22_X2 inst_1550 ( .B2(net_3405), .A2(net_3360), .ZN(net_3355), .A1(net_3277), .B1(net_420) );
CLKBUF_X2 inst_14353 ( .A(net_12243), .Z(net_14315) );
CLKBUF_X2 inst_14288 ( .A(net_14249), .Z(net_14250) );
SDFF_X2 inst_910 ( .Q(net_7147), .D(net_7147), .SE(net_3903), .SI(net_3809), .CK(net_11583) );
NAND2_X2 inst_4097 ( .A1(net_6528), .A2(net_1645), .ZN(net_955) );
SDFF_X2 inst_693 ( .Q(net_6730), .D(net_6730), .SE(net_3815), .SI(net_3799), .CK(net_11098) );
AOI222_X2 inst_7586 ( .A1(net_7234), .ZN(net_5365), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_328), .C2(net_326) );
CLKBUF_X2 inst_10134 ( .A(net_10095), .Z(net_10096) );
CLKBUF_X2 inst_13080 ( .A(net_13041), .Z(net_13042) );
CLKBUF_X2 inst_8772 ( .A(net_8733), .Z(net_8734) );
CLKBUF_X2 inst_12494 ( .A(net_8753), .Z(net_12456) );
AOI222_X2 inst_7562 ( .A1(net_7242), .ZN(net_5337), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_336), .C2(net_334) );
CLKBUF_X2 inst_12344 ( .A(net_12305), .Z(net_12306) );
CLKBUF_X2 inst_11515 ( .A(net_11476), .Z(net_11477) );
CLKBUF_X2 inst_10119 ( .A(net_9555), .Z(net_10081) );
CLKBUF_X2 inst_8920 ( .A(net_8881), .Z(net_8882) );
DFF_X2 inst_6217 ( .QN(net_7683), .D(net_3860), .CK(net_10792) );
AOI22_X2 inst_7383 ( .A2(net_5916), .B2(net_2957), .ZN(net_2937), .B1(net_2667), .A1(net_856) );
AOI22_X2 inst_7401 ( .B1(net_5939), .A2(net_2838), .ZN(net_2837), .A1(net_479), .B2(net_203) );
SDFF_X2 inst_937 ( .SI(net_7179), .Q(net_7179), .SE(net_3817), .D(net_3785), .CK(net_7909) );
AOI22_X2 inst_7390 ( .B1(net_5939), .A2(net_5916), .ZN(net_2929), .A1(net_838), .B2(net_194) );
CLKBUF_X2 inst_8303 ( .A(net_8264), .Z(net_8265) );
SDFF_X2 inst_908 ( .Q(net_7144), .D(net_7144), .SE(net_3903), .SI(net_3811), .CK(net_7857) );
SDFF_X2 inst_355 ( .SI(net_7613), .Q(net_7613), .D(net_4802), .SE(net_3870), .CK(net_10279) );
CLKBUF_X2 inst_11690 ( .A(net_10560), .Z(net_11652) );
CLKBUF_X2 inst_13731 ( .A(net_13044), .Z(net_13693) );
CLKBUF_X2 inst_9259 ( .A(net_8727), .Z(net_9221) );
CLKBUF_X2 inst_9227 ( .A(net_8434), .Z(net_9189) );
SDFF_X2 inst_218 ( .Q(net_6336), .SI(net_6335), .D(net_3653), .SE(net_392), .CK(net_14057) );
DFF_X1 inst_6584 ( .QN(net_7554), .D(net_5066), .CK(net_10313) );
NAND2_X2 inst_3647 ( .A1(net_7064), .ZN(net_1816), .A2(net_791) );
NAND2_X2 inst_3498 ( .ZN(net_2620), .A2(net_2424), .A1(net_653) );
DFF_X1 inst_6753 ( .QN(net_7649), .D(net_4840), .CK(net_10288) );
CLKBUF_X2 inst_11865 ( .A(net_9305), .Z(net_11827) );
CLKBUF_X2 inst_11098 ( .A(net_11059), .Z(net_11060) );
CLKBUF_X2 inst_8226 ( .A(net_8102), .Z(net_8188) );
CLKBUF_X2 inst_10706 ( .A(net_10667), .Z(net_10668) );
DFF_X2 inst_6228 ( .QN(net_6963), .D(net_3719), .CK(net_8569) );
NAND2_X2 inst_3693 ( .A2(net_1798), .ZN(net_1750), .A1(net_1749) );
CLKBUF_X2 inst_11309 ( .A(net_10558), .Z(net_11271) );
AOI21_X2 inst_7655 ( .B2(net_3439), .ZN(net_3390), .A(net_3216), .B1(net_755) );
DFF_X1 inst_6806 ( .D(net_3459), .CK(net_10421), .Q(x397) );
NAND2_X2 inst_3769 ( .A1(net_7171), .A2(net_1637), .ZN(net_1576) );
NAND2_X2 inst_4053 ( .A1(net_6792), .A2(net_1651), .ZN(net_999) );
OAI21_X2 inst_1747 ( .ZN(net_5521), .A(net_4820), .B2(net_4153), .B1(net_1074) );
INV_X4 inst_5236 ( .A(net_839), .ZN(net_455) );
CLKBUF_X2 inst_10477 ( .A(net_10044), .Z(net_10439) );
CLKBUF_X2 inst_9066 ( .A(net_9027), .Z(net_9028) );
INV_X4 inst_5109 ( .A(net_7814), .ZN(net_3836) );
CLKBUF_X2 inst_11834 ( .A(net_8698), .Z(net_11796) );
INV_X4 inst_5357 ( .A(net_6086), .ZN(net_3489) );
CLKBUF_X2 inst_12992 ( .A(net_9054), .Z(net_12954) );
CLKBUF_X2 inst_11978 ( .A(net_11939), .Z(net_11940) );
CLKBUF_X2 inst_14204 ( .A(net_14165), .Z(net_14166) );
CLKBUF_X2 inst_13026 ( .A(net_12987), .Z(net_12988) );
CLKBUF_X2 inst_13352 ( .A(net_9962), .Z(net_13314) );
NAND2_X2 inst_3917 ( .ZN(net_1387), .A2(net_1386), .A1(net_1079) );
CLKBUF_X2 inst_14104 ( .A(net_11026), .Z(net_14066) );
CLKBUF_X2 inst_13243 ( .A(net_13204), .Z(net_13205) );
CLKBUF_X2 inst_9467 ( .A(net_8494), .Z(net_9429) );
CLKBUF_X2 inst_9419 ( .A(net_9380), .Z(net_9381) );
AOI222_X2 inst_7601 ( .A1(net_7238), .ZN(net_5345), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_332), .C2(net_330) );
CLKBUF_X2 inst_12231 ( .A(net_12192), .Z(net_12193) );
NAND3_X2 inst_2682 ( .ZN(net_3204), .A2(net_2937), .A3(net_2844), .A1(net_2776) );
NAND3_X2 inst_2574 ( .ZN(net_5765), .A1(net_5660), .A2(net_5284), .A3(net_4234) );
CLKBUF_X2 inst_8517 ( .A(net_8478), .Z(net_8479) );
CLKBUF_X2 inst_12434 ( .A(net_12395), .Z(net_12396) );
INV_X4 inst_4699 ( .A(net_5976), .ZN(net_3364) );
NOR2_X4 inst_2229 ( .ZN(net_5669), .A1(net_5531), .A2(net_4499) );
CLKBUF_X2 inst_10023 ( .A(net_9984), .Z(net_9985) );
CLKBUF_X2 inst_11456 ( .A(net_11417), .Z(net_11418) );
DFF_X2 inst_6252 ( .QN(net_7763), .D(net_3057), .CK(net_9504) );
INV_X4 inst_4749 ( .ZN(net_2631), .A(net_226) );
SDFF_X2 inst_964 ( .Q(net_6443), .D(net_6443), .SE(net_3820), .SI(net_3807), .CK(net_8856) );
NAND2_X2 inst_3372 ( .ZN(net_3502), .A1(net_3501), .A2(net_3223) );
SDFF_X2 inst_1245 ( .SI(net_6540), .Q(net_6540), .D(net_3805), .SE(net_3756), .CK(net_8400) );
CLKBUF_X2 inst_7940 ( .A(net_7901), .Z(net_7902) );
CLKBUF_X2 inst_10165 ( .A(net_10126), .Z(net_10127) );
NOR2_X2 inst_2313 ( .A2(net_6201), .A1(net_5843), .ZN(net_5828) );
CLKBUF_X2 inst_12560 ( .A(net_8493), .Z(net_12522) );
DFF_X1 inst_6422 ( .QN(net_6177), .D(net_5748), .CK(net_8744) );
CLKBUF_X2 inst_10649 ( .A(net_10610), .Z(net_10611) );
CLKBUF_X2 inst_12660 ( .A(net_11622), .Z(net_12622) );
INV_X4 inst_5409 ( .A(net_7682), .ZN(net_1199) );
NAND2_X2 inst_3788 ( .A1(net_7164), .A2(net_1637), .ZN(net_1557) );
CLKBUF_X2 inst_12629 ( .A(net_12590), .Z(net_12591) );
CLKBUF_X2 inst_14030 ( .A(net_13991), .Z(net_13992) );
CLKBUF_X2 inst_12965 ( .A(net_12926), .Z(net_12927) );
INV_X2 inst_6114 ( .ZN(net_5929), .A(net_5925) );
NAND2_X2 inst_3663 ( .ZN(net_1800), .A1(net_1799), .A2(net_1798) );
CLKBUF_X2 inst_11977 ( .A(net_11938), .Z(net_11939) );
DFF_X2 inst_6193 ( .QN(net_7229), .D(net_5053), .CK(net_9371) );
NAND2_X2 inst_3001 ( .ZN(net_5010), .A2(net_4331), .A1(net_2257) );
CLKBUF_X2 inst_14111 ( .A(net_14072), .Z(net_14073) );
CLKBUF_X2 inst_13741 ( .A(net_13702), .Z(net_13703) );
NAND3_X2 inst_2818 ( .ZN(net_2280), .A3(net_1604), .A1(net_1404), .A2(net_941) );
NAND2_X2 inst_3008 ( .A1(net_6886), .A2(net_5006), .ZN(net_5001) );
INV_X4 inst_5515 ( .A(net_7268), .ZN(net_2047) );
NAND2_X2 inst_3198 ( .ZN(net_4728), .A2(net_3986), .A1(net_1855) );
INV_X2 inst_5900 ( .A(net_5994), .ZN(net_2601) );
CLKBUF_X2 inst_8234 ( .A(net_8195), .Z(net_8196) );
CLKBUF_X2 inst_7979 ( .A(net_7940), .Z(net_7941) );
NAND2_X4 inst_2904 ( .A2(net_2916), .ZN(net_2711), .A1(net_2626) );
CLKBUF_X2 inst_10075 ( .A(net_10036), .Z(net_10037) );
NOR2_X2 inst_2383 ( .A1(net_5778), .ZN(net_4597), .A2(net_4170) );
OAI21_X2 inst_1701 ( .ZN(net_5593), .A(net_5267), .B2(net_4477), .B1(net_4228) );
CLKBUF_X2 inst_12853 ( .A(net_12814), .Z(net_12815) );
CLKBUF_X2 inst_10640 ( .A(net_8726), .Z(net_10602) );
CLKBUF_X2 inst_13853 ( .A(net_13814), .Z(net_13815) );
CLKBUF_X2 inst_10401 ( .A(net_9926), .Z(net_10363) );
CLKBUF_X2 inst_13614 ( .A(net_12326), .Z(net_13576) );
CLKBUF_X2 inst_8738 ( .A(net_8584), .Z(net_8700) );
NAND2_X2 inst_4071 ( .A1(net_6806), .A2(net_1651), .ZN(net_981) );
CLKBUF_X2 inst_13577 ( .A(net_8698), .Z(net_13539) );
CLKBUF_X2 inst_11363 ( .A(net_11324), .Z(net_11325) );
INV_X4 inst_4987 ( .ZN(net_745), .A(net_703) );
CLKBUF_X2 inst_8249 ( .A(net_8210), .Z(net_8211) );
CLKBUF_X2 inst_9667 ( .A(net_8656), .Z(net_9629) );
NOR2_X2 inst_2469 ( .A2(net_5778), .ZN(net_2669), .A1(net_418) );
CLKBUF_X2 inst_12262 ( .A(net_8247), .Z(net_12224) );
CLKBUF_X2 inst_9287 ( .A(net_9248), .Z(net_9249) );
CLKBUF_X2 inst_7868 ( .A(net_7829), .Z(net_7830) );
CLKBUF_X2 inst_9838 ( .A(net_9799), .Z(net_9800) );
CLKBUF_X2 inst_9627 ( .A(net_9588), .Z(net_9589) );
CLKBUF_X2 inst_9163 ( .A(net_8050), .Z(net_9125) );
CLKBUF_X2 inst_13405 ( .A(net_13366), .Z(net_13367) );
CLKBUF_X2 inst_8593 ( .A(net_8554), .Z(net_8555) );
CLKBUF_X2 inst_13230 ( .A(net_8849), .Z(net_13192) );
INV_X4 inst_4736 ( .A(net_5962), .ZN(net_3878) );
CLKBUF_X2 inst_14442 ( .A(net_14403), .Z(net_14404) );
CLKBUF_X2 inst_12503 ( .A(net_12464), .Z(net_12465) );
CLKBUF_X2 inst_8437 ( .A(net_8398), .Z(net_8399) );
CLKBUF_X2 inst_9671 ( .A(net_9197), .Z(net_9633) );
SDFF_X2 inst_1135 ( .SI(net_6658), .Q(net_6658), .D(net_3892), .SE(net_3471), .CK(net_10043) );
DFF_X2 inst_6259 ( .QN(net_5963), .D(net_2736), .CK(net_10728) );
CLKBUF_X2 inst_10330 ( .A(net_10291), .Z(net_10292) );
DFFR_X2 inst_6983 ( .QN(net_6016), .D(net_3446), .CK(net_11445), .RN(x1822) );
NAND2_X2 inst_3715 ( .A1(net_6500), .A2(net_1642), .ZN(net_1631) );
CLKBUF_X2 inst_10929 ( .A(net_10890), .Z(net_10891) );
CLKBUF_X2 inst_8333 ( .A(net_8294), .Z(net_8295) );
CLKBUF_X2 inst_11871 ( .A(net_11832), .Z(net_11833) );
CLKBUF_X2 inst_14419 ( .A(net_11223), .Z(net_14381) );
NAND2_X2 inst_3127 ( .ZN(net_4836), .A2(net_4153), .A1(net_2205) );
NAND2_X2 inst_3042 ( .A1(net_6993), .A2(net_4977), .ZN(net_4965) );
CLKBUF_X2 inst_10945 ( .A(net_10906), .Z(net_10907) );
CLKBUF_X2 inst_8822 ( .A(net_8783), .Z(net_8784) );
NAND2_X2 inst_3243 ( .A1(net_7767), .ZN(net_4304), .A2(net_4145) );
CLKBUF_X2 inst_14039 ( .A(net_14000), .Z(net_14001) );
CLKBUF_X2 inst_8605 ( .A(net_8566), .Z(net_8567) );
CLKBUF_X2 inst_10564 ( .A(net_10525), .Z(net_10526) );
SDFF_X2 inst_981 ( .Q(net_6456), .D(net_6456), .SE(net_3904), .SI(net_3792), .CK(net_11550) );
CLKBUF_X2 inst_11940 ( .A(net_11901), .Z(net_11902) );
AOI21_X2 inst_7735 ( .B1(net_6600), .ZN(net_4028), .B2(net_2583), .A(net_2290) );
CLKBUF_X2 inst_8815 ( .A(net_8776), .Z(net_8777) );
SDFF_X2 inst_1266 ( .Q(net_6556), .D(net_3420), .SI(net_3419), .SE(net_2244), .CK(net_10700) );
CLKBUF_X2 inst_8904 ( .A(net_8439), .Z(net_8866) );
DFF_X2 inst_6189 ( .QN(net_6960), .D(net_5076), .CK(net_11370) );
CLKBUF_X2 inst_12260 ( .A(net_12221), .Z(net_12222) );
CLKBUF_X2 inst_12064 ( .A(net_12025), .Z(net_12026) );
OAI21_X2 inst_2094 ( .B2(net_4447), .ZN(net_4322), .B1(net_4080), .A(net_3570) );
INV_X4 inst_5102 ( .A(net_7808), .ZN(net_3810) );
INV_X4 inst_4872 ( .ZN(net_1268), .A(net_639) );
DFF_X2 inst_6287 ( .D(net_2394), .QN(net_263), .CK(net_10782) );
NAND2_X1 inst_4317 ( .ZN(net_4547), .A2(net_3870), .A1(net_1513) );
CLKBUF_X2 inst_13310 ( .A(net_11191), .Z(net_13272) );
DFF_X2 inst_6279 ( .QN(net_6184), .D(net_2617), .CK(net_7929) );
NAND2_X2 inst_3417 ( .A2(net_5893), .ZN(net_3333), .A1(net_626) );
CLKBUF_X2 inst_13347 ( .A(net_10781), .Z(net_13309) );
DFFR_X2 inst_7090 ( .QN(net_7724), .D(net_2791), .CK(net_10740), .RN(x1822) );
DFF_X1 inst_6794 ( .D(net_3944), .CK(net_12619), .Q(x494) );
CLKBUF_X2 inst_14337 ( .A(net_14298), .Z(net_14299) );
CLKBUF_X2 inst_11379 ( .A(net_11340), .Z(net_11341) );
INV_X4 inst_5406 ( .ZN(net_418), .A(net_288) );
DFF_X2 inst_6292 ( .QN(net_6401), .D(net_1837), .CK(net_12965) );
CLKBUF_X2 inst_13959 ( .A(net_13887), .Z(net_13921) );
INV_X4 inst_5324 ( .A(net_6418), .ZN(net_896) );
NAND2_X2 inst_3491 ( .ZN(net_2648), .A1(net_2647), .A2(net_2646) );
NOR2_X2 inst_2393 ( .A2(net_3996), .ZN(net_3995), .A1(net_2452) );
OAI21_X2 inst_1838 ( .B1(net_5365), .ZN(net_5334), .A(net_4375), .B2(net_3853) );
XNOR2_X2 inst_71 ( .B(net_6421), .ZN(net_1703), .A(net_1071) );
CLKBUF_X2 inst_9414 ( .A(net_9375), .Z(net_9376) );
OAI22_X2 inst_1454 ( .B2(net_5899), .B1(net_4650), .ZN(net_4615), .A2(net_4614), .A1(net_4066) );
CLKBUF_X2 inst_9438 ( .A(net_9399), .Z(net_9400) );
CLKBUF_X2 inst_10114 ( .A(net_9614), .Z(net_10076) );
NAND2_X2 inst_4079 ( .A1(net_6665), .A2(net_1655), .ZN(net_973) );
NAND2_X2 inst_3231 ( .ZN(net_4524), .A2(net_4292), .A1(net_1734) );
NAND2_X2 inst_3147 ( .ZN(net_4816), .A2(net_4153), .A1(net_2071) );
CLKBUF_X2 inst_9084 ( .A(net_9045), .Z(net_9046) );
OAI21_X2 inst_1945 ( .B1(net_5232), .ZN(net_5080), .A(net_4732), .B2(net_3986) );
INV_X4 inst_5564 ( .A(net_7431), .ZN(net_2093) );
NAND3_X2 inst_2657 ( .ZN(net_3943), .A3(net_3440), .A2(net_2933), .A1(net_2823) );
CLKBUF_X2 inst_12884 ( .A(net_12845), .Z(net_12846) );
CLKBUF_X2 inst_14407 ( .A(net_9283), .Z(net_14369) );
INV_X2 inst_5722 ( .ZN(net_4006), .A(net_3916) );
SDFF_X2 inst_336 ( .SI(net_7458), .Q(net_7458), .D(net_5094), .SE(net_3993), .CK(net_9760) );
CLKBUF_X2 inst_12129 ( .A(net_12090), .Z(net_12091) );
AOI21_X2 inst_7720 ( .B1(net_6594), .ZN(net_5903), .B2(net_2583), .A(net_2279) );
CLKBUF_X2 inst_13239 ( .A(net_13200), .Z(net_13201) );
CLKBUF_X2 inst_13043 ( .A(net_12624), .Z(net_13005) );
CLKBUF_X2 inst_12930 ( .A(net_12891), .Z(net_12892) );
SDFF_X2 inst_376 ( .SI(net_7671), .Q(net_7671), .D(net_4790), .SE(net_3866), .CK(net_7984) );
DFF_X1 inst_6479 ( .QN(net_7401), .D(net_5573), .CK(net_9819) );
CLKBUF_X2 inst_10816 ( .A(net_10777), .Z(net_10778) );
INV_X4 inst_5157 ( .ZN(net_557), .A(net_556) );
OAI21_X2 inst_1939 ( .B1(net_5542), .ZN(net_5096), .A(net_4738), .B2(net_3988) );
NAND2_X2 inst_3268 ( .ZN(net_3710), .A1(net_3709), .A2(net_3226) );
NAND2_X4 inst_2902 ( .ZN(net_3392), .A1(net_3240), .A2(net_3222) );
AND2_X4 inst_7844 ( .A2(net_6409), .A1(net_6408), .ZN(net_1823) );
CLKBUF_X2 inst_14066 ( .A(net_11481), .Z(net_14028) );
CLKBUF_X2 inst_8726 ( .A(net_8687), .Z(net_8688) );
CLKBUF_X2 inst_11676 ( .A(net_11637), .Z(net_11638) );
CLKBUF_X2 inst_12167 ( .A(net_12075), .Z(net_12129) );
CLKBUF_X2 inst_8508 ( .A(net_8469), .Z(net_8470) );
INV_X4 inst_5174 ( .A(net_650), .ZN(net_533) );
CLKBUF_X2 inst_13450 ( .A(net_13411), .Z(net_13412) );
CLKBUF_X2 inst_9553 ( .A(net_9514), .Z(net_9515) );
AND2_X2 inst_7856 ( .ZN(net_3015), .A2(net_2817), .A1(net_2254) );
CLKBUF_X2 inst_10991 ( .A(net_10952), .Z(net_10953) );
CLKBUF_X2 inst_11736 ( .A(net_8213), .Z(net_11698) );
CLKBUF_X2 inst_8897 ( .A(net_8858), .Z(net_8859) );
DFF_X2 inst_6299 ( .QN(net_5977), .D(net_1661), .CK(net_12525) );
CLKBUF_X2 inst_8263 ( .A(net_7969), .Z(net_8225) );
CLKBUF_X2 inst_12627 ( .A(net_12588), .Z(net_12589) );
INV_X2 inst_5870 ( .A(net_892), .ZN(net_488) );
CLKBUF_X2 inst_13251 ( .A(net_10699), .Z(net_13213) );
CLKBUF_X2 inst_10852 ( .A(net_10813), .Z(net_10814) );
CLKBUF_X2 inst_9951 ( .A(net_9912), .Z(net_9913) );
NAND2_X2 inst_3880 ( .A1(net_7115), .A2(net_1675), .ZN(net_1440) );
NAND2_X2 inst_3100 ( .ZN(net_4903), .A2(net_4327), .A1(net_2245) );
CLKBUF_X2 inst_8359 ( .A(net_7883), .Z(net_8321) );
INV_X2 inst_5998 ( .A(net_7628), .ZN(net_1895) );
NAND2_X2 inst_4052 ( .A1(net_6537), .A2(net_1645), .ZN(net_1000) );
CLKBUF_X2 inst_8552 ( .A(net_8513), .Z(net_8514) );
NAND2_X1 inst_4251 ( .ZN(net_4675), .A2(net_3988), .A1(net_2218) );
INV_X8 inst_4487 ( .ZN(net_4666), .A(net_3412) );
OAI22_X2 inst_1596 ( .A1(net_3289), .B2(net_3200), .A2(net_3187), .ZN(net_3141), .B1(net_740) );
NAND2_X1 inst_4364 ( .ZN(net_4363), .A2(net_3853), .A1(net_2004) );
DFF_X1 inst_6400 ( .QN(net_6139), .D(net_5688), .CK(net_11533) );
NAND2_X2 inst_3752 ( .A1(net_7035), .A2(net_1975), .ZN(net_1593) );
DFFR_X2 inst_7078 ( .QN(net_7748), .D(net_2796), .CK(net_8580), .RN(x1822) );
CLKBUF_X2 inst_10174 ( .A(net_10135), .Z(net_10136) );
NOR2_X4 inst_2265 ( .ZN(net_5621), .A1(net_5466), .A2(net_4417) );
SDFF_X2 inst_284 ( .D(net_6397), .SE(net_6052), .SI(net_322), .Q(net_322), .CK(net_13827) );
CLKBUF_X2 inst_13494 ( .A(net_13455), .Z(net_13456) );
OAI22_X2 inst_1555 ( .B2(net_3405), .A2(net_3360), .ZN(net_3350), .A1(net_3131), .B1(net_423) );
CLKBUF_X2 inst_13809 ( .A(net_9501), .Z(net_13771) );
SDFF_X2 inst_1293 ( .D(net_3812), .SE(net_3256), .SI(net_142), .Q(net_142), .CK(net_10683) );
NAND2_X2 inst_3805 ( .A1(net_6633), .A2(net_1624), .ZN(net_1540) );
NAND3_X2 inst_2579 ( .ZN(net_5760), .A1(net_5655), .A2(net_5277), .A3(net_4305) );
SDFF_X2 inst_280 ( .Q(net_6366), .SI(net_6365), .D(net_3556), .SE(net_392), .CK(net_13610) );
CLKBUF_X2 inst_11249 ( .A(net_11210), .Z(net_11211) );
CLKBUF_X2 inst_12668 ( .A(net_12629), .Z(net_12630) );
NAND2_X2 inst_3157 ( .ZN(net_4806), .A2(net_4805), .A1(net_4257) );
OAI21_X2 inst_1713 ( .ZN(net_5581), .A(net_5126), .B2(net_4416), .B1(net_4030) );
DFFR_X2 inst_6970 ( .QN(net_6015), .D(net_4004), .CK(net_10455), .RN(x1822) );
INV_X4 inst_5650 ( .A(net_7232), .ZN(net_598) );
CLKBUF_X2 inst_9888 ( .A(net_8199), .Z(net_9850) );
INV_X8 inst_4527 ( .ZN(net_3756), .A(net_3113) );
CLKBUF_X2 inst_11657 ( .A(net_10918), .Z(net_11619) );
CLKBUF_X2 inst_9532 ( .A(net_9202), .Z(net_9494) );
NAND2_X2 inst_3137 ( .ZN(net_4826), .A2(net_4153), .A1(net_2081) );
CLKBUF_X2 inst_13648 ( .A(net_13609), .Z(net_13610) );
INV_X4 inst_4676 ( .ZN(net_3462), .A(net_3461) );
CLKBUF_X2 inst_11668 ( .A(net_9270), .Z(net_11630) );
CLKBUF_X2 inst_14071 ( .A(net_14032), .Z(net_14033) );
INV_X4 inst_5437 ( .A(net_6088), .ZN(net_3485) );
AOI222_X2 inst_7544 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1874), .A1(net_1873), .B1(net_1872), .C1(net_1871) );
CLKBUF_X2 inst_8110 ( .A(net_8071), .Z(net_8072) );
CLKBUF_X2 inst_11556 ( .A(net_9127), .Z(net_11518) );
CLKBUF_X2 inst_10344 ( .A(net_10305), .Z(net_10306) );
INV_X8 inst_4496 ( .ZN(net_3903), .A(net_3110) );
AOI22_X2 inst_7357 ( .B2(net_3105), .ZN(net_3092), .A2(net_2712), .A1(net_1131), .B1(net_760) );
DFF_X1 inst_6344 ( .QN(net_6187), .D(net_5841), .CK(net_13644) );
SDFF_X2 inst_951 ( .SI(net_7194), .Q(net_7194), .SE(net_3819), .D(net_3800), .CK(net_10622) );
CLKBUF_X2 inst_12565 ( .A(net_11354), .Z(net_12527) );
DFF_X1 inst_6586 ( .QN(net_7556), .D(net_5064), .CK(net_13085) );
CLKBUF_X2 inst_9836 ( .A(net_9724), .Z(net_9798) );
AOI21_X2 inst_7727 ( .B1(net_6462), .ZN(net_4439), .B2(net_2580), .A(net_2379) );
CLKBUF_X2 inst_11188 ( .A(net_9079), .Z(net_11150) );
INV_X2 inst_5831 ( .A(net_1300), .ZN(net_907) );
NAND2_X1 inst_4393 ( .ZN(net_4334), .A2(net_3859), .A1(net_2208) );
CLKBUF_X2 inst_10268 ( .A(net_8738), .Z(net_10230) );
CLKBUF_X2 inst_8299 ( .A(net_8260), .Z(net_8261) );
CLKBUF_X2 inst_11253 ( .A(net_9857), .Z(net_11215) );
CLKBUF_X2 inst_12743 ( .A(net_12704), .Z(net_12705) );
CLKBUF_X2 inst_8938 ( .A(net_8899), .Z(net_8900) );
SDFFR_X2 inst_1359 ( .SI(net_6035), .Q(net_6035), .D(net_3883), .SE(net_3087), .CK(net_9972), .RN(x1822) );
CLKBUF_X2 inst_10345 ( .A(net_10306), .Z(net_10307) );
AOI222_X2 inst_7499 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2076), .A1(net_2075), .B1(net_2074), .C1(net_2073) );
NAND2_X2 inst_3188 ( .ZN(net_4745), .A2(net_3941), .A1(net_2212) );
AOI22_X2 inst_7358 ( .B2(net_3105), .ZN(net_3091), .A2(net_2712), .A1(net_1109), .B1(net_694) );
CLKBUF_X2 inst_11545 ( .A(net_10790), .Z(net_11507) );
AOI22_X2 inst_7435 ( .B1(net_7079), .A1(net_7047), .ZN(net_1976), .A2(net_1975), .B2(net_791) );
AOI22_X2 inst_7351 ( .B2(net_3105), .ZN(net_3099), .A2(net_2712), .A1(net_1111), .B1(net_452) );
NAND2_X2 inst_3129 ( .ZN(net_4834), .A2(net_4153), .A1(net_2085) );
CLKBUF_X2 inst_12590 ( .A(net_12551), .Z(net_12552) );
INV_X4 inst_4674 ( .ZN(net_3467), .A(net_3466) );
CLKBUF_X2 inst_11328 ( .A(net_11289), .Z(net_11290) );
NAND2_X2 inst_3797 ( .A1(net_6499), .A2(net_1642), .ZN(net_1548) );
XNOR2_X2 inst_100 ( .ZN(net_2257), .A(net_1150), .B(net_1144) );
INV_X4 inst_5581 ( .A(net_6009), .ZN(net_2968) );
NAND2_X1 inst_4352 ( .ZN(net_4375), .A2(net_3853), .A1(net_2161) );
SDFF_X2 inst_921 ( .Q(net_7159), .D(net_7159), .SE(net_3903), .SI(net_3793), .CK(net_8079) );
SDFF_X2 inst_279 ( .D(net_6398), .SE(net_6052), .SI(net_323), .Q(net_323), .CK(net_13828) );
CLKBUF_X2 inst_14202 ( .A(net_14163), .Z(net_14164) );
CLKBUF_X2 inst_10772 ( .A(net_9302), .Z(net_10734) );
AOI21_X4 inst_7618 ( .B2(net_5945), .B1(net_5944), .ZN(net_5610), .A(x1062) );
AOI22_X2 inst_7425 ( .A1(net_2970), .B1(net_2772), .ZN(net_2767), .A2(net_236), .B2(net_162) );
NAND2_X2 inst_3970 ( .ZN(net_1310), .A2(net_1107), .A1(net_811) );
NAND2_X2 inst_3387 ( .ZN(net_3456), .A2(net_3455), .A1(net_3375) );
CLKBUF_X2 inst_11683 ( .A(net_11644), .Z(net_11645) );
CLKBUF_X2 inst_11014 ( .A(net_10975), .Z(net_10976) );
CLKBUF_X2 inst_8271 ( .A(net_7877), .Z(net_8233) );
XNOR2_X2 inst_81 ( .ZN(net_1647), .A(net_1646), .B(net_826) );
CLKBUF_X2 inst_11499 ( .A(net_10572), .Z(net_11461) );
INV_X2 inst_5806 ( .ZN(net_1277), .A(net_689) );
CLKBUF_X2 inst_13424 ( .A(net_13385), .Z(net_13386) );
CLKBUF_X2 inst_9761 ( .A(net_9722), .Z(net_9723) );
DFF_X1 inst_6395 ( .QN(net_6134), .D(net_5693), .CK(net_10974) );
DFFR_X2 inst_7087 ( .QN(net_7747), .D(net_2797), .CK(net_8579), .RN(x1822) );
CLKBUF_X2 inst_9471 ( .A(net_9432), .Z(net_9433) );
CLKBUF_X2 inst_8825 ( .A(net_8786), .Z(net_8787) );
CLKBUF_X2 inst_14411 ( .A(net_14372), .Z(net_14373) );
CLKBUF_X2 inst_12040 ( .A(net_10777), .Z(net_12002) );
SDFF_X2 inst_790 ( .SI(net_6920), .Q(net_6920), .SE(net_3887), .D(net_3789), .CK(net_8134) );
CLKBUF_X2 inst_10515 ( .A(net_10476), .Z(net_10477) );
SDFF_X2 inst_1009 ( .SI(net_6501), .Q(net_6501), .SE(net_3886), .D(net_3811), .CK(net_11650) );
CLKBUF_X2 inst_8931 ( .A(net_8892), .Z(net_8893) );
CLKBUF_X2 inst_8024 ( .A(net_7985), .Z(net_7986) );
NAND2_X2 inst_2954 ( .ZN(net_5486), .A1(net_4941), .A2(net_4940) );
CLKBUF_X2 inst_9711 ( .A(net_9037), .Z(net_9673) );
CLKBUF_X2 inst_13217 ( .A(net_13178), .Z(net_13179) );
CLKBUF_X2 inst_12045 ( .A(net_12006), .Z(net_12007) );
CLKBUF_X2 inst_11844 ( .A(net_8222), .Z(net_11806) );
NOR3_X2 inst_2197 ( .ZN(net_3879), .A1(net_3378), .A3(net_1263), .A2(net_782) );
CLKBUF_X2 inst_7995 ( .A(net_7956), .Z(net_7957) );
SDFF_X2 inst_733 ( .Q(net_6849), .D(net_6849), .SE(net_3893), .SI(net_3805), .CK(net_10905) );
INV_X2 inst_5885 ( .A(net_7653), .ZN(net_1986) );
CLKBUF_X2 inst_13064 ( .A(net_8478), .Z(net_13026) );
OAI21_X2 inst_1959 ( .B1(net_5200), .ZN(net_5061), .A(net_4706), .B2(net_3986) );
NAND3_X2 inst_2582 ( .ZN(net_5757), .A1(net_5652), .A2(net_5274), .A3(net_4312) );
SDFF_X2 inst_142 ( .Q(net_6236), .SI(net_6235), .SE(net_392), .D(net_142), .CK(net_13619) );
CLKBUF_X2 inst_14294 ( .A(net_12279), .Z(net_14256) );
XNOR2_X2 inst_78 ( .ZN(net_1934), .B(net_676), .A(net_639) );
CLKBUF_X2 inst_13182 ( .A(net_13143), .Z(net_13144) );
CLKBUF_X2 inst_8020 ( .A(net_7935), .Z(net_7982) );
CLKBUF_X2 inst_7896 ( .A(net_7844), .Z(net_7858) );
NAND3_X2 inst_2813 ( .ZN(net_2285), .A3(net_1582), .A1(net_1375), .A2(net_1038) );
SDFF_X2 inst_177 ( .Q(net_6277), .SI(net_6276), .D(net_3501), .SE(net_392), .CK(net_13485) );
CLKBUF_X2 inst_7892 ( .A(net_7853), .Z(net_7854) );
SDFF_X2 inst_783 ( .SI(net_6912), .Q(net_6912), .D(net_3807), .SE(net_3781), .CK(net_11723) );
DFF_X1 inst_6416 ( .QN(net_6163), .D(net_5754), .CK(net_11039) );
CLKBUF_X2 inst_7910 ( .A(net_7871), .Z(net_7872) );
CLKBUF_X2 inst_8450 ( .A(net_8411), .Z(net_8412) );
INV_X4 inst_5696 ( .A(net_6087), .ZN(net_3487) );
OAI21_X2 inst_2014 ( .B2(net_4497), .ZN(net_4494), .B1(net_4110), .A(net_3658) );
INV_X8 inst_4471 ( .ZN(net_5244), .A(net_4277) );
INV_X16 inst_6122 ( .ZN(net_4977), .A(net_4265) );
CLKBUF_X2 inst_10144 ( .A(net_10105), .Z(net_10106) );
SDFF_X2 inst_615 ( .Q(net_6593), .D(net_6593), .SE(net_3830), .SI(net_3802), .CK(net_12910) );
CLKBUF_X2 inst_12182 ( .A(net_12143), .Z(net_12144) );
CLKBUF_X2 inst_12597 ( .A(net_12558), .Z(net_12559) );
CLKBUF_X2 inst_12821 ( .A(net_11813), .Z(net_12783) );
CLKBUF_X2 inst_9999 ( .A(net_8062), .Z(net_9961) );
CLKBUF_X2 inst_9157 ( .A(net_9118), .Z(net_9119) );
CLKBUF_X2 inst_8456 ( .A(net_8008), .Z(net_8418) );
NAND3_X2 inst_2822 ( .A2(net_3849), .ZN(net_1829), .A3(net_1828), .A1(net_657) );
NOR2_X2 inst_2467 ( .A2(net_2729), .ZN(net_2728), .A1(net_2727) );
CLKBUF_X2 inst_7906 ( .A(net_7867), .Z(net_7868) );
DFF_X2 inst_6176 ( .Q(net_6398), .D(net_6397), .CK(net_14189) );
NAND2_X2 inst_3843 ( .A2(net_1696), .ZN(net_1495), .A1(net_1494) );
CLKBUF_X2 inst_11583 ( .A(net_10631), .Z(net_11545) );
CLKBUF_X2 inst_10621 ( .A(net_10582), .Z(net_10583) );
CLKBUF_X2 inst_10335 ( .A(net_10296), .Z(net_10297) );
CLKBUF_X2 inst_8656 ( .A(net_8617), .Z(net_8618) );
OAI21_X2 inst_2031 ( .B2(net_4476), .ZN(net_4472), .B1(net_4173), .A(net_3602) );
NAND2_X1 inst_4386 ( .ZN(net_4341), .A2(net_3859), .A1(net_2037) );
CLKBUF_X2 inst_13632 ( .A(net_9409), .Z(net_13594) );
INV_X4 inst_5593 ( .A(net_6064), .ZN(net_3585) );
CLKBUF_X2 inst_11282 ( .A(net_11243), .Z(net_11244) );
CLKBUF_X2 inst_10255 ( .A(net_10216), .Z(net_10217) );
CLKBUF_X2 inst_11527 ( .A(net_11488), .Z(net_11489) );
CLKBUF_X2 inst_8525 ( .A(net_8486), .Z(net_8487) );
INV_X4 inst_4941 ( .ZN(net_749), .A(net_748) );
AND2_X4 inst_7835 ( .ZN(net_2924), .A1(net_2704), .A2(net_264) );
DFFR_X2 inst_7095 ( .QN(net_7720), .D(net_2593), .CK(net_9599), .RN(x1822) );
INV_X4 inst_5133 ( .ZN(net_3152), .A(net_587) );
CLKBUF_X2 inst_9986 ( .A(net_9947), .Z(net_9948) );
SDFF_X2 inst_338 ( .SI(net_7527), .Q(net_7527), .D(net_5097), .SE(net_3988), .CK(net_12438) );
INV_X4 inst_5577 ( .A(net_7699), .ZN(net_438) );
NOR2_X2 inst_2412 ( .A1(net_6019), .ZN(net_3411), .A2(net_3404) );
INV_X4 inst_4928 ( .ZN(net_1656), .A(net_625) );
NAND2_X2 inst_4005 ( .ZN(net_1279), .A1(net_686), .A2(net_630) );
CLKBUF_X2 inst_10384 ( .A(net_10345), .Z(net_10346) );
INV_X4 inst_5424 ( .A(net_5995), .ZN(net_551) );
NAND2_X1 inst_4323 ( .ZN(net_4541), .A2(net_3870), .A1(net_1398) );
NOR3_X2 inst_2214 ( .ZN(net_2224), .A1(net_1916), .A3(net_1682), .A2(net_871) );
DFF_X1 inst_6468 ( .QN(net_6169), .D(net_5591), .CK(net_7967) );
CLKBUF_X2 inst_10018 ( .A(net_9979), .Z(net_9980) );
NOR2_X2 inst_2474 ( .A2(net_5778), .ZN(net_2608), .A1(net_2607) );
CLKBUF_X2 inst_14051 ( .A(net_14012), .Z(net_14013) );
SDFF_X2 inst_579 ( .Q(net_6576), .D(net_6576), .SE(net_3823), .SI(net_3808), .CK(net_12188) );
INV_X4 inst_5247 ( .ZN(net_1728), .A(net_886) );
NOR2_X2 inst_2495 ( .ZN(net_1748), .A2(net_1747), .A1(net_1072) );
NAND2_X2 inst_4019 ( .A1(net_6669), .A2(net_1655), .ZN(net_1033) );
DFF_X1 inst_6902 ( .D(net_2493), .Q(net_183), .CK(net_9938) );
CLKBUF_X2 inst_11265 ( .A(net_11226), .Z(net_11227) );
AOI222_X2 inst_7462 ( .ZN(net_2206), .A1(net_2205), .A2(net_2204), .B1(net_2203), .B2(net_2202), .C1(net_2201), .C2(net_2200) );
CLKBUF_X2 inst_11697 ( .A(net_11658), .Z(net_11659) );
CLKBUF_X2 inst_11219 ( .A(net_8815), .Z(net_11181) );
NAND2_X2 inst_3236 ( .ZN(net_4279), .A2(net_4278), .A1(net_1975) );
SDFF_X2 inst_698 ( .SI(net_6758), .Q(net_6758), .SE(net_3816), .D(net_3792), .CK(net_8280) );
CLKBUF_X2 inst_14378 ( .A(net_14339), .Z(net_14340) );
CLKBUF_X2 inst_11096 ( .A(net_11057), .Z(net_11058) );
CLKBUF_X2 inst_10474 ( .A(net_10435), .Z(net_10436) );
NAND2_X2 inst_3964 ( .A1(net_6433), .A2(net_1677), .ZN(net_1318) );
NAND2_X2 inst_3944 ( .A1(net_6979), .A2(net_1833), .ZN(net_1347) );
NAND2_X2 inst_3394 ( .ZN(net_3757), .A2(net_3363), .A1(net_2887) );
NAND2_X2 inst_3408 ( .ZN(net_3340), .A1(net_3339), .A2(net_435) );
XNOR2_X2 inst_88 ( .ZN(net_1917), .A(net_724), .B(net_600) );
INV_X2 inst_5978 ( .A(net_7661), .ZN(net_1901) );
INV_X2 inst_6054 ( .ZN(net_1261), .A(net_121) );
CLKBUF_X2 inst_10397 ( .A(net_9615), .Z(net_10359) );
NAND2_X4 inst_2863 ( .ZN(net_4288), .A1(net_4280), .A2(net_1654) );
CLKBUF_X2 inst_10356 ( .A(net_9902), .Z(net_10318) );
CLKBUF_X2 inst_8401 ( .A(net_8362), .Z(net_8363) );
CLKBUF_X2 inst_12882 ( .A(net_10729), .Z(net_12844) );
CLKBUF_X2 inst_11190 ( .A(net_11151), .Z(net_11152) );
SDFF_X2 inst_360 ( .SI(net_7608), .Q(net_7608), .D(net_4789), .SE(net_3870), .CK(net_10278) );
NAND2_X2 inst_3897 ( .A1(net_7109), .A2(net_1675), .ZN(net_1417) );
INV_X4 inst_5534 ( .A(net_6131), .ZN(net_3631) );
DFF_X1 inst_6604 ( .QN(net_7511), .D(net_5404), .CK(net_9235) );
CLKBUF_X2 inst_11458 ( .A(net_11419), .Z(net_11420) );
CLKBUF_X2 inst_10876 ( .A(net_10837), .Z(net_10838) );
CLKBUF_X2 inst_11693 ( .A(net_11385), .Z(net_11655) );
NAND2_X2 inst_3908 ( .A1(net_7112), .A2(net_1675), .ZN(net_1402) );
NAND2_X2 inst_3754 ( .A1(net_7045), .A2(net_1975), .ZN(net_1591) );
INV_X1 inst_6160 ( .A(net_5853), .ZN(x96) );
CLKBUF_X2 inst_12574 ( .A(net_12535), .Z(net_12536) );
DFF_X1 inst_6797 ( .D(net_3943), .CK(net_9567), .Q(x699) );
SDFF_X2 inst_1129 ( .SI(net_6680), .Q(net_6680), .D(net_3898), .SE(net_3471), .CK(net_11998) );
CLKBUF_X2 inst_10229 ( .A(net_10190), .Z(net_10191) );
CLKBUF_X2 inst_8922 ( .A(net_8883), .Z(net_8884) );
SDFF_X2 inst_837 ( .Q(net_7016), .D(net_7016), .SE(net_3899), .SI(net_3805), .CK(net_9031) );
INV_X2 inst_5716 ( .ZN(net_4250), .A(net_4121) );
SDFF_X2 inst_744 ( .Q(net_6833), .D(net_6833), .SE(net_3893), .SI(net_3799), .CK(net_11813) );
CLKBUF_X2 inst_13116 ( .A(net_13077), .Z(net_13078) );
CLKBUF_X2 inst_13375 ( .A(net_13336), .Z(net_13337) );
NAND2_X2 inst_3827 ( .A1(net_6839), .A2(net_1521), .ZN(net_1516) );
CLKBUF_X2 inst_14425 ( .A(net_14386), .Z(net_14387) );
CLKBUF_X2 inst_8956 ( .A(net_8917), .Z(net_8918) );
CLKBUF_X2 inst_12385 ( .A(net_12346), .Z(net_12347) );
DFF_X1 inst_6509 ( .QN(net_7431), .D(net_5514), .CK(net_12488) );
INV_X4 inst_5457 ( .A(net_6069), .ZN(net_3621) );
CLKBUF_X2 inst_13492 ( .A(net_11714), .Z(net_13454) );
NAND2_X2 inst_4112 ( .A1(net_6660), .A2(net_1655), .ZN(net_940) );
DFFR_X2 inst_7025 ( .D(net_3292), .QN(net_279), .CK(net_9616), .RN(x1822) );
CLKBUF_X2 inst_8785 ( .A(net_8746), .Z(net_8747) );
AND3_X4 inst_7798 ( .ZN(net_2587), .A1(net_2389), .A3(net_2229), .A2(net_1709) );
CLKBUF_X2 inst_10497 ( .A(net_10458), .Z(net_10459) );
AOI21_X2 inst_7664 ( .B2(net_5927), .ZN(net_3312), .A(net_3311), .B1(net_1214) );
CLKBUF_X2 inst_11002 ( .A(net_10963), .Z(net_10964) );
XNOR2_X2 inst_65 ( .ZN(net_2480), .A(net_1077), .B(net_559) );
CLKBUF_X2 inst_12443 ( .A(net_12404), .Z(net_12405) );
SDFF_X2 inst_536 ( .Q(net_7240), .D(net_7240), .SE(net_3822), .SI(net_336), .CK(net_12679) );
CLKBUF_X2 inst_9563 ( .A(net_9524), .Z(net_9525) );
CLKBUF_X2 inst_12711 ( .A(net_12672), .Z(net_12673) );
NAND2_X2 inst_3592 ( .ZN(net_2408), .A2(net_1888), .A1(net_1445) );
DFF_X1 inst_6822 ( .QN(net_5972), .D(net_3016), .CK(net_8571) );
INV_X4 inst_5121 ( .A(net_601), .ZN(net_596) );
NAND2_X2 inst_3732 ( .A1(net_6912), .A2(net_1639), .ZN(net_1613) );
CLKBUF_X2 inst_11032 ( .A(net_10993), .Z(net_10994) );
INV_X8 inst_4503 ( .ZN(net_3816), .A(net_3262) );
CLKBUF_X2 inst_9658 ( .A(net_9619), .Z(net_9620) );
CLKBUF_X2 inst_8146 ( .A(net_8107), .Z(net_8108) );
INV_X4 inst_4907 ( .A(net_3810), .ZN(net_3198) );
OAI21_X2 inst_2027 ( .ZN(net_4478), .B1(net_4477), .B2(net_4476), .A(net_3612) );
INV_X2 inst_5882 ( .ZN(net_3073), .A(net_279) );
NAND2_X2 inst_2926 ( .ZN(net_5529), .A1(net_5003), .A2(net_5002) );
AOI222_X2 inst_7487 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2116), .A1(net_2115), .B1(net_2114), .C1(net_2113) );
SDFF_X2 inst_416 ( .D(net_6392), .SE(net_5799), .SI(net_377), .Q(net_377), .CK(net_13894) );
CLKBUF_X2 inst_9169 ( .A(net_9130), .Z(net_9131) );
SDFF_X2 inst_1158 ( .SI(net_6821), .Q(net_6821), .D(net_3800), .SE(net_3729), .CK(net_11375) );
CLKBUF_X2 inst_9059 ( .A(net_9020), .Z(net_9021) );
OAI21_X2 inst_1870 ( .ZN(net_5241), .B1(net_5240), .A(net_4593), .B2(net_3867) );
CLKBUF_X2 inst_13445 ( .A(net_13406), .Z(net_13407) );
CLKBUF_X2 inst_10871 ( .A(net_10832), .Z(net_10833) );
DFFR_X2 inst_7038 ( .QN(net_5984), .D(net_3129), .CK(net_10347), .RN(x1822) );
OR2_X2 inst_1406 ( .A1(net_6417), .A2(net_6416), .ZN(x30) );
CLKBUF_X2 inst_8396 ( .A(net_8357), .Z(net_8358) );
INV_X4 inst_5500 ( .A(net_5986), .ZN(net_440) );
INV_X4 inst_5330 ( .A(net_6032), .ZN(net_572) );
INV_X4 inst_5270 ( .ZN(net_1145), .A(net_421) );
NAND2_X1 inst_4319 ( .ZN(net_4545), .A2(net_3870), .A1(net_1372) );
CLKBUF_X2 inst_10943 ( .A(net_10904), .Z(net_10905) );
CLKBUF_X2 inst_9520 ( .A(net_9481), .Z(net_9482) );
CLKBUF_X2 inst_8436 ( .A(net_8221), .Z(net_8398) );
CLKBUF_X2 inst_8046 ( .A(net_7975), .Z(net_8008) );
NOR2_X2 inst_2445 ( .A2(net_5967), .ZN(net_3154), .A1(net_2999) );
NAND2_X1 inst_4432 ( .A1(net_7613), .A2(net_2131), .ZN(net_1420) );
CLKBUF_X2 inst_11039 ( .A(net_8778), .Z(net_11001) );
CLKBUF_X2 inst_13014 ( .A(net_9647), .Z(net_12976) );
NAND2_X2 inst_3039 ( .A1(net_7024), .A2(net_4979), .ZN(net_4968) );
INV_X4 inst_5477 ( .A(net_7558), .ZN(net_2091) );
SDFF_X2 inst_973 ( .Q(net_6426), .D(net_6426), .SE(net_3820), .SI(net_3802), .CK(net_8855) );
CLKBUF_X2 inst_13374 ( .A(net_10819), .Z(net_13336) );
NAND2_X2 inst_3058 ( .A1(net_7156), .A2(net_4954), .ZN(net_4947) );
SDFF_X2 inst_461 ( .SI(net_6918), .Q(net_6918), .D(net_3898), .SE(net_3887), .CK(net_11520) );
INV_X2 inst_6092 ( .ZN(net_3080), .A(net_290) );
CLKBUF_X2 inst_11258 ( .A(net_11219), .Z(net_11220) );
CLKBUF_X2 inst_11884 ( .A(net_11845), .Z(net_11846) );
CLKBUF_X2 inst_8291 ( .A(net_8061), .Z(net_8253) );
CLKBUF_X2 inst_11771 ( .A(net_9839), .Z(net_11733) );
DFF_X1 inst_6387 ( .QN(net_6118), .D(net_5701), .CK(net_11202) );
OAI21_X2 inst_1973 ( .B1(net_4868), .ZN(net_4863), .A(net_4374), .B2(net_3856) );
NAND2_X2 inst_3089 ( .A1(net_6452), .A2(net_4925), .ZN(net_4914) );
NAND2_X2 inst_3051 ( .ZN(net_4956), .A2(net_4329), .A1(net_2253) );
CLKBUF_X2 inst_8326 ( .A(net_8287), .Z(net_8288) );
NAND3_X2 inst_2668 ( .ZN(net_3961), .A2(net_3875), .A3(net_3737), .A1(net_2239) );
SDFF_X2 inst_1122 ( .SI(net_6672), .Q(net_6672), .D(net_3776), .SE(net_3465), .CK(net_12140) );
CLKBUF_X2 inst_12170 ( .A(net_12131), .Z(net_12132) );
NAND2_X2 inst_3324 ( .ZN(net_3598), .A1(net_3597), .A2(net_3228) );
CLKBUF_X2 inst_14447 ( .A(net_14408), .Z(net_14409) );
CLKBUF_X2 inst_14238 ( .A(net_11342), .Z(net_14200) );
CLKBUF_X2 inst_7987 ( .A(net_7948), .Z(net_7949) );
AOI222_X2 inst_7478 ( .ZN(net_2149), .A1(net_2148), .B1(net_2147), .C1(net_2146), .A2(net_2135), .B2(net_2133), .C2(net_2131) );
INV_X2 inst_5742 ( .ZN(net_3723), .A(net_3421) );
CLKBUF_X2 inst_14351 ( .A(net_14312), .Z(net_14313) );
INV_X2 inst_5775 ( .ZN(net_2876), .A(net_2808) );
INV_X4 inst_4808 ( .ZN(net_4786), .A(net_1174) );
INV_X4 inst_4657 ( .ZN(net_5879), .A(net_4141) );
NAND2_X2 inst_2981 ( .A1(net_6750), .A2(net_5033), .ZN(net_5030) );
OAI221_X2 inst_1669 ( .C2(net_5903), .ZN(net_4638), .B1(net_4637), .B2(net_4403), .C1(net_4030), .A(net_3488) );
AOI22_X2 inst_7456 ( .A2(net_7743), .B2(net_7741), .A1(net_7714), .B1(net_7712), .ZN(net_658) );
INV_X4 inst_4998 ( .A(net_7814), .ZN(net_3900) );
CLKBUF_X2 inst_9240 ( .A(net_9201), .Z(net_9202) );
INV_X4 inst_5390 ( .A(net_7572), .ZN(net_1838) );
NAND2_X1 inst_4406 ( .A2(net_3087), .ZN(net_2912), .A1(net_2911) );
CLKBUF_X2 inst_12195 ( .A(net_12156), .Z(net_12157) );
HA_X1 inst_6169 ( .S(net_1693), .CO(net_895), .A(net_894), .B(net_705) );
DFF_X1 inst_6696 ( .QN(net_7294), .D(net_5379), .CK(net_10176) );
NAND2_X2 inst_3162 ( .ZN(net_4771), .A2(net_3941), .A1(net_2033) );
NAND2_X2 inst_3956 ( .A1(net_6842), .A2(net_1521), .ZN(net_1329) );
XNOR2_X2 inst_90 ( .ZN(net_1202), .B(net_1201), .A(net_778) );
CLKBUF_X2 inst_11166 ( .A(net_11127), .Z(net_11128) );
CLKBUF_X2 inst_10850 ( .A(net_10811), .Z(net_10812) );
DFF_X1 inst_6858 ( .D(net_2551), .Q(net_224), .CK(net_12824) );
CLKBUF_X2 inst_8860 ( .A(net_8821), .Z(net_8822) );
INV_X4 inst_4650 ( .ZN(net_4614), .A(net_4276) );
OAI21_X2 inst_1801 ( .ZN(net_5389), .A(net_4716), .B2(net_3986), .B1(net_1167) );
CLKBUF_X2 inst_12777 ( .A(net_12738), .Z(net_12739) );
INV_X4 inst_5093 ( .A(net_7804), .ZN(net_3813) );
AOI21_X4 inst_7625 ( .B1(net_6998), .ZN(net_4624), .A(net_2462), .B2(net_1100) );
CLKBUF_X2 inst_9964 ( .A(net_9925), .Z(net_9926) );
NAND2_X2 inst_3833 ( .A1(net_6974), .A2(net_1833), .ZN(net_1506) );
SDFF_X2 inst_720 ( .D(net_7799), .SI(net_6764), .Q(net_6764), .SE(net_3872), .CK(net_11088) );
SDFF_X2 inst_958 ( .Q(net_6435), .D(net_6435), .SE(net_3820), .SI(net_3813), .CK(net_8651) );
CLKBUF_X2 inst_8457 ( .A(net_8418), .Z(net_8419) );
NOR2_X2 inst_2460 ( .A2(net_6184), .ZN(net_2907), .A1(net_637) );
SDFF_X2 inst_1217 ( .SI(net_7207), .Q(net_7207), .D(net_3812), .SE(net_3750), .CK(net_12132) );
CLKBUF_X2 inst_12412 ( .A(net_12373), .Z(net_12374) );
CLKBUF_X2 inst_10468 ( .A(net_8504), .Z(net_10430) );
CLKBUF_X2 inst_13465 ( .A(net_13426), .Z(net_13427) );
SDFF_X2 inst_368 ( .SI(net_7639), .Q(net_7639), .D(net_4790), .SE(net_3867), .CK(net_7992) );
CLKBUF_X2 inst_10832 ( .A(net_9564), .Z(net_10794) );
OAI21_X2 inst_1697 ( .ZN(net_5597), .A(net_5285), .B2(net_4498), .B1(net_4105) );
CLKBUF_X2 inst_10788 ( .A(net_10749), .Z(net_10750) );
CLKBUF_X2 inst_10285 ( .A(net_10246), .Z(net_10247) );
DFFR_X2 inst_6995 ( .QN(net_7704), .D(net_3358), .CK(net_10365), .RN(x1822) );
DFF_X1 inst_6938 ( .D(net_2396), .Q(net_252), .CK(net_13263) );
DFFR_X1 inst_7126 ( .Q(net_6014), .D(net_4798), .CK(net_10460), .RN(x1822) );
CLKBUF_X2 inst_10187 ( .A(net_10148), .Z(net_10149) );
INV_X2 inst_5907 ( .A(net_7473), .ZN(net_2096) );
NAND2_X2 inst_3027 ( .A1(net_7018), .ZN(net_4982), .A2(net_4979) );
NAND2_X2 inst_3689 ( .A1(net_7344), .A2(net_1798), .ZN(net_1756) );
CLKBUF_X2 inst_8614 ( .A(net_8575), .Z(net_8576) );
NAND2_X2 inst_3556 ( .ZN(net_2511), .A2(net_2052), .A1(net_1779) );
CLKBUF_X2 inst_14059 ( .A(net_14020), .Z(net_14021) );
CLKBUF_X2 inst_14016 ( .A(net_13127), .Z(net_13978) );
CLKBUF_X2 inst_10235 ( .A(net_10196), .Z(net_10197) );
AOI222_X2 inst_7480 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2143), .A1(net_2142), .B1(net_2141), .C1(net_2140) );
XNOR2_X2 inst_68 ( .ZN(net_2482), .A(net_1082), .B(net_588) );
CLKBUF_X2 inst_8811 ( .A(net_8160), .Z(net_8773) );
CLKBUF_X2 inst_8029 ( .A(net_7990), .Z(net_7991) );
OAI21_X2 inst_1966 ( .B1(net_5399), .ZN(net_5039), .A(net_4694), .B2(net_3989) );
NAND2_X2 inst_3914 ( .A1(net_6432), .A2(net_1677), .ZN(net_1392) );
SDFF_X2 inst_1253 ( .SI(net_6522), .Q(net_6522), .D(net_3802), .SE(net_3756), .CK(net_11619) );
CLKBUF_X2 inst_10913 ( .A(net_8592), .Z(net_10875) );
CLKBUF_X2 inst_11943 ( .A(net_8397), .Z(net_11905) );
CLKBUF_X2 inst_10689 ( .A(net_10650), .Z(net_10651) );
INV_X4 inst_4716 ( .ZN(net_3119), .A(net_3041) );
DFF_X1 inst_6838 ( .D(net_2509), .Q(net_179), .CK(net_12782) );
NAND3_X2 inst_2793 ( .ZN(net_2307), .A3(net_1561), .A1(net_1502), .A2(net_992) );
OAI21_X2 inst_1884 ( .ZN(net_5199), .B1(net_5198), .A(net_4574), .B2(net_3867) );
OAI21_X2 inst_2018 ( .B2(net_4497), .ZN(net_4490), .B1(net_4097), .A(net_3650) );
NOR2_X2 inst_2435 ( .ZN(net_3434), .A1(net_3050), .A2(net_3049) );
DFF_X1 inst_6488 ( .QN(net_7419), .D(net_5564), .CK(net_12127) );
CLKBUF_X2 inst_13172 ( .A(net_13133), .Z(net_13134) );
CLKBUF_X2 inst_8540 ( .A(net_8501), .Z(net_8502) );
CLKBUF_X2 inst_14078 ( .A(net_14039), .Z(net_14040) );
OAI21_X2 inst_1690 ( .B2(net_5904), .ZN(net_5604), .A(net_5306), .B1(net_4132) );
CLKBUF_X2 inst_10101 ( .A(net_8179), .Z(net_10063) );
DFF_X1 inst_6413 ( .QN(net_6160), .D(net_5757), .CK(net_11048) );
OAI221_X2 inst_1678 ( .ZN(net_3371), .A(net_3182), .B2(net_2981), .C2(net_2905), .C1(net_2861), .B1(net_1972) );
CLKBUF_X2 inst_9815 ( .A(net_9776), .Z(net_9777) );
INV_X4 inst_5312 ( .A(net_6083), .ZN(net_3538) );
CLKBUF_X2 inst_9540 ( .A(net_9501), .Z(net_9502) );
CLKBUF_X2 inst_11602 ( .A(net_7990), .Z(net_11564) );
CLKBUF_X2 inst_10839 ( .A(net_9318), .Z(net_10801) );
CLKBUF_X2 inst_13015 ( .A(net_12976), .Z(net_12977) );
SDFF_X2 inst_1287 ( .D(net_3799), .SE(net_3256), .SI(net_134), .Q(net_134), .CK(net_8471) );
NOR2_X4 inst_2233 ( .ZN(net_5665), .A1(net_5524), .A2(net_4493) );
NAND2_X1 inst_4231 ( .ZN(net_4696), .A2(net_3989), .A1(net_2165) );
AOI22_X2 inst_7266 ( .B1(net_6945), .A1(net_6913), .A2(net_5298), .B2(net_5297), .ZN(net_5284) );
CLKBUF_X2 inst_13939 ( .A(net_13900), .Z(net_13901) );
INV_X2 inst_5826 ( .ZN(net_928), .A(net_927) );
NAND2_X1 inst_4266 ( .ZN(net_4653), .A2(net_3993), .A1(net_1421) );
SDFF_X2 inst_1169 ( .D(net_7807), .SI(net_6939), .Q(net_6939), .SE(net_3734), .CK(net_8621) );
CLKBUF_X2 inst_13870 ( .A(net_13831), .Z(net_13832) );
NAND2_X2 inst_3483 ( .ZN(net_2671), .A1(net_2670), .A2(net_2669) );
INV_X4 inst_5704 ( .ZN(net_5942), .A(net_5941) );
CLKBUF_X2 inst_9440 ( .A(net_9401), .Z(net_9402) );
CLKBUF_X2 inst_8634 ( .A(net_8536), .Z(net_8596) );
SDFF_X2 inst_396 ( .SI(net_7337), .Q(net_7337), .D(net_4781), .SE(net_3856), .CK(net_12755) );
NAND2_X2 inst_3382 ( .ZN(net_3482), .A1(net_3481), .A2(net_3223) );
CLKBUF_X2 inst_12251 ( .A(net_12212), .Z(net_12213) );
NAND2_X2 inst_3377 ( .ZN(net_3492), .A1(net_3491), .A2(net_3225) );
NAND2_X4 inst_2877 ( .A1(net_4274), .ZN(net_4262), .A2(net_1677) );
CLKBUF_X2 inst_12908 ( .A(net_12869), .Z(net_12870) );
INV_X4 inst_5128 ( .ZN(net_588), .A(net_587) );
DFF_X1 inst_6514 ( .QN(net_7445), .D(net_5443), .CK(net_9296) );
CLKBUF_X2 inst_11221 ( .A(net_9168), .Z(net_11183) );
AOI222_X2 inst_7502 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2064), .A1(net_2063), .B1(net_2062), .C1(net_2061) );
CLKBUF_X2 inst_14330 ( .A(net_14291), .Z(net_14292) );
CLKBUF_X2 inst_11709 ( .A(net_11670), .Z(net_11671) );
CLKBUF_X2 inst_10371 ( .A(net_10332), .Z(net_10333) );
CLKBUF_X2 inst_11894 ( .A(net_11570), .Z(net_11856) );
CLKBUF_X2 inst_12062 ( .A(net_8257), .Z(net_12024) );
CLKBUF_X2 inst_9095 ( .A(net_9056), .Z(net_9057) );
NAND2_X4 inst_2845 ( .ZN(net_5478), .A1(net_4928), .A2(net_4926) );
OR2_X2 inst_1418 ( .ZN(net_2858), .A2(net_787), .A1(net_520) );
CLKBUF_X2 inst_14124 ( .A(net_14085), .Z(net_14086) );
CLKBUF_X2 inst_10171 ( .A(net_10132), .Z(net_10133) );
AOI21_X2 inst_7760 ( .B1(net_7134), .ZN(net_5899), .B2(net_2582), .A(net_2361) );
OAI21_X2 inst_1740 ( .ZN(net_5538), .B1(net_5537), .A(net_4807), .B2(net_4153) );
NAND2_X2 inst_2977 ( .A1(net_6748), .ZN(net_5036), .A2(net_5033) );
INV_X4 inst_5663 ( .A(net_6120), .ZN(net_3691) );
SDFF_X2 inst_1092 ( .SI(net_6951), .Q(net_6951), .D(net_3790), .SE(net_3741), .CK(net_8129) );
CLKBUF_X2 inst_11181 ( .A(net_9575), .Z(net_11143) );
CLKBUF_X2 inst_9843 ( .A(net_9804), .Z(net_9805) );
AOI222_X2 inst_7492 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2098), .A1(net_2097), .B1(net_2096), .C1(net_2095) );
CLKBUF_X2 inst_11176 ( .A(net_9383), .Z(net_11138) );
AND2_X4 inst_7822 ( .ZN(net_3118), .A2(net_3049), .A1(net_1253) );
INV_X4 inst_4836 ( .ZN(net_5102), .A(net_1074) );
OAI21_X2 inst_2001 ( .B2(net_4518), .ZN(net_4512), .B1(net_4126), .A(net_3618) );
CLKBUF_X2 inst_11784 ( .A(net_11745), .Z(net_11746) );
CLKBUF_X2 inst_10011 ( .A(net_7960), .Z(net_9973) );
CLKBUF_X2 inst_10321 ( .A(net_10282), .Z(net_10283) );
OAI221_X2 inst_1657 ( .ZN(net_4796), .A(net_4573), .C2(net_3973), .B2(net_3962), .C1(net_3764), .B1(net_1961) );
CLKBUF_X2 inst_14231 ( .A(net_14192), .Z(net_14193) );
CLKBUF_X2 inst_14385 ( .A(net_14346), .Z(net_14347) );
CLKBUF_X2 inst_12982 ( .A(net_12943), .Z(net_12944) );
CLKBUF_X2 inst_10085 ( .A(net_10046), .Z(net_10047) );
OAI21_X2 inst_2077 ( .B2(net_4415), .ZN(net_4413), .B1(net_4028), .A(net_3510) );
CLKBUF_X2 inst_12729 ( .A(net_12028), .Z(net_12691) );
CLKBUF_X2 inst_11356 ( .A(net_11317), .Z(net_11318) );
CLKBUF_X2 inst_8078 ( .A(net_8039), .Z(net_8040) );
AOI21_X2 inst_7780 ( .B1(net_6607), .ZN(net_4018), .B2(net_2583), .A(net_2316) );
INV_X4 inst_4592 ( .ZN(net_4306), .A(net_4174) );
SDFF_X2 inst_451 ( .D(net_6390), .SE(net_6050), .SI(net_300), .Q(net_300), .CK(net_14210) );
INV_X4 inst_5478 ( .A(net_6422), .ZN(net_1938) );
OAI211_X2 inst_2166 ( .B(net_2724), .ZN(net_2722), .C1(net_2299), .A(net_1671), .C2(net_1670) );
CLKBUF_X2 inst_13704 ( .A(net_13665), .Z(net_13666) );
CLKBUF_X2 inst_13930 ( .A(net_13891), .Z(net_13892) );
DFF_X1 inst_6656 ( .QN(net_7663), .D(net_5189), .CK(net_10554) );
CLKBUF_X2 inst_9910 ( .A(net_9871), .Z(net_9872) );
CLKBUF_X2 inst_12179 ( .A(net_10049), .Z(net_12141) );
SDFF_X2 inst_797 ( .SI(net_6898), .Q(net_6898), .SE(net_3887), .D(net_3798), .CK(net_8923) );
OAI22_X2 inst_1495 ( .B1(net_4666), .B2(net_4519), .A1(net_4132), .A2(net_4130), .ZN(net_4112) );
INV_X4 inst_5546 ( .ZN(net_565), .A(net_272) );
INV_X4 inst_5051 ( .ZN(net_3852), .A(net_3224) );
AOI222_X2 inst_7471 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2167), .A1(net_2166), .B1(net_2165), .C1(net_2164) );
CLKBUF_X2 inst_9310 ( .A(net_8245), .Z(net_9272) );
NAND2_X2 inst_3032 ( .A1(net_6988), .A2(net_4977), .ZN(net_4975) );
INV_X4 inst_5295 ( .A(net_6826), .ZN(net_571) );
NAND2_X2 inst_3657 ( .A1(net_7074), .ZN(net_1806), .A2(net_791) );
CLKBUF_X2 inst_8882 ( .A(net_7966), .Z(net_8844) );
AOI22_X2 inst_7319 ( .ZN(net_4573), .B2(net_3974), .A2(net_3382), .A1(net_1740), .B1(net_932) );
DFF_X1 inst_6896 ( .D(net_2512), .QN(net_176), .CK(net_12779) );
CLKBUF_X2 inst_12069 ( .A(net_8993), .Z(net_12031) );
OAI21_X2 inst_1998 ( .B2(net_4518), .ZN(net_4515), .B1(net_4135), .A(net_3474) );
DFF_X1 inst_6856 ( .D(net_2558), .Q(net_207), .CK(net_9232) );
CLKBUF_X2 inst_13195 ( .A(net_13156), .Z(net_13157) );
DFF_X1 inst_6787 ( .Q(net_7779), .D(net_4296), .CK(net_9548) );
NAND2_X2 inst_3302 ( .ZN(net_3642), .A1(net_3641), .A2(net_3229) );
CLKBUF_X2 inst_11157 ( .A(net_9581), .Z(net_11119) );
NAND2_X4 inst_2870 ( .A1(net_5882), .ZN(net_4269), .A2(net_2582) );
NAND2_X2 inst_3583 ( .ZN(net_2426), .A2(net_2425), .A1(net_868) );
CLKBUF_X2 inst_13242 ( .A(net_13203), .Z(net_13204) );
CLKBUF_X2 inst_8446 ( .A(net_8407), .Z(net_8408) );
INV_X4 inst_4933 ( .ZN(net_761), .A(net_760) );
SDFF_X2 inst_1115 ( .Q(net_7096), .D(net_3426), .SI(net_3425), .SE(net_2252), .CK(net_9326) );
DFF_X2 inst_6234 ( .Q(net_6391), .D(net_6390), .CK(net_14178) );
SDFF_X2 inst_874 ( .SI(net_7032), .Q(net_7032), .SE(net_3818), .D(net_3799), .CK(net_11935) );
NAND2_X2 inst_2976 ( .ZN(net_5037), .A2(net_4332), .A1(net_2242) );
SDFF_X2 inst_1021 ( .SI(net_6517), .Q(net_6517), .SE(net_3889), .D(net_3821), .CK(net_11234) );
OAI221_X2 inst_1681 ( .C1(net_5940), .ZN(net_3254), .B1(net_3252), .A(net_3037), .C2(net_217), .B2(net_180) );
CLKBUF_X2 inst_10222 ( .A(net_8085), .Z(net_10184) );
CLKBUF_X2 inst_9140 ( .A(net_9101), .Z(net_9102) );
NAND2_X2 inst_4204 ( .A2(net_6010), .ZN(net_1157), .A1(net_592) );
CLKBUF_X2 inst_12095 ( .A(net_12056), .Z(net_12057) );
CLKBUF_X2 inst_9173 ( .A(net_9134), .Z(net_9135) );
OAI221_X2 inst_1652 ( .ZN(net_4857), .B1(net_4855), .C2(net_4624), .B2(net_4600), .C1(net_4228), .A(net_3592) );
CLKBUF_X2 inst_9391 ( .A(net_9352), .Z(net_9353) );
INV_X4 inst_4827 ( .A(net_2853), .ZN(net_2804) );
SDFF_X2 inst_572 ( .SI(net_6513), .Q(net_6513), .D(net_3898), .SE(net_3886), .CK(net_11265) );
OAI22_X2 inst_1622 ( .B1(net_5942), .A1(net_2784), .ZN(net_2782), .B2(net_214), .A2(net_177) );
CLKBUF_X2 inst_13965 ( .A(net_9320), .Z(net_13927) );
CLKBUF_X2 inst_12699 ( .A(net_12660), .Z(net_12661) );
CLKBUF_X2 inst_12392 ( .A(net_12353), .Z(net_12354) );
OAI21_X2 inst_1735 ( .ZN(net_5552), .B1(net_5551), .A(net_4812), .B2(net_4153) );
INV_X4 inst_5036 ( .A(net_7800), .ZN(net_3890) );
SDFF_X2 inst_257 ( .Q(net_6377), .SI(net_6376), .D(net_3707), .SE(net_392), .CK(net_13509) );
OAI21_X2 inst_2050 ( .B2(net_4457), .ZN(net_4450), .B1(net_4072), .A(net_3496) );
CLKBUF_X2 inst_9516 ( .A(net_9477), .Z(net_9478) );
CLKBUF_X2 inst_12971 ( .A(net_12286), .Z(net_12933) );
INV_X4 inst_5458 ( .A(net_6094), .ZN(net_3515) );
INV_X8 inst_4555 ( .ZN(net_2200), .A(net_790) );
SDFF_X2 inst_485 ( .Q(net_6967), .D(net_6967), .SI(net_3892), .SE(net_3891), .CK(net_9127) );
CLKBUF_X2 inst_10684 ( .A(net_10645), .Z(net_10646) );
CLKBUF_X2 inst_8681 ( .A(net_8642), .Z(net_8643) );
SDFF_X2 inst_1189 ( .SI(net_7060), .Q(net_7060), .D(net_3792), .SE(net_3742), .CK(net_9063) );
SDFF_X2 inst_1205 ( .SI(net_7089), .Q(net_7089), .D(net_3821), .SE(net_3747), .CK(net_8182) );
NOR2_X2 inst_2360 ( .ZN(net_5304), .A2(net_4633), .A1(net_4505) );
CLKBUF_X2 inst_11052 ( .A(net_11013), .Z(net_11014) );
INV_X4 inst_5085 ( .A(net_7794), .ZN(net_3778) );
CLKBUF_X2 inst_11048 ( .A(net_8718), .Z(net_11010) );
XNOR2_X2 inst_33 ( .ZN(net_2477), .A(net_2476), .B(net_912) );
OAI21_X2 inst_2107 ( .ZN(net_3970), .A(net_3969), .B2(net_3873), .B1(net_884) );
CLKBUF_X2 inst_12756 ( .A(net_10694), .Z(net_12718) );
SDFF_X2 inst_232 ( .Q(net_6322), .SI(net_6321), .D(net_3641), .SE(net_392), .CK(net_14013) );
DFF_X2 inst_6253 ( .QN(net_7765), .D(net_3006), .CK(net_8015) );
CLKBUF_X2 inst_8310 ( .A(net_8271), .Z(net_8272) );
AOI222_X2 inst_7575 ( .A1(net_7246), .ZN(net_5359), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_340), .C2(net_338) );
CLKBUF_X2 inst_8641 ( .A(net_8602), .Z(net_8603) );
INV_X4 inst_4628 ( .ZN(net_4194), .A(net_4048) );
CLKBUF_X2 inst_14409 ( .A(net_14370), .Z(net_14371) );
NAND2_X2 inst_3794 ( .A1(net_7036), .A2(net_1975), .ZN(net_1551) );
CLKBUF_X2 inst_9648 ( .A(net_9137), .Z(net_9610) );
DFF_X1 inst_6929 ( .D(net_2407), .Q(net_257), .CK(net_10806) );
NAND2_X2 inst_3716 ( .A1(net_6769), .A2(net_1635), .ZN(net_1630) );
SDFF_X2 inst_253 ( .Q(net_6341), .SI(net_6340), .D(net_3593), .SE(net_392), .CK(net_13495) );
CLKBUF_X2 inst_9608 ( .A(net_9569), .Z(net_9570) );
AOI21_X2 inst_7730 ( .B1(net_6593), .ZN(net_5902), .B2(net_2583), .A(net_2280) );
CLKBUF_X2 inst_14080 ( .A(net_13269), .Z(net_14042) );
CLKBUF_X2 inst_13945 ( .A(net_13906), .Z(net_13907) );
NAND2_X2 inst_3652 ( .A1(net_7076), .ZN(net_1811), .A2(net_791) );
SDFF_X2 inst_589 ( .Q(net_6588), .D(net_6588), .SE(net_3823), .SI(net_3821), .CK(net_12031) );
INV_X4 inst_5229 ( .ZN(net_785), .A(net_467) );
CLKBUF_X2 inst_12428 ( .A(net_12389), .Z(net_12390) );
INV_X4 inst_4868 ( .ZN(net_1077), .A(net_630) );
CLKBUF_X2 inst_11969 ( .A(net_7957), .Z(net_11931) );
CLKBUF_X2 inst_10176 ( .A(net_10137), .Z(net_10138) );
INV_X4 inst_5043 ( .A(net_2887), .ZN(net_782) );
NAND2_X1 inst_4273 ( .ZN(net_4640), .A2(net_3993), .A1(net_1327) );
CLKBUF_X2 inst_9829 ( .A(net_9790), .Z(net_9791) );
CLKBUF_X2 inst_13751 ( .A(net_11880), .Z(net_13713) );
CLKBUF_X2 inst_9822 ( .A(net_9783), .Z(net_9784) );
DFF_X1 inst_6907 ( .D(net_2492), .Q(net_187), .CK(net_12399) );
CLKBUF_X2 inst_9331 ( .A(net_8133), .Z(net_9293) );
SDFF_X2 inst_602 ( .Q(net_6606), .D(net_6606), .SE(net_3830), .SI(net_3810), .CK(net_12172) );
XNOR2_X2 inst_59 ( .B(net_3985), .ZN(net_1926), .A(net_1685) );
OAI21_X2 inst_1877 ( .ZN(net_5223), .B1(net_5222), .A(net_4585), .B2(net_3867) );
NOR2_X2 inst_2367 ( .ZN(net_5269), .A2(net_4623), .A1(net_4466) );
CLKBUF_X2 inst_9182 ( .A(net_9143), .Z(net_9144) );
SDFF_X2 inst_135 ( .Q(net_6215), .SI(net_6214), .SE(net_392), .D(net_149), .CK(net_14233) );
CLKBUF_X2 inst_10533 ( .A(net_9733), .Z(net_10495) );
CLKBUF_X2 inst_10091 ( .A(net_9205), .Z(net_10053) );
NAND2_X2 inst_3256 ( .A2(net_3869), .ZN(net_3867), .A1(net_3861) );
CLKBUF_X2 inst_12867 ( .A(net_12828), .Z(net_12829) );
CLKBUF_X2 inst_11711 ( .A(net_11672), .Z(net_11673) );
CLKBUF_X2 inst_9050 ( .A(net_9011), .Z(net_9012) );
AOI21_X2 inst_7673 ( .B1(net_7008), .ZN(net_4227), .A(net_2467), .B2(net_1100) );
OAI21_X2 inst_1865 ( .ZN(net_5249), .B1(net_5204), .A(net_4534), .B2(net_3870) );
CLKBUF_X2 inst_11960 ( .A(net_11783), .Z(net_11922) );
DFF_X1 inst_6390 ( .QN(net_6121), .D(net_5698), .CK(net_8385) );
XNOR2_X2 inst_37 ( .ZN(net_2451), .A(net_1690), .B(net_426) );
OAI221_X2 inst_1664 ( .C2(net_5898), .ZN(net_4654), .B1(net_4650), .B2(net_4447), .C1(net_4080), .A(net_3531) );
CLKBUF_X2 inst_10037 ( .A(net_8000), .Z(net_9999) );
OAI22_X2 inst_1447 ( .B2(net_5907), .B1(net_4660), .A2(net_4629), .ZN(net_4627), .A1(net_4087) );
CLKBUF_X2 inst_9321 ( .A(net_9282), .Z(net_9283) );
NAND2_X2 inst_3117 ( .A1(net_6621), .A2(net_4899), .ZN(net_4884) );
INV_X2 inst_6072 ( .A(net_7759), .ZN(net_5873) );
NAND2_X2 inst_3770 ( .A1(net_7173), .A2(net_1637), .ZN(net_1575) );
CLKBUF_X2 inst_8157 ( .A(net_8118), .Z(net_8119) );
CLKBUF_X2 inst_9601 ( .A(net_9562), .Z(net_9563) );
CLKBUF_X2 inst_13863 ( .A(net_8059), .Z(net_13825) );
NAND3_X2 inst_2709 ( .ZN(net_2468), .A2(net_1805), .A3(net_1567), .A1(net_1415) );
SDFF_X2 inst_224 ( .Q(net_6330), .SI(net_6329), .D(net_3665), .SE(net_392), .CK(net_14036) );
CLKBUF_X2 inst_14003 ( .A(net_12445), .Z(net_13965) );
CLKBUF_X2 inst_9661 ( .A(net_8430), .Z(net_9623) );
INV_X4 inst_4730 ( .A(net_3200), .ZN(net_3144) );
NAND2_X2 inst_3635 ( .ZN(net_1948), .A1(net_1290), .A2(net_1132) );
INV_X4 inst_5399 ( .A(net_6071), .ZN(net_3647) );
NAND2_X2 inst_3075 ( .A1(net_6478), .ZN(net_4930), .A2(net_4927) );
INV_X4 inst_5058 ( .A(net_7819), .ZN(net_3790) );
NAND3_X2 inst_2800 ( .ZN(net_2298), .A3(net_1576), .A1(net_1330), .A2(net_982) );
CLKBUF_X2 inst_9487 ( .A(net_9448), .Z(net_9449) );
CLKBUF_X2 inst_14297 ( .A(net_14258), .Z(net_14259) );
NOR2_X2 inst_2406 ( .A2(net_7771), .A1(net_5930), .ZN(net_4001) );
SDFF_X2 inst_766 ( .Q(net_6890), .D(net_6890), .SE(net_3901), .SI(net_3821), .CK(net_11470) );
CLKBUF_X2 inst_8796 ( .A(net_8665), .Z(net_8758) );
NAND2_X2 inst_3270 ( .ZN(net_3706), .A1(net_3705), .A2(net_3225) );
OAI21_X2 inst_1908 ( .B1(net_5353), .ZN(net_5160), .A(net_4761), .B2(net_3941) );
NAND2_X2 inst_3273 ( .ZN(net_3700), .A1(net_3699), .A2(net_3231) );
SDFF_X2 inst_801 ( .Q(net_6964), .D(net_6964), .SE(net_3891), .SI(net_3797), .CK(net_9038) );
CLKBUF_X2 inst_10617 ( .A(net_7858), .Z(net_10579) );
CLKBUF_X2 inst_9943 ( .A(net_9107), .Z(net_9905) );
INV_X16 inst_6139 ( .ZN(net_1497), .A(net_786) );
SDFF_X2 inst_870 ( .SI(net_7057), .Q(net_7057), .D(net_3821), .SE(net_3777), .CK(net_8211) );
CLKBUF_X2 inst_12544 ( .A(net_10976), .Z(net_12506) );
CLKBUF_X2 inst_14282 ( .A(net_14243), .Z(net_14244) );
CLKBUF_X2 inst_9660 ( .A(net_8572), .Z(net_9622) );
XNOR2_X2 inst_11 ( .A(net_4142), .ZN(net_3825), .B(net_758) );
DFF_X1 inst_6552 ( .Q(net_7777), .D(net_5605), .CK(net_9985) );
OAI22_X2 inst_1619 ( .B1(net_5937), .ZN(net_2787), .A1(net_2786), .B2(net_210), .A2(net_173) );
NAND2_X2 inst_3110 ( .A1(net_6585), .A2(net_4897), .ZN(net_4891) );
SDFF_X2 inst_441 ( .Q(net_7393), .D(net_7393), .SE(net_3994), .SI(net_358), .CK(net_12063) );
CLKBUF_X2 inst_13468 ( .A(net_13429), .Z(net_13430) );
AOI21_X2 inst_7688 ( .B1(net_7136), .ZN(net_5909), .B2(net_2582), .A(net_2376) );
NOR2_X4 inst_2276 ( .ZN(net_3847), .A1(net_3406), .A2(net_3241) );
CLKBUF_X2 inst_8425 ( .A(net_8386), .Z(net_8387) );
DFF_X2 inst_6201 ( .QN(net_6822), .D(net_4397), .CK(net_11412) );
CLKBUF_X2 inst_11414 ( .A(net_9475), .Z(net_11376) );
CLKBUF_X2 inst_8892 ( .A(net_8490), .Z(net_8854) );
INV_X4 inst_5228 ( .A(net_841), .ZN(net_461) );
NOR2_X2 inst_2301 ( .A2(net_6186), .ZN(net_5841), .A1(net_5840) );
SDFF_X2 inst_808 ( .Q(net_6981), .D(net_6981), .SE(net_3891), .SI(net_3808), .CK(net_8083) );
CLKBUF_X2 inst_8202 ( .A(net_8000), .Z(net_8164) );
SDFF_X2 inst_557 ( .Q(net_6434), .D(net_6434), .SI(net_3894), .SE(net_3820), .CK(net_8658) );
CLKBUF_X2 inst_13639 ( .A(net_10437), .Z(net_13601) );
NAND2_X2 inst_3859 ( .A1(net_6430), .A2(net_1677), .ZN(net_1474) );
CLKBUF_X2 inst_9683 ( .A(net_9644), .Z(net_9645) );
CLKBUF_X2 inst_14300 ( .A(net_14261), .Z(net_14262) );
CLKBUF_X2 inst_11154 ( .A(net_11115), .Z(net_11116) );
OR2_X4 inst_1383 ( .ZN(net_2901), .A2(net_2752), .A1(net_289) );
NAND2_X2 inst_3279 ( .ZN(net_3688), .A1(net_3687), .A2(net_3231) );
SDFF_X2 inst_823 ( .Q(net_6969), .D(net_6969), .SE(net_3891), .SI(net_3798), .CK(net_11961) );
OAI22_X2 inst_1461 ( .B2(net_5903), .B1(net_4637), .ZN(net_4606), .A2(net_4605), .A1(net_4016) );
CLKBUF_X2 inst_8809 ( .A(net_8770), .Z(net_8771) );
INV_X1 inst_6153 ( .A(net_5857), .ZN(x124) );
NAND2_X4 inst_2838 ( .ZN(net_5550), .A1(net_5022), .A2(net_5021) );
NAND2_X2 inst_3773 ( .A1(net_7042), .A2(net_1975), .ZN(net_1572) );
NAND2_X2 inst_3423 ( .A2(net_5914), .ZN(net_3325), .A1(net_649) );
NAND2_X4 inst_2833 ( .ZN(net_5561), .A1(net_5034), .A2(net_5032) );
INV_X4 inst_4767 ( .ZN(net_2433), .A(net_1934) );
OAI21_X2 inst_2042 ( .ZN(net_4461), .B1(net_4460), .B2(net_4457), .A(net_3569) );
CLKBUF_X2 inst_10608 ( .A(net_10569), .Z(net_10570) );
CLKBUF_X2 inst_8383 ( .A(net_8344), .Z(net_8345) );
CLKBUF_X2 inst_8248 ( .A(net_8209), .Z(net_8210) );
CLKBUF_X2 inst_13154 ( .A(net_10280), .Z(net_13116) );
INV_X4 inst_5620 ( .A(net_6157), .ZN(net_3605) );
CLKBUF_X2 inst_11409 ( .A(net_9914), .Z(net_11371) );
DFFR_X2 inst_7104 ( .D(net_1959), .QN(net_126), .CK(net_12316), .RN(x1822) );
CLKBUF_X2 inst_13361 ( .A(net_13322), .Z(net_13323) );
AOI21_X2 inst_7746 ( .B1(net_6742), .ZN(net_4120), .B2(net_2581), .A(net_2315) );
INV_X4 inst_5156 ( .ZN(net_559), .A(net_558) );
CLKBUF_X2 inst_10758 ( .A(net_7962), .Z(net_10720) );
INV_X2 inst_6107 ( .A(net_7631), .ZN(net_1899) );
CLKBUF_X2 inst_9976 ( .A(net_9937), .Z(net_9938) );
CLKBUF_X2 inst_8342 ( .A(net_8303), .Z(net_8304) );
NAND3_X2 inst_2796 ( .ZN(net_2304), .A3(net_1539), .A1(net_1340), .A2(net_1032) );
CLKBUF_X2 inst_14084 ( .A(net_14045), .Z(net_14046) );
CLKBUF_X2 inst_10587 ( .A(net_10548), .Z(net_10549) );
NAND3_X2 inst_2729 ( .ZN(net_2372), .A3(net_1615), .A1(net_1467), .A2(net_1027) );
OR2_X2 inst_1413 ( .ZN(net_3767), .A2(net_795), .A1(net_446) );
CLKBUF_X2 inst_8364 ( .A(net_7885), .Z(net_8326) );
CLKBUF_X2 inst_8842 ( .A(net_8803), .Z(net_8804) );
CLKBUF_X2 inst_13320 ( .A(net_13281), .Z(net_13282) );
OAI21_X2 inst_1815 ( .ZN(net_5373), .B1(net_5347), .A(net_4340), .B2(net_3859) );
NAND2_X2 inst_3993 ( .A2(net_1910), .ZN(net_1198), .A1(net_1197) );
DFF_X1 inst_6926 ( .D(net_2398), .Q(net_238), .CK(net_10285) );
CLKBUF_X2 inst_13187 ( .A(net_13148), .Z(net_13149) );
INV_X4 inst_5267 ( .A(net_855), .ZN(net_423) );
CLKBUF_X2 inst_11140 ( .A(net_10283), .Z(net_11102) );
CLKBUF_X2 inst_10422 ( .A(net_10383), .Z(net_10384) );
CLKBUF_X2 inst_13272 ( .A(net_13233), .Z(net_13234) );
DFFR_X2 inst_7010 ( .D(net_3274), .QN(net_280), .CK(net_12650), .RN(x1822) );
OAI211_X2 inst_2169 ( .B(net_2724), .ZN(net_2713), .C2(net_2652), .A(net_2222), .C1(net_1666) );
CLKBUF_X2 inst_12379 ( .A(net_11322), .Z(net_12341) );
CLKBUF_X2 inst_11903 ( .A(net_10582), .Z(net_11865) );
SDFF_X2 inst_1326 ( .D(net_6381), .SE(net_5800), .SI(net_346), .Q(net_346), .CK(net_14134) );
CLKBUF_X2 inst_8960 ( .A(net_8921), .Z(net_8922) );
DFF_X1 inst_6708 ( .QN(net_7314), .D(net_5366), .CK(net_12710) );
CLKBUF_X2 inst_10840 ( .A(net_10801), .Z(net_10802) );
CLKBUF_X2 inst_8191 ( .A(net_8152), .Z(net_8153) );
CLKBUF_X2 inst_11920 ( .A(net_11881), .Z(net_11882) );
CLKBUF_X2 inst_10319 ( .A(net_7953), .Z(net_10281) );
INV_X4 inst_5442 ( .A(net_7406), .ZN(net_2115) );
NAND2_X1 inst_4238 ( .ZN(net_4689), .A2(net_3989), .A1(net_2120) );
CLKBUF_X2 inst_9496 ( .A(net_9457), .Z(net_9458) );
INV_X4 inst_5275 ( .ZN(net_612), .A(net_417) );
INV_X4 inst_4758 ( .ZN(net_2626), .A(net_2488) );
CLKBUF_X2 inst_9857 ( .A(net_9818), .Z(net_9819) );
NAND2_X2 inst_3875 ( .A1(net_6829), .A2(net_1521), .ZN(net_1446) );
NAND3_X2 inst_2629 ( .ZN(net_5700), .A1(net_5677), .A2(net_5311), .A3(net_4251) );
CLKBUF_X2 inst_8989 ( .A(net_8950), .Z(net_8951) );
CLKBUF_X2 inst_13658 ( .A(net_8188), .Z(net_13620) );
CLKBUF_X2 inst_9732 ( .A(net_8545), .Z(net_9694) );
CLKBUF_X2 inst_14342 ( .A(net_14303), .Z(net_14304) );
CLKBUF_X2 inst_9595 ( .A(net_9556), .Z(net_9557) );
CLKBUF_X2 inst_9197 ( .A(net_9158), .Z(net_9159) );
INV_X16 inst_6127 ( .ZN(net_4497), .A(net_3846) );
SDFFR_X2 inst_1341 ( .Q(net_7708), .D(net_7708), .SI(net_3808), .SE(net_3405), .CK(net_13191), .RN(x1822) );
OAI21_X2 inst_2154 ( .B1(net_3919), .ZN(net_2698), .A(net_2622), .B2(net_1680) );
SDFF_X2 inst_587 ( .Q(net_6586), .D(net_6586), .SE(net_3823), .SI(net_3789), .CK(net_9124) );
SDFF_X2 inst_666 ( .Q(net_6725), .D(net_6725), .SE(net_3871), .SI(net_3800), .CK(net_11392) );
CLKBUF_X2 inst_10798 ( .A(net_10759), .Z(net_10760) );
INV_X4 inst_4602 ( .ZN(net_4242), .A(net_4102) );
INV_X2 inst_5937 ( .A(net_7329), .ZN(net_1793) );
NAND3_X2 inst_2602 ( .ZN(net_5737), .A1(net_5632), .A2(net_5181), .A3(net_4197) );
OAI21_X2 inst_1829 ( .ZN(net_5352), .B1(net_5351), .A(net_4389), .B2(net_3856) );
XNOR2_X2 inst_109 ( .A(net_2567), .ZN(net_834), .B(net_833) );
SDFF_X2 inst_1182 ( .SI(net_6955), .Q(net_6955), .D(net_3801), .SE(net_3741), .CK(net_8114) );
DFF_X1 inst_6875 ( .D(net_2498), .Q(net_163), .CK(net_12238) );
DFF_X1 inst_6446 ( .QN(net_6097), .D(net_5724), .CK(net_12061) );
NAND2_X2 inst_3983 ( .ZN(net_1287), .A1(net_885), .A2(net_311) );
CLKBUF_X2 inst_9868 ( .A(net_9829), .Z(net_9830) );
AOI22_X2 inst_7368 ( .B1(net_7737), .A1(net_7708), .A2(net_5916), .B2(net_2957), .ZN(net_2954) );
CLKBUF_X2 inst_12376 ( .A(net_12337), .Z(net_12338) );
CLKBUF_X2 inst_12275 ( .A(net_12236), .Z(net_12237) );
CLKBUF_X2 inst_11019 ( .A(net_10481), .Z(net_10981) );
INV_X2 inst_5984 ( .A(net_7298), .ZN(net_2073) );
OAI22_X2 inst_1444 ( .B2(net_5896), .B1(net_4660), .ZN(net_4631), .A2(net_4629), .A1(net_4093) );
INV_X4 inst_5252 ( .ZN(net_2959), .A(net_438) );
CLKBUF_X2 inst_11993 ( .A(net_11954), .Z(net_11955) );
CLKBUF_X2 inst_11217 ( .A(net_11178), .Z(net_11179) );
AOI222_X2 inst_7594 ( .A1(net_7393), .ZN(net_5539), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_356), .C2(net_354) );
INV_X4 inst_5490 ( .A(net_7553), .ZN(net_2101) );
SDFF_X2 inst_1231 ( .SI(net_7225), .Q(net_7225), .D(net_3801), .SE(net_3751), .CK(net_10605) );
CLKBUF_X2 inst_11939 ( .A(net_11900), .Z(net_11901) );
CLKBUF_X2 inst_12210 ( .A(net_12171), .Z(net_12172) );
CLKBUF_X2 inst_13547 ( .A(net_13508), .Z(net_13509) );
SDFF_X2 inst_904 ( .SI(net_7802), .Q(net_7108), .D(net_7108), .SE(net_3888), .CK(net_13363) );
NAND2_X2 inst_3315 ( .ZN(net_3616), .A1(net_3615), .A2(net_3228) );
AOI22_X2 inst_7347 ( .B2(net_3105), .ZN(net_3103), .A2(net_2712), .A1(net_1117), .B1(net_629) );
CLKBUF_X2 inst_12100 ( .A(net_11092), .Z(net_12062) );
CLKBUF_X2 inst_10628 ( .A(net_10589), .Z(net_10590) );
CLKBUF_X2 inst_13147 ( .A(net_13108), .Z(net_13109) );
OAI21_X2 inst_2159 ( .A(net_2232), .B1(net_1920), .ZN(net_1681), .B2(net_1231) );
AOI21_X2 inst_7753 ( .B1(net_6469), .ZN(net_4051), .B2(net_2580), .A(net_2320) );
DFFR_X2 inst_7051 ( .QN(net_6022), .D(net_3135), .CK(net_8586), .RN(x1822) );
DFF_X2 inst_6266 ( .QN(net_5978), .D(net_2637), .CK(net_12530) );
NAND2_X2 inst_3923 ( .A1(net_6977), .A2(net_1833), .ZN(net_1379) );
CLKBUF_X2 inst_13094 ( .A(net_11448), .Z(net_13056) );
CLKBUF_X2 inst_11652 ( .A(net_11613), .Z(net_11614) );
INV_X4 inst_4831 ( .A(net_2704), .ZN(net_2703) );
SDFF_X2 inst_757 ( .Q(net_6880), .D(net_6880), .SE(net_3901), .SI(net_3807), .CK(net_11732) );
CLKBUF_X2 inst_10431 ( .A(net_10392), .Z(net_10393) );
SDFF_X2 inst_343 ( .SI(net_7343), .Q(net_7343), .D(net_4876), .SE(net_3856), .CK(net_9415) );
OAI22_X2 inst_1627 ( .A2(net_2820), .B2(net_2718), .ZN(net_2697), .A1(net_2274), .B1(net_579) );
INV_X4 inst_4739 ( .A(net_3087), .ZN(net_3084) );
CLKBUF_X2 inst_12670 ( .A(net_10295), .Z(net_12632) );
SDFF_X2 inst_543 ( .SI(net_6496), .Q(net_6496), .SE(net_3889), .D(net_3814), .CK(net_11270) );
SDFF_X2 inst_1106 ( .D(net_7802), .SI(net_6664), .Q(net_6664), .SE(net_3465), .CK(net_9144) );
CLKBUF_X2 inst_12131 ( .A(net_12092), .Z(net_12093) );
CLKBUF_X2 inst_14194 ( .A(net_14155), .Z(net_14156) );
CLKBUF_X2 inst_13557 ( .A(net_13518), .Z(net_13519) );
CLKBUF_X2 inst_12994 ( .A(net_12955), .Z(net_12956) );
CLKBUF_X2 inst_13122 ( .A(net_11925), .Z(net_13084) );
DFF_X1 inst_6882 ( .D(net_2526), .Q(net_232), .CK(net_12231) );
NAND2_X2 inst_3817 ( .A1(net_6641), .A2(net_1624), .ZN(net_1528) );
AOI21_X2 inst_7697 ( .B1(net_6741), .ZN(net_4122), .B2(net_2581), .A(net_2314) );
OAI21_X2 inst_2070 ( .B1(net_5900), .B2(net_4436), .ZN(net_4423), .A(net_3682) );
INV_X4 inst_5065 ( .A(net_3004), .ZN(net_716) );
SDFF_X2 inst_1256 ( .SI(net_6524), .Q(net_6524), .D(net_3799), .SE(net_3756), .CK(net_8822) );
INV_X2 inst_5765 ( .ZN(net_3023), .A(net_3022) );
NAND2_X4 inst_2890 ( .ZN(net_4080), .A2(net_3326), .A1(net_2911) );
CLKBUF_X2 inst_13858 ( .A(net_13819), .Z(net_13820) );
CLKBUF_X2 inst_9549 ( .A(net_9510), .Z(net_9511) );
CLKBUF_X2 inst_12538 ( .A(net_12499), .Z(net_12500) );
DFF_X2 inst_6337 ( .QN(net_7820), .CK(net_8233), .D(x1374) );
AOI222_X2 inst_7555 ( .A1(net_7544), .ZN(net_5198), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_376), .C2(net_374) );
OAI21_X2 inst_1903 ( .B1(net_5363), .ZN(net_5166), .A(net_4766), .B2(net_3941) );
CLKBUF_X2 inst_14254 ( .A(net_14215), .Z(net_14216) );
CLKBUF_X2 inst_9503 ( .A(net_9464), .Z(net_9465) );
CLKBUF_X2 inst_8347 ( .A(net_8010), .Z(net_8309) );
CLKBUF_X2 inst_11230 ( .A(net_11191), .Z(net_11192) );
CLKBUF_X2 inst_13716 ( .A(net_13677), .Z(net_13678) );
NAND2_X1 inst_4304 ( .ZN(net_4562), .A2(net_3866), .A1(net_1860) );
NOR2_X2 inst_2554 ( .A2(net_6034), .A1(net_6028), .ZN(net_2885) );
DFF_X1 inst_6848 ( .D(net_2561), .QN(net_214), .CK(net_9541) );
CLKBUF_X2 inst_13810 ( .A(net_13771), .Z(net_13772) );
NAND3_X2 inst_2745 ( .ZN(net_2356), .A3(net_1556), .A1(net_1444), .A2(net_1036) );
CLKBUF_X2 inst_9423 ( .A(net_9384), .Z(net_9385) );
CLKBUF_X2 inst_14422 ( .A(net_14383), .Z(net_14384) );
NAND3_X2 inst_2604 ( .ZN(net_5735), .A1(net_5630), .A2(net_5173), .A3(net_4195) );
CLKBUF_X2 inst_11802 ( .A(net_11763), .Z(net_11764) );
AOI22_X2 inst_7253 ( .B1(net_6821), .A1(net_6789), .A2(net_5316), .B2(net_5315), .ZN(net_5307) );
CLKBUF_X2 inst_13125 ( .A(net_13086), .Z(net_13087) );
CLKBUF_X2 inst_11297 ( .A(net_9063), .Z(net_11259) );
CLKBUF_X2 inst_12452 ( .A(net_12413), .Z(net_12414) );
NAND2_X1 inst_4410 ( .A2(net_5982), .A1(net_5981), .ZN(net_2882) );
SDFF_X2 inst_1244 ( .SI(net_6539), .Q(net_6539), .D(net_3807), .SE(net_3756), .CK(net_8756) );
CLKBUF_X2 inst_8134 ( .A(net_8095), .Z(net_8096) );
NAND2_X2 inst_3248 ( .ZN(net_5383), .A1(net_3857), .A2(net_3467) );
SDFF_X2 inst_582 ( .Q(net_6579), .D(net_6579), .SE(net_3823), .SI(net_3805), .CK(net_12179) );
INV_X8 inst_4515 ( .ZN(net_3815), .A(net_3176) );
CLKBUF_X2 inst_12329 ( .A(net_11156), .Z(net_12291) );
OAI21_X2 inst_2110 ( .ZN(net_3744), .B1(net_3441), .B2(net_2751), .A(net_419) );
OAI21_X2 inst_1850 ( .B1(net_5341), .ZN(net_5322), .A(net_4362), .B2(net_3853) );
NAND2_X2 inst_3477 ( .ZN(net_2860), .A2(net_2705), .A1(net_2630) );
CLKBUF_X2 inst_9774 ( .A(net_7846), .Z(net_9736) );
OAI21_X2 inst_1950 ( .B1(net_5220), .ZN(net_5070), .A(net_4727), .B2(net_3986) );
CLKBUF_X2 inst_12057 ( .A(net_12018), .Z(net_12019) );
CLKBUF_X2 inst_13896 ( .A(net_9717), .Z(net_13858) );
AOI222_X2 inst_7463 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2199), .A1(net_2198), .B1(net_2197), .C1(net_2196) );
INV_X4 inst_5287 ( .A(net_6690), .ZN(net_823) );
CLKBUF_X2 inst_9402 ( .A(net_9363), .Z(net_9364) );
AOI21_X2 inst_7690 ( .B1(net_6732), .ZN(net_4521), .B2(net_2581), .A(net_2375) );
AOI22_X2 inst_7292 ( .B1(net_6542), .A1(net_6510), .ZN(net_5186), .A2(net_5184), .B2(net_5183) );
CLKBUF_X2 inst_12914 ( .A(net_12875), .Z(net_12876) );
CLKBUF_X2 inst_12673 ( .A(net_12193), .Z(net_12635) );
OAI21_X2 inst_2057 ( .B1(net_5909), .B2(net_4457), .ZN(net_4441), .A(net_3526) );
CLKBUF_X2 inst_13408 ( .A(net_13369), .Z(net_13370) );
SDFF_X2 inst_843 ( .Q(net_7024), .D(net_7024), .SE(net_3899), .SI(net_3788), .CK(net_10864) );
OAI21_X2 inst_1779 ( .ZN(net_5415), .B1(net_5414), .A(net_4693), .B2(net_3989) );
CLKBUF_X2 inst_10710 ( .A(net_8948), .Z(net_10672) );
AOI22_X2 inst_7299 ( .B1(net_6549), .A1(net_6517), .A2(net_5184), .B2(net_5183), .ZN(net_5170) );
OAI21_X2 inst_2115 ( .ZN(net_3300), .B1(net_3299), .B2(net_3297), .A(net_3083) );
INV_X4 inst_5146 ( .ZN(net_570), .A(net_569) );
NAND2_X2 inst_3251 ( .ZN(net_5057), .A1(net_3854), .A2(net_3714) );
XNOR2_X2 inst_112 ( .ZN(net_2389), .A(net_1201), .B(net_826) );
OAI21_X2 inst_1728 ( .ZN(net_5566), .B1(net_5434), .A(net_4831), .B2(net_4153) );
SDFF_X2 inst_916 ( .Q(net_7153), .D(net_7153), .SE(net_3903), .SI(net_3804), .CK(net_11576) );
OAI21_X2 inst_1722 ( .ZN(net_5572), .B1(net_5446), .A(net_4837), .B2(net_4153) );
CLKBUF_X2 inst_11161 ( .A(net_10042), .Z(net_11123) );
INV_X4 inst_5570 ( .A(net_6068), .ZN(net_3709) );
CLKBUF_X2 inst_13799 ( .A(net_13760), .Z(net_13761) );
CLKBUF_X2 inst_9824 ( .A(net_9785), .Z(net_9786) );
CLKBUF_X2 inst_9523 ( .A(net_9484), .Z(net_9485) );
CLKBUF_X2 inst_8754 ( .A(net_8158), .Z(net_8716) );
AOI22_X2 inst_7300 ( .B1(net_6550), .A1(net_6518), .A2(net_5184), .B2(net_5183), .ZN(net_5169) );
DFF_X1 inst_6409 ( .QN(net_6156), .D(net_5761), .CK(net_9054) );
NAND2_X2 inst_3665 ( .A2(net_1798), .ZN(net_1796), .A1(net_1795) );
CLKBUF_X2 inst_8376 ( .A(net_8337), .Z(net_8338) );
AOI22_X2 inst_7441 ( .ZN(net_5414), .A2(net_1225), .B1(net_1223), .B2(net_365), .A1(net_353) );
NAND3_X2 inst_2724 ( .ZN(net_2377), .A3(net_1636), .A1(net_1491), .A2(net_1030) );
NOR2_X2 inst_2525 ( .ZN(net_2705), .A2(net_273), .A1(net_267) );
CLKBUF_X2 inst_9353 ( .A(net_9314), .Z(net_9315) );
NAND2_X2 inst_2968 ( .ZN(net_5459), .A1(net_4884), .A2(net_4883) );
CLKBUF_X2 inst_12010 ( .A(net_9594), .Z(net_11972) );
CLKBUF_X2 inst_11334 ( .A(net_11295), .Z(net_11296) );
DFFR_X2 inst_7067 ( .QN(net_6029), .D(net_3061), .CK(net_12850), .RN(x1822) );
CLKBUF_X2 inst_12875 ( .A(net_10483), .Z(net_12837) );
CLKBUF_X2 inst_7916 ( .A(net_7877), .Z(net_7878) );
NAND2_X2 inst_2964 ( .ZN(net_5463), .A1(net_4892), .A2(net_4891) );
CLKBUF_X2 inst_11760 ( .A(net_11721), .Z(net_11722) );
NAND2_X2 inst_3721 ( .A1(net_6638), .ZN(net_1625), .A2(net_1624) );
NOR2_X2 inst_2349 ( .ZN(net_5655), .A1(net_5507), .A2(net_4474) );
CLKBUF_X2 inst_8855 ( .A(net_8816), .Z(net_8817) );
SDFF_X2 inst_646 ( .SI(net_6631), .Q(net_6631), .SE(net_3851), .D(net_3814), .CK(net_12895) );
INV_X2 inst_5751 ( .ZN(net_3911), .A(net_3738) );
INV_X4 inst_5076 ( .A(net_2893), .ZN(net_793) );
DFF_X1 inst_6667 ( .QN(net_7261), .D(net_5165), .CK(net_10193) );
NAND2_X2 inst_4032 ( .A1(net_6928), .A2(net_1654), .ZN(net_1020) );
CLKBUF_X2 inst_8062 ( .A(net_7921), .Z(net_8024) );
CLKBUF_X2 inst_14310 ( .A(net_14271), .Z(net_14272) );
CLKBUF_X2 inst_10213 ( .A(net_10174), .Z(net_10175) );
NAND2_X2 inst_3169 ( .ZN(net_4764), .A2(net_3941), .A1(net_2079) );
CLKBUF_X2 inst_9387 ( .A(net_9348), .Z(net_9349) );
SDFF_X2 inst_382 ( .SI(net_7670), .Q(net_7670), .D(net_4791), .SE(net_3866), .CK(net_13235) );
CLKBUF_X2 inst_13278 ( .A(net_13239), .Z(net_13240) );
CLKBUF_X2 inst_9841 ( .A(net_9802), .Z(net_9803) );
INV_X4 inst_5344 ( .A(net_6175), .ZN(net_3711) );
NOR2_X2 inst_2329 ( .A2(net_6289), .A1(net_5840), .ZN(net_5812) );
CLKBUF_X2 inst_11119 ( .A(net_9081), .Z(net_11081) );
INV_X2 inst_6101 ( .A(net_7502), .ZN(net_2113) );
CLKBUF_X2 inst_10361 ( .A(net_10192), .Z(net_10323) );
CLKBUF_X2 inst_14248 ( .A(net_14209), .Z(net_14210) );
CLKBUF_X2 inst_9799 ( .A(net_9483), .Z(net_9761) );
INV_X2 inst_6067 ( .A(net_7757), .ZN(net_5871) );
NAND3_X2 inst_2788 ( .ZN(net_2312), .A3(net_1570), .A1(net_1423), .A2(net_974) );
CLKBUF_X2 inst_10560 ( .A(net_10521), .Z(net_10522) );
INV_X2 inst_6015 ( .A(net_7440), .ZN(net_1448) );
CLKBUF_X2 inst_11891 ( .A(net_11852), .Z(net_11853) );
DFF_X1 inst_6565 ( .QN(net_7501), .D(net_5109), .CK(net_9257) );
CLKBUF_X2 inst_10415 ( .A(net_10376), .Z(net_10377) );
SDFF_X2 inst_1049 ( .Q(net_7236), .D(net_7236), .SE(net_3822), .SI(net_332), .CK(net_12661) );
CLKBUF_X2 inst_10194 ( .A(net_10155), .Z(net_10156) );
CLKBUF_X2 inst_8418 ( .A(net_8072), .Z(net_8380) );
SDFF_X2 inst_168 ( .Q(net_6246), .SI(net_6245), .D(net_3681), .SE(net_392), .CK(net_13530) );
CLKBUF_X2 inst_9139 ( .A(net_9100), .Z(net_9101) );
INV_X4 inst_5116 ( .ZN(net_638), .A(net_601) );
CLKBUF_X2 inst_8085 ( .A(net_7833), .Z(net_8047) );
INV_X4 inst_4575 ( .ZN(net_5784), .A(net_5783) );
INV_X2 inst_6037 ( .A(net_7597), .ZN(net_1372) );
CLKBUF_X2 inst_13819 ( .A(net_13780), .Z(net_13781) );
CLKBUF_X2 inst_8688 ( .A(net_8649), .Z(net_8650) );
CLKBUF_X2 inst_10547 ( .A(net_10508), .Z(net_10509) );
SDFF_X2 inst_991 ( .Q(net_6478), .D(net_6478), .SE(net_3904), .SI(net_3804), .CK(net_8413) );
CLKBUF_X2 inst_12258 ( .A(net_12219), .Z(net_12220) );
CLKBUF_X2 inst_10642 ( .A(net_10603), .Z(net_10604) );
INV_X4 inst_5613 ( .A(net_6179), .ZN(net_3705) );
CLKBUF_X2 inst_9643 ( .A(net_9604), .Z(net_9605) );
CLKBUF_X2 inst_9249 ( .A(net_9210), .Z(net_9211) );
SDFF_X2 inst_580 ( .Q(net_6578), .D(net_6578), .SE(net_3823), .SI(net_3807), .CK(net_12184) );
SDFF_X2 inst_170 ( .Q(net_6244), .SI(net_6243), .D(net_3709), .SE(net_392), .CK(net_13972) );
CLKBUF_X2 inst_13533 ( .A(net_13494), .Z(net_13495) );
CLKBUF_X2 inst_9160 ( .A(net_9121), .Z(net_9122) );
NAND2_X2 inst_3691 ( .A1(net_7334), .A2(net_1798), .ZN(net_1753) );
CLKBUF_X2 inst_13159 ( .A(net_9990), .Z(net_13121) );
AND2_X4 inst_7823 ( .ZN(net_3117), .A2(net_3047), .A1(net_1251) );
OAI21_X2 inst_1857 ( .ZN(net_5261), .B1(net_5232), .A(net_4546), .B2(net_3870) );
CLKBUF_X2 inst_12647 ( .A(net_10576), .Z(net_12609) );
CLKBUF_X2 inst_11536 ( .A(net_11497), .Z(net_11498) );
AOI22_X2 inst_7336 ( .B2(net_3439), .ZN(net_3306), .A2(net_2712), .B1(net_1965), .A1(net_146) );
CLKBUF_X2 inst_11304 ( .A(net_10454), .Z(net_11266) );
SDFF_X2 inst_468 ( .Q(net_7547), .D(net_7547), .SE(net_3896), .SI(net_381), .CK(net_13129) );
SDFF_X2 inst_1099 ( .SI(net_6813), .Q(net_6813), .D(net_3803), .SE(net_3729), .CK(net_11314) );
DFF_X1 inst_6611 ( .QN(net_7572), .D(net_5396), .CK(net_13286) );
CLKBUF_X2 inst_9103 ( .A(net_9064), .Z(net_9065) );
CLKBUF_X2 inst_8746 ( .A(net_8665), .Z(net_8708) );
NAND2_X1 inst_4428 ( .A1(net_7605), .A2(net_2131), .ZN(net_1450) );
NAND2_X2 inst_3616 ( .ZN(net_2266), .A2(net_1936), .A1(net_1304) );
INV_X4 inst_4889 ( .A(net_2382), .ZN(net_878) );
CLKBUF_X2 inst_13842 ( .A(net_13803), .Z(net_13804) );
NOR3_X2 inst_2190 ( .ZN(net_5952), .A2(net_3952), .A3(net_3880), .A1(net_3762) );
SDFF_X2 inst_429 ( .SI(net_7756), .Q(net_7756), .SE(net_5925), .D(net_3909), .CK(net_10390) );
NAND3_X2 inst_2692 ( .ZN(net_3110), .A2(net_3109), .A3(net_3041), .A1(net_3000) );
CLKBUF_X2 inst_13580 ( .A(net_13541), .Z(net_13542) );
OAI22_X2 inst_1599 ( .A1(net_3282), .B2(net_3200), .A2(net_3144), .ZN(net_3137), .B1(net_761) );
CLKBUF_X2 inst_10298 ( .A(net_10259), .Z(net_10260) );
AND2_X4 inst_7808 ( .ZN(net_3844), .A2(net_3843), .A1(net_1140) );
INV_X4 inst_5026 ( .A(net_6688), .ZN(net_664) );
NAND2_X2 inst_3565 ( .ZN(net_2502), .A2(net_2010), .A1(net_1771) );
AOI22_X2 inst_7348 ( .B1(net_3849), .B2(net_3105), .ZN(net_3102), .A2(net_2712), .A1(net_1133) );
INV_X2 inst_5995 ( .A(net_7479), .ZN(net_2185) );
CLKBUF_X2 inst_8055 ( .A(net_8016), .Z(net_8017) );
CLKBUF_X2 inst_14141 ( .A(net_13464), .Z(net_14103) );
CLKBUF_X2 inst_7922 ( .A(net_7846), .Z(net_7884) );
INV_X4 inst_5687 ( .A(net_6070), .ZN(net_3681) );
CLKBUF_X2 inst_13824 ( .A(net_13785), .Z(net_13786) );
CLKBUF_X2 inst_13567 ( .A(net_13528), .Z(net_13529) );
DFFR_X2 inst_6960 ( .QN(net_7722), .D(net_5777), .CK(net_10378), .RN(x1822) );
CLKBUF_X2 inst_8629 ( .A(net_8590), .Z(net_8591) );
NAND2_X2 inst_3977 ( .ZN(net_1293), .A1(net_885), .A2(net_318) );
NAND2_X2 inst_3467 ( .A2(net_2957), .ZN(net_2758), .A1(net_2757) );
NAND3_X2 inst_2593 ( .ZN(net_5746), .A1(net_5641), .A2(net_5224), .A3(net_4205) );
NAND2_X2 inst_3064 ( .A1(net_7159), .A2(net_4954), .ZN(net_4941) );
CLKBUF_X2 inst_11717 ( .A(net_11678), .Z(net_11679) );
NAND2_X2 inst_3676 ( .A1(net_7340), .A2(net_1798), .ZN(net_1780) );
CLKBUF_X2 inst_9850 ( .A(net_8522), .Z(net_9812) );
INV_X4 inst_5021 ( .ZN(net_876), .A(net_792) );
CLKBUF_X2 inst_13550 ( .A(net_13511), .Z(net_13512) );
SDFF_X2 inst_318 ( .SI(net_7461), .Q(net_7461), .D(net_5100), .SE(net_3993), .CK(net_9707) );
CLKBUF_X2 inst_7948 ( .A(net_7908), .Z(net_7910) );
NAND2_X2 inst_4033 ( .A1(net_6793), .A2(net_1651), .ZN(net_1019) );
CLKBUF_X2 inst_14210 ( .A(net_14171), .Z(net_14172) );
CLKBUF_X2 inst_8538 ( .A(net_8499), .Z(net_8500) );
INV_X4 inst_5044 ( .A(net_3234), .ZN(net_649) );
NAND2_X4 inst_2899 ( .A1(net_5914), .ZN(net_3403), .A2(net_462) );
NAND2_X2 inst_4065 ( .A1(net_6671), .A2(net_1655), .ZN(net_987) );
CLKBUF_X2 inst_13790 ( .A(net_13751), .Z(net_13752) );
OAI22_X2 inst_1486 ( .B1(net_4666), .B2(net_4135), .A1(net_4132), .ZN(net_4129), .A2(net_4128) );
CLKBUF_X2 inst_13449 ( .A(net_13410), .Z(net_13411) );
NOR2_X4 inst_2281 ( .ZN(net_3837), .A1(net_3399), .A2(net_3243) );
SDFF_X2 inst_1175 ( .SI(net_6946), .Q(net_6946), .D(net_3836), .SE(net_3741), .CK(net_8124) );
CLKBUF_X2 inst_12666 ( .A(net_9288), .Z(net_12628) );
CLKBUF_X2 inst_13929 ( .A(net_13890), .Z(net_13891) );
CLKBUF_X2 inst_14222 ( .A(net_10702), .Z(net_14184) );
INV_X2 inst_5877 ( .A(net_6016), .ZN(net_2612) );
INV_X4 inst_5256 ( .ZN(net_633), .A(net_435) );
NAND2_X2 inst_4096 ( .A1(net_6663), .A2(net_1655), .ZN(net_956) );
CLKBUF_X2 inst_12208 ( .A(net_10756), .Z(net_12170) );
CLKBUF_X2 inst_12164 ( .A(net_12125), .Z(net_12126) );
CLKBUF_X2 inst_8305 ( .A(net_7857), .Z(net_8267) );
CLKBUF_X2 inst_8962 ( .A(net_7995), .Z(net_8924) );
INV_X8 inst_4509 ( .ZN(net_3889), .A(net_3257) );
SDFF_X2 inst_395 ( .SI(net_7336), .Q(net_7336), .D(net_4782), .SE(net_3856), .CK(net_9914) );
CLKBUF_X2 inst_14106 ( .A(net_14067), .Z(net_14068) );
CLKBUF_X2 inst_10927 ( .A(net_10149), .Z(net_10889) );
DFF_X1 inst_6808 ( .D(net_3754), .CK(net_10418), .Q(x315) );
SDFF_X2 inst_841 ( .Q(net_7022), .D(net_7022), .SE(net_3899), .SI(net_3790), .CK(net_11000) );
NAND2_X2 inst_3963 ( .A1(net_6835), .A2(net_1521), .ZN(net_1319) );
CLKBUF_X2 inst_13682 ( .A(net_13643), .Z(net_13644) );
CLKBUF_X2 inst_12508 ( .A(net_12469), .Z(net_12470) );
AOI22_X2 inst_7328 ( .A2(net_3435), .B2(net_3434), .ZN(net_3418), .B1(net_2565), .A1(net_1254) );
SDFF_X2 inst_689 ( .Q(net_6755), .D(net_6755), .SI(net_3821), .SE(net_3815), .CK(net_11332) );
CLKBUF_X2 inst_13412 ( .A(net_13201), .Z(net_13374) );
NAND2_X1 inst_4453 ( .A2(net_1256), .ZN(net_1124), .A1(net_1123) );
NAND3_X2 inst_2689 ( .ZN(net_3153), .A2(net_3152), .A3(net_3049), .A1(net_2999) );
CLKBUF_X2 inst_13538 ( .A(net_12133), .Z(net_13500) );
DFF_X1 inst_6361 ( .QN(net_6221), .D(net_5823), .CK(net_14122) );
INV_X4 inst_4895 ( .A(net_3852), .ZN(net_3042) );
NAND2_X2 inst_3896 ( .A1(net_6428), .A2(net_1677), .ZN(net_1418) );
CLKBUF_X2 inst_9622 ( .A(net_9583), .Z(net_9584) );
OAI22_X2 inst_1558 ( .B2(net_3405), .A2(net_3360), .ZN(net_3347), .A1(net_3282), .B1(net_436) );
NAND2_X2 inst_3679 ( .A2(net_1798), .ZN(net_1775), .A1(net_1774) );
CLKBUF_X2 inst_14212 ( .A(net_14173), .Z(net_14174) );
CLKBUF_X2 inst_12630 ( .A(net_12591), .Z(net_12592) );
NAND2_X4 inst_2906 ( .ZN(net_1864), .A2(net_1672), .A1(net_1657) );
DFF_X2 inst_6272 ( .QN(net_5920), .D(net_390), .CK(net_12772) );
INV_X2 inst_5848 ( .ZN(net_701), .A(net_700) );
CLKBUF_X2 inst_14206 ( .A(net_14167), .Z(net_14168) );
CLKBUF_X2 inst_13398 ( .A(net_13359), .Z(net_13360) );
CLKBUF_X2 inst_12836 ( .A(net_9038), .Z(net_12798) );
NAND2_X2 inst_3886 ( .A1(net_6697), .A2(net_1497), .ZN(net_1433) );
CLKBUF_X2 inst_13587 ( .A(net_13548), .Z(net_13549) );
CLKBUF_X2 inst_9072 ( .A(net_8251), .Z(net_9034) );
CLKBUF_X2 inst_8797 ( .A(net_8344), .Z(net_8759) );
CLKBUF_X2 inst_8685 ( .A(net_8012), .Z(net_8647) );
OAI22_X2 inst_1615 ( .A1(net_3275), .A2(net_3087), .B2(net_3084), .ZN(net_3056), .B1(net_3055) );
CLKBUF_X2 inst_13201 ( .A(net_11438), .Z(net_13163) );
CLKBUF_X2 inst_9148 ( .A(net_9109), .Z(net_9110) );
CLKBUF_X2 inst_11692 ( .A(net_11653), .Z(net_11654) );
CLKBUF_X2 inst_11434 ( .A(net_11395), .Z(net_11396) );
CLKBUF_X2 inst_9505 ( .A(net_8338), .Z(net_9467) );
AOI222_X2 inst_7503 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2060), .A1(net_2059), .B1(net_2058), .C1(net_2057) );
CLKBUF_X2 inst_10643 ( .A(net_8815), .Z(net_10605) );
CLKBUF_X2 inst_12406 ( .A(net_8270), .Z(net_12368) );
CLKBUF_X2 inst_11510 ( .A(net_11471), .Z(net_11472) );
CLKBUF_X2 inst_13760 ( .A(net_13721), .Z(net_13722) );
CLKBUF_X2 inst_9890 ( .A(net_9851), .Z(net_9852) );
CLKBUF_X2 inst_8313 ( .A(net_7929), .Z(net_8275) );
OAI21_X2 inst_2145 ( .B1(net_5778), .ZN(net_2799), .A(net_2674), .B2(net_2672) );
SDFF_X2 inst_709 ( .SI(net_6781), .Q(net_6781), .SE(net_3872), .D(net_3780), .CK(net_11326) );
NOR2_X2 inst_2375 ( .ZN(net_5154), .A2(net_4609), .A1(net_4425) );
CLKBUF_X2 inst_12127 ( .A(net_9190), .Z(net_12089) );
INV_X2 inst_5725 ( .ZN(net_4003), .A(net_3910) );
SDFF_X2 inst_920 ( .Q(net_7158), .D(net_7158), .SE(net_3903), .SI(net_3794), .CK(net_8702) );
NAND2_X2 inst_3454 ( .A2(net_5925), .ZN(net_2918), .A1(net_1826) );
DFF_X2 inst_6298 ( .QN(net_5969), .D(net_1663), .CK(net_11404) );
INV_X2 inst_5741 ( .ZN(net_3724), .A(net_3424) );
CLKBUF_X2 inst_13400 ( .A(net_13361), .Z(net_13362) );
DFF_X1 inst_6571 ( .QN(net_7552), .D(net_5083), .CK(net_12274) );
CLKBUF_X2 inst_12080 ( .A(net_11127), .Z(net_12042) );
CLKBUF_X2 inst_9956 ( .A(net_9917), .Z(net_9918) );
CLKBUF_X2 inst_12517 ( .A(net_8189), .Z(net_12479) );
CLKBUF_X2 inst_12331 ( .A(net_12292), .Z(net_12293) );
CLKBUF_X2 inst_12106 ( .A(net_12067), .Z(net_12068) );
AOI22_X2 inst_7389 ( .A2(net_5916), .B2(net_2957), .ZN(net_2930), .B1(net_2647), .A1(net_713) );
INV_X4 inst_4610 ( .ZN(net_4234), .A(net_4086) );
CLKBUF_X2 inst_13350 ( .A(net_13311), .Z(net_13312) );
CLKBUF_X2 inst_11629 ( .A(net_9929), .Z(net_11591) );
INV_X2 inst_6116 ( .A(net_5932), .ZN(net_5931) );
NAND2_X1 inst_4403 ( .A2(net_3297), .ZN(net_3074), .A1(net_3073) );
CLKBUF_X2 inst_13797 ( .A(net_9471), .Z(net_13759) );
CLKBUF_X2 inst_14203 ( .A(net_14164), .Z(net_14165) );
NAND2_X4 inst_2889 ( .ZN(net_4057), .A2(net_3328), .A1(net_3093) );
CLKBUF_X2 inst_11432 ( .A(net_7911), .Z(net_11394) );
CLKBUF_X2 inst_11380 ( .A(net_10247), .Z(net_11342) );
CLKBUF_X2 inst_10109 ( .A(net_7909), .Z(net_10071) );
CLKBUF_X2 inst_9885 ( .A(net_9846), .Z(net_9847) );
CLKBUF_X2 inst_13743 ( .A(net_13704), .Z(net_13705) );
CLKBUF_X2 inst_8034 ( .A(net_7995), .Z(net_7996) );
NOR3_X2 inst_2189 ( .ZN(net_5950), .A2(net_3953), .A3(net_3881), .A1(net_3765) );
INV_X4 inst_5448 ( .A(net_6097), .ZN(net_3509) );
NAND2_X2 inst_4198 ( .A2(net_5936), .ZN(net_2735), .A1(net_769) );
SDFF_X2 inst_315 ( .SI(net_7457), .Q(net_7457), .D(net_5103), .SE(net_3993), .CK(net_12449) );
NAND2_X2 inst_2935 ( .ZN(net_5512), .A1(net_4985), .A2(net_4984) );
CLKBUF_X2 inst_13176 ( .A(net_13137), .Z(net_13138) );
AOI21_X2 inst_7653 ( .B2(net_3439), .ZN(net_3393), .A(net_3209), .B1(net_3075) );
SDFF_X2 inst_216 ( .Q(net_6338), .SI(net_6337), .D(net_3649), .SE(net_392), .CK(net_14062) );
NAND2_X2 inst_3369 ( .ZN(net_3508), .A1(net_3507), .A2(net_3223) );
CLKBUF_X2 inst_8992 ( .A(net_8536), .Z(net_8954) );
CLKBUF_X2 inst_13612 ( .A(net_13573), .Z(net_13574) );
CLKBUF_X2 inst_10924 ( .A(net_10885), .Z(net_10886) );
CLKBUF_X2 inst_14444 ( .A(net_10827), .Z(net_14406) );
CLKBUF_X2 inst_13099 ( .A(net_9730), .Z(net_13061) );
CLKBUF_X2 inst_12987 ( .A(net_12948), .Z(net_12949) );
CLKBUF_X2 inst_9202 ( .A(net_9163), .Z(net_9164) );
OAI21_X2 inst_2060 ( .B2(net_4436), .ZN(net_4435), .B1(net_4061), .A(net_3551) );
CLKBUF_X2 inst_10179 ( .A(net_10140), .Z(net_10141) );
CLKBUF_X2 inst_8771 ( .A(net_8662), .Z(net_8733) );
NAND3_X2 inst_2680 ( .ZN(net_3335), .A3(net_3102), .A1(net_2854), .A2(net_2769) );
SDFF_X2 inst_415 ( .D(net_6392), .SE(net_5801), .SI(net_337), .Q(net_337), .CK(net_14314) );
CLKBUF_X2 inst_10592 ( .A(net_10539), .Z(net_10554) );
AOI22_X2 inst_7321 ( .ZN(net_4550), .B2(net_3970), .A2(net_3377), .A1(net_1264), .B1(net_928) );
CLKBUF_X2 inst_9225 ( .A(net_9156), .Z(net_9187) );
CLKBUF_X2 inst_12005 ( .A(net_7887), .Z(net_11967) );
CLKBUF_X2 inst_7866 ( .A(net_7825), .Z(net_7828) );
OAI21_X2 inst_1795 ( .ZN(net_5395), .A(net_4722), .B2(net_3986), .B1(net_1265) );
AOI21_X2 inst_7652 ( .B2(net_3439), .ZN(net_3394), .A(net_3214), .B1(net_285) );
AOI22_X2 inst_7291 ( .B1(net_7216), .A1(net_7184), .A2(net_5244), .B2(net_5243), .ZN(net_5210) );
SDFF_X2 inst_828 ( .Q(net_7007), .D(net_7007), .SE(net_3899), .SI(net_3813), .CK(net_10867) );
INV_X4 inst_4697 ( .A(net_5968), .ZN(net_3366) );
CLKBUF_X2 inst_9074 ( .A(net_9035), .Z(net_9036) );
DFF_X2 inst_6278 ( .D(net_2614), .QN(net_266), .CK(net_10783) );
CLKBUF_X2 inst_13522 ( .A(net_13483), .Z(net_13484) );
NAND2_X2 inst_4164 ( .ZN(net_931), .A1(net_514), .A2(net_439) );
CLKBUF_X2 inst_10869 ( .A(net_9423), .Z(net_10831) );
CLKBUF_X2 inst_14185 ( .A(net_14146), .Z(net_14147) );
CLKBUF_X2 inst_10408 ( .A(net_8664), .Z(net_10370) );
OAI22_X2 inst_1561 ( .B2(net_3405), .A2(net_3360), .ZN(net_3344), .A1(net_3111), .B1(net_512) );
CLKBUF_X2 inst_8899 ( .A(net_8860), .Z(net_8861) );
CLKBUF_X2 inst_13919 ( .A(net_9731), .Z(net_13881) );
OAI21_X2 inst_2104 ( .ZN(net_3976), .A(net_3975), .B2(net_3876), .B1(net_725) );
CLKBUF_X2 inst_12190 ( .A(net_12151), .Z(net_12152) );
CLKBUF_X2 inst_8052 ( .A(net_8013), .Z(net_8014) );
CLKBUF_X2 inst_12437 ( .A(net_12398), .Z(net_12399) );
CLKBUF_X2 inst_10854 ( .A(net_7954), .Z(net_10816) );
CLKBUF_X2 inst_9530 ( .A(net_9491), .Z(net_9492) );
NAND3_X2 inst_2573 ( .ZN(net_5766), .A1(net_5661), .A2(net_5289), .A3(net_4235) );
CLKBUF_X2 inst_8762 ( .A(net_8723), .Z(net_8724) );
AOI21_X2 inst_7733 ( .B1(net_6460), .ZN(net_5910), .B2(net_2580), .A(net_2306) );
AOI22_X2 inst_7382 ( .A2(net_5916), .B2(net_2957), .ZN(net_2939), .B1(net_2938), .A1(net_859) );
DFF_X2 inst_6182 ( .QN(net_6553), .D(net_5450), .CK(net_7936) );
CLKBUF_X2 inst_8749 ( .A(net_8710), .Z(net_8711) );
DFF_X2 inst_6233 ( .QN(net_6063), .D(net_3456), .CK(net_13205) );
DFF_X2 inst_6240 ( .QN(net_7531), .D(net_3034), .CK(net_9509) );
CLKBUF_X2 inst_11426 ( .A(net_9006), .Z(net_11388) );
CLKBUF_X2 inst_9629 ( .A(net_8128), .Z(net_9591) );
CLKBUF_X2 inst_10127 ( .A(net_10088), .Z(net_10089) );
CLKBUF_X2 inst_10794 ( .A(net_8918), .Z(net_10756) );
CLKBUF_X2 inst_9137 ( .A(net_9098), .Z(net_9099) );
OAI21_X2 inst_2096 ( .B2(net_4426), .ZN(net_4320), .B1(net_4057), .A(net_3586) );
CLKBUF_X2 inst_10169 ( .A(net_10130), .Z(net_10131) );
SDFF_X2 inst_552 ( .SI(net_7807), .Q(net_6438), .D(net_6438), .SE(net_3820), .CK(net_8661) );
CLKBUF_X2 inst_10951 ( .A(net_10912), .Z(net_10913) );
NAND2_X2 inst_3050 ( .A1(net_6985), .A2(net_4977), .ZN(net_4957) );
INV_X4 inst_4793 ( .ZN(net_4782), .A(net_1267) );
CLKBUF_X2 inst_11349 ( .A(net_11310), .Z(net_11311) );
INV_X4 inst_4997 ( .A(net_784), .ZN(net_694) );
CLKBUF_X2 inst_13916 ( .A(net_13877), .Z(net_13878) );
CLKBUF_X2 inst_8491 ( .A(net_8452), .Z(net_8453) );
CLKBUF_X2 inst_12483 ( .A(net_12444), .Z(net_12445) );
NAND2_X2 inst_3913 ( .A1(net_6844), .A2(net_1521), .ZN(net_1393) );
OAI22_X2 inst_1564 ( .A2(net_3297), .ZN(net_3290), .A1(net_3289), .B2(net_3286), .B1(net_749) );
INV_X2 inst_5807 ( .A(net_1692), .ZN(net_1210) );
DFFR_X2 inst_6985 ( .QN(net_6038), .D(net_3444), .CK(net_12566), .RN(x1822) );
CLKBUF_X2 inst_12625 ( .A(net_12586), .Z(net_12587) );
CLKBUF_X2 inst_10995 ( .A(net_10956), .Z(net_10957) );
AOI222_X2 inst_7484 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2126), .A1(net_2125), .B1(net_2124), .C1(net_2123) );
OAI21_X2 inst_1941 ( .B1(net_5537), .ZN(net_5092), .A(net_4736), .B2(net_3988) );
DFF_X1 inst_6477 ( .QN(net_6090), .D(net_5582), .CK(net_12953) );
DFF_X2 inst_6247 ( .QN(net_7751), .D(net_3027), .CK(net_12538) );
CLKBUF_X2 inst_8064 ( .A(net_8005), .Z(net_8026) );
XNOR2_X2 inst_9 ( .A(net_4144), .ZN(net_3827), .B(net_747) );
CLKBUF_X2 inst_9492 ( .A(net_9453), .Z(net_9454) );
SDFF_X2 inst_356 ( .SI(net_7609), .Q(net_7609), .D(net_4797), .SE(net_3870), .CK(net_13259) );
CLKBUF_X2 inst_9311 ( .A(net_9272), .Z(net_9273) );
NAND2_X2 inst_3358 ( .ZN(net_3529), .A1(net_3528), .A2(net_3226) );
DFF_X1 inst_6719 ( .QN(net_7320), .D(net_5342), .CK(net_10142) );
INV_X4 inst_5587 ( .A(net_7552), .ZN(net_2129) );
CLKBUF_X2 inst_10735 ( .A(net_10696), .Z(net_10697) );
DFF_X1 inst_6884 ( .D(net_2511), .QN(net_173), .CK(net_9952) );
OAI22_X2 inst_1594 ( .A1(net_3293), .B2(net_3200), .ZN(net_3145), .A2(net_3144), .B1(net_607) );
CLKBUF_X2 inst_9267 ( .A(net_9228), .Z(net_9229) );
SDFF_X2 inst_902 ( .SI(net_7799), .Q(net_7105), .D(net_7105), .SE(net_3888), .CK(net_8712) );
CLKBUF_X2 inst_9105 ( .A(net_8707), .Z(net_9067) );
CLKBUF_X2 inst_12224 ( .A(net_12185), .Z(net_12186) );
NAND2_X2 inst_3489 ( .A2(net_2724), .ZN(net_2653), .A1(net_2652) );
SDFF_X2 inst_778 ( .SI(net_6906), .Q(net_6906), .SE(net_3887), .D(net_3811), .CK(net_8872) );
NAND2_X1 inst_4286 ( .ZN(net_4581), .A2(net_3867), .A1(net_1186) );
CLKBUF_X2 inst_10118 ( .A(net_9361), .Z(net_10080) );
OAI21_X2 inst_1935 ( .B1(net_5554), .ZN(net_5110), .A(net_4742), .B2(net_3988) );
INV_X2 inst_6032 ( .ZN(net_400), .A(x940) );
CLKBUF_X2 inst_9332 ( .A(net_9293), .Z(net_9294) );
CLKBUF_X2 inst_7912 ( .A(net_7873), .Z(net_7874) );
CLKBUF_X2 inst_8678 ( .A(net_8639), .Z(net_8640) );
CLKBUF_X2 inst_8235 ( .A(net_8196), .Z(net_8197) );
CLKBUF_X2 inst_11486 ( .A(net_11447), .Z(net_11448) );
CLKBUF_X2 inst_13884 ( .A(net_13845), .Z(net_13846) );
CLKBUF_X2 inst_8845 ( .A(net_8806), .Z(net_8807) );
AND2_X4 inst_7810 ( .ZN(net_3840), .A2(net_3839), .A1(net_1146) );
OAI21_X2 inst_2140 ( .A(net_5924), .ZN(net_2808), .B1(net_2807), .B2(net_2806) );
CLKBUF_X2 inst_8353 ( .A(net_8314), .Z(net_8315) );
CLKBUF_X2 inst_9641 ( .A(net_9602), .Z(net_9603) );
CLKBUF_X2 inst_12855 ( .A(net_12816), .Z(net_12817) );
CLKBUF_X2 inst_13895 ( .A(net_13856), .Z(net_13857) );
SDFF_X2 inst_781 ( .SI(net_6909), .Q(net_6909), .SE(net_3887), .D(net_3786), .CK(net_8497) );
CLKBUF_X2 inst_11386 ( .A(net_10725), .Z(net_11348) );
CLKBUF_X2 inst_12033 ( .A(net_11994), .Z(net_11995) );
CLKBUF_X2 inst_12368 ( .A(net_11177), .Z(net_12330) );
NAND2_X2 inst_4042 ( .A1(net_6944), .A2(net_1654), .ZN(net_1010) );
CLKBUF_X2 inst_13409 ( .A(net_13370), .Z(net_13371) );
AOI21_X2 inst_7629 ( .ZN(net_4259), .A(net_4258), .B1(net_4257), .B2(net_4001) );
CLKBUF_X2 inst_9450 ( .A(net_9411), .Z(net_9412) );
NAND2_X2 inst_3696 ( .ZN(net_1734), .A1(net_1282), .A2(net_1095) );
CLKBUF_X2 inst_9499 ( .A(net_9460), .Z(net_9461) );
CLKBUF_X2 inst_13120 ( .A(net_13081), .Z(net_13082) );
CLKBUF_X2 inst_9971 ( .A(net_9932), .Z(net_9933) );
DFFR_X2 inst_7053 ( .QN(net_6023), .D(net_3197), .CK(net_8583), .RN(x1822) );
OAI22_X2 inst_1559 ( .B2(net_3405), .A2(net_3360), .ZN(net_3346), .A1(net_3280), .B1(net_521) );
OAI21_X2 inst_1928 ( .ZN(net_5117), .A(net_4753), .B2(net_3941), .B1(net_1168) );
OAI21_X2 inst_1967 ( .ZN(net_4873), .B1(net_4872), .A(net_4343), .B2(net_3859) );
CLKBUF_X2 inst_8830 ( .A(net_8791), .Z(net_8792) );
CLKBUF_X2 inst_13733 ( .A(net_10903), .Z(net_13695) );
DFF_X1 inst_6752 ( .QN(net_7667), .D(net_4841), .CK(net_8325) );
INV_X8 inst_4485 ( .ZN(net_4272), .A(net_3923) );
SDFF_X2 inst_927 ( .Q(net_7136), .D(net_7136), .SE(net_3903), .SI(net_3798), .CK(net_13348) );
CLKBUF_X2 inst_12944 ( .A(net_12905), .Z(net_12906) );
AOI21_X2 inst_7659 ( .ZN(net_5958), .B2(net_3439), .A(net_3212), .B1(net_1220) );
CLKBUF_X2 inst_13304 ( .A(net_13265), .Z(net_13266) );
AOI22_X2 inst_7420 ( .A1(net_2970), .ZN(net_2773), .B1(net_2772), .A2(net_238), .B2(net_164) );
CLKBUF_X2 inst_13258 ( .A(net_13219), .Z(net_13220) );
CLKBUF_X2 inst_10967 ( .A(net_10928), .Z(net_10929) );
XNOR2_X2 inst_73 ( .ZN(net_1935), .B(net_670), .A(net_666) );
OAI22_X2 inst_1488 ( .B1(net_4666), .A1(net_4132), .B2(net_4128), .ZN(net_4125), .A2(net_4124) );
OAI21_X2 inst_1719 ( .ZN(net_5575), .B1(net_5539), .A(net_4685), .B2(net_3989) );
OAI21_X2 inst_1947 ( .B1(net_5227), .ZN(net_5073), .A(net_4730), .B2(net_3986) );
CLKBUF_X2 inst_8030 ( .A(net_7991), .Z(net_7992) );
AOI22_X2 inst_7318 ( .ZN(net_4590), .B2(net_3976), .A2(net_3384), .A1(net_1158), .B1(net_926) );
DFF_X2 inst_6285 ( .D(net_2415), .QN(net_226), .CK(net_12594) );
INV_X4 inst_4690 ( .ZN(net_4144), .A(net_3331) );
CLKBUF_X2 inst_9236 ( .A(net_9197), .Z(net_9198) );
SDFF_X2 inst_890 ( .Q(net_7121), .D(net_7121), .SE(net_3888), .SI(net_3804), .CK(net_11590) );
CLKBUF_X2 inst_12510 ( .A(net_12471), .Z(net_12472) );
CLKBUF_X2 inst_12352 ( .A(net_12313), .Z(net_12314) );
OAI21_X2 inst_1851 ( .B1(net_5339), .ZN(net_5321), .A(net_4361), .B2(net_3853) );
INV_X2 inst_5911 ( .A(net_7297), .ZN(net_2053) );
INV_X4 inst_4585 ( .A(net_5040), .ZN(net_4327) );
CLKBUF_X2 inst_12896 ( .A(net_12857), .Z(net_12858) );
CLKBUF_X2 inst_8105 ( .A(net_8066), .Z(net_8067) );
INV_X8 inst_4514 ( .ZN(net_3888), .A(net_3207) );
DFF_X1 inst_6903 ( .D(net_2506), .QN(net_184), .CK(net_12411) );
CLKBUF_X2 inst_9539 ( .A(net_9500), .Z(net_9501) );
CLKBUF_X2 inst_9126 ( .A(net_8447), .Z(net_9088) );
SDFF_X2 inst_1168 ( .SI(net_6938), .Q(net_6938), .D(net_3811), .SE(net_3734), .CK(net_8622) );
CLKBUF_X2 inst_12963 ( .A(net_12924), .Z(net_12925) );
CLKBUF_X2 inst_11294 ( .A(net_11255), .Z(net_11256) );
AOI222_X2 inst_7573 ( .A1(net_7546), .ZN(net_5237), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_378), .C2(net_376) );
SDFF_X2 inst_659 ( .Q(net_6717), .D(net_6717), .SE(net_3871), .SI(net_3782), .CK(net_11752) );
AOI21_X2 inst_7681 ( .B1(net_7014), .ZN(net_4216), .A(net_2458), .B2(net_1100) );
DFF_X1 inst_6890 ( .D(net_2525), .Q(net_233), .CK(net_9428) );
CLKBUF_X2 inst_12868 ( .A(net_11369), .Z(net_12830) );
CLKBUF_X2 inst_11747 ( .A(net_10665), .Z(net_11709) );
CLKBUF_X2 inst_12883 ( .A(net_12844), .Z(net_12845) );
NAND2_X1 inst_4363 ( .ZN(net_4364), .A2(net_3853), .A1(net_2008) );
SDFF_X2 inst_1161 ( .D(net_7799), .SI(net_6796), .Q(net_6796), .SE(net_3729), .CK(net_11062) );
NAND2_X2 inst_3362 ( .ZN(net_3522), .A1(net_3521), .A2(net_3225) );
INV_X4 inst_5273 ( .ZN(net_707), .A(net_608) );
CLKBUF_X2 inst_8094 ( .A(net_8055), .Z(net_8056) );
INV_X4 inst_5505 ( .A(net_6040), .ZN(net_2839) );
CLKBUF_X2 inst_10289 ( .A(net_9718), .Z(net_10251) );
NAND2_X2 inst_3199 ( .ZN(net_4727), .A2(net_3986), .A1(net_1845) );
DFF_X2 inst_6178 ( .QN(net_6688), .D(net_5455), .CK(net_9730) );
NAND2_X2 inst_3612 ( .ZN(net_2270), .A2(net_1932), .A1(net_1306) );
OAI22_X2 inst_1581 ( .B2(net_3200), .ZN(net_3199), .A1(net_3198), .A2(net_3196), .B1(net_443) );
CLKBUF_X2 inst_14096 ( .A(net_13992), .Z(net_14058) );
CLKBUF_X2 inst_10703 ( .A(net_10664), .Z(net_10665) );
NOR2_X2 inst_2388 ( .ZN(net_4292), .A1(net_4142), .A2(net_4141) );
NOR2_X2 inst_2312 ( .A2(net_6202), .A1(net_5843), .ZN(net_5829) );
INV_X4 inst_5633 ( .A(net_5988), .ZN(net_427) );
INV_X4 inst_5336 ( .A(net_6042), .ZN(net_2911) );
NAND2_X1 inst_4309 ( .ZN(net_4557), .A2(net_3866), .A1(net_1978) );
CLKBUF_X2 inst_11642 ( .A(net_11603), .Z(net_11604) );
NAND2_X2 inst_3500 ( .A2(net_2714), .ZN(net_2618), .A1(net_405) );
NAND3_X2 inst_2634 ( .ZN(net_5695), .A1(net_5672), .A2(net_5302), .A3(net_4246) );
CLKBUF_X2 inst_10526 ( .A(net_10487), .Z(net_10488) );
DFF_X1 inst_6381 ( .QN(net_6281), .D(net_5803), .CK(net_13638) );
NAND2_X2 inst_3711 ( .A1(net_6758), .ZN(net_1636), .A2(net_1635) );
DFFR_X2 inst_7103 ( .D(net_1943), .QN(net_128), .CK(net_12320), .RN(x1822) );
CLKBUF_X2 inst_13419 ( .A(net_13380), .Z(net_13381) );
NOR2_X4 inst_2241 ( .ZN(net_5645), .A1(net_5491), .A2(net_4459) );
CLKBUF_X2 inst_8165 ( .A(net_7969), .Z(net_8127) );
AOI222_X2 inst_7568 ( .ZN(net_5351), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_344), .C2(net_342), .A1(net_330) );
NOR4_X2 inst_2182 ( .ZN(net_2424), .A3(net_1674), .A4(net_1673), .A1(net_1234), .A2(net_1230) );
CLKBUF_X2 inst_8334 ( .A(net_8295), .Z(net_8296) );
SDFF_X2 inst_650 ( .Q(net_6706), .D(net_6706), .SE(net_3871), .SI(net_3812), .CK(net_8298) );
SDFF_X2 inst_289 ( .D(net_6396), .SE(net_6050), .SI(net_303), .Q(net_303), .CK(net_14219) );
NAND3_X2 inst_2667 ( .ZN(net_3963), .A2(net_3876), .A3(net_3738), .A1(net_2235) );
CLKBUF_X2 inst_8674 ( .A(net_7989), .Z(net_8636) );
NAND2_X2 inst_4194 ( .ZN(net_899), .A1(net_888), .A2(net_395) );
SDFF_X2 inst_987 ( .Q(net_6473), .D(net_6473), .SE(net_3904), .SI(net_3808), .CK(net_8778) );
CLKBUF_X2 inst_12467 ( .A(net_11522), .Z(net_12429) );
CLKBUF_X2 inst_8701 ( .A(net_8662), .Z(net_8663) );
CLKBUF_X2 inst_9376 ( .A(net_9337), .Z(net_9338) );
CLKBUF_X2 inst_8643 ( .A(net_8604), .Z(net_8605) );
SDFF_X2 inst_679 ( .Q(net_6743), .D(net_6743), .SE(net_3815), .SI(net_3808), .CK(net_11341) );
INV_X4 inst_5627 ( .A(net_7432), .ZN(net_2154) );
NAND2_X2 inst_3006 ( .A1(net_6885), .A2(net_5006), .ZN(net_5003) );
CLKBUF_X2 inst_12532 ( .A(net_10309), .Z(net_12494) );
CLKBUF_X2 inst_9703 ( .A(net_8560), .Z(net_9665) );
AOI21_X2 inst_7689 ( .B1(net_6726), .ZN(net_4508), .B2(net_2581), .A(net_2377) );
NAND2_X2 inst_3364 ( .ZN(net_3518), .A1(net_3517), .A2(net_3223) );
SDFFR_X2 inst_1351 ( .D(net_3800), .SE(net_3256), .SI(net_153), .Q(net_153), .CK(net_10398), .RN(x1822) );
CLKBUF_X2 inst_10443 ( .A(net_10404), .Z(net_10405) );
XNOR2_X2 inst_44 ( .B(net_6690), .ZN(net_2445), .A(net_1239) );
NAND2_X1 inst_4433 ( .A2(net_2131), .ZN(net_1414), .A1(net_1413) );
SDFF_X2 inst_371 ( .SI(net_7643), .Q(net_7643), .D(net_4787), .SE(net_3867), .CK(net_8311) );
CLKBUF_X2 inst_13994 ( .A(net_13955), .Z(net_13956) );
CLKBUF_X2 inst_12805 ( .A(net_9830), .Z(net_12767) );
SDFF_X2 inst_435 ( .Q(net_7387), .D(net_7387), .SE(net_3994), .SI(net_352), .CK(net_9641) );
DFF_X1 inst_6498 ( .QN(net_7410), .D(net_5538), .CK(net_9300) );
INV_X4 inst_4962 ( .ZN(net_3277), .A(net_718) );
CLKBUF_X2 inst_11563 ( .A(net_8309), .Z(net_11525) );
CLKBUF_X2 inst_10768 ( .A(net_10729), .Z(net_10730) );
CLKBUF_X2 inst_10791 ( .A(net_10752), .Z(net_10753) );
CLKBUF_X2 inst_10305 ( .A(net_10266), .Z(net_10267) );
INV_X4 inst_4619 ( .ZN(net_4203), .A(net_4067) );
CLKBUF_X2 inst_13474 ( .A(net_13435), .Z(net_13436) );
NAND2_X2 inst_3787 ( .A1(net_7044), .A2(net_1975), .ZN(net_1558) );
AOI222_X2 inst_7470 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2171), .A1(net_2170), .B1(net_2169), .C1(net_2168) );
INV_X4 inst_4982 ( .A(net_772), .ZN(net_724) );
SDFF_X2 inst_628 ( .SI(net_6639), .Q(net_6639), .SE(net_3850), .D(net_3785), .CK(net_10660) );
NAND2_X2 inst_3684 ( .A2(net_1798), .ZN(net_1765), .A1(net_1764) );
CLKBUF_X2 inst_13633 ( .A(net_13594), .Z(net_13595) );
OAI21_X2 inst_1923 ( .ZN(net_5122), .A(net_4756), .B2(net_3941), .B1(net_1141) );
NAND3_X2 inst_2748 ( .ZN(net_2353), .A3(net_1598), .A1(net_1522), .A2(net_1037) );
NAND2_X2 inst_3013 ( .A1(net_6856), .A2(net_5004), .ZN(net_4996) );
CLKBUF_X2 inst_9201 ( .A(net_8968), .Z(net_9163) );
INV_X4 inst_4744 ( .A(net_2754), .ZN(net_2748) );
NAND2_X2 inst_3642 ( .ZN(net_2230), .A2(net_1919), .A1(net_1691) );
CLKBUF_X2 inst_11873 ( .A(net_11834), .Z(net_11835) );
INV_X4 inst_5087 ( .A(net_7809), .ZN(net_3786) );
CLKBUF_X2 inst_9130 ( .A(net_9091), .Z(net_9092) );
AOI222_X2 inst_7563 ( .A1(net_7244), .ZN(net_5363), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_338), .C2(net_336) );
NAND2_X2 inst_3092 ( .A1(net_6486), .A2(net_4927), .ZN(net_4911) );
CLKBUF_X2 inst_14162 ( .A(net_12842), .Z(net_14124) );
DFF_X1 inst_6587 ( .QN(net_7557), .D(net_5063), .CK(net_13168) );
CLKBUF_X2 inst_11127 ( .A(net_10418), .Z(net_11089) );
CLKBUF_X2 inst_13931 ( .A(net_12526), .Z(net_13893) );
NAND3_X2 inst_2734 ( .ZN(net_2367), .A3(net_1555), .A1(net_1339), .A2(net_1025) );
INV_X4 inst_4920 ( .A(net_3894), .ZN(net_3273) );
NAND2_X2 inst_3395 ( .ZN(net_4300), .A2(net_3441), .A1(net_2855) );
SDFF_X2 inst_1130 ( .SI(net_6681), .Q(net_6681), .D(net_3790), .SE(net_3471), .CK(net_11997) );
CLKBUF_X2 inst_11608 ( .A(net_11569), .Z(net_11570) );
CLKBUF_X2 inst_9300 ( .A(net_9261), .Z(net_9262) );
DFF_X1 inst_6518 ( .QN(net_7449), .D(net_5435), .CK(net_9677) );
SDFF_X2 inst_855 ( .SI(net_7040), .Q(net_7040), .D(net_3812), .SE(net_3777), .CK(net_8220) );
OAI21_X2 inst_2039 ( .B1(net_4621), .B2(net_4476), .ZN(net_4464), .A(net_3582) );
CLKBUF_X2 inst_12706 ( .A(net_12667), .Z(net_12668) );
DFF_X2 inst_6304 ( .QN(net_7690), .D(net_837), .CK(net_9487) );
NAND2_X2 inst_3233 ( .ZN(net_4303), .A2(net_4164), .A1(net_663) );
AND2_X2 inst_7851 ( .A1(net_7770), .ZN(net_4002), .A2(net_4001) );
CLKBUF_X2 inst_8996 ( .A(net_8474), .Z(net_8958) );
CLKBUF_X2 inst_11823 ( .A(net_10087), .Z(net_11785) );
INV_X2 inst_5866 ( .A(net_826), .ZN(net_536) );
INV_X4 inst_5466 ( .A(net_6130), .ZN(net_3633) );
AOI222_X2 inst_7588 ( .A1(net_7385), .ZN(net_5448), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_348), .C2(net_346) );
INV_X4 inst_5425 ( .A(net_5996), .ZN(net_629) );
CLKBUF_X2 inst_10160 ( .A(net_10121), .Z(net_10122) );
CLKBUF_X2 inst_9304 ( .A(net_9265), .Z(net_9266) );
NAND2_X1 inst_4295 ( .ZN(net_4571), .A2(net_3866), .A1(net_2128) );
SDFF_X2 inst_518 ( .Q(net_6751), .D(net_6751), .SI(net_3898), .SE(net_3815), .CK(net_8378) );
SDFFR_X2 inst_1363 ( .SI(net_7738), .Q(net_7738), .D(net_4596), .SE(net_2608), .CK(net_10331), .RN(x1822) );
INV_X4 inst_4851 ( .ZN(net_1056), .A(net_1055) );
INV_X2 inst_5894 ( .A(net_7363), .ZN(net_2050) );
CLKBUF_X2 inst_8242 ( .A(net_8032), .Z(net_8204) );
NAND2_X2 inst_3863 ( .A1(net_6983), .A2(net_1833), .ZN(net_1469) );
NOR2_X2 inst_2345 ( .A2(net_6014), .A1(net_5778), .ZN(net_5706) );
CLKBUF_X2 inst_8059 ( .A(net_8020), .Z(net_8021) );
CLKBUF_X2 inst_12157 ( .A(net_12118), .Z(net_12119) );
DFF_X1 inst_6538 ( .QN(net_7470), .D(net_5578), .CK(net_9267) );
NAND2_X2 inst_3602 ( .ZN(net_2398), .A2(net_1843), .A1(net_1364) );
CLKBUF_X2 inst_9614 ( .A(net_9575), .Z(net_9576) );
CLKBUF_X2 inst_12388 ( .A(net_8010), .Z(net_12350) );
CLKBUF_X2 inst_14291 ( .A(net_11570), .Z(net_14253) );
AOI222_X2 inst_7582 ( .A1(net_7536), .ZN(net_5240), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_368), .C2(net_366) );
INV_X4 inst_5260 ( .ZN(net_432), .A(net_431) );
CLKBUF_X2 inst_12637 ( .A(net_9255), .Z(net_12599) );
CLKBUF_X2 inst_11815 ( .A(net_11776), .Z(net_11777) );
CLKBUF_X2 inst_11372 ( .A(net_8850), .Z(net_11334) );
CLKBUF_X2 inst_12336 ( .A(net_12297), .Z(net_12298) );
INV_X4 inst_5190 ( .A(net_844), .ZN(net_513) );
SDFFR_X2 inst_1354 ( .D(net_3804), .SE(net_3256), .SI(net_152), .Q(net_152), .CK(net_8544), .RN(x1822) );
CLKBUF_X2 inst_11806 ( .A(net_10719), .Z(net_11768) );
SDFF_X2 inst_970 ( .Q(net_6450), .D(net_6450), .SE(net_3820), .SI(net_3790), .CK(net_8415) );
CLKBUF_X2 inst_11992 ( .A(net_11953), .Z(net_11954) );
DFF_X1 inst_6731 ( .QN(net_7350), .D(net_5324), .CK(net_10123) );
SDFF_X2 inst_1278 ( .D(net_3798), .SE(net_3256), .SI(net_135), .Q(net_135), .CK(net_8481) );
NAND2_X2 inst_3763 ( .A1(net_6911), .A2(net_1639), .ZN(net_1582) );
CLKBUF_X2 inst_10136 ( .A(net_10097), .Z(net_10098) );
SDFF_X2 inst_749 ( .Q(net_6861), .D(net_6861), .SE(net_3901), .SI(net_3792), .CK(net_8937) );
CLKBUF_X2 inst_11975 ( .A(net_11936), .Z(net_11937) );
DFF_X1 inst_6688 ( .QN(net_7277), .D(net_5123), .CK(net_9960) );
SDFF_X2 inst_1030 ( .Q(net_7536), .D(net_7536), .SE(net_3896), .SI(net_370), .CK(net_9393) );
OAI21_X2 inst_2127 ( .ZN(net_3005), .B1(net_2997), .A(net_2873), .B2(net_2623) );
CLKBUF_X2 inst_13689 ( .A(net_11986), .Z(net_13651) );
CLKBUF_X2 inst_13626 ( .A(net_13587), .Z(net_13588) );
CLKBUF_X2 inst_10611 ( .A(net_10572), .Z(net_10573) );
NAND3_X2 inst_2649 ( .ZN(net_4153), .A1(net_4152), .A3(net_3992), .A2(net_1730) );
CLKBUF_X2 inst_11441 ( .A(net_11402), .Z(net_11403) );
OR2_X4 inst_1373 ( .ZN(net_3448), .A2(net_3249), .A1(net_2601) );
NOR2_X4 inst_2268 ( .ZN(net_5618), .A1(net_5463), .A2(net_4412) );
NOR2_X2 inst_2458 ( .ZN(net_2994), .A1(net_2805), .A2(net_227) );
NAND2_X2 inst_3828 ( .A1(net_6838), .A2(net_1521), .ZN(net_1515) );
AOI22_X2 inst_7285 ( .B1(net_7222), .A1(net_7190), .A2(net_5244), .B2(net_5243), .ZN(net_5224) );
CLKBUF_X2 inst_14303 ( .A(net_14264), .Z(net_14265) );
CLKBUF_X2 inst_8474 ( .A(net_8246), .Z(net_8436) );
INV_X2 inst_5841 ( .ZN(net_765), .A(net_624) );
CLKBUF_X2 inst_9923 ( .A(net_9884), .Z(net_9885) );
DFF_X1 inst_6898 ( .D(net_2510), .QN(net_178), .CK(net_9948) );
NAND2_X2 inst_3155 ( .ZN(net_4808), .A2(net_4153), .A1(net_2097) );
INV_X4 inst_5481 ( .A(net_6002), .ZN(net_442) );
NAND2_X2 inst_3134 ( .ZN(net_4829), .A2(net_4153), .A1(net_2170) );
SDFF_X2 inst_1006 ( .SI(net_6488), .Q(net_6488), .SE(net_3889), .D(net_3792), .CK(net_8772) );
OAI21_X2 inst_1985 ( .B1(net_4849), .ZN(net_4844), .A(net_4581), .B2(net_3867) );
AOI22_X2 inst_7311 ( .B1(net_6684), .A1(net_6652), .A2(net_5139), .B2(net_5138), .ZN(net_5132) );
CLKBUF_X2 inst_13519 ( .A(net_13480), .Z(net_13481) );
CLKBUF_X2 inst_11787 ( .A(net_8875), .Z(net_11749) );
DFF_X1 inst_6710 ( .QN(net_7326), .D(net_5360), .CK(net_10153) );
NAND2_X2 inst_4043 ( .A1(net_6796), .A2(net_1651), .ZN(net_1009) );
CLKBUF_X2 inst_10473 ( .A(net_10434), .Z(net_10435) );
CLKBUF_X2 inst_9817 ( .A(net_9778), .Z(net_9779) );
INV_X4 inst_5134 ( .ZN(net_3918), .A(net_803) );
CLKBUF_X2 inst_8407 ( .A(net_8017), .Z(net_8369) );
CLKBUF_X2 inst_11999 ( .A(net_11960), .Z(net_11961) );
INV_X2 inst_5755 ( .A(net_3404), .ZN(net_3330) );
CLKBUF_X2 inst_11933 ( .A(net_11894), .Z(net_11895) );
CLKBUF_X2 inst_8691 ( .A(net_8652), .Z(net_8653) );
INV_X4 inst_4753 ( .ZN(net_2622), .A(net_392) );
CLKBUF_X2 inst_10960 ( .A(net_10921), .Z(net_10922) );
CLKBUF_X2 inst_8122 ( .A(net_8008), .Z(net_8084) );
CLKBUF_X2 inst_11885 ( .A(net_7827), .Z(net_11847) );
CLKBUF_X2 inst_10082 ( .A(net_8575), .Z(net_10044) );
CLKBUF_X2 inst_11957 ( .A(net_11918), .Z(net_11919) );
INV_X4 inst_4947 ( .ZN(net_738), .A(net_737) );
CLKBUF_X2 inst_13435 ( .A(net_12706), .Z(net_13397) );
CLKBUF_X2 inst_8915 ( .A(net_8876), .Z(net_8877) );
CLKBUF_X2 inst_11671 ( .A(net_11632), .Z(net_11633) );
CLKBUF_X2 inst_12349 ( .A(net_12310), .Z(net_12311) );
INV_X2 inst_5783 ( .ZN(net_2446), .A(net_2445) );
CLKBUF_X2 inst_12490 ( .A(net_8892), .Z(net_12452) );
CLKBUF_X2 inst_12755 ( .A(net_12716), .Z(net_12717) );
DFF_X1 inst_6457 ( .QN(net_6110), .D(net_5602), .CK(net_11175) );
INV_X4 inst_4588 ( .ZN(net_4314), .A(net_4226) );
CLKBUF_X2 inst_13746 ( .A(net_13707), .Z(net_13708) );
CLKBUF_X2 inst_9099 ( .A(net_9060), .Z(net_9061) );
CLKBUF_X2 inst_9898 ( .A(net_9859), .Z(net_9860) );
NAND2_X2 inst_4184 ( .ZN(net_1046), .A2(net_481), .A1(net_427) );
NAND2_X2 inst_4049 ( .A1(net_6934), .A2(net_1654), .ZN(net_1003) );
INV_X4 inst_5067 ( .A(net_3230), .ZN(net_1216) );
NAND3_X2 inst_2702 ( .A1(net_5932), .ZN(net_2645), .A3(net_2644), .A2(net_689) );
CLKBUF_X2 inst_12820 ( .A(net_12781), .Z(net_12782) );
DFF_X1 inst_6531 ( .QN(net_7478), .D(net_5420), .CK(net_9271) );
NAND2_X2 inst_2910 ( .ZN(net_5785), .A2(net_5771), .A1(net_414) );
CLKBUF_X2 inst_11517 ( .A(net_11478), .Z(net_11479) );
INV_X4 inst_4670 ( .ZN(net_3541), .A(net_3540) );
INV_X4 inst_5701 ( .A(net_5939), .ZN(net_5938) );
NAND2_X2 inst_3238 ( .ZN(net_4275), .A1(net_4274), .A2(net_1642) );
SDFF_X2 inst_145 ( .Q(net_6233), .SI(net_6232), .SE(net_392), .D(net_139), .CK(net_14114) );
CLKBUF_X2 inst_13703 ( .A(net_11084), .Z(net_13665) );
NAND2_X4 inst_2854 ( .ZN(net_5469), .A1(net_4907), .A2(net_4906) );
NAND2_X2 inst_3030 ( .A1(net_6987), .ZN(net_4978), .A2(net_4977) );
AOI21_X2 inst_7717 ( .B1(net_6864), .ZN(net_5897), .B2(net_2579), .A(net_2343) );
INV_X4 inst_4594 ( .ZN(net_5090), .A(net_4295) );
NOR2_X4 inst_2230 ( .ZN(net_5668), .A1(net_5529), .A2(net_4496) );
CLKBUF_X2 inst_9689 ( .A(net_8824), .Z(net_9651) );
INV_X4 inst_5355 ( .A(net_6037), .ZN(net_2597) );
INV_X4 inst_5630 ( .A(net_6143), .ZN(net_3645) );
CLKBUF_X2 inst_13028 ( .A(net_12989), .Z(net_12990) );
DFF_X2 inst_6214 ( .D(net_4002), .QN(net_154), .CK(net_12383) );
CLKBUF_X2 inst_10199 ( .A(net_10160), .Z(net_10161) );
CLKBUF_X2 inst_10511 ( .A(net_10472), .Z(net_10473) );
CLKBUF_X2 inst_12240 ( .A(net_12201), .Z(net_12202) );
INV_X4 inst_5345 ( .A(net_7784), .ZN(net_888) );
OAI22_X2 inst_1437 ( .B1(net_5852), .ZN(net_5686), .A2(net_5498), .B2(net_5497), .A1(net_5258) );
CLKBUF_X2 inst_13820 ( .A(net_11686), .Z(net_13782) );
CLKBUF_X2 inst_10481 ( .A(net_10442), .Z(net_10443) );
CLKBUF_X2 inst_9292 ( .A(net_9253), .Z(net_9254) );
CLKBUF_X2 inst_9119 ( .A(net_8200), .Z(net_9081) );
CLKBUF_X2 inst_14174 ( .A(net_14135), .Z(net_14136) );
CLKBUF_X2 inst_10557 ( .A(net_8268), .Z(net_10519) );
CLKBUF_X2 inst_13661 ( .A(net_13622), .Z(net_13623) );
INV_X8 inst_4477 ( .ZN(net_4979), .A(net_4266) );
NOR2_X2 inst_2533 ( .ZN(net_1646), .A2(net_703), .A1(net_488) );
NOR2_X2 inst_2391 ( .ZN(net_3998), .A2(net_3996), .A1(net_1203) );
AOI222_X2 inst_7606 ( .A1(net_7237), .ZN(net_5347), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_331), .C2(net_329) );
NOR2_X4 inst_2239 ( .ZN(net_5659), .A1(net_5512), .A2(net_4481) );
XNOR2_X2 inst_27 ( .ZN(net_2568), .B(net_2567), .A(net_2440) );
CLKBUF_X2 inst_10027 ( .A(net_9988), .Z(net_9989) );
CLKBUF_X2 inst_10741 ( .A(net_10702), .Z(net_10703) );
CLKBUF_X2 inst_8790 ( .A(net_8386), .Z(net_8752) );
DFF_X2 inst_6335 ( .QN(net_7812), .CK(net_8432), .D(x1443) );
OAI222_X2 inst_1639 ( .C2(net_4107), .ZN(net_4009), .A2(net_4008), .B2(net_4007), .A1(net_2444), .B1(net_1650), .C1(net_430) );
NAND2_X1 inst_4446 ( .ZN(net_1258), .A1(net_1257), .A2(net_1256) );
CLKBUF_X2 inst_13645 ( .A(net_11273), .Z(net_13607) );
CLKBUF_X2 inst_11468 ( .A(net_11429), .Z(net_11430) );
CLKBUF_X2 inst_10717 ( .A(net_10678), .Z(net_10679) );
CLKBUF_X2 inst_11761 ( .A(net_11722), .Z(net_11723) );
CLKBUF_X2 inst_10063 ( .A(net_9348), .Z(net_10025) );
INV_X4 inst_5155 ( .A(net_565), .ZN(net_560) );
CLKBUF_X2 inst_10365 ( .A(net_8084), .Z(net_10327) );
CLKBUF_X2 inst_11071 ( .A(net_10918), .Z(net_11033) );
CLKBUF_X2 inst_9756 ( .A(net_9717), .Z(net_9718) );
AOI22_X2 inst_7403 ( .B1(net_5939), .A2(net_2838), .ZN(net_2835), .A1(net_2834), .B2(net_207) );
DFF_X1 inst_6420 ( .QN(net_6175), .D(net_5750), .CK(net_8748) );
INV_X4 inst_5230 ( .ZN(net_1666), .A(net_460) );
CLKBUF_X2 inst_9045 ( .A(net_9006), .Z(net_9007) );
SDFF_X2 inst_639 ( .SI(net_6652), .Q(net_6652), .SE(net_3851), .D(net_3821), .CK(net_12011) );
SDFF_X2 inst_155 ( .QN(net_6259), .SI(net_6258), .D(net_3538), .SE(net_392), .CK(net_14001) );
INV_X4 inst_4858 ( .ZN(net_1670), .A(net_1042) );
CLKBUF_X2 inst_10170 ( .A(net_10131), .Z(net_10132) );
NAND2_X2 inst_3939 ( .A1(net_7116), .A2(net_1675), .ZN(net_1354) );
INV_X2 inst_6043 ( .A(net_7379), .ZN(net_399) );
INV_X4 inst_5309 ( .A(net_7532), .ZN(net_435) );
XNOR2_X2 inst_55 ( .ZN(net_2246), .A(net_2245), .B(net_2244) );
OAI211_X2 inst_2167 ( .B(net_2724), .ZN(net_2721), .A(net_1922), .C2(net_1921), .C1(net_1057) );
NOR2_X4 inst_2280 ( .ZN(net_3841), .A1(net_3400), .A2(net_3236) );
DFFR_X2 inst_7008 ( .D(net_3281), .QN(net_272), .CK(net_12343), .RN(x1822) );
CLKBUF_X2 inst_12193 ( .A(net_11597), .Z(net_12155) );
AOI22_X2 inst_7412 ( .B1(net_5939), .A2(net_2838), .ZN(net_2823), .A1(net_742), .B2(net_197) );
DFF_X2 inst_6328 ( .QN(net_7821), .CK(net_8241), .D(x1366) );
CLKBUF_X2 inst_9872 ( .A(net_9833), .Z(net_9834) );
DFFR_X2 inst_7097 ( .D(net_1956), .QN(net_116), .CK(net_9594), .RN(x1822) );
CLKBUF_X2 inst_12561 ( .A(net_9871), .Z(net_12523) );
NAND2_X1 inst_4248 ( .ZN(net_4678), .A2(net_3988), .A1(net_2184) );
OAI221_X2 inst_1651 ( .ZN(net_5044), .C2(net_5043), .B2(net_5040), .A(net_4523), .B1(net_2429), .C1(net_1088) );
CLKBUF_X2 inst_12176 ( .A(net_12137), .Z(net_12138) );
CLKBUF_X2 inst_9758 ( .A(net_8431), .Z(net_9720) );
CLKBUF_X2 inst_8281 ( .A(net_8242), .Z(net_8243) );
NAND2_X2 inst_4127 ( .A2(net_1225), .ZN(net_1190), .A1(net_364) );
CLKBUF_X2 inst_11634 ( .A(net_11595), .Z(net_11596) );
CLKBUF_X2 inst_11159 ( .A(net_11120), .Z(net_11121) );
DFF_X1 inst_6451 ( .QN(net_6102), .D(net_5719), .CK(net_9215) );
SDFF_X2 inst_1137 ( .D(net_7799), .SI(net_6661), .Q(net_6661), .SE(net_3465), .CK(net_12889) );
SDFF_X2 inst_323 ( .SI(net_7488), .Q(net_7488), .D(net_5104), .SE(net_3989), .CK(net_12070) );
OR2_X4 inst_1389 ( .A2(net_7782), .A1(net_7781), .ZN(net_768) );
CLKBUF_X2 inst_9032 ( .A(net_8207), .Z(net_8994) );
CLKBUF_X2 inst_14043 ( .A(net_14004), .Z(net_14005) );
NAND2_X2 inst_3065 ( .A1(net_7127), .A2(net_4950), .ZN(net_4940) );
SDFF_X2 inst_715 ( .SI(net_6760), .Q(net_6760), .SE(net_3816), .D(net_3802), .CK(net_8959) );
OAI22_X2 inst_1494 ( .B1(net_4666), .B2(net_4521), .A2(net_4134), .A1(net_4132), .ZN(net_4113) );
INV_X4 inst_5206 ( .ZN(net_2999), .A(net_492) );
AOI22_X2 inst_7333 ( .A2(net_3420), .B2(net_3419), .ZN(net_3413), .B1(net_2571), .A1(net_1244) );
DFF_X1 inst_6354 ( .QN(net_6204), .D(net_5830), .CK(net_13701) );
CLKBUF_X2 inst_8941 ( .A(net_8902), .Z(net_8903) );
INV_X4 inst_5213 ( .A(net_3093), .ZN(net_482) );
CLKBUF_X2 inst_14113 ( .A(net_14074), .Z(net_14075) );
NAND2_X2 inst_3525 ( .ZN(net_2542), .A2(net_2126), .A1(net_1472) );
CLKBUF_X2 inst_12734 ( .A(net_11635), .Z(net_12696) );
CLKBUF_X2 inst_10479 ( .A(net_10440), .Z(net_10441) );
NAND2_X2 inst_3449 ( .A2(net_5925), .ZN(net_2923), .A1(net_1828) );
OAI221_X2 inst_1682 ( .C1(net_5940), .ZN(net_3253), .B1(net_3252), .A(net_3038), .C2(net_221), .B2(net_184) );
INV_X4 inst_5077 ( .A(net_7813), .ZN(net_3783) );
SDFFR_X2 inst_1340 ( .Q(net_7710), .D(net_7710), .SI(net_3807), .SE(net_3405), .CK(net_10716), .RN(x1822) );
OAI22_X2 inst_1481 ( .A1(net_4855), .B1(net_4228), .B2(net_4222), .A2(net_4173), .ZN(net_4172) );
CLKBUF_X2 inst_14275 ( .A(net_14236), .Z(net_14237) );
CLKBUF_X2 inst_13778 ( .A(net_11489), .Z(net_13740) );
CLKBUF_X2 inst_10630 ( .A(net_10291), .Z(net_10592) );
CLKBUF_X2 inst_13194 ( .A(net_13155), .Z(net_13156) );
CLKBUF_X2 inst_10191 ( .A(net_9418), .Z(net_10153) );
AND4_X2 inst_7794 ( .ZN(net_837), .A3(net_836), .A2(x1155), .A1(x1126), .A4(x1101) );
CLKBUF_X2 inst_13349 ( .A(net_13310), .Z(net_13311) );
XNOR2_X2 inst_31 ( .ZN(net_2481), .A(net_2480), .B(net_935) );
NAND2_X2 inst_3505 ( .ZN(net_2562), .A2(net_2199), .A1(net_1489) );
CLKBUF_X2 inst_9355 ( .A(net_8512), .Z(net_9317) );
CLKBUF_X2 inst_8788 ( .A(net_8749), .Z(net_8750) );
CLKBUF_X2 inst_10128 ( .A(net_9435), .Z(net_10090) );
AOI21_X2 inst_7707 ( .B1(net_6867), .ZN(net_4500), .B2(net_2579), .A(net_2357) );
CLKBUF_X2 inst_10204 ( .A(net_10165), .Z(net_10166) );
NAND2_X2 inst_3217 ( .ZN(net_4709), .A2(net_3986), .A1(net_1979) );
CLKBUF_X2 inst_9556 ( .A(net_9517), .Z(net_9518) );
CLKBUF_X2 inst_10937 ( .A(net_8651), .Z(net_10899) );
DFF_X1 inst_6440 ( .QN(net_6083), .D(net_5730), .CK(net_11677) );
CLKBUF_X2 inst_12730 ( .A(net_12691), .Z(net_12692) );
CLKBUF_X2 inst_9787 ( .A(net_8045), .Z(net_9749) );
NAND2_X1 inst_4376 ( .ZN(net_4351), .A2(net_3859), .A1(net_2065) );
NAND2_X2 inst_3537 ( .ZN(net_2530), .A2(net_2163), .A1(net_1786) );
CLKBUF_X2 inst_12606 ( .A(net_12567), .Z(net_12568) );
INV_X8 inst_4556 ( .ZN(net_2133), .A(net_779) );
CLKBUF_X2 inst_14449 ( .A(net_14410), .Z(net_14411) );
CLKBUF_X2 inst_11778 ( .A(net_11739), .Z(net_11740) );
INV_X2 inst_6023 ( .ZN(net_401), .A(x906) );
OAI21_X2 inst_1833 ( .ZN(net_5344), .B1(net_5343), .A(net_4357), .B2(net_3856) );
CLKBUF_X2 inst_8160 ( .A(net_8121), .Z(net_8122) );
INV_X4 inst_5301 ( .A(net_6822), .ZN(net_574) );
OAI21_X2 inst_2122 ( .B1(net_3299), .B2(net_3087), .ZN(net_3086), .A(net_2909) );
NAND2_X2 inst_3044 ( .A1(net_6994), .A2(net_4977), .ZN(net_4963) );
INV_X4 inst_5443 ( .A(net_6118), .ZN(net_3473) );
NAND2_X2 inst_3520 ( .ZN(net_2547), .A2(net_2122), .A1(net_1508) );
CLKBUF_X2 inst_11601 ( .A(net_11562), .Z(net_11563) );
CLKBUF_X2 inst_9809 ( .A(net_9770), .Z(net_9771) );
CLKBUF_X2 inst_13041 ( .A(net_13002), .Z(net_13003) );
CLKBUF_X2 inst_11914 ( .A(net_11875), .Z(net_11876) );
NAND2_X2 inst_3573 ( .ZN(net_2494), .A2(net_2056), .A1(net_1794) );
CLKBUF_X2 inst_13453 ( .A(net_12943), .Z(net_13415) );
CLKBUF_X2 inst_12324 ( .A(net_12285), .Z(net_12286) );
CLKBUF_X2 inst_11306 ( .A(net_10492), .Z(net_11268) );
SDFF_X2 inst_623 ( .SI(net_6623), .Q(net_6623), .SE(net_3851), .D(net_3797), .CK(net_9694) );
SDFF_X2 inst_1072 ( .SI(net_6536), .Q(net_6536), .D(net_3786), .SE(net_3755), .CK(net_8758) );
CLKBUF_X2 inst_8557 ( .A(net_8518), .Z(net_8519) );
OAI22_X2 inst_1621 ( .B1(net_5938), .A1(net_2786), .ZN(net_2783), .B2(net_213), .A2(net_176) );
OAI21_X2 inst_1993 ( .ZN(net_4599), .B2(net_4598), .B1(net_4228), .A(net_3594) );
CLKBUF_X2 inst_10373 ( .A(net_10334), .Z(net_10335) );
CLKBUF_X2 inst_14193 ( .A(net_14154), .Z(net_14155) );
CLKBUF_X2 inst_9791 ( .A(net_9752), .Z(net_9753) );
NAND2_X2 inst_3226 ( .A2(net_7780), .ZN(net_5253), .A1(net_4297) );
DFF_X1 inst_6671 ( .QN(net_7266), .D(net_5159), .CK(net_9890) );
CLKBUF_X2 inst_10674 ( .A(net_10635), .Z(net_10636) );
CLKBUF_X2 inst_8435 ( .A(net_8396), .Z(net_8397) );
CLKBUF_X2 inst_9609 ( .A(net_9570), .Z(net_9571) );
CLKBUF_X2 inst_13224 ( .A(net_13185), .Z(net_13186) );
DFF_X1 inst_6470 ( .QN(net_6171), .D(net_5589), .CK(net_7957) );
NAND2_X2 inst_3617 ( .ZN(net_2265), .A2(net_1940), .A1(net_1308) );
CLKBUF_X2 inst_10893 ( .A(net_10854), .Z(net_10855) );
OR2_X4 inst_1377 ( .ZN(net_3444), .A2(net_3251), .A1(net_2609) );
NAND2_X2 inst_3125 ( .ZN(net_4838), .A2(net_4153), .A1(net_2174) );
CLKBUF_X2 inst_10571 ( .A(net_10532), .Z(net_10533) );
NOR3_X2 inst_2201 ( .ZN(net_3173), .A1(net_2979), .A3(net_1743), .A2(net_1103) );
CLKBUF_X2 inst_14130 ( .A(net_9686), .Z(net_14092) );
CLKBUF_X2 inst_10581 ( .A(net_10542), .Z(net_10543) );
CLKBUF_X2 inst_10750 ( .A(net_10711), .Z(net_10712) );
CLKBUF_X2 inst_10562 ( .A(net_10523), .Z(net_10524) );
SDFF_X2 inst_760 ( .Q(net_6883), .D(net_6883), .SE(net_3901), .SI(net_3804), .CK(net_10894) );
CLKBUF_X2 inst_14144 ( .A(net_9598), .Z(net_14106) );
CLKBUF_X2 inst_12842 ( .A(net_12803), .Z(net_12804) );
CLKBUF_X2 inst_10814 ( .A(net_10775), .Z(net_10776) );
CLKBUF_X2 inst_8867 ( .A(net_8828), .Z(net_8829) );
INV_X4 inst_5671 ( .A(net_7789), .ZN(net_1928) );
OAI21_X2 inst_1696 ( .ZN(net_5598), .A(net_5286), .B2(net_4500), .B1(net_4105) );
CLKBUF_X2 inst_9347 ( .A(net_9308), .Z(net_9309) );
INV_X4 inst_4911 ( .A(net_3883), .ZN(net_3111) );
INV_X8 inst_4525 ( .ZN(net_3751), .A(net_3114) );
NAND2_X2 inst_4115 ( .A2(net_1225), .ZN(net_1178), .A1(net_359) );
CLKBUF_X2 inst_13264 ( .A(net_13225), .Z(net_13226) );
CLKBUF_X2 inst_9831 ( .A(net_9357), .Z(net_9793) );
CLKBUF_X2 inst_8174 ( .A(net_8135), .Z(net_8136) );
NAND2_X2 inst_3727 ( .A1(net_7165), .A2(net_1637), .ZN(net_1618) );
CLKBUF_X2 inst_12237 ( .A(net_12198), .Z(net_12199) );
CLKBUF_X2 inst_10812 ( .A(net_9741), .Z(net_10774) );
CLKBUF_X2 inst_8417 ( .A(net_8113), .Z(net_8379) );
INV_X4 inst_5591 ( .A(net_7733), .ZN(net_2679) );
AOI22_X2 inst_7258 ( .B1(net_6949), .A1(net_6917), .A2(net_5298), .B2(net_5297), .ZN(net_5296) );
OAI21_X2 inst_1687 ( .B1(net_5778), .ZN(net_5777), .A(net_5711), .B2(net_5710) );
OAI21_X2 inst_1970 ( .ZN(net_4867), .B1(net_4866), .A(net_4352), .B2(net_3859) );
NAND2_X2 inst_3989 ( .A1(net_6425), .A2(net_1677), .ZN(net_1275) );
CLKBUF_X2 inst_12211 ( .A(net_8579), .Z(net_12173) );
CLKBUF_X2 inst_10000 ( .A(net_8527), .Z(net_9962) );
CLKBUF_X2 inst_12934 ( .A(net_8317), .Z(net_12896) );
DFF_X1 inst_6790 ( .D(net_3933), .CK(net_13215), .Q(x447) );
CLKBUF_X2 inst_14100 ( .A(net_14061), .Z(net_14062) );
CLKBUF_X2 inst_10256 ( .A(net_9268), .Z(net_10218) );
NAND2_X2 inst_3569 ( .ZN(net_2498), .A2(net_1998), .A1(net_1800) );
AOI22_X2 inst_7268 ( .B1(net_7082), .A1(net_7050), .ZN(net_5282), .A2(net_5280), .B2(net_5279) );
NAND2_X2 inst_3411 ( .ZN(net_4157), .A2(net_3321), .A1(net_2853) );
CLKBUF_X2 inst_10436 ( .A(net_10397), .Z(net_10398) );
AOI22_X2 inst_7417 ( .B1(net_5939), .A1(net_2777), .ZN(net_2776), .B2(net_220), .A2(net_183) );
CLKBUF_X2 inst_12576 ( .A(net_12537), .Z(net_12538) );
NOR2_X2 inst_2524 ( .ZN(net_3833), .A2(net_892), .A1(net_703) );
CLKBUF_X2 inst_9486 ( .A(net_9447), .Z(net_9448) );
OAI22_X2 inst_1446 ( .B2(net_5906), .B1(net_4660), .A2(net_4629), .ZN(net_4628), .A1(net_4089) );
SDFF_X2 inst_390 ( .SI(net_7310), .Q(net_7310), .D(net_4784), .SE(net_3859), .CK(net_12360) );
NOR2_X2 inst_2421 ( .A2(net_5890), .ZN(net_3229), .A1(net_617) );
INV_X4 inst_4842 ( .ZN(net_5876), .A(net_2997) );
CLKBUF_X2 inst_8181 ( .A(net_8142), .Z(net_8143) );
SDFF_X2 inst_1062 ( .Q(net_6868), .D(net_6868), .SE(net_3901), .SI(net_3890), .CK(net_11706) );
CLKBUF_X2 inst_13757 ( .A(net_9622), .Z(net_13719) );
CLKBUF_X2 inst_7996 ( .A(net_7949), .Z(net_7958) );
NAND3_X2 inst_2663 ( .ZN(net_3933), .A3(net_3394), .A2(net_2948), .A1(net_2833) );
NAND2_X2 inst_3289 ( .ZN(net_3668), .A1(net_3667), .A2(net_3229) );
AOI222_X2 inst_7477 ( .C1(net_7521), .B1(net_7489), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2151), .A1(net_2150) );
CLKBUF_X2 inst_12814 ( .A(net_12775), .Z(net_12776) );
CLKBUF_X2 inst_7930 ( .A(net_7891), .Z(net_7892) );
CLKBUF_X2 inst_14361 ( .A(net_13248), .Z(net_14323) );
CLKBUF_X2 inst_12650 ( .A(net_12611), .Z(net_12612) );
CLKBUF_X2 inst_12116 ( .A(net_11647), .Z(net_12078) );
CLKBUF_X2 inst_10508 ( .A(net_10469), .Z(net_10470) );
CLKBUF_X2 inst_12087 ( .A(net_12048), .Z(net_12049) );
CLKBUF_X2 inst_10277 ( .A(net_10238), .Z(net_10239) );
SDFF_X2 inst_401 ( .SI(net_7344), .Q(net_7344), .D(net_4777), .SE(net_3856), .CK(net_9403) );
CLKBUF_X2 inst_8086 ( .A(net_8047), .Z(net_8048) );
NAND2_X2 inst_3210 ( .ZN(net_4716), .A2(net_3986), .A1(net_1881) );
CLKBUF_X2 inst_12440 ( .A(net_12401), .Z(net_12402) );
DFFR_X2 inst_7063 ( .QN(net_6041), .D(net_3067), .CK(net_12642), .RN(x1822) );
CLKBUF_X2 inst_12539 ( .A(net_12500), .Z(net_12501) );
INV_X4 inst_5200 ( .ZN(net_663), .A(net_500) );
NAND3_X2 inst_2642 ( .ZN(net_5687), .A1(net_5664), .A2(net_5292), .A3(net_4238) );
INV_X16 inst_6145 ( .ZN(net_1637), .A(net_821) );
INV_X4 inst_4653 ( .ZN(net_4622), .A(net_4278) );
INV_X2 inst_6087 ( .A(net_7287), .ZN(net_2003) );
CLKBUF_X2 inst_12028 ( .A(net_9086), .Z(net_11990) );
INV_X8 inst_4465 ( .ZN(net_5243), .A(net_4286) );
CLKBUF_X2 inst_14394 ( .A(net_14355), .Z(net_14356) );
CLKBUF_X2 inst_13107 ( .A(net_13068), .Z(net_13069) );
CLKBUF_X2 inst_12281 ( .A(net_12242), .Z(net_12243) );
INV_X4 inst_4865 ( .A(net_2709), .ZN(net_1105) );
CLKBUF_X2 inst_13479 ( .A(net_13440), .Z(net_13441) );
CLKBUF_X2 inst_8548 ( .A(net_8509), .Z(net_8510) );
INV_X4 inst_5250 ( .ZN(net_441), .A(net_440) );
SDFF_X2 inst_123 ( .QN(net_6199), .SI(net_6198), .D(net_3374), .SE(net_392), .CK(net_14247) );
SDFF_X2 inst_930 ( .SI(net_7802), .Q(net_7140), .D(net_7140), .SE(net_3903), .CK(net_13343) );
AOI21_X2 inst_7634 ( .ZN(net_3956), .B2(net_3772), .B1(net_2894), .A(net_1046) );
CLKBUF_X2 inst_11908 ( .A(net_11869), .Z(net_11870) );
DFF_X1 inst_6801 ( .D(net_3935), .CK(net_9566), .Q(x589) );
OAI21_X2 inst_2160 ( .ZN(net_2806), .A(net_303), .B2(net_300), .B1(net_290) );
CLKBUF_X2 inst_8494 ( .A(net_8171), .Z(net_8456) );
INV_X4 inst_5181 ( .ZN(net_631), .A(net_522) );
CLKBUF_X2 inst_10981 ( .A(net_10897), .Z(net_10943) );
NOR2_X2 inst_2298 ( .A2(net_6189), .ZN(net_5845), .A1(net_5840) );
CLKBUF_X2 inst_10453 ( .A(net_9639), .Z(net_10415) );
CLKBUF_X2 inst_14355 ( .A(net_14316), .Z(net_14317) );
DFF_X1 inst_6622 ( .QN(net_7583), .D(net_5385), .CK(net_13437) );
CLKBUF_X2 inst_11660 ( .A(net_11621), .Z(net_11622) );
SDFF_X2 inst_167 ( .Q(net_6247), .SI(net_6246), .D(net_3647), .SE(net_392), .CK(net_13531) );
CLKBUF_X2 inst_13138 ( .A(net_13099), .Z(net_13100) );
CLKBUF_X2 inst_11354 ( .A(net_10119), .Z(net_11316) );
CLKBUF_X2 inst_13650 ( .A(net_13611), .Z(net_13612) );
INV_X4 inst_4913 ( .A(net_3798), .ZN(net_3280) );
NAND2_X2 inst_3874 ( .A1(net_7117), .A2(net_1675), .ZN(net_1447) );
CLKBUF_X2 inst_8524 ( .A(net_8485), .Z(net_8486) );
CLKBUF_X2 inst_9168 ( .A(net_9129), .Z(net_9130) );
SDFF_X2 inst_1251 ( .SI(net_6548), .Q(net_6548), .D(net_3793), .SE(net_3756), .CK(net_11624) );
CLKBUF_X2 inst_12245 ( .A(net_12206), .Z(net_12207) );
INV_X4 inst_4874 ( .ZN(net_1270), .A(net_906) );
NOR2_X2 inst_2475 ( .A2(net_5778), .ZN(net_2606), .A1(net_2605) );
AOI22_X2 inst_7360 ( .ZN(net_2995), .A2(net_2994), .B2(net_2993), .A1(net_1155), .B1(net_636) );
DFF_X1 inst_6824 ( .QN(net_5980), .D(net_3014), .CK(net_10519) );
CLKBUF_X2 inst_13033 ( .A(net_12994), .Z(net_12995) );
CLKBUF_X2 inst_9195 ( .A(net_9156), .Z(net_9157) );
CLKBUF_X2 inst_13131 ( .A(net_13092), .Z(net_13093) );
CLKBUF_X2 inst_12488 ( .A(net_11914), .Z(net_12450) );
SDFF_X2 inst_331 ( .SI(net_7517), .Q(net_7517), .D(net_5098), .SE(net_3988), .CK(net_9765) );
CLKBUF_X2 inst_10300 ( .A(net_10261), .Z(net_10262) );
CLKBUF_X2 inst_10270 ( .A(net_10231), .Z(net_10232) );
AOI22_X2 inst_7433 ( .A1(net_2970), .B1(net_2772), .ZN(net_2759), .A2(net_235), .B2(net_161) );
CLKBUF_X2 inst_10691 ( .A(net_10287), .Z(net_10653) );
CLKBUF_X2 inst_9937 ( .A(net_7856), .Z(net_9899) );
CLKBUF_X2 inst_13312 ( .A(net_12516), .Z(net_13274) );
CLKBUF_X2 inst_14317 ( .A(net_14278), .Z(net_14279) );
CLKBUF_X2 inst_8948 ( .A(net_8909), .Z(net_8910) );
AOI22_X2 inst_7369 ( .A1(net_7691), .A2(net_5916), .B2(net_2957), .ZN(net_2953), .B1(net_916) );
NOR4_X2 inst_2172 ( .ZN(net_3249), .A4(net_3120), .A1(net_2632), .A3(net_2474), .A2(net_832) );
CLKBUF_X2 inst_11227 ( .A(net_9500), .Z(net_11189) );
NOR2_X2 inst_2353 ( .ZN(net_5651), .A1(net_5503), .A2(net_4470) );
CLKBUF_X2 inst_11921 ( .A(net_11882), .Z(net_11883) );
CLKBUF_X2 inst_8005 ( .A(net_7966), .Z(net_7967) );
SDFF_X2 inst_667 ( .Q(net_6698), .D(net_6698), .SE(net_3871), .SI(net_3799), .CK(net_11109) );
CLKBUF_X2 inst_13483 ( .A(net_13444), .Z(net_13445) );
NAND3_X2 inst_2762 ( .ZN(net_2339), .A1(net_1426), .A3(net_1274), .A2(net_1013) );
CLKBUF_X2 inst_12646 ( .A(net_12607), .Z(net_12608) );
CLKBUF_X2 inst_8870 ( .A(net_8831), .Z(net_8832) );
NAND2_X4 inst_2896 ( .A1(net_5917), .ZN(net_3406), .A2(net_516) );
SDFF_X2 inst_997 ( .Q(net_6485), .D(net_6485), .SE(net_3904), .SI(net_3821), .CK(net_8406) );
SDFF_X2 inst_857 ( .D(net_7807), .SI(net_7042), .Q(net_7042), .SE(net_3777), .CK(net_10857) );
CLKBUF_X2 inst_8732 ( .A(net_8693), .Z(net_8694) );
INV_X4 inst_4824 ( .ZN(net_1088), .A(net_1087) );
NAND3_X2 inst_2691 ( .ZN(net_3148), .A2(net_3147), .A3(net_3045), .A1(net_3002) );
CLKBUF_X2 inst_14401 ( .A(net_14362), .Z(net_14363) );
DFF_X2 inst_6311 ( .QN(net_7814), .CK(net_10888), .D(x1424) );
OAI22_X2 inst_1511 ( .B1(net_4650), .A1(net_4080), .B2(net_4079), .ZN(net_4075), .A2(net_4074) );
DFF_X1 inst_6403 ( .QN(net_6142), .D(net_5767), .CK(net_8167) );
AOI222_X2 inst_7543 ( .C1(net_7678), .A1(net_7646), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1876), .B1(net_1875) );
CLKBUF_X2 inst_10777 ( .A(net_10738), .Z(net_10739) );
NAND2_X2 inst_4179 ( .A2(net_6823), .ZN(net_771), .A1(net_450) );
CLKBUF_X2 inst_12721 ( .A(net_12682), .Z(net_12683) );
INV_X2 inst_5951 ( .A(net_7769), .ZN(net_407) );
CLKBUF_X2 inst_8977 ( .A(net_8938), .Z(net_8939) );
CLKBUF_X2 inst_7988 ( .A(net_7915), .Z(net_7950) );
DFF_X1 inst_6645 ( .QN(net_7619), .D(net_5209), .CK(net_10298) );
NAND2_X2 inst_4006 ( .ZN(net_1278), .A2(net_666), .A1(net_613) );
NAND2_X1 inst_4243 ( .ZN(net_4684), .A2(net_3989), .A1(net_2189) );
NAND2_X2 inst_3203 ( .ZN(net_4723), .A2(net_3986), .A1(net_1838) );
CLKBUF_X2 inst_14344 ( .A(net_14305), .Z(net_14306) );
CLKBUF_X2 inst_13659 ( .A(net_12887), .Z(net_13621) );
INV_X4 inst_5073 ( .A(net_6553), .ZN(net_1153) );
OAI22_X2 inst_1504 ( .B1(net_4660), .A1(net_4105), .B2(net_4093), .ZN(net_4090), .A2(net_4089) );
NAND2_X2 inst_3403 ( .A2(net_5929), .ZN(net_3375), .A1(net_3374) );
CLKBUF_X2 inst_13951 ( .A(net_13912), .Z(net_13913) );
INV_X2 inst_5830 ( .A(net_1306), .ZN(net_908) );
SDFF_X2 inst_1310 ( .D(net_6386), .SE(net_5799), .SI(net_371), .Q(net_371), .CK(net_13873) );
NAND2_X2 inst_3280 ( .ZN(net_3686), .A1(net_3685), .A2(net_3231) );
CLKBUF_X2 inst_9802 ( .A(net_9763), .Z(net_9764) );
INV_X8 inst_4491 ( .ZN(net_4650), .A(net_3408) );
CLKBUF_X2 inst_9006 ( .A(net_8840), .Z(net_8968) );
AOI222_X2 inst_7518 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2016), .A1(net_2015), .B1(net_2014), .C1(net_2013) );
AOI22_X2 inst_7397 ( .A2(net_3105), .B1(net_2970), .ZN(net_2844), .A1(net_2843), .B2(net_257) );
CLKBUF_X2 inst_11594 ( .A(net_11555), .Z(net_11556) );
NAND3_X2 inst_2823 ( .A2(net_3857), .ZN(net_1827), .A3(net_1826), .A1(net_654) );
CLKBUF_X2 inst_13981 ( .A(net_13942), .Z(net_13943) );
NAND2_X2 inst_3807 ( .A1(net_6632), .A2(net_1624), .ZN(net_1538) );
CLKBUF_X2 inst_13413 ( .A(net_10626), .Z(net_13375) );
SDFF_X2 inst_1069 ( .SI(net_6547), .Q(net_6547), .D(net_3794), .SE(net_3756), .CK(net_11227) );
CLKBUF_X2 inst_12719 ( .A(net_12680), .Z(net_12681) );
CLKBUF_X2 inst_11327 ( .A(net_8194), .Z(net_11289) );
CLKBUF_X2 inst_14153 ( .A(net_8812), .Z(net_14115) );
SDFF_X2 inst_136 ( .Q(net_6214), .SI(net_6213), .SE(net_392), .D(net_148), .CK(net_14228) );
CLKBUF_X2 inst_13083 ( .A(net_10408), .Z(net_13045) );
CLKBUF_X2 inst_11733 ( .A(net_11694), .Z(net_11695) );
CLKBUF_X2 inst_10326 ( .A(net_10287), .Z(net_10288) );
INV_X2 inst_5839 ( .ZN(net_783), .A(net_782) );
NAND2_X2 inst_3541 ( .ZN(net_2526), .A2(net_2149), .A1(net_1198) );
CLKBUF_X2 inst_13837 ( .A(net_13798), .Z(net_13799) );
OAI22_X2 inst_1526 ( .B1(net_4644), .A1(net_4057), .B2(net_4047), .ZN(net_4044), .A2(net_4043) );
CLKBUF_X2 inst_11503 ( .A(net_11464), .Z(net_11465) );
CLKBUF_X2 inst_13825 ( .A(net_8078), .Z(net_13787) );
NOR2_X2 inst_2547 ( .A2(net_7232), .ZN(net_1247), .A1(net_445) );
INV_X4 inst_4637 ( .ZN(net_4185), .A(net_4031) );
SDFF_X2 inst_1047 ( .Q(net_7248), .D(net_7248), .SE(net_3822), .SI(net_344), .CK(net_12664) );
DFF_X1 inst_6860 ( .D(net_2547), .Q(net_197), .CK(net_12077) );
INV_X4 inst_5167 ( .ZN(net_543), .A(net_542) );
NAND2_X2 inst_3850 ( .A1(net_6709), .A2(net_1497), .ZN(net_1486) );
CLKBUF_X2 inst_12582 ( .A(net_10285), .Z(net_12544) );
CLKBUF_X2 inst_8507 ( .A(net_8468), .Z(net_8469) );
CLKBUF_X2 inst_11768 ( .A(net_11729), .Z(net_11730) );
CLKBUF_X2 inst_14368 ( .A(net_11626), .Z(net_14330) );
CLKBUF_X2 inst_12432 ( .A(net_12393), .Z(net_12394) );
CLKBUF_X2 inst_10972 ( .A(net_10933), .Z(net_10934) );
DFF_X1 inst_6744 ( .QN(net_7618), .D(net_4843), .CK(net_12244) );
NAND2_X2 inst_3700 ( .A1(net_7460), .ZN(net_1704), .A2(net_1696) );
OAI21_X2 inst_1858 ( .ZN(net_5260), .B1(net_5230), .A(net_4545), .B2(net_3870) );
OAI21_X2 inst_1786 ( .B1(net_5440), .ZN(net_5405), .A(net_4679), .B2(net_3988) );
CLKBUF_X2 inst_13668 ( .A(net_13629), .Z(net_13630) );
NAND2_X2 inst_3846 ( .A1(net_6694), .A2(net_1497), .ZN(net_1491) );
SDFFR_X2 inst_1334 ( .SI(net_7743), .Q(net_7743), .D(net_4596), .SE(net_3930), .CK(net_13197), .RN(x1822) );
SDFF_X2 inst_496 ( .Q(net_7120), .D(net_7120), .SI(net_3900), .SE(net_3888), .CK(net_8797) );
CLKBUF_X2 inst_10639 ( .A(net_10600), .Z(net_10601) );
CLKBUF_X2 inst_12356 ( .A(net_12317), .Z(net_12318) );
CLKBUF_X2 inst_10304 ( .A(net_8680), .Z(net_10266) );
INV_X4 inst_5369 ( .A(net_7721), .ZN(net_2847) );
INV_X2 inst_5944 ( .A(net_7317), .ZN(net_1770) );
CLKBUF_X2 inst_9011 ( .A(net_8972), .Z(net_8973) );
INV_X2 inst_5733 ( .ZN(net_3958), .A(net_3957) );
DFF_X1 inst_6867 ( .D(net_2548), .QN(net_211), .CK(net_12609) );
INV_X16 inst_6129 ( .ZN(net_4457), .A(net_3842) );
INV_X4 inst_5383 ( .A(net_7384), .ZN(net_826) );
NAND2_X2 inst_3749 ( .A1(net_6909), .A2(net_1639), .ZN(net_1596) );
CLKBUF_X2 inst_12130 ( .A(net_10736), .Z(net_12092) );
AOI22_X2 inst_7273 ( .B1(net_7087), .A1(net_7055), .A2(net_5280), .B2(net_5279), .ZN(net_5275) );
NAND3_X2 inst_2620 ( .ZN(net_5719), .A1(net_5614), .A2(net_5131), .A3(net_4178) );
OAI222_X2 inst_1633 ( .A1(net_5865), .C2(net_5077), .ZN(net_5076), .A2(net_5075), .B2(net_5074), .B1(net_2439), .C1(net_585) );
CLKBUF_X2 inst_12425 ( .A(net_12386), .Z(net_12387) );
CLKBUF_X2 inst_11453 ( .A(net_11414), .Z(net_11415) );
SDFF_X2 inst_1262 ( .D(net_6389), .SE(net_5801), .SI(net_334), .Q(net_334), .CK(net_14304) );
INV_X4 inst_5303 ( .A(net_7581), .ZN(net_1877) );
CLKBUF_X2 inst_9364 ( .A(net_8628), .Z(net_9326) );
SDFF_X2 inst_265 ( .Q(net_6369), .SI(net_6368), .D(net_3525), .SE(net_392), .CK(net_14073) );
CLKBUF_X2 inst_8048 ( .A(net_7971), .Z(net_8010) );
OAI21_X2 inst_2055 ( .B1(net_5899), .B2(net_4457), .ZN(net_4443), .A(net_3555) );
CLKBUF_X2 inst_11702 ( .A(net_11663), .Z(net_11664) );
DFF_X1 inst_6799 ( .D(net_3938), .CK(net_12830), .Q(x786) );
NAND2_X2 inst_3856 ( .A1(net_6699), .A2(net_1497), .ZN(net_1479) );
CLKBUF_X2 inst_12453 ( .A(net_12414), .Z(net_12415) );
AOI21_X2 inst_7783 ( .B1(net_6595), .ZN(net_5912), .B2(net_2583), .A(net_2362) );
INV_X4 inst_5091 ( .ZN(net_2299), .A(net_861) );
INV_X4 inst_5554 ( .A(net_6961), .ZN(net_451) );
CLKBUF_X2 inst_14169 ( .A(net_8799), .Z(net_14131) );
CLKBUF_X2 inst_11650 ( .A(net_11545), .Z(net_11612) );
NAND2_X2 inst_3262 ( .ZN(net_4143), .A1(net_3855), .A2(net_3540) );
CLKBUF_X2 inst_12577 ( .A(net_9155), .Z(net_12539) );
CLKBUF_X2 inst_11482 ( .A(net_11443), .Z(net_11444) );
DFF_X1 inst_6432 ( .QN(net_6075), .D(net_5738), .CK(net_8113) );
INV_X8 inst_4566 ( .ZN(net_1645), .A(net_490) );
CLKBUF_X2 inst_10716 ( .A(net_7866), .Z(net_10678) );
CLKBUF_X2 inst_12993 ( .A(net_11714), .Z(net_12955) );
CLKBUF_X2 inst_10653 ( .A(net_10614), .Z(net_10615) );
DFF_X2 inst_6301 ( .D(net_1692), .QN(net_191), .CK(net_12286) );
SDFF_X2 inst_1077 ( .SI(net_7213), .Q(net_7213), .D(net_3897), .SE(net_3750), .CK(net_7902) );
CLKBUF_X2 inst_7975 ( .A(net_7869), .Z(net_7937) );
AOI22_X2 inst_7249 ( .B1(net_6817), .A1(net_6785), .A2(net_5316), .B2(net_5315), .ZN(net_5311) );
CLKBUF_X2 inst_12956 ( .A(net_12917), .Z(net_12918) );
NAND2_X2 inst_3954 ( .A1(net_6569), .A2(net_1705), .ZN(net_1331) );
CLKBUF_X2 inst_9367 ( .A(net_9328), .Z(net_9329) );
DFF_X1 inst_6461 ( .QN(net_6130), .D(net_5598), .CK(net_10958) );
NAND3_X2 inst_2757 ( .ZN(net_2344), .A3(net_1602), .A1(net_1500), .A2(net_1031) );
SDFF_X2 inst_222 ( .Q(net_6332), .SI(net_6331), .D(net_3661), .SE(net_392), .CK(net_14044) );
OAI21_X2 inst_1932 ( .ZN(net_5113), .A(net_4750), .B2(net_3941), .B1(net_1086) );
CLKBUF_X2 inst_10822 ( .A(net_8859), .Z(net_10784) );
CLKBUF_X2 inst_9733 ( .A(net_8773), .Z(net_9695) );
DFF_X1 inst_6372 ( .QN(net_6290), .D(net_5812), .CK(net_14275) );
CLKBUF_X2 inst_7884 ( .A(net_7830), .Z(net_7846) );
INV_X2 inst_6073 ( .A(net_7288), .ZN(net_1999) );
NAND2_X2 inst_3704 ( .ZN(net_5943), .A2(net_1672), .A1(net_531) );
CLKBUF_X2 inst_13903 ( .A(net_11011), .Z(net_13865) );
CLKBUF_X2 inst_13166 ( .A(net_13127), .Z(net_13128) );
CLKBUF_X2 inst_12218 ( .A(net_9156), .Z(net_12180) );
CLKBUF_X2 inst_11828 ( .A(net_8156), .Z(net_11790) );
DFF_X1 inst_6728 ( .QN(net_7362), .D(net_5327), .CK(net_12701) );
SDFF_X2 inst_1052 ( .Q(net_7241), .D(net_7241), .SE(net_3822), .SI(net_337), .CK(net_9823) );
SDFF_X2 inst_1280 ( .D(net_3894), .SE(net_3256), .SI(net_140), .Q(net_140), .CK(net_8536) );
SDFF_X2 inst_1302 ( .SI(net_7766), .Q(net_7766), .SE(net_5923), .D(net_2746), .CK(net_10772) );
CLKBUF_X2 inst_12740 ( .A(net_8198), .Z(net_12702) );
DFF_X1 inst_6435 ( .QN(net_6078), .D(net_5735), .CK(net_8440) );
INV_X4 inst_5362 ( .A(net_6121), .ZN(net_3617) );
CLKBUF_X2 inst_13904 ( .A(net_13865), .Z(net_13866) );
CLKBUF_X2 inst_9578 ( .A(net_8815), .Z(net_9540) );
INV_X2 inst_6112 ( .A(net_5922), .ZN(net_5921) );
CLKBUF_X2 inst_10609 ( .A(net_10570), .Z(net_10571) );
OAI221_X2 inst_1648 ( .ZN(net_5078), .C2(net_5077), .B2(net_5074), .A(net_4526), .B1(net_2433), .C1(net_1269) );
CLKBUF_X2 inst_13958 ( .A(net_13919), .Z(net_13920) );
INV_X2 inst_5847 ( .A(net_1151), .ZN(net_721) );
SDFF_X2 inst_1079 ( .SI(net_7195), .Q(net_7195), .D(net_3792), .SE(net_3750), .CK(net_10319) );
CLKBUF_X2 inst_13833 ( .A(net_13794), .Z(net_13795) );
DFF_X2 inst_6200 ( .QN(net_6687), .D(net_4398), .CK(net_9719) );
NAND2_X2 inst_3925 ( .A1(net_6847), .A2(net_1521), .ZN(net_1375) );
NAND3_X2 inst_2606 ( .ZN(net_5733), .A1(net_5628), .A2(net_5171), .A3(net_4193) );
CLKBUF_X2 inst_9837 ( .A(net_9158), .Z(net_9799) );
NAND2_X1 inst_4314 ( .ZN(net_4552), .A2(net_3866), .A1(net_1867) );
NOR2_X2 inst_2523 ( .A1(net_6406), .ZN(net_1042), .A2(net_938) );
SDFF_X2 inst_506 ( .SI(net_6765), .Q(net_6765), .D(net_3890), .SE(net_3816), .CK(net_11756) );
CLKBUF_X2 inst_13569 ( .A(net_10150), .Z(net_13531) );
CLKBUF_X2 inst_10662 ( .A(net_10623), .Z(net_10624) );
CLKBUF_X2 inst_11782 ( .A(net_11743), .Z(net_11744) );
CLKBUF_X2 inst_8572 ( .A(net_8330), .Z(net_8534) );
SDFF_X2 inst_134 ( .Q(net_6216), .SI(net_6215), .SE(net_392), .D(net_150), .CK(net_14235) );
NOR2_X2 inst_2409 ( .ZN(net_3730), .A2(net_3335), .A1(net_3031) );
NAND2_X2 inst_3322 ( .ZN(net_3602), .A1(net_3601), .A2(net_3228) );
CLKBUF_X2 inst_10835 ( .A(net_10796), .Z(net_10797) );
SDFF_X2 inst_1085 ( .SI(net_7082), .Q(net_7082), .D(net_3775), .SE(net_3747), .CK(net_8193) );
SDFF_X2 inst_1323 ( .D(net_6384), .SE(net_5801), .SI(net_329), .Q(net_329), .CK(net_14288) );
NAND2_X2 inst_3425 ( .A2(net_5892), .ZN(net_3323), .A1(net_644) );
CLKBUF_X2 inst_14048 ( .A(net_14009), .Z(net_14010) );
NOR2_X2 inst_2328 ( .A2(net_6290), .A1(net_5843), .ZN(net_5813) );
CLKBUF_X2 inst_10464 ( .A(net_10420), .Z(net_10426) );
CLKBUF_X2 inst_8791 ( .A(net_8752), .Z(net_8753) );
CLKBUF_X2 inst_8060 ( .A(net_8016), .Z(net_8022) );
NAND3_X2 inst_2655 ( .ZN(net_3945), .A3(net_3389), .A2(net_2947), .A1(net_2825) );
SDFF_X2 inst_160 ( .Q(net_6254), .SI(net_6253), .D(net_3575), .SE(net_392), .CK(net_13536) );
OAI21_X2 inst_1720 ( .ZN(net_5574), .B1(net_5537), .A(net_4684), .B2(net_3989) );
CLKBUF_X2 inst_8889 ( .A(net_8779), .Z(net_8851) );
INV_X2 inst_5779 ( .ZN(net_2896), .A(net_266) );
CLKBUF_X2 inst_14420 ( .A(net_14381), .Z(net_14382) );
CLKBUF_X2 inst_13541 ( .A(net_9867), .Z(net_13503) );
NAND2_X2 inst_2912 ( .ZN(net_5781), .A2(net_5769), .A1(net_401) );
CLKBUF_X2 inst_9243 ( .A(net_8162), .Z(net_9205) );
AOI22_X2 inst_7450 ( .A2(net_2949), .B2(net_2679), .ZN(net_843), .A1(net_842), .B1(net_841) );
SDFF_X2 inst_762 ( .Q(net_6885), .D(net_6885), .SE(net_3901), .SI(net_3796), .CK(net_8873) );
SDFF_X2 inst_370 ( .SI(net_7642), .Q(net_7642), .D(net_4788), .SE(net_3867), .CK(net_13391) );
CLKBUF_X2 inst_10414 ( .A(net_10375), .Z(net_10376) );
AND2_X4 inst_7825 ( .ZN(net_3115), .A2(net_3045), .A1(net_1245) );
NAND2_X2 inst_3025 ( .A1(net_6850), .A2(net_5004), .ZN(net_4984) );
SDFF_X2 inst_1265 ( .Q(net_7231), .D(net_3423), .SI(net_3422), .SE(net_2249), .CK(net_10468) );
CLKBUF_X2 inst_10669 ( .A(net_10630), .Z(net_10631) );
AOI222_X2 inst_7530 ( .B2(net_2135), .C2(net_2133), .ZN(net_1915), .A1(net_1914), .B1(net_1913), .C1(net_1912), .A2(net_1910) );
CLKBUF_X2 inst_10434 ( .A(net_10395), .Z(net_10396) );
CLKBUF_X2 inst_8371 ( .A(net_8332), .Z(net_8333) );
INV_X8 inst_4530 ( .ZN(net_3439), .A(net_2645) );
CLKBUF_X2 inst_11882 ( .A(net_11843), .Z(net_11844) );
CLKBUF_X2 inst_8176 ( .A(net_8137), .Z(net_8138) );
CLKBUF_X2 inst_11288 ( .A(net_10250), .Z(net_11250) );
SDFF_X2 inst_1321 ( .D(net_6385), .SE(net_6052), .SI(net_310), .Q(net_310), .CK(net_13804) );
SDFF_X2 inst_1012 ( .SI(net_6505), .Q(net_6505), .SE(net_3886), .D(net_3776), .CK(net_8850) );
CLKBUF_X2 inst_12768 ( .A(net_12729), .Z(net_12730) );
INV_X4 inst_5255 ( .ZN(net_3920), .A(net_1679) );
CLKBUF_X2 inst_13843 ( .A(net_13475), .Z(net_13805) );
CLKBUF_X2 inst_8341 ( .A(net_8302), .Z(net_8303) );
OAI21_X2 inst_1956 ( .B1(net_5206), .ZN(net_5064), .A(net_4709), .B2(net_3986) );
CLKBUF_X2 inst_8378 ( .A(net_8339), .Z(net_8340) );
NAND2_X2 inst_3492 ( .ZN(net_2733), .A2(net_2628), .A1(net_2585) );
CLKBUF_X2 inst_10687 ( .A(net_7838), .Z(net_10649) );
CLKBUF_X2 inst_10935 ( .A(net_10896), .Z(net_10897) );
SDFF_X2 inst_751 ( .Q(net_6873), .D(net_6873), .SE(net_3901), .SI(net_3812), .CK(net_11485) );
CLKBUF_X2 inst_14032 ( .A(net_13993), .Z(net_13994) );
CLKBUF_X2 inst_9015 ( .A(net_7972), .Z(net_8977) );
NAND2_X2 inst_3149 ( .ZN(net_4814), .A2(net_4153), .A1(net_2154) );
NAND2_X1 inst_4283 ( .ZN(net_4584), .A2(net_3867), .A1(net_1846) );
NOR2_X2 inst_2471 ( .A2(net_5778), .ZN(net_2681), .A1(net_2611) );
NAND2_X2 inst_4034 ( .A1(net_6538), .A2(net_1645), .ZN(net_1018) );
CLKBUF_X2 inst_13570 ( .A(net_8252), .Z(net_13532) );
SDFF_X2 inst_377 ( .SI(net_7672), .Q(net_7672), .D(net_4789), .SE(net_3866), .CK(net_13240) );
DFFR_X2 inst_6993 ( .QN(net_7703), .D(net_3359), .CK(net_10367), .RN(x1822) );
CLKBUF_X2 inst_10157 ( .A(net_10076), .Z(net_10119) );
INV_X4 inst_4760 ( .ZN(net_2872), .A(net_2786) );
NAND2_X2 inst_3946 ( .A1(net_6841), .A2(net_1521), .ZN(net_1342) );
NAND2_X2 inst_3244 ( .ZN(net_3993), .A2(net_3992), .A1(net_3983) );
DFFS_X2 inst_6953 ( .QN(net_6408), .D(net_2721), .CK(net_14399), .SN(x1822) );
NAND2_X2 inst_3920 ( .A1(net_7099), .A2(net_1675), .ZN(net_1383) );
DFF_X1 inst_6920 ( .D(net_2408), .Q(net_255), .CK(net_13270) );
NAND2_X2 inst_3821 ( .A1(net_7169), .A2(net_1637), .ZN(net_1524) );
AOI22_X2 inst_7443 ( .ZN(net_5399), .A2(net_1225), .B1(net_1223), .B2(net_364), .A1(net_352) );
INV_X2 inst_5981 ( .ZN(net_1135), .A(net_125) );
NAND2_X2 inst_3018 ( .A1(net_6891), .A2(net_5006), .ZN(net_4991) );
CLKBUF_X2 inst_13750 ( .A(net_13711), .Z(net_13712) );
NAND2_X2 inst_3078 ( .A1(net_6447), .ZN(net_4926), .A2(net_4925) );
CLKBUF_X2 inst_12779 ( .A(net_12740), .Z(net_12741) );
INV_X2 inst_5792 ( .A(net_5961), .ZN(net_2236) );
CLKBUF_X2 inst_12675 ( .A(net_12636), .Z(net_12637) );
CLKBUF_X2 inst_13579 ( .A(net_13540), .Z(net_13541) );
CLKBUF_X2 inst_13330 ( .A(net_11976), .Z(net_13292) );
CLKBUF_X2 inst_9731 ( .A(net_9692), .Z(net_9693) );
INV_X4 inst_4623 ( .ZN(net_4199), .A(net_4059) );
INV_X2 inst_5926 ( .A(net_7346), .ZN(net_2161) );
INV_X4 inst_5054 ( .A(net_7815), .ZN(net_3775) );
NAND2_X2 inst_3835 ( .A1(net_7110), .A2(net_1675), .ZN(net_1504) );
INV_X4 inst_4627 ( .ZN(net_4195), .A(net_4050) );
CLKBUF_X2 inst_14429 ( .A(net_14390), .Z(net_14391) );
CLKBUF_X2 inst_13559 ( .A(net_13520), .Z(net_13521) );
CLKBUF_X2 inst_12414 ( .A(net_12258), .Z(net_12376) );
CLKBUF_X2 inst_14191 ( .A(net_14152), .Z(net_14153) );
XNOR2_X2 inst_107 ( .B(net_6420), .ZN(net_1039), .A(net_807) );
OAI21_X2 inst_2117 ( .B2(net_3297), .ZN(net_3296), .A(net_3079), .B1(net_3071) );
SDFF_X2 inst_990 ( .Q(net_6476), .D(net_6476), .SE(net_3904), .SI(net_3805), .CK(net_10843) );
CLKBUF_X2 inst_12381 ( .A(net_11560), .Z(net_12343) );
CLKBUF_X2 inst_10412 ( .A(net_10373), .Z(net_10374) );
NAND2_X2 inst_3140 ( .ZN(net_4823), .A2(net_4153), .A1(net_2152) );
INV_X4 inst_4710 ( .ZN(net_2979), .A(net_2978) );
CLKBUF_X2 inst_13812 ( .A(net_8887), .Z(net_13774) );
CLKBUF_X2 inst_12035 ( .A(net_11996), .Z(net_11997) );
NAND2_X2 inst_3628 ( .ZN(net_1955), .A1(net_1289), .A2(net_1120) );
CLKBUF_X2 inst_11941 ( .A(net_10577), .Z(net_11903) );
CLKBUF_X2 inst_12308 ( .A(net_11250), .Z(net_12270) );
CLKBUF_X2 inst_10093 ( .A(net_10054), .Z(net_10055) );
NOR2_X2 inst_2366 ( .ZN(net_5270), .A2(net_4625), .A1(net_4467) );
CLKBUF_X2 inst_11200 ( .A(net_10473), .Z(net_11162) );
INV_X4 inst_4642 ( .ZN(net_4180), .A(net_4019) );
AOI22_X2 inst_7340 ( .B2(net_3439), .ZN(net_3302), .B1(net_3077), .A2(net_2712), .A1(net_152) );
INV_X4 inst_5049 ( .A(net_6958), .ZN(net_1148) );
NAND2_X2 inst_3316 ( .ZN(net_3614), .A1(net_3613), .A2(net_3228) );
CLKBUF_X2 inst_9385 ( .A(net_8521), .Z(net_9347) );
CLKBUF_X2 inst_11343 ( .A(net_11304), .Z(net_11305) );
CLKBUF_X2 inst_14155 ( .A(net_14116), .Z(net_14117) );
NAND2_X1 inst_4411 ( .A2(net_5962), .A1(net_5961), .ZN(net_2881) );
CLKBUF_X2 inst_11471 ( .A(net_11432), .Z(net_11433) );
CLKBUF_X2 inst_13998 ( .A(net_10175), .Z(net_13960) );
AOI21_X2 inst_7772 ( .B1(net_7142), .ZN(net_4079), .B2(net_2582), .A(net_2323) );
NAND2_X2 inst_4014 ( .A1(net_6943), .A2(net_1654), .ZN(net_1038) );
INV_X4 inst_4605 ( .ZN(net_4239), .A(net_4096) );
NAND2_X2 inst_3694 ( .ZN(net_1736), .A1(net_1278), .A2(net_1098) );
INV_X4 inst_4882 ( .A(net_3048), .ZN(net_1079) );
CLKBUF_X2 inst_11207 ( .A(net_11168), .Z(net_11169) );
CLKBUF_X2 inst_10351 ( .A(net_9578), .Z(net_10313) );
NAND3_X2 inst_2698 ( .ZN(net_2694), .A3(net_2570), .A2(net_2432), .A1(net_2268) );
SDFF_X2 inst_1237 ( .SI(net_6530), .Q(net_6530), .D(net_3894), .SE(net_3755), .CK(net_8619) );
CLKBUF_X2 inst_12873 ( .A(net_12834), .Z(net_12835) );
CLKBUF_X2 inst_9908 ( .A(net_9869), .Z(net_9870) );
NOR2_X2 inst_2518 ( .ZN(net_1062), .A2(net_667), .A1(net_611) );
NAND2_X2 inst_3460 ( .A2(net_5966), .ZN(net_2892), .A1(net_2891) );
INV_X4 inst_5152 ( .A(net_894), .ZN(net_564) );
INV_X4 inst_5544 ( .A(net_7251), .ZN(net_2039) );
OAI21_X2 inst_2075 ( .ZN(net_4417), .B1(net_4416), .B2(net_4415), .A(net_3514) );
NAND2_X2 inst_3062 ( .A1(net_7158), .A2(net_4954), .ZN(net_4943) );
NAND2_X2 inst_3310 ( .ZN(net_3626), .A1(net_3625), .A2(net_3231) );
OAI21_X2 inst_1911 ( .ZN(net_5157), .B1(net_4872), .A(net_4759), .B2(net_3941) );
DFF_X2 inst_6267 ( .QN(net_5962), .D(net_2633), .CK(net_10727) );
INV_X4 inst_5689 ( .ZN(net_530), .A(net_293) );
CLKBUF_X2 inst_14249 ( .A(net_9249), .Z(net_14211) );
CLKBUF_X2 inst_10841 ( .A(net_8509), .Z(net_10803) );
CLKBUF_X2 inst_13459 ( .A(net_13420), .Z(net_13421) );
SDFF_X2 inst_585 ( .Q(net_6583), .D(net_6583), .SE(net_3823), .SI(net_3791), .CK(net_10668) );
INV_X4 inst_5100 ( .ZN(net_2419), .A(net_618) );
CLKBUF_X2 inst_8536 ( .A(net_8076), .Z(net_8498) );
CLKBUF_X2 inst_8816 ( .A(net_8777), .Z(net_8778) );
CLKBUF_X2 inst_13967 ( .A(net_13928), .Z(net_13929) );
INV_X4 inst_5435 ( .A(net_6171), .ZN(net_3554) );
INV_X4 inst_5107 ( .A(net_1726), .ZN(net_814) );
INV_X2 inst_6013 ( .A(net_7603), .ZN(net_1413) );
INV_X2 inst_5763 ( .ZN(net_3030), .A(net_2926) );
CLKBUF_X2 inst_11171 ( .A(net_10818), .Z(net_11133) );
SDFF_X2 inst_383 ( .SI(net_7678), .Q(net_7678), .D(net_4785), .SE(net_3866), .CK(net_10269) );
CLKBUF_X2 inst_12137 ( .A(net_12098), .Z(net_12099) );
DFF_X1 inst_6453 ( .QN(net_6092), .D(net_5717), .CK(net_9207) );
NOR2_X2 inst_2428 ( .ZN(net_3432), .A2(net_3122), .A1(net_3048) );
CLKBUF_X2 inst_11793 ( .A(net_11754), .Z(net_11755) );
CLKBUF_X2 inst_13561 ( .A(net_13522), .Z(net_13523) );
INV_X4 inst_5115 ( .ZN(net_691), .A(net_602) );
CLKBUF_X2 inst_14382 ( .A(net_14343), .Z(net_14344) );
AOI21_X2 inst_7670 ( .B1(net_7004), .ZN(net_4230), .A(net_2470), .B2(net_1100) );
DFFR_X2 inst_7031 ( .QN(net_5988), .D(net_3137), .CK(net_13224), .RN(x1822) );
NAND2_X2 inst_4132 ( .ZN(net_1267), .A2(net_1222), .A1(net_336) );
AOI21_X2 inst_7679 ( .B1(net_6996), .ZN(net_4600), .A(net_2472), .B2(net_1100) );
CLKBUF_X2 inst_9765 ( .A(net_8603), .Z(net_9727) );
AOI222_X2 inst_7553 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1843), .A1(net_1842), .B1(net_1841), .C1(net_1840) );
SDFF_X2 inst_1124 ( .SI(net_6674), .Q(net_6674), .D(net_3784), .SE(net_3471), .CK(net_12135) );
NAND2_X2 inst_4086 ( .A1(net_6791), .A2(net_1651), .ZN(net_966) );
CLKBUF_X2 inst_11091 ( .A(net_11052), .Z(net_11053) );
CLKBUF_X2 inst_11801 ( .A(net_10141), .Z(net_11763) );
INV_X4 inst_5372 ( .A(net_6103), .ZN(net_3497) );
NOR2_X2 inst_2555 ( .A1(net_6045), .A2(net_6039), .ZN(net_2887) );
NAND2_X2 inst_3375 ( .ZN(net_3496), .A1(net_3495), .A2(net_3225) );
SDFF_X2 inst_234 ( .SI(net_6359), .Q(net_6320), .D(net_3667), .SE(net_392), .CK(net_14003) );
CLKBUF_X2 inst_13922 ( .A(net_11138), .Z(net_13884) );
DFFR_X2 inst_6966 ( .QN(net_7781), .D(net_5918), .CK(net_10250), .RN(x1822) );
INV_X4 inst_5293 ( .A(net_6018), .ZN(net_645) );
CLKBUF_X2 inst_13447 ( .A(net_13408), .Z(net_13409) );
INV_X4 inst_5240 ( .ZN(net_630), .A(net_450) );
CLKBUF_X2 inst_12450 ( .A(net_9969), .Z(net_12412) );
INV_X4 inst_5343 ( .A(net_6091), .ZN(net_3519) );
CLKBUF_X2 inst_12398 ( .A(net_12359), .Z(net_12360) );
NAND2_X2 inst_3714 ( .A1(net_6768), .A2(net_1635), .ZN(net_1632) );
CLKBUF_X2 inst_12317 ( .A(net_12278), .Z(net_12279) );
CLKBUF_X2 inst_12269 ( .A(net_8205), .Z(net_12231) );
INV_X4 inst_5285 ( .A(net_7410), .ZN(net_2190) );
CLKBUF_X2 inst_13975 ( .A(net_13621), .Z(net_13937) );
DFF_X1 inst_6658 ( .QN(net_7665), .D(net_5187), .CK(net_13273) );
INV_X4 inst_5611 ( .A(net_6074), .ZN(net_3607) );
SDFF_X2 inst_1304 ( .SE(net_7378), .Q(net_7378), .D(net_2991), .SI(net_2990), .CK(net_9471) );
NAND2_X2 inst_3429 ( .ZN(net_3219), .A2(net_3103), .A1(net_2771) );
SDFFR_X2 inst_1328 ( .SI(net_7737), .Q(net_7737), .SE(net_5683), .D(net_4596), .CK(net_10333), .RN(x1822) );
CLKBUF_X2 inst_9027 ( .A(net_8988), .Z(net_8989) );
CLKBUF_X2 inst_8429 ( .A(net_8390), .Z(net_8391) );
DFF_X1 inst_6815 ( .D(net_3204), .CK(net_10819), .Q(x217) );
NAND2_X2 inst_3292 ( .ZN(net_3662), .A1(net_3661), .A2(net_3229) );
CLKBUF_X2 inst_8575 ( .A(net_8227), .Z(net_8537) );
OAI21_X2 inst_1776 ( .B1(net_5436), .ZN(net_5418), .A(net_4697), .B2(net_3989) );
AOI21_X2 inst_7751 ( .B1(net_6873), .ZN(net_4101), .B2(net_2579), .A(net_2352) );
INV_X4 inst_5024 ( .A(net_7228), .ZN(net_665) );
NOR2_X2 inst_2335 ( .A2(net_6283), .A1(net_5843), .ZN(net_5806) );
AOI21_X2 inst_7715 ( .B1(net_6862), .ZN(net_4485), .B2(net_2579), .A(net_2345) );
CLKBUF_X2 inst_13157 ( .A(net_9693), .Z(net_13119) );
SDFF_X2 inst_919 ( .Q(net_7157), .D(net_7157), .SE(net_3903), .SI(net_3795), .CK(net_8704) );
CLKBUF_X2 inst_10530 ( .A(net_10491), .Z(net_10492) );
CLKBUF_X2 inst_12772 ( .A(net_12733), .Z(net_12734) );
SDFF_X2 inst_598 ( .Q(net_6591), .D(net_6591), .SE(net_3830), .SI(net_3792), .CK(net_12914) );
OAI21_X2 inst_1916 ( .B1(net_5345), .ZN(net_5148), .A(net_4748), .B2(net_3941) );
CLKBUF_X2 inst_9705 ( .A(net_9666), .Z(net_9667) );
OAI22_X2 inst_1624 ( .B1(net_6421), .A2(net_2820), .ZN(net_2738), .B2(net_2718), .A1(net_1703) );
CLKBUF_X2 inst_14057 ( .A(net_14018), .Z(net_14019) );
CLKBUF_X2 inst_10595 ( .A(net_10556), .Z(net_10557) );
CLKBUF_X2 inst_12403 ( .A(net_12364), .Z(net_12365) );
OAI21_X2 inst_1797 ( .ZN(net_5393), .A(net_4721), .B2(net_3986), .B1(net_1075) );
CLKBUF_X2 inst_10728 ( .A(net_10689), .Z(net_10690) );
NAND2_X2 inst_3167 ( .ZN(net_4766), .A2(net_3941), .A1(net_2067) );
CLKBUF_X2 inst_13501 ( .A(net_13462), .Z(net_13463) );
NAND2_X1 inst_4408 ( .A2(net_3087), .ZN(net_2909), .A1(net_2834) );
NAND3_X2 inst_2708 ( .ZN(net_2469), .A2(net_1817), .A3(net_1593), .A1(net_1408) );
CLKBUF_X2 inst_14029 ( .A(net_8600), .Z(net_13991) );
DFF_X2 inst_6197 ( .Q(net_6395), .D(net_6394), .CK(net_13848) );
CLKBUF_X2 inst_9866 ( .A(net_9827), .Z(net_9828) );
NAND2_X2 inst_3530 ( .ZN(net_2537), .A2(net_2104), .A1(net_1374) );
INV_X4 inst_5009 ( .A(net_7820), .ZN(net_3794) );
INV_X4 inst_4785 ( .ZN(net_2640), .A(net_1658) );
CLKBUF_X2 inst_13552 ( .A(net_9072), .Z(net_13514) );
AOI21_X2 inst_7785 ( .B1(net_7071), .ZN(net_4173), .A(net_2336), .B2(net_791) );
NAND3_X2 inst_2592 ( .ZN(net_5747), .A1(net_5642), .A2(net_5229), .A3(net_4206) );
SDFF_X2 inst_325 ( .SI(net_7490), .Q(net_7490), .D(net_5094), .SE(net_3989), .CK(net_9777) );
DFF_X1 inst_6502 ( .QN(net_7424), .D(net_5528), .CK(net_12116) );
CLKBUF_X2 inst_12752 ( .A(net_12339), .Z(net_12714) );
CLKBUF_X2 inst_8858 ( .A(net_8812), .Z(net_8820) );
INV_X4 inst_4769 ( .ZN(net_2435), .A(net_1932) );
AOI22_X2 inst_7331 ( .A2(net_3426), .B2(net_3425), .ZN(net_3415), .B1(net_2569), .A1(net_1246) );
SDFF_X2 inst_1197 ( .SI(net_7061), .Q(net_7061), .D(net_3806), .SE(net_3742), .CK(net_11846) );
NAND2_X2 inst_3116 ( .A1(net_6588), .A2(net_4897), .ZN(net_4885) );
NAND2_X1 inst_4378 ( .ZN(net_4349), .A2(net_3859), .A1(net_2077) );
CLKBUF_X2 inst_10544 ( .A(net_10505), .Z(net_10506) );
CLKBUF_X2 inst_9682 ( .A(net_9643), .Z(net_9644) );
DFFR_X2 inst_6958 ( .QN(net_7728), .D(net_5775), .CK(net_9620), .RN(x1822) );
SDFF_X2 inst_955 ( .SI(net_7171), .Q(net_7171), .SE(net_3819), .D(net_3814), .CK(net_10486) );
XNOR2_X2 inst_114 ( .ZN(net_2393), .B(net_1199), .A(net_820) );
CLKBUF_X2 inst_11767 ( .A(net_11728), .Z(net_11729) );
DFFR_X1 inst_7116 ( .QN(net_5854), .D(net_5794), .CK(net_9466), .RN(x1822) );
NOR2_X4 inst_2278 ( .ZN(net_3843), .A1(net_3403), .A2(net_3234) );
CLKBUF_X2 inst_11041 ( .A(net_11002), .Z(net_11003) );
INV_X4 inst_4866 ( .A(net_2708), .ZN(net_1103) );
CLKBUF_X2 inst_11415 ( .A(net_11376), .Z(net_11377) );
CLKBUF_X2 inst_7924 ( .A(net_7885), .Z(net_7886) );
AND3_X2 inst_7800 ( .ZN(net_3334), .A3(net_3096), .A2(net_2929), .A1(net_2928) );
CLKBUF_X2 inst_9519 ( .A(net_9480), .Z(net_9481) );
NAND2_X2 inst_4150 ( .A2(net_1225), .ZN(net_1074), .A1(net_360) );
CLKBUF_X2 inst_9630 ( .A(net_8947), .Z(net_9592) );
INV_X2 inst_5851 ( .ZN(net_676), .A(net_675) );
CLKBUF_X2 inst_12371 ( .A(net_8124), .Z(net_12333) );
SDFF_X2 inst_534 ( .SI(net_7807), .Q(net_6605), .D(net_6605), .SE(net_3830), .CK(net_12932) );
CLKBUF_X2 inst_12422 ( .A(net_9399), .Z(net_12384) );
DFF_X1 inst_6665 ( .QN(net_7250), .D(net_5167), .CK(net_12731) );
CLKBUF_X2 inst_8636 ( .A(net_8597), .Z(net_8598) );
CLKBUF_X2 inst_13816 ( .A(net_13777), .Z(net_13778) );
CLKBUF_X2 inst_12502 ( .A(net_9269), .Z(net_12464) );
CLKBUF_X2 inst_9033 ( .A(net_8401), .Z(net_8995) );
CLKBUF_X2 inst_10682 ( .A(net_10643), .Z(net_10644) );
DFFR_X1 inst_7117 ( .QN(net_5853), .D(net_5793), .CK(net_12811), .RN(x1822) );
INV_X4 inst_5618 ( .A(net_7728), .ZN(net_2757) );
CLKBUF_X2 inst_13663 ( .A(net_13624), .Z(net_13625) );
CLKBUF_X2 inst_11142 ( .A(net_11103), .Z(net_11104) );
NAND2_X4 inst_2842 ( .ZN(net_5536), .A1(net_5014), .A2(net_5013) );
INV_X2 inst_5711 ( .ZN(net_4255), .A(net_4133) );
INV_X4 inst_5193 ( .ZN(net_1694), .A(net_510) );
OAI21_X2 inst_2084 ( .B2(net_4415), .ZN(net_4406), .B1(net_4405), .A(net_3486) );
NAND2_X4 inst_2836 ( .ZN(net_5556), .A1(net_5026), .A2(net_5025) );
NAND2_X2 inst_3792 ( .A1(net_6498), .A2(net_1642), .ZN(net_1553) );
NAND2_X1 inst_4336 ( .ZN(net_4391), .A2(net_3853), .A1(net_2020) );
CLKBUF_X2 inst_12310 ( .A(net_11855), .Z(net_12272) );
CLKBUF_X2 inst_11534 ( .A(net_8918), .Z(net_11496) );
CLKBUF_X2 inst_8203 ( .A(net_8032), .Z(net_8165) );
CLKBUF_X2 inst_10424 ( .A(net_10385), .Z(net_10386) );
NAND3_X2 inst_2770 ( .ZN(net_2330), .A3(net_1584), .A1(net_1483), .A2(net_989) );
CLKBUF_X2 inst_11735 ( .A(net_11696), .Z(net_11697) );
CLKBUF_X2 inst_9184 ( .A(net_9145), .Z(net_9146) );
INV_X4 inst_4573 ( .ZN(net_5788), .A(net_5787) );
NAND2_X2 inst_3444 ( .ZN(net_3160), .A1(net_3159), .A2(net_3158) );
AOI22_X2 inst_7284 ( .B1(net_7221), .A1(net_7189), .A2(net_5244), .B2(net_5243), .ZN(net_5229) );
CLKBUF_X2 inst_10848 ( .A(net_10809), .Z(net_10810) );
SDFF_X2 inst_803 ( .Q(net_6976), .D(net_6976), .SE(net_3891), .SI(net_3812), .CK(net_8224) );
CLKBUF_X2 inst_12011 ( .A(net_9099), .Z(net_11973) );
CLKBUF_X2 inst_9295 ( .A(net_9256), .Z(net_9257) );
INV_X4 inst_4732 ( .A(net_3200), .ZN(net_3196) );
NOR2_X2 inst_2348 ( .ZN(net_5656), .A1(net_5508), .A2(net_4475) );
NAND2_X2 inst_4021 ( .A1(net_6927), .A2(net_1654), .ZN(net_1031) );
CLKBUF_X2 inst_10312 ( .A(net_10273), .Z(net_10274) );
CLKBUF_X2 inst_11936 ( .A(net_11897), .Z(net_11898) );
CLKBUF_X2 inst_11059 ( .A(net_11020), .Z(net_11021) );
SDFF_X2 inst_662 ( .Q(net_6721), .D(net_6721), .SE(net_3871), .SI(net_3789), .CK(net_11352) );
OAI22_X2 inst_1533 ( .B1(net_4637), .ZN(net_4031), .A1(net_4030), .A2(net_4029), .B2(net_4028) );
NAND2_X2 inst_3495 ( .A2(net_2644), .ZN(net_2624), .A1(net_623) );
CLKBUF_X2 inst_9827 ( .A(net_9467), .Z(net_9789) );
AOI21_X2 inst_7741 ( .B1(net_7145), .ZN(net_4072), .B2(net_2582), .A(net_2321) );
CLKBUF_X2 inst_8290 ( .A(net_8251), .Z(net_8252) );
CLKBUF_X2 inst_11046 ( .A(net_11007), .Z(net_11008) );
CLKBUF_X2 inst_11114 ( .A(net_11075), .Z(net_11076) );
CLKBUF_X2 inst_12491 ( .A(net_12452), .Z(net_12453) );
AOI21_X2 inst_7713 ( .B1(net_6878), .ZN(net_4091), .B2(net_2579), .A(net_2348) );
INV_X4 inst_5080 ( .ZN(net_3854), .A(net_3227) );
INV_X4 inst_4666 ( .ZN(net_3996), .A(net_3745) );
CLKBUF_X2 inst_14115 ( .A(net_14076), .Z(net_14077) );
OAI22_X2 inst_1465 ( .B2(net_5087), .ZN(net_4397), .A1(net_4148), .A2(net_3828), .B1(net_1181) );
CLKBUF_X2 inst_12653 ( .A(net_9076), .Z(net_12615) );
INV_X4 inst_5030 ( .ZN(net_760), .A(net_662) );
XNOR2_X2 inst_53 ( .ZN(net_2248), .A(net_1919), .B(net_887) );
INV_X4 inst_5265 ( .A(net_826), .ZN(net_425) );
CLKBUF_X2 inst_13009 ( .A(net_10605), .Z(net_12971) );
DFF_X1 inst_6550 ( .Q(net_7775), .D(net_5607), .CK(net_10425) );
NAND3_X2 inst_2614 ( .ZN(net_5725), .A1(net_5620), .A2(net_5137), .A3(net_4184) );
NAND2_X2 inst_3337 ( .ZN(net_3572), .A1(net_3571), .A2(net_3225) );
CLKBUF_X2 inst_10513 ( .A(net_10474), .Z(net_10475) );
NAND2_X2 inst_4215 ( .A2(net_6411), .A1(net_6410), .ZN(net_2275) );
NAND2_X2 inst_4090 ( .A1(net_7213), .A2(net_1648), .ZN(net_962) );
SDFF_X2 inst_999 ( .Q(net_6486), .D(net_6486), .SE(net_3904), .SI(net_3801), .CK(net_8060) );
AND2_X4 inst_7805 ( .A1(net_7767), .ZN(net_4805), .A2(net_4304) );
CLKBUF_X2 inst_12378 ( .A(net_12339), .Z(net_12340) );
CLKBUF_X2 inst_8083 ( .A(net_8044), .Z(net_8045) );
OAI21_X2 inst_2111 ( .ZN(net_3457), .B2(net_3455), .A(net_3373), .B1(net_402) );
OAI21_X2 inst_1846 ( .B1(net_5349), .ZN(net_5326), .A(net_4367), .B2(net_3853) );
CLKBUF_X2 inst_8419 ( .A(net_8380), .Z(net_8381) );
CLKBUF_X2 inst_13943 ( .A(net_11191), .Z(net_13905) );
OAI21_X2 inst_2139 ( .ZN(net_2811), .A(net_506), .B1(net_264), .B2(net_262) );
NAND2_X1 inst_4278 ( .ZN(net_4589), .A2(net_3867), .A1(net_1895) );
OAI22_X2 inst_1463 ( .B2(net_5913), .B1(net_4637), .A2(net_4605), .ZN(net_4603), .A1(net_4012) );
CLKBUF_X2 inst_14242 ( .A(net_14203), .Z(net_14204) );
CLKBUF_X2 inst_10236 ( .A(net_10127), .Z(net_10198) );
SDFF_X2 inst_186 ( .Q(net_6268), .SI(net_6267), .D(net_3479), .SE(net_392), .CK(net_13914) );
CLKBUF_X2 inst_9665 ( .A(net_9626), .Z(net_9627) );
NAND2_X1 inst_4271 ( .ZN(net_4643), .A2(net_3993), .A1(net_1409) );
CLKBUF_X2 inst_13463 ( .A(net_11733), .Z(net_13425) );
CLKBUF_X2 inst_10756 ( .A(net_9364), .Z(net_10718) );
SDFF_X2 inst_759 ( .Q(net_6881), .D(net_6881), .SE(net_3901), .SI(net_3805), .CK(net_10898) );
CLKBUF_X2 inst_11655 ( .A(net_11220), .Z(net_11617) );
CLKBUF_X2 inst_9820 ( .A(net_9616), .Z(net_9782) );
NAND2_X2 inst_3071 ( .A1(net_7151), .A2(net_4954), .ZN(net_4934) );
CLKBUF_X2 inst_10395 ( .A(net_10356), .Z(net_10357) );
CLKBUF_X2 inst_13192 ( .A(net_12686), .Z(net_13154) );
CLKBUF_X2 inst_11963 ( .A(net_11924), .Z(net_11925) );
CLKBUF_X2 inst_13536 ( .A(net_13497), .Z(net_13498) );
CLKBUF_X2 inst_8283 ( .A(net_8244), .Z(net_8245) );
SDFF_X2 inst_863 ( .SI(net_7048), .Q(net_7048), .D(net_3783), .SE(net_3777), .CK(net_9018) );
CLKBUF_X2 inst_8669 ( .A(net_8630), .Z(net_8631) );
DFF_X2 inst_6315 ( .Q(net_7799), .CK(net_10949), .D(x1550) );
OR2_X4 inst_1385 ( .A2(net_6184), .ZN(net_3087), .A1(net_1701) );
DFF_X1 inst_6513 ( .QN(net_7444), .D(net_5445), .CK(net_10092) );
INV_X2 inst_5921 ( .A(net_7445), .ZN(net_1381) );
INV_X2 inst_5770 ( .ZN(net_2985), .A(net_2984) );
OAI22_X2 inst_1573 ( .A2(net_3297), .B2(net_3286), .ZN(net_3274), .A1(net_3273), .B1(net_576) );
DFF_X1 inst_6596 ( .QN(net_7598), .D(net_5259), .CK(net_13083) );
INV_X4 inst_5521 ( .A(net_6162), .ZN(net_3597) );
CLKBUF_X2 inst_8394 ( .A(net_8355), .Z(net_8356) );
OR2_X4 inst_1390 ( .A2(net_7764), .ZN(net_2899), .A1(net_278) );
CLKBUF_X2 inst_9274 ( .A(net_8640), .Z(net_9236) );
NAND2_X2 inst_3586 ( .ZN(net_2416), .A2(net_1896), .A1(net_1429) );
CLKBUF_X2 inst_13652 ( .A(net_11178), .Z(net_13614) );
SDFF_X2 inst_229 ( .Q(net_6325), .SI(net_6324), .D(net_3635), .SE(net_392), .CK(net_14021) );
CLKBUF_X2 inst_9124 ( .A(net_9085), .Z(net_9086) );
AOI21_X2 inst_7744 ( .B1(net_7147), .ZN(net_4068), .B2(net_2582), .A(net_2335) );
CLKBUF_X2 inst_9974 ( .A(net_9935), .Z(net_9936) );
NOR2_X4 inst_2282 ( .ZN(net_5892), .A2(net_5874), .A1(net_3028) );
CLKBUF_X2 inst_12920 ( .A(net_8220), .Z(net_12882) );
CLKBUF_X2 inst_9596 ( .A(net_9557), .Z(net_9558) );
INV_X4 inst_4992 ( .ZN(net_2382), .A(net_681) );
INV_X4 inst_4689 ( .ZN(net_4151), .A(net_3333) );
CLKBUF_X2 inst_11719 ( .A(net_8276), .Z(net_11681) );
INV_X1 inst_6151 ( .ZN(net_3029), .A(net_3028) );
CLKBUF_X2 inst_9187 ( .A(net_9148), .Z(net_9149) );
OAI21_X2 inst_2131 ( .ZN(net_2904), .A(net_2903), .B2(net_2897), .B1(net_909) );
INV_X2 inst_5718 ( .ZN(net_4248), .A(net_4117) );
CLKBUF_X2 inst_12007 ( .A(net_10895), .Z(net_11969) );
CLKBUF_X2 inst_9949 ( .A(net_9910), .Z(net_9911) );
AOI22_X2 inst_7297 ( .B1(net_6547), .A1(net_6515), .A2(net_5184), .B2(net_5183), .ZN(net_5172) );
CLKBUF_X2 inst_8804 ( .A(net_8765), .Z(net_8766) );
SDFF_X2 inst_169 ( .Q(net_6245), .SI(net_6244), .D(net_3621), .SE(net_392), .CK(net_13982) );
CLKBUF_X2 inst_9453 ( .A(net_9414), .Z(net_9415) );
INV_X1 inst_6158 ( .A(net_5856), .ZN(x114) );
SDFF_X2 inst_421 ( .D(net_6391), .SE(net_5801), .SI(net_336), .Q(net_336), .CK(net_14309) );
CLKBUF_X2 inst_12880 ( .A(net_12841), .Z(net_12842) );
CLKBUF_X2 inst_11263 ( .A(net_11224), .Z(net_11225) );
CLKBUF_X2 inst_11748 ( .A(net_11709), .Z(net_11710) );
CLKBUF_X2 inst_8014 ( .A(net_7888), .Z(net_7976) );
SDFF_X2 inst_555 ( .Q(net_6442), .D(net_6442), .SI(net_3897), .SE(net_3820), .CK(net_8890) );
DFFR_X2 inst_7016 ( .D(net_3298), .QN(net_290), .CK(net_12423), .RN(x1822) );
SDFF_X2 inst_816 ( .Q(net_6991), .D(net_6991), .SE(net_3891), .SI(net_3794), .CK(net_8420) );
CLKBUF_X2 inst_11000 ( .A(net_9376), .Z(net_10962) );
CLKBUF_X2 inst_12911 ( .A(net_12872), .Z(net_12873) );
CLKBUF_X2 inst_10293 ( .A(net_9816), .Z(net_10255) );
CLKBUF_X2 inst_12978 ( .A(net_12939), .Z(net_12940) );
NAND3_X2 inst_2798 ( .ZN(net_2302), .A3(net_1543), .A1(net_1462), .A2(net_949) );
SDFF_X2 inst_1184 ( .SI(net_6928), .Q(net_6928), .D(net_3892), .SE(net_3741), .CK(net_8908) );
CLKBUF_X2 inst_12903 ( .A(net_11624), .Z(net_12865) );
CLKBUF_X2 inst_12692 ( .A(net_12653), .Z(net_12654) );
CLKBUF_X2 inst_9352 ( .A(net_9313), .Z(net_9314) );
INV_X4 inst_4685 ( .ZN(net_3738), .A(net_3366) );
CLKBUF_X2 inst_14325 ( .A(net_14286), .Z(net_14287) );
CLKBUF_X2 inst_13694 ( .A(net_13655), .Z(net_13656) );
INV_X1 inst_6157 ( .A(net_5854), .ZN(x101) );
AOI222_X2 inst_7596 ( .A1(net_7248), .ZN(net_5355), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_342), .C2(net_340) );
CLKBUF_X2 inst_12523 ( .A(net_12484), .Z(net_12485) );
CLKBUF_X2 inst_8197 ( .A(net_8158), .Z(net_8159) );
AND3_X4 inst_7796 ( .ZN(net_2589), .A1(net_2414), .A3(net_2227), .A2(net_1711) );
SDFF_X2 inst_1108 ( .SI(net_6525), .Q(net_6525), .D(net_3798), .SE(net_3756), .CK(net_11628) );
DFF_X1 inst_6580 ( .QN(net_7626), .D(net_5238), .CK(net_10591) );
CLKBUF_X2 inst_11863 ( .A(net_11824), .Z(net_11825) );
CLKBUF_X2 inst_9480 ( .A(net_9441), .Z(net_9442) );
INV_X4 inst_5148 ( .ZN(net_703), .A(net_568) );
INV_X4 inst_5140 ( .A(net_871), .ZN(net_684) );
CLKBUF_X2 inst_11578 ( .A(net_7901), .Z(net_11540) );
CLKBUF_X2 inst_8756 ( .A(net_8717), .Z(net_8718) );
CLKBUF_X2 inst_12273 ( .A(net_12234), .Z(net_12235) );
INV_X8 inst_4534 ( .ZN(net_5843), .A(net_392) );
CLKBUF_X2 inst_8952 ( .A(net_8913), .Z(net_8914) );
AOI222_X2 inst_7521 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2006), .A1(net_2005), .B1(net_2004), .C1(net_2003) );
CLKBUF_X2 inst_12931 ( .A(net_12892), .Z(net_12893) );
NAND2_X2 inst_3991 ( .ZN(net_1921), .A2(net_1042), .A1(net_484) );
CLKBUF_X2 inst_8286 ( .A(net_8247), .Z(net_8248) );
CLKBUF_X2 inst_13620 ( .A(net_8144), .Z(net_13582) );
CLKBUF_X2 inst_9546 ( .A(net_9412), .Z(net_9508) );
CLKBUF_X2 inst_11422 ( .A(net_11383), .Z(net_11384) );
CLKBUF_X2 inst_8604 ( .A(net_8565), .Z(net_8566) );
DFF_X2 inst_6203 ( .QN(net_7092), .D(net_4395), .CK(net_9369) );
CLKBUF_X2 inst_8617 ( .A(net_8578), .Z(net_8579) );
NAND2_X2 inst_3343 ( .ZN(net_3561), .A1(net_3560), .A2(net_3225) );
CLKBUF_X2 inst_9718 ( .A(net_9679), .Z(net_9680) );
NAND2_X2 inst_4140 ( .A2(net_1228), .ZN(net_1094), .A1(net_384) );
CLKBUF_X2 inst_13340 ( .A(net_13301), .Z(net_13302) );
OAI22_X2 inst_1543 ( .B1(net_4637), .B2(net_4416), .A1(net_4030), .A2(net_4028), .ZN(net_4010) );
CLKBUF_X2 inst_13892 ( .A(net_13853), .Z(net_13854) );
AOI22_X2 inst_7290 ( .B1(net_7215), .A1(net_7183), .A2(net_5244), .B2(net_5243), .ZN(net_5211) );
NAND2_X1 inst_4219 ( .ZN(net_4741), .A2(net_3988), .A1(net_2119) );
NAND3_X2 inst_2801 ( .ZN(net_2297), .A3(net_1554), .A1(net_1370), .A2(net_985) );
SDFF_X2 inst_1118 ( .SI(net_6666), .Q(net_6666), .D(net_3813), .SE(net_3465), .CK(net_9325) );
CLKBUF_X2 inst_9153 ( .A(net_9114), .Z(net_9115) );
NOR2_X2 inst_2303 ( .A2(net_6219), .A1(net_5843), .ZN(net_5838) );
CLKBUF_X2 inst_13714 ( .A(net_8025), .Z(net_13676) );
DFFR_X2 inst_6978 ( .QN(net_7785), .D(net_3990), .CK(net_13025), .RN(x1822) );
INV_X2 inst_6109 ( .A(net_7434), .ZN(net_1421) );
CLKBUF_X2 inst_8090 ( .A(net_7951), .Z(net_8052) );
CLKBUF_X2 inst_10948 ( .A(net_10909), .Z(net_10910) );
SDFF_X2 inst_473 ( .Q(net_7149), .D(net_7149), .SE(net_3903), .SI(net_3897), .CK(net_7926) );
CLKBUF_X2 inst_10140 ( .A(net_8777), .Z(net_10102) );
NOR3_X2 inst_2211 ( .ZN(net_2276), .A3(net_2275), .A2(net_1920), .A1(net_1836) );
NAND2_X2 inst_3771 ( .A1(net_7170), .A2(net_1637), .ZN(net_1574) );
NAND2_X2 inst_3083 ( .A1(net_6449), .A2(net_4925), .ZN(net_4920) );
CLKBUF_X2 inst_9170 ( .A(net_9131), .Z(net_9132) );
OAI21_X2 inst_1695 ( .B2(net_5907), .ZN(net_5599), .A(net_5287), .B1(net_4105) );
INV_X4 inst_5557 ( .A(net_7258), .ZN(net_1993) );
CLKBUF_X2 inst_12609 ( .A(net_12570), .Z(net_12571) );
CLKBUF_X2 inst_8954 ( .A(net_8915), .Z(net_8916) );
CLKBUF_X2 inst_9917 ( .A(net_9059), .Z(net_9879) );
CLKBUF_X2 inst_12942 ( .A(net_12903), .Z(net_12904) );
CLKBUF_X2 inst_9724 ( .A(net_9685), .Z(net_9686) );
CLKBUF_X2 inst_11034 ( .A(net_10995), .Z(net_10996) );
OR2_X2 inst_1404 ( .ZN(net_3066), .A2(net_3065), .A1(net_2876) );
NAND2_X2 inst_2989 ( .A1(net_6754), .A2(net_5033), .ZN(net_5022) );
INV_X2 inst_5880 ( .A(net_6023), .ZN(net_412) );
NAND2_X2 inst_3479 ( .ZN(net_2683), .A1(net_2682), .A2(net_2681) );
SDFFR_X2 inst_1339 ( .Q(net_7714), .D(net_7714), .SI(net_3782), .SE(net_3405), .CK(net_10717), .RN(x1822) );
CLKBUF_X2 inst_11235 ( .A(net_11196), .Z(net_11197) );
NAND2_X1 inst_4284 ( .ZN(net_4583), .A2(net_3867), .A1(net_1862) );
INV_X4 inst_4971 ( .ZN(net_695), .A(net_694) );
INV_X4 inst_4704 ( .ZN(net_3321), .A(net_3240) );
INV_X4 inst_4724 ( .A(net_5963), .ZN(net_3051) );
CLKBUF_X2 inst_13512 ( .A(net_11376), .Z(net_13474) );
INV_X8 inst_4467 ( .ZN(net_5138), .A(net_4284) );
NAND2_X2 inst_3575 ( .ZN(net_2492), .A2(net_2012), .A1(net_1797) );
CLKBUF_X2 inst_9238 ( .A(net_8012), .Z(net_9200) );
INV_X8 inst_4493 ( .ZN(net_3823), .A(net_3155) );
NAND2_X2 inst_3654 ( .A1(net_7065), .ZN(net_1809), .A2(net_791) );
SDFF_X2 inst_977 ( .Q(net_6429), .D(net_6429), .SE(net_3820), .SI(net_3798), .CK(net_11668) );
CLKBUF_X2 inst_8484 ( .A(net_8445), .Z(net_8446) );
CLKBUF_X2 inst_10180 ( .A(net_10141), .Z(net_10142) );
AOI22_X2 inst_7251 ( .B1(net_6819), .A1(net_6787), .A2(net_5316), .B2(net_5315), .ZN(net_5309) );
DFF_X1 inst_6901 ( .D(net_2527), .Q(net_182), .CK(net_9940) );
INV_X4 inst_5669 ( .A(net_7681), .ZN(net_522) );
INV_X4 inst_4802 ( .ZN(net_5097), .A(net_1190) );
CLKBUF_X2 inst_10941 ( .A(net_10902), .Z(net_10903) );
SDFF_X2 inst_297 ( .D(net_6394), .SE(net_5801), .SI(net_339), .Q(net_339), .CK(net_14317) );
OR2_X4 inst_1395 ( .A2(net_7530), .ZN(net_790), .A1(net_705) );
NOR2_X2 inst_2477 ( .A2(net_5778), .ZN(net_2603), .A1(net_542) );
CLKBUF_X2 inst_13933 ( .A(net_13192), .Z(net_13895) );
CLKBUF_X2 inst_13145 ( .A(net_13106), .Z(net_13107) );
CLKBUF_X2 inst_11728 ( .A(net_11689), .Z(net_11690) );
INV_X4 inst_5460 ( .A(net_7272), .ZN(net_2033) );
CLKBUF_X2 inst_11424 ( .A(net_11385), .Z(net_11386) );
CLKBUF_X2 inst_8322 ( .A(net_8283), .Z(net_8284) );
INV_X4 inst_4838 ( .A(net_2853), .ZN(net_1072) );
NOR3_X2 inst_2188 ( .ZN(net_5948), .A2(net_3954), .A3(net_3882), .A1(net_3768) );
NAND2_X2 inst_3436 ( .ZN(net_3212), .A2(net_3094), .A1(net_2761) );
OAI21_X2 inst_1875 ( .ZN(net_5228), .B1(net_5227), .A(net_4587), .B2(net_3867) );
NAND2_X2 inst_3351 ( .ZN(net_3545), .A1(net_3544), .A2(net_3226) );
CLKBUF_X2 inst_13057 ( .A(net_11197), .Z(net_13019) );
CLKBUF_X2 inst_10466 ( .A(net_10427), .Z(net_10428) );
CLKBUF_X2 inst_10005 ( .A(net_9966), .Z(net_9967) );
NAND2_X2 inst_3190 ( .ZN(net_4738), .A2(net_3988), .A1(net_2105) );
SDFF_X2 inst_162 ( .Q(net_6252), .SI(net_6251), .D(net_3550), .SE(net_392), .CK(net_13988) );
CLKBUF_X2 inst_8459 ( .A(net_7882), .Z(net_8421) );
NAND2_X2 inst_3308 ( .ZN(net_3630), .A1(net_3629), .A2(net_3229) );
CLKBUF_X2 inst_10873 ( .A(net_10834), .Z(net_10835) );
NAND2_X2 inst_3397 ( .ZN(net_3713), .A2(net_3325), .A1(net_3235) );
AOI22_X2 inst_7373 ( .A2(net_5916), .B2(net_2957), .ZN(net_2948), .B1(net_2676), .A1(net_848) );
CLKBUF_X2 inst_13286 ( .A(net_10803), .Z(net_13248) );
AOI22_X2 inst_7302 ( .B1(net_6540), .A1(net_6508), .A2(net_5184), .B2(net_5183), .ZN(net_5149) );
INV_X4 inst_5484 ( .A(net_5848), .ZN(net_4257) );
CLKBUF_X2 inst_13387 ( .A(net_11378), .Z(net_13349) );
CLKBUF_X2 inst_11544 ( .A(net_11505), .Z(net_11506) );
NAND2_X1 inst_4421 ( .A2(net_2131), .ZN(net_1514), .A1(net_1513) );
NAND3_X2 inst_2829 ( .A2(net_3852), .ZN(net_1212), .A3(net_1211), .A1(net_656) );
NAND2_X2 inst_3819 ( .A1(net_6624), .A2(net_1624), .ZN(net_1526) );
CLKBUF_X2 inst_11383 ( .A(net_11344), .Z(net_11345) );
CLKBUF_X2 inst_8448 ( .A(net_7892), .Z(net_8410) );
NAND2_X1 inst_4233 ( .ZN(net_4694), .A2(net_3989), .A1(net_2169) );
NAND2_X2 inst_3668 ( .A1(net_7343), .A2(net_1798), .ZN(net_1791) );
DFFR_X1 inst_7128 ( .D(net_3370), .Q(net_286), .CK(net_12349), .RN(x1822) );
INV_X2 inst_5905 ( .A(net_7497), .ZN(net_2172) );
NAND2_X2 inst_3968 ( .A1(net_6576), .A2(net_1705), .ZN(net_1312) );
CLKBUF_X2 inst_8208 ( .A(net_8031), .Z(net_8170) );
CLKBUF_X2 inst_13010 ( .A(net_10874), .Z(net_12972) );
CLKBUF_X2 inst_12086 ( .A(net_12047), .Z(net_12048) );
INV_X4 inst_4633 ( .ZN(net_4189), .A(net_4038) );
CLKBUF_X2 inst_8143 ( .A(net_8016), .Z(net_8105) );
SDFF_X2 inst_1098 ( .D(net_7802), .SI(net_6799), .Q(net_6799), .SE(net_3729), .CK(net_11080) );
DFFR_X2 inst_7077 ( .QN(net_6419), .D(net_2849), .CK(net_10240), .RN(x1822) );
NAND2_X2 inst_4149 ( .A2(net_1228), .ZN(net_1075), .A1(net_377) );
CLKBUF_X2 inst_8113 ( .A(net_8074), .Z(net_8075) );
CLKBUF_X2 inst_10051 ( .A(net_8951), .Z(net_10013) );
NOR2_X2 inst_2443 ( .A2(net_5963), .ZN(net_3158), .A1(net_3001) );
DFF_X1 inst_6660 ( .QN(net_7652), .D(net_5180), .CK(net_13146) );
CLKBUF_X2 inst_10915 ( .A(net_10876), .Z(net_10877) );
CLKBUF_X2 inst_8027 ( .A(net_7882), .Z(net_7989) );
DFF_X1 inst_6411 ( .QN(net_6158), .D(net_5759), .CK(net_8252) );
SDFF_X2 inst_723 ( .Q(net_6829), .D(net_6829), .SE(net_3893), .SI(net_3797), .CK(net_8953) );
CLKBUF_X2 inst_10990 ( .A(net_10951), .Z(net_10952) );
CLKBUF_X2 inst_9525 ( .A(net_9486), .Z(net_9487) );
CLKBUF_X2 inst_8921 ( .A(net_8882), .Z(net_8883) );
CLKBUF_X2 inst_8769 ( .A(net_8730), .Z(net_8731) );
SDFF_X2 inst_618 ( .Q(net_6595), .D(net_6595), .SE(net_3830), .SI(net_3799), .CK(net_12906) );
NOR2_X2 inst_2444 ( .A2(net_5983), .ZN(net_3169), .A1(net_3000) );
CLKBUF_X2 inst_11980 ( .A(net_11941), .Z(net_11942) );
NAND2_X2 inst_3893 ( .A1(net_6440), .A2(net_1677), .ZN(net_1423) );
CLKBUF_X2 inst_11616 ( .A(net_11577), .Z(net_11578) );
CLKBUF_X2 inst_11055 ( .A(net_11016), .Z(net_11017) );
NAND2_X2 inst_3057 ( .A1(net_7123), .A2(net_4950), .ZN(net_4948) );
CLKBUF_X2 inst_13274 ( .A(net_10246), .Z(net_13236) );
INV_X2 inst_5777 ( .ZN(net_2897), .A(net_229) );
NOR2_X2 inst_2462 ( .ZN(net_2737), .A1(net_2735), .A2(net_2729) );
DFF_X1 inst_6706 ( .QN(net_7290), .D(net_5368), .CK(net_10162) );
SDFF_X2 inst_474 ( .Q(net_6850), .D(net_6850), .SI(net_3900), .SE(net_3893), .CK(net_10937) );
CLKBUF_X2 inst_7894 ( .A(net_7855), .Z(net_7856) );
OAI21_X2 inst_2067 ( .B2(net_4436), .ZN(net_4428), .B1(net_4047), .A(net_3539) );
INV_X4 inst_5561 ( .A(net_7427), .ZN(net_2138) );
SDFF_X2 inst_626 ( .SI(net_6636), .Q(net_6636), .SE(net_3850), .D(net_3811), .CK(net_9335) );
CLKBUF_X2 inst_13075 ( .A(net_7942), .Z(net_13037) );
CLKBUF_X2 inst_8268 ( .A(net_8229), .Z(net_8230) );
CLKBUF_X2 inst_11539 ( .A(net_11500), .Z(net_11501) );
CLKBUF_X2 inst_9879 ( .A(net_9840), .Z(net_9841) );
AOI222_X2 inst_7476 ( .C1(net_7520), .B1(net_7488), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2153), .A1(net_2152) );
NAND3_X2 inst_2777 ( .ZN(net_2323), .A3(net_1546), .A1(net_1504), .A2(net_960) );
CLKBUF_X2 inst_12283 ( .A(net_12211), .Z(net_12245) );
DFF_X1 inst_6830 ( .D(net_2587), .QN(net_188), .CK(net_12302) );
DFF_X1 inst_6784 ( .QN(net_6065), .D(net_4319), .CK(net_8102) );
CLKBUF_X2 inst_10247 ( .A(net_9544), .Z(net_10209) );
NOR2_X2 inst_2446 ( .A2(net_5920), .ZN(net_3057), .A1(net_508) );
CLKBUF_X2 inst_13602 ( .A(net_13563), .Z(net_13564) );
INV_X4 inst_5046 ( .A(net_2885), .ZN(net_776) );
CLKBUF_X2 inst_8880 ( .A(net_8841), .Z(net_8842) );
CLKBUF_X2 inst_8452 ( .A(net_8305), .Z(net_8414) );
AND2_X4 inst_7840 ( .ZN(net_1386), .A2(net_795), .A1(net_646) );
CLKBUF_X2 inst_14128 ( .A(net_10867), .Z(net_14090) );
CLKBUF_X2 inst_11457 ( .A(net_8384), .Z(net_11419) );
CLKBUF_X2 inst_13070 ( .A(net_10583), .Z(net_13032) );
CLKBUF_X2 inst_12641 ( .A(net_12602), .Z(net_12603) );
SDFF_X2 inst_798 ( .D(net_7799), .SI(net_6899), .Q(net_6899), .SE(net_3887), .CK(net_11790) );
CLKBUF_X2 inst_14260 ( .A(net_14221), .Z(net_14222) );
CLKBUF_X2 inst_12648 ( .A(net_9168), .Z(net_12610) );
INV_X4 inst_5210 ( .ZN(net_1726), .A(net_892) );
DFF_X1 inst_6613 ( .QN(net_7574), .D(net_5394), .CK(net_8037) );
NAND2_X1 inst_4340 ( .ZN(net_4387), .A2(net_3856), .A1(net_1781) );
CLKBUF_X2 inst_12767 ( .A(net_12728), .Z(net_12729) );
OAI22_X2 inst_1434 ( .B1(net_5855), .ZN(net_5795), .A2(net_5786), .B2(net_5785), .A1(net_5771) );
CLKBUF_X2 inst_12727 ( .A(net_12688), .Z(net_12689) );
INV_X4 inst_5464 ( .A(net_6076), .ZN(net_3550) );
OAI21_X2 inst_1886 ( .B1(net_5240), .ZN(net_5195), .A(net_4571), .B2(net_3866) );
CLKBUF_X2 inst_14089 ( .A(net_14050), .Z(net_14051) );
CLKBUF_X2 inst_10211 ( .A(net_9578), .Z(net_10173) );
CLKBUF_X2 inst_12889 ( .A(net_12521), .Z(net_12851) );
CLKBUF_X2 inst_8831 ( .A(net_8792), .Z(net_8793) );
CLKBUF_X2 inst_8778 ( .A(net_8739), .Z(net_8740) );
NAND2_X1 inst_4349 ( .ZN(net_4378), .A2(net_3856), .A1(net_1761) );
OAI22_X2 inst_1457 ( .B2(net_5900), .B1(net_4644), .ZN(net_4611), .A2(net_4610), .A1(net_4045) );
CLKBUF_X2 inst_8366 ( .A(net_8327), .Z(net_8328) );
CLKBUF_X2 inst_8627 ( .A(net_8588), .Z(net_8589) );
DFFR_X2 inst_7110 ( .D(net_1953), .QN(net_123), .CK(net_9578), .RN(x1822) );
OAI21_X2 inst_1818 ( .ZN(net_5370), .B1(net_5341), .A(net_4337), .B2(net_3859) );
CLKBUF_X2 inst_10552 ( .A(net_10513), .Z(net_10514) );
CLKBUF_X2 inst_10705 ( .A(net_10666), .Z(net_10667) );
CLKBUF_X2 inst_13244 ( .A(net_12928), .Z(net_13206) );
CLKBUF_X2 inst_10264 ( .A(net_10225), .Z(net_10226) );
CLKBUF_X2 inst_8209 ( .A(net_8170), .Z(net_8171) );
CLKBUF_X2 inst_11254 ( .A(net_11215), .Z(net_11216) );
NAND2_X2 inst_3662 ( .A1(net_7338), .ZN(net_1801), .A2(net_1798) );
OAI21_X2 inst_1766 ( .B1(net_5545), .ZN(net_5428), .A(net_4643), .B2(net_3993) );
NAND3_X2 inst_2670 ( .ZN(net_3957), .A2(net_3873), .A3(net_3735), .A1(net_2238) );
CLKBUF_X2 inst_13888 ( .A(net_13849), .Z(net_13850) );
CLKBUF_X2 inst_10983 ( .A(net_10944), .Z(net_10945) );
CLKBUF_X2 inst_8380 ( .A(net_8341), .Z(net_8342) );
CLKBUF_X2 inst_8216 ( .A(net_7945), .Z(net_8178) );
NAND2_X2 inst_2974 ( .ZN(net_5493), .A2(net_5253), .A1(net_398) );
OAI21_X2 inst_1895 ( .B1(net_5208), .ZN(net_5182), .A(net_4558), .B2(net_3866) );
CLKBUF_X2 inst_9639 ( .A(net_9600), .Z(net_9601) );
CLKBUF_X2 inst_8476 ( .A(net_8437), .Z(net_8438) );
NAND3_X2 inst_2730 ( .ZN(net_2371), .A3(net_1580), .A1(net_1480), .A2(net_997) );
INV_X8 inst_4548 ( .ZN(net_2204), .A(net_706) );
SDFF_X2 inst_737 ( .Q(net_6855), .D(net_6855), .SE(net_3893), .SI(net_3790), .CK(net_8148) );
CLKBUF_X2 inst_11725 ( .A(net_11686), .Z(net_11687) );
SDFF_X2 inst_876 ( .D(net_7799), .SI(net_7034), .Q(net_7034), .SE(net_3818), .CK(net_11932) );
CLKBUF_X2 inst_11178 ( .A(net_11139), .Z(net_11140) );
NAND2_X2 inst_2979 ( .A1(net_6749), .ZN(net_5034), .A2(net_5033) );
CLKBUF_X2 inst_8990 ( .A(net_8951), .Z(net_8952) );
INV_X4 inst_4727 ( .A(net_5975), .ZN(net_3043) );
SDFF_X2 inst_545 ( .Q(net_7239), .D(net_7239), .SE(net_3822), .SI(net_335), .CK(net_12674) );
CLKBUF_X2 inst_8373 ( .A(net_8334), .Z(net_8335) );
CLKBUF_X2 inst_10189 ( .A(net_8768), .Z(net_10151) );
CLKBUF_X2 inst_8132 ( .A(net_8024), .Z(net_8094) );
NOR2_X2 inst_2433 ( .A1(net_3128), .ZN(net_3069), .A2(net_3068) );
DFF_X1 inst_6854 ( .D(net_2541), .Q(net_223), .CK(net_12541) );
CLKBUF_X2 inst_11665 ( .A(net_11626), .Z(net_11627) );
CLKBUF_X2 inst_12188 ( .A(net_10697), .Z(net_12150) );
CLKBUF_X2 inst_11751 ( .A(net_11712), .Z(net_11713) );
DFF_X1 inst_6682 ( .QN(net_7270), .D(net_5122), .CK(net_9888) );
CLKBUF_X2 inst_13595 ( .A(net_12978), .Z(net_13557) );
CLKBUF_X2 inst_9845 ( .A(net_9806), .Z(net_9807) );
SDFF_X2 inst_562 ( .SI(net_7184), .Q(net_7184), .D(net_3836), .SE(net_3817), .CK(net_11591) );
NOR2_X2 inst_2480 ( .A2(net_5778), .ZN(net_2663), .A1(net_2601) );
AND2_X4 inst_7832 ( .ZN(net_3012), .A2(net_2814), .A1(net_2243) );
CLKBUF_X2 inst_8917 ( .A(net_8656), .Z(net_8879) );
CLKBUF_X2 inst_8624 ( .A(net_8585), .Z(net_8586) );
INV_X2 inst_5878 ( .A(net_7327), .ZN(net_1757) );
CLKBUF_X2 inst_14383 ( .A(net_12466), .Z(net_14345) );
CLKBUF_X2 inst_11445 ( .A(net_11406), .Z(net_11407) );
DFF_X1 inst_6385 ( .QN(net_6116), .D(net_5703), .CK(net_11206) );
AOI221_X2 inst_7615 ( .C2(net_3105), .B1(net_2970), .ZN(net_2964), .A(net_2787), .C1(net_650), .B2(net_247) );
CLKBUF_X2 inst_8910 ( .A(net_8871), .Z(net_8872) );
CLKBUF_X2 inst_8277 ( .A(net_8153), .Z(net_8239) );
INV_X4 inst_4953 ( .ZN(net_731), .A(net_730) );
CLKBUF_X2 inst_12404 ( .A(net_12365), .Z(net_12366) );
CLKBUF_X2 inst_9589 ( .A(net_9550), .Z(net_9551) );
CLKBUF_X2 inst_13356 ( .A(net_13317), .Z(net_13318) );
NAND2_X2 inst_3659 ( .A1(net_7077), .ZN(net_1804), .A2(net_791) );
AOI222_X2 inst_7465 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2191), .A1(net_2190), .B1(net_2189), .C1(net_2188) );
DFF_X1 inst_6573 ( .QN(net_7563), .D(net_5081), .CK(net_10594) );
NAND2_X2 inst_3604 ( .ZN(net_2396), .A2(net_1892), .A1(net_1451) );
CLKBUF_X2 inst_13067 ( .A(net_13028), .Z(net_13029) );
CLKBUF_X2 inst_12347 ( .A(net_12308), .Z(net_12309) );
DFF_X1 inst_6487 ( .QN(net_7418), .D(net_5565), .CK(net_9686) );
SDFF_X2 inst_1109 ( .SI(net_6685), .Q(net_6685), .D(net_3801), .SE(net_3471), .CK(net_9083) );
CLKBUF_X2 inst_12054 ( .A(net_12015), .Z(net_12016) );
CLKBUF_X2 inst_10559 ( .A(net_10520), .Z(net_10521) );
CLKBUF_X2 inst_13879 ( .A(net_13840), .Z(net_13841) );
NAND2_X1 inst_4415 ( .A2(net_5970), .A1(net_5969), .ZN(net_2877) );
NAND2_X2 inst_4209 ( .A2(net_5987), .A1(net_5986), .ZN(net_3232) );
NAND2_X2 inst_3037 ( .A1(net_7023), .A2(net_4979), .ZN(net_4970) );
CLKBUF_X2 inst_10266 ( .A(net_10227), .Z(net_10228) );
DFF_X1 inst_6635 ( .QN(net_7591), .D(net_5247), .CK(net_13432) );
CLKBUF_X2 inst_10275 ( .A(net_8893), .Z(net_10237) );
CLKBUF_X2 inst_11522 ( .A(net_11483), .Z(net_11484) );
CLKBUF_X2 inst_8561 ( .A(net_7879), .Z(net_8523) );
CLKBUF_X2 inst_8972 ( .A(net_8112), .Z(net_8934) );
CLKBUF_X2 inst_7956 ( .A(net_7917), .Z(net_7918) );
SDFF_X2 inst_1314 ( .D(net_6384), .SE(net_5799), .SI(net_369), .Q(net_369), .CK(net_14296) );
CLKBUF_X2 inst_12072 ( .A(net_12033), .Z(net_12034) );
INV_X2 inst_5828 ( .ZN(net_924), .A(net_923) );
NAND2_X1 inst_4260 ( .ZN(net_4662), .A2(net_3993), .A1(net_1395) );
CLKBUF_X2 inst_10218 ( .A(net_10179), .Z(net_10180) );
INV_X4 inst_5533 ( .A(net_6099), .ZN(net_3505) );
SDFF_X2 inst_1156 ( .SI(net_6819), .Q(net_6819), .D(net_3821), .SE(net_3722), .CK(net_11379) );
CLKBUF_X2 inst_8072 ( .A(net_7853), .Z(net_8034) );
NAND2_X2 inst_3378 ( .ZN(net_3490), .A1(net_3489), .A2(net_3223) );
CLKBUF_X2 inst_11466 ( .A(net_9839), .Z(net_11428) );
INV_X2 inst_5993 ( .A(net_7300), .ZN(net_2045) );
CLKBUF_X2 inst_12512 ( .A(net_12473), .Z(net_12474) );
NAND2_X2 inst_3484 ( .ZN(net_2668), .A1(net_2667), .A2(net_2666) );
CLKBUF_X2 inst_13868 ( .A(net_13829), .Z(net_13830) );
CLKBUF_X2 inst_13676 ( .A(net_13637), .Z(net_13638) );
SDFF_X2 inst_942 ( .SI(net_7185), .Q(net_7185), .SE(net_3819), .D(net_3804), .CK(net_11560) );
CLKBUF_X2 inst_14259 ( .A(net_14220), .Z(net_14221) );
AOI21_X2 inst_7755 ( .B1(net_6472), .ZN(net_4045), .B2(net_2580), .A(net_2312) );
CLKBUF_X2 inst_12077 ( .A(net_12038), .Z(net_12039) );
CLKBUF_X2 inst_8269 ( .A(net_8230), .Z(net_8231) );
SDFF_X2 inst_1295 ( .D(net_6387), .SE(net_5799), .SI(net_372), .Q(net_372), .CK(net_13880) );
OAI21_X2 inst_1880 ( .ZN(net_5207), .B1(net_5206), .A(net_4578), .B2(net_3867) );
CLKBUF_X2 inst_13174 ( .A(net_13135), .Z(net_13136) );
AOI22_X2 inst_7457 ( .A2(net_7738), .B2(net_7737), .A1(net_7709), .B1(net_7708), .ZN(net_628) );
SDFF_X2 inst_262 ( .Q(net_6372), .SI(net_6371), .D(net_3566), .SE(net_392), .CK(net_14083) );
DFF_X1 inst_6603 ( .QN(net_7510), .D(net_5405), .CK(net_9240) );
NAND2_X2 inst_3630 ( .ZN(net_1953), .A1(net_1296), .A2(net_1118) );
CLKBUF_X2 inst_10333 ( .A(net_10294), .Z(net_10295) );
AOI22_X2 inst_7338 ( .B2(net_3439), .ZN(net_3304), .A2(net_2712), .B1(net_1226), .A1(net_149) );
INV_X4 inst_4675 ( .ZN(net_3464), .A(net_3463) );
AOI22_X2 inst_7353 ( .B2(net_3105), .ZN(net_3097), .A2(net_2712), .A1(net_1119), .B1(net_469) );
INV_X8 inst_4501 ( .ZN(net_3777), .A(net_3263) );
NAND2_X1 inst_4252 ( .ZN(net_4674), .A2(net_3988), .A1(net_2168) );
SDFF_X2 inst_1035 ( .Q(net_7537), .D(net_7537), .SE(net_3896), .SI(net_371), .CK(net_9388) );
CLKBUF_X2 inst_7942 ( .A(net_7903), .Z(net_7904) );
CLKBUF_X2 inst_11758 ( .A(net_11719), .Z(net_11720) );
NAND2_X2 inst_3637 ( .ZN(net_1946), .A1(net_1283), .A2(net_1114) );
CLKBUF_X2 inst_11490 ( .A(net_9541), .Z(net_11452) );
DFF_X1 inst_6356 ( .QN(net_6202), .D(net_5828), .CK(net_14284) );
OAI21_X2 inst_1883 ( .ZN(net_5201), .B1(net_5200), .A(net_4575), .B2(net_3867) );
CLKBUF_X2 inst_12863 ( .A(net_8912), .Z(net_12825) );
CLKBUF_X2 inst_9580 ( .A(net_8525), .Z(net_9542) );
CLKBUF_X2 inst_8258 ( .A(net_8219), .Z(net_8220) );
NAND2_X2 inst_3621 ( .ZN(net_1966), .A1(net_1965), .A2(net_1964) );
INV_X4 inst_5451 ( .A(net_7378), .ZN(net_891) );
DFF_X1 inst_6393 ( .QN(net_6112), .D(net_5695), .CK(net_11188) );
SDFF_X2 inst_864 ( .SI(net_7050), .Q(net_7050), .SE(net_3777), .D(net_3775), .CK(net_8215) );
SDFF_X2 inst_418 ( .D(net_6392), .SE(net_6051), .SI(net_309), .Q(net_309), .CK(net_13741) );
XNOR2_X2 inst_86 ( .B(net_2259), .ZN(net_1303), .A(net_1302) );
SDFF_X2 inst_949 ( .SI(net_7165), .Q(net_7165), .SE(net_3819), .D(net_3802), .CK(net_13335) );
NAND2_X2 inst_3283 ( .ZN(net_3680), .A1(net_3679), .A2(net_3231) );
NAND2_X2 inst_3961 ( .A1(net_6439), .A2(net_1677), .ZN(net_1323) );
CLKBUF_X2 inst_12580 ( .A(net_10348), .Z(net_12542) );
CLKBUF_X2 inst_13294 ( .A(net_13255), .Z(net_13256) );
CLKBUF_X2 inst_9526 ( .A(net_8603), .Z(net_9488) );
NAND2_X2 inst_3730 ( .A1(net_6765), .A2(net_1635), .ZN(net_1615) );
CLKBUF_X2 inst_10342 ( .A(net_10303), .Z(net_10304) );
NAND2_X2 inst_3598 ( .ZN(net_2402), .A2(net_1847), .A1(net_1399) );
CLKBUF_X2 inst_11851 ( .A(net_11570), .Z(net_11813) );
INV_X2 inst_5871 ( .A(net_886), .ZN(net_448) );
CLKBUF_X2 inst_10016 ( .A(net_9977), .Z(net_9978) );
CLKBUF_X2 inst_12140 ( .A(net_12101), .Z(net_12102) );
OAI21_X2 inst_1826 ( .ZN(net_5358), .B1(net_5357), .A(net_4381), .B2(net_3856) );
OAI21_X2 inst_2109 ( .ZN(net_3835), .B1(net_3834), .B2(net_3833), .A(net_3470) );
INV_X4 inst_5395 ( .A(net_6101), .ZN(net_3501) );
DFF_X2 inst_6192 ( .QN(net_7095), .D(net_5056), .CK(net_9374) );
OAI21_X2 inst_2020 ( .B2(net_4497), .ZN(net_4488), .B1(net_4487), .A(net_3638) );
NAND2_X1 inst_4361 ( .ZN(net_4366), .A2(net_3853), .A1(net_2046) );
CLKBUF_X2 inst_13957 ( .A(net_13918), .Z(net_13919) );
SDFF_X2 inst_1177 ( .SI(net_6949), .Q(net_6949), .D(net_3779), .SE(net_3734), .CK(net_11690) );
CLKBUF_X2 inst_13721 ( .A(net_13682), .Z(net_13683) );
NAND3_X2 inst_2820 ( .ZN(net_2278), .A3(net_1589), .A1(net_1490), .A2(net_940) );
NOR2_X2 inst_2548 ( .A2(net_6692), .ZN(net_1253), .A1(net_492) );
CLKBUF_X2 inst_14417 ( .A(net_14378), .Z(net_14379) );
NOR2_X2 inst_2404 ( .ZN(net_3762), .A1(net_3761), .A2(net_3760) );
CLKBUF_X2 inst_14075 ( .A(net_8737), .Z(net_14037) );
CLKBUF_X2 inst_11494 ( .A(net_11455), .Z(net_11456) );
CLKBUF_X2 inst_7994 ( .A(net_7955), .Z(net_7956) );
INV_X4 inst_5127 ( .ZN(net_687), .A(net_589) );
CLKBUF_X2 inst_8022 ( .A(net_7893), .Z(net_7984) );
OAI22_X2 inst_1578 ( .A2(net_3297), .B2(net_3286), .ZN(net_3266), .A1(net_3265), .B1(net_464) );
CLKBUF_X2 inst_12587 ( .A(net_12548), .Z(net_12549) );
CLKBUF_X2 inst_9051 ( .A(net_7873), .Z(net_9013) );
AND2_X4 inst_7849 ( .ZN(net_1665), .A2(net_861), .A1(net_681) );
OAI221_X2 inst_1666 ( .C2(net_5900), .ZN(net_4647), .B1(net_4644), .B2(net_4426), .C1(net_4057), .A(net_3535) );
AOI21_X2 inst_7662 ( .B2(net_5926), .ZN(net_3316), .A(net_3315), .B1(net_1217) );
SDFF_X2 inst_735 ( .Q(net_6852), .D(net_6852), .SE(net_3893), .SI(net_3782), .CK(net_11748) );
OAI22_X2 inst_1529 ( .B1(net_4644), .B2(net_4439), .A2(net_4061), .A1(net_4057), .ZN(net_4038) );
CLKBUF_X2 inst_9053 ( .A(net_9014), .Z(net_9015) );
CLKBUF_X2 inst_12445 ( .A(net_9528), .Z(net_12407) );
INV_X4 inst_4612 ( .ZN(net_4210), .A(net_4084) );
CLKBUF_X2 inst_10426 ( .A(net_10387), .Z(net_10388) );
CLKBUF_X2 inst_7890 ( .A(net_7851), .Z(net_7852) );
OAI221_X2 inst_1653 ( .ZN(net_4856), .B1(net_4855), .C2(net_4621), .B2(net_4598), .C1(net_4228), .A(net_3590) );
CLKBUF_X2 inst_9598 ( .A(net_9559), .Z(net_9560) );
CLKBUF_X2 inst_11398 ( .A(net_11359), .Z(net_11360) );
CLKBUF_X2 inst_13376 ( .A(net_13337), .Z(net_13338) );
CLKBUF_X2 inst_8820 ( .A(net_8435), .Z(net_8782) );
CLKBUF_X2 inst_11627 ( .A(net_11588), .Z(net_11589) );
NAND2_X2 inst_2984 ( .A1(net_6719), .A2(net_5031), .ZN(net_5027) );
SDFF_X2 inst_175 ( .Q(net_6279), .SI(net_6278), .D(net_3497), .SE(net_392), .CK(net_13930) );
NAND2_X2 inst_3258 ( .ZN(net_3859), .A2(net_3858), .A1(net_3834) );
CLKBUF_X2 inst_13002 ( .A(net_12963), .Z(net_12964) );
CLKBUF_X2 inst_11989 ( .A(net_9276), .Z(net_11951) );
CLKBUF_X2 inst_12150 ( .A(net_12111), .Z(net_12112) );
CLKBUF_X2 inst_10491 ( .A(net_8157), .Z(net_10453) );
INV_X4 inst_5010 ( .A(net_7822), .ZN(net_3821) );
CLKBUF_X2 inst_10895 ( .A(net_10856), .Z(net_10857) );
OAI21_X2 inst_1737 ( .ZN(net_5546), .B1(net_5545), .A(net_4810), .B2(net_4153) );
CLKBUF_X2 inst_8594 ( .A(net_8011), .Z(net_8556) );
OAI21_X2 inst_1805 ( .ZN(net_5385), .A(net_4711), .B2(net_3986), .B1(net_1183) );
NAND2_X2 inst_2995 ( .A1(net_6757), .A2(net_5033), .ZN(net_5016) );
NAND2_X2 inst_3563 ( .ZN(net_2504), .A2(net_2022), .A1(net_1796) );
CLKBUF_X2 inst_9675 ( .A(net_7961), .Z(net_9637) );
DFFR_X2 inst_7081 ( .QN(net_7733), .D(net_2801), .CK(net_7975), .RN(x1822) );
INV_X4 inst_5513 ( .A(net_5987), .ZN(net_3093) );
CLKBUF_X2 inst_8231 ( .A(net_8192), .Z(net_8193) );
INV_X8 inst_4541 ( .ZN(net_2579), .A(net_1281) );
CLKBUF_X2 inst_8936 ( .A(net_8895), .Z(net_8898) );
NAND3_X2 inst_2752 ( .ZN(net_2349), .A3(net_1596), .A1(net_1403), .A2(net_1044) );
CLKBUF_X2 inst_10095 ( .A(net_8057), .Z(net_10057) );
CLKBUF_X2 inst_14073 ( .A(net_14034), .Z(net_14035) );
SDFF_X2 inst_1149 ( .SI(net_6810), .Q(net_6810), .D(net_3805), .SE(net_3722), .CK(net_8346) );
CLKBUF_X2 inst_10146 ( .A(net_9187), .Z(net_10108) );
CLKBUF_X2 inst_14354 ( .A(net_14315), .Z(net_14316) );
SDFF_X2 inst_1281 ( .D(net_3813), .SE(net_3256), .SI(net_141), .Q(net_141), .CK(net_8535) );
OAI22_X2 inst_1509 ( .B1(net_4650), .ZN(net_4081), .A1(net_4080), .A2(net_4079), .B2(net_4078) );
INV_X4 inst_5640 ( .A(net_7401), .ZN(net_2174) );
NAND2_X2 inst_3088 ( .A1(net_6484), .A2(net_4927), .ZN(net_4915) );
CLKBUF_X2 inst_10386 ( .A(net_9847), .Z(net_10348) );
CLKBUF_X2 inst_9000 ( .A(net_8961), .Z(net_8962) );
CLKBUF_X2 inst_11475 ( .A(net_11436), .Z(net_11437) );
CLKBUF_X2 inst_9696 ( .A(net_9657), .Z(net_9658) );
NAND2_X2 inst_3782 ( .A1(net_6760), .A2(net_1635), .ZN(net_1563) );
INV_X4 inst_4719 ( .ZN(net_3024), .A(net_2866) );
AOI222_X2 inst_7486 ( .B1(net_7372), .C1(net_7308), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2118), .A1(net_2117) );
DFF_X1 inst_6630 ( .QN(net_7601), .D(net_5254), .CK(net_13278) );
INV_X2 inst_6003 ( .A(net_7755), .ZN(net_5872) );
NAND2_X1 inst_4353 ( .ZN(net_4374), .A2(net_3856), .A1(net_1764) );
CLKBUF_X2 inst_9285 ( .A(net_9246), .Z(net_9247) );
NAND2_X2 inst_3934 ( .A1(net_6981), .A2(net_1833), .ZN(net_1360) );
CLKBUF_X2 inst_9716 ( .A(net_9006), .Z(net_9678) );
CLKBUF_X2 inst_13302 ( .A(net_12220), .Z(net_13264) );
CLKBUF_X2 inst_12475 ( .A(net_12436), .Z(net_12437) );
CLKBUF_X2 inst_8054 ( .A(net_7987), .Z(net_8016) );
INV_X2 inst_5809 ( .A(net_1691), .ZN(net_1208) );
SDFF_X2 inst_948 ( .SI(net_7191), .Q(net_7191), .SE(net_3817), .D(net_3793), .CK(net_10629) );
SDFF_X2 inst_1140 ( .SI(net_6790), .Q(net_6790), .D(net_3797), .SE(net_3729), .CK(net_11076) );
CLKBUF_X2 inst_9251 ( .A(net_9212), .Z(net_9213) );
INV_X16 inst_6140 ( .ZN(net_1677), .A(net_780) );
OAI21_X2 inst_1800 ( .ZN(net_5390), .A(net_4717), .B2(net_3986), .B1(net_1165) );
INV_X4 inst_4773 ( .ZN(net_1722), .A(net_1721) );
CLKBUF_X2 inst_8463 ( .A(net_8424), .Z(net_8425) );
CLKBUF_X2 inst_11087 ( .A(net_10982), .Z(net_11049) );
DFF_X1 inst_6644 ( .QN(net_7633), .D(net_5221), .CK(net_13275) );
SDFF_X2 inst_448 ( .D(net_6390), .SE(net_5800), .SI(net_355), .Q(net_355), .CK(net_14145) );
INV_X2 inst_5966 ( .A(net_7470), .ZN(net_2114) );
CLKBUF_X2 inst_13493 ( .A(net_13454), .Z(net_13455) );
CLKBUF_X2 inst_11407 ( .A(net_11368), .Z(net_11369) );
CLKBUF_X2 inst_11275 ( .A(net_11236), .Z(net_11237) );
INV_X4 inst_5680 ( .A(net_7379), .ZN(net_417) );
CLKBUF_X2 inst_10253 ( .A(net_10214), .Z(net_10215) );
CLKBUF_X2 inst_8039 ( .A(net_7856), .Z(net_8001) );
INV_X2 inst_6056 ( .ZN(net_1111), .A(net_128) );
INV_X4 inst_4921 ( .A(net_3778), .ZN(net_3071) );
CLKBUF_X2 inst_14367 ( .A(net_14328), .Z(net_14329) );
CLKBUF_X2 inst_11647 ( .A(net_11608), .Z(net_11609) );
CLKBUF_X2 inst_9966 ( .A(net_8421), .Z(net_9928) );
CLKBUF_X2 inst_9374 ( .A(net_8296), .Z(net_9336) );
INV_X4 inst_5444 ( .A(net_7230), .ZN(net_833) );
INV_X2 inst_6030 ( .ZN(net_2927), .A(net_268) );
NAND2_X1 inst_4380 ( .ZN(net_4347), .A2(net_3859), .A1(net_2057) );
OAI21_X2 inst_2002 ( .B2(net_4518), .ZN(net_4511), .B1(net_4124), .A(net_3690) );
CLKBUF_X2 inst_10862 ( .A(net_9885), .Z(net_10824) );
CLKBUF_X2 inst_10053 ( .A(net_8595), .Z(net_10015) );
CLKBUF_X2 inst_13017 ( .A(net_9570), .Z(net_12979) );
CLKBUF_X2 inst_10471 ( .A(net_10432), .Z(net_10433) );
CLKBUF_X2 inst_8430 ( .A(net_8391), .Z(net_8392) );
CLKBUF_X2 inst_8212 ( .A(net_8173), .Z(net_8174) );
SDFF_X2 inst_608 ( .Q(net_6613), .D(net_6613), .SE(net_3830), .SI(net_3804), .CK(net_9170) );
SDFFR_X2 inst_1343 ( .Q(net_7711), .D(net_7711), .SI(net_3805), .SE(net_3405), .CK(net_13190), .RN(x1822) );
CLKBUF_X2 inst_9068 ( .A(net_8542), .Z(net_9030) );
CLKBUF_X2 inst_8050 ( .A(net_7864), .Z(net_8012) );
SDFF_X2 inst_834 ( .Q(net_7013), .D(net_7013), .SE(net_3899), .SI(net_3808), .CK(net_11898) );
CLKBUF_X2 inst_11183 ( .A(net_7961), .Z(net_11145) );
CLKBUF_X2 inst_8729 ( .A(net_8690), .Z(net_8691) );
AOI222_X2 inst_7536 ( .C1(net_7670), .A1(net_7638), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1892), .B1(net_1891) );
NAND2_X2 inst_2920 ( .A2(net_7774), .ZN(net_5772), .A1(net_5608) );
NAND2_X2 inst_4054 ( .A1(net_6809), .A2(net_1651), .ZN(net_998) );
AND2_X4 inst_7813 ( .ZN(net_3994), .A2(net_3339), .A1(net_633) );
DFF_X1 inst_6713 ( .QN(net_7329), .D(net_5354), .CK(net_12250) );
SDFF_X2 inst_966 ( .Q(net_6444), .D(net_6444), .SE(net_3820), .SI(net_3805), .CK(net_10853) );
CLKBUF_X2 inst_11833 ( .A(net_11794), .Z(net_11795) );
CLKBUF_X2 inst_8924 ( .A(net_8885), .Z(net_8886) );
SDFF_X2 inst_1246 ( .SI(net_6541), .Q(net_6541), .D(net_3900), .SE(net_3756), .CK(net_8046) );
NAND2_X2 inst_2961 ( .ZN(net_5466), .A1(net_4900), .A2(net_4898) );
NAND2_X2 inst_3185 ( .ZN(net_4748), .A2(net_3941), .A1(net_2216) );
INV_X4 inst_4679 ( .ZN(net_3385), .A(net_3384) );
NOR2_X2 inst_2506 ( .ZN(net_1238), .A2(net_675), .A1(net_639) );
CLKBUF_X2 inst_13214 ( .A(net_8328), .Z(net_13176) );
CLKBUF_X2 inst_11699 ( .A(net_11660), .Z(net_11661) );
CLKBUF_X2 inst_11269 ( .A(net_11230), .Z(net_11231) );
INV_X2 inst_5836 ( .ZN(net_810), .A(net_809) );
CLKBUF_X2 inst_13163 ( .A(net_8025), .Z(net_13125) );
INV_X2 inst_5976 ( .A(net_7630), .ZN(net_1852) );
INV_X4 inst_5647 ( .A(net_7705), .ZN(net_842) );
CLKBUF_X2 inst_10623 ( .A(net_10327), .Z(net_10585) );
INV_X4 inst_5245 ( .A(net_1824), .ZN(net_1232) );
INV_X4 inst_5580 ( .A(net_6409), .ZN(net_529) );
INV_X4 inst_5575 ( .A(net_6125), .ZN(net_3643) );
INV_X8 inst_4557 ( .ZN(net_2209), .A(net_778) );
CLKBUF_X2 inst_12180 ( .A(net_12141), .Z(net_12142) );
NAND2_X2 inst_3607 ( .ZN(net_2391), .A2(net_1849), .A1(net_1510) );
CLKBUF_X2 inst_8568 ( .A(net_8529), .Z(net_8530) );
OAI21_X2 inst_2029 ( .B2(net_4476), .ZN(net_4474), .B1(net_4211), .A(net_3606) );
CLKBUF_X2 inst_10632 ( .A(net_10593), .Z(net_10594) );
CLKBUF_X2 inst_12812 ( .A(net_12773), .Z(net_12774) );
CLKBUF_X2 inst_8583 ( .A(net_7904), .Z(net_8545) );
CLKBUF_X2 inst_10498 ( .A(net_10459), .Z(net_10460) );
CLKBUF_X2 inst_8779 ( .A(net_8740), .Z(net_8741) );
INV_X4 inst_4936 ( .A(net_2299), .ZN(net_757) );
CLKBUF_X2 inst_13324 ( .A(net_13285), .Z(net_13286) );
NAND2_X2 inst_3160 ( .ZN(net_4773), .A2(net_3941), .A1(net_2051) );
CLKBUF_X2 inst_14022 ( .A(net_11582), .Z(net_13984) );
NAND2_X4 inst_2861 ( .A1(net_5880), .ZN(net_5040), .A2(net_4138) );
XNOR2_X2 inst_66 ( .ZN(net_2476), .A(net_1055), .B(net_489) );
INV_X4 inst_4814 ( .ZN(net_4789), .A(net_1164) );
CLKBUF_X2 inst_11139 ( .A(net_11100), .Z(net_11101) );
CLKBUF_X2 inst_11012 ( .A(net_10973), .Z(net_10974) );
CLKBUF_X2 inst_10604 ( .A(net_10565), .Z(net_10566) );
CLKBUF_X2 inst_7920 ( .A(net_7881), .Z(net_7882) );
CLKBUF_X2 inst_8807 ( .A(net_8334), .Z(net_8769) );
CLKBUF_X2 inst_12297 ( .A(net_8422), .Z(net_12259) );
SDFF_X2 inst_273 ( .D(net_6399), .SE(net_5800), .SI(net_364), .Q(net_364), .CK(net_13683) );
CLKBUF_X2 inst_13443 ( .A(net_8068), .Z(net_13405) );
OAI21_X2 inst_1965 ( .B1(net_5410), .ZN(net_5045), .A(net_4652), .B2(net_3993) );
NAND2_X2 inst_3915 ( .A1(net_6438), .A2(net_1677), .ZN(net_1391) );
INV_X4 inst_5419 ( .A(net_7231), .ZN(net_445) );
SDFF_X2 inst_366 ( .SI(net_7636), .Q(net_7636), .D(net_4792), .SE(net_3867), .CK(net_13253) );
NOR2_X2 inst_2418 ( .A2(net_7768), .ZN(net_4258), .A1(net_3341) );
CLKBUF_X2 inst_8144 ( .A(net_8105), .Z(net_8106) );
DFFR_X2 inst_7019 ( .D(net_3284), .QN(net_294), .CK(net_10452), .RN(x1822) );
INV_X2 inst_5743 ( .ZN(net_3721), .A(net_3418) );
INV_X4 inst_5422 ( .A(net_7260), .ZN(net_2067) );
CLKBUF_X2 inst_12542 ( .A(net_12503), .Z(net_12504) );
CLKBUF_X2 inst_9565 ( .A(net_9526), .Z(net_9527) );
CLKBUF_X2 inst_9397 ( .A(net_9358), .Z(net_9359) );
CLKBUF_X2 inst_7964 ( .A(net_7925), .Z(net_7926) );
AOI22_X2 inst_7313 ( .B1(net_6686), .A1(net_6654), .A2(net_5139), .B2(net_5138), .ZN(net_5130) );
NAND2_X2 inst_3285 ( .ZN(net_3676), .A1(net_3675), .A2(net_3231) );
DFFS_X2 inst_6948 ( .QN(net_6411), .D(net_2725), .CK(net_14416), .SN(x1822) );
DFF_X1 inst_6492 ( .QN(net_7404), .D(net_5555), .CK(net_12505) );
INV_X2 inst_5896 ( .A(net_7331), .ZN(net_1778) );
INV_X4 inst_4746 ( .ZN(net_2753), .A(net_2631) );
CLKBUF_X2 inst_7950 ( .A(net_7911), .Z(net_7912) );
CLKBUF_X2 inst_14091 ( .A(net_14052), .Z(net_14053) );
SDFF_X2 inst_1025 ( .SI(net_6493), .Q(net_6493), .SE(net_3886), .D(net_3798), .CK(net_11633) );
SDFF_X2 inst_707 ( .SI(net_6778), .Q(net_6778), .SE(net_3816), .D(net_3783), .CK(net_10910) );
INV_X4 inst_4655 ( .ZN(net_5877), .A(net_4150) );
CLKBUF_X2 inst_11931 ( .A(net_8521), .Z(net_11893) );
CLKBUF_X2 inst_11790 ( .A(net_11609), .Z(net_11752) );
AOI222_X2 inst_7566 ( .A1(net_7245), .ZN(net_5361), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_339), .C2(net_337) );
NAND2_X2 inst_3670 ( .A2(net_1798), .ZN(net_1789), .A1(net_1788) );
CLKBUF_X2 inst_11568 ( .A(net_11529), .Z(net_11530) );
NAND2_X1 inst_4460 ( .A2(net_1256), .ZN(net_1110), .A1(net_1109) );
CLKBUF_X2 inst_8336 ( .A(net_8297), .Z(net_8298) );
AOI222_X2 inst_7570 ( .ZN(net_5434), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_364), .C2(net_362), .A1(net_350) );
INV_X4 inst_5635 ( .A(net_7724), .ZN(net_2664) );
CLKBUF_X2 inst_12559 ( .A(net_12520), .Z(net_12521) );
AND2_X4 inst_7834 ( .ZN(net_2990), .A1(net_2853), .A2(net_190) );
CLKBUF_X2 inst_11681 ( .A(net_11642), .Z(net_11643) );
DFFR_X2 inst_7002 ( .QN(net_7719), .D(net_3350), .CK(net_8600), .RN(x1822) );
NAND3_X2 inst_2804 ( .ZN(net_2294), .A3(net_1638), .A1(net_1493), .A2(net_957) );
INV_X4 inst_5542 ( .A(net_7533), .ZN(net_894) );
CLKBUF_X2 inst_8654 ( .A(net_8615), .Z(net_8616) );
INV_X4 inst_5131 ( .A(net_1221), .ZN(net_584) );
CLKBUF_X2 inst_10080 ( .A(net_10041), .Z(net_10042) );
CLKBUF_X2 inst_13710 ( .A(net_13671), .Z(net_13672) );
CLKBUF_X2 inst_13654 ( .A(net_13615), .Z(net_13616) );
AOI22_X2 inst_7269 ( .B1(net_7083), .A1(net_7051), .ZN(net_5281), .A2(net_5280), .B2(net_5279) );
NAND3_X2 inst_2576 ( .ZN(net_5763), .A1(net_5658), .A2(net_5282), .A3(net_4316) );
NAND3_X2 inst_2631 ( .ZN(net_5698), .A1(net_5675), .A2(net_5309), .A3(net_4249) );
SDFF_X2 inst_772 ( .SI(net_7799), .Q(net_6867), .D(net_6867), .SE(net_3901), .CK(net_11805) );
NAND2_X2 inst_3810 ( .A1(net_6636), .A2(net_1624), .ZN(net_1535) );
CLKBUF_X2 inst_8453 ( .A(net_8237), .Z(net_8415) );
DFF_X1 inst_6738 ( .QN(net_7364), .D(net_4861), .CK(net_12694) );
CLKBUF_X2 inst_13261 ( .A(net_13222), .Z(net_13223) );
NAND2_X2 inst_3682 ( .A2(net_1798), .ZN(net_1769), .A1(net_1768) );
INV_X4 inst_4940 ( .ZN(net_751), .A(net_750) );
INV_X8 inst_4523 ( .ZN(net_3747), .A(net_3115) );
DFFR_X2 inst_7073 ( .D(net_2813), .QN(net_276), .CK(net_12331), .RN(x1822) );
INV_X4 inst_4583 ( .A(net_5054), .ZN(net_4329) );
NAND3_X2 inst_2636 ( .ZN(net_5693), .A1(net_5670), .A2(net_5300), .A3(net_4244) );
CLKBUF_X2 inst_13282 ( .A(net_13243), .Z(net_13244) );
DFF_X2 inst_6198 ( .QN(net_7227), .D(net_4394), .CK(net_10518) );
CLKBUF_X2 inst_10525 ( .A(net_8999), .Z(net_10487) );
AOI222_X2 inst_7579 ( .A1(net_7549), .ZN(net_5230), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_381), .C2(net_379) );
CLKBUF_X2 inst_14396 ( .A(net_14357), .Z(net_14358) );
CLKBUF_X2 inst_11561 ( .A(net_11522), .Z(net_11523) );
INV_X4 inst_4870 ( .ZN(net_3849), .A(net_687) );
CLKBUF_X2 inst_13618 ( .A(net_13579), .Z(net_13580) );
CLKBUF_X2 inst_12961 ( .A(net_12922), .Z(net_12923) );
SDFF_X2 inst_445 ( .Q(net_7400), .D(net_7400), .SE(net_3994), .SI(net_365), .CK(net_9622) );
INV_X4 inst_5454 ( .A(net_7271), .ZN(net_2087) );
INV_X4 inst_5192 ( .A(net_858), .ZN(net_511) );
DFF_X2 inst_6224 ( .QN(net_7232), .D(net_3724), .CK(net_9366) );
CLKBUF_X2 inst_11566 ( .A(net_11527), .Z(net_11528) );
CLKBUF_X2 inst_11400 ( .A(net_11361), .Z(net_11362) );
DFF_X1 inst_6761 ( .QN(net_7347), .D(net_4859), .CK(net_12793) );
SDFF_X2 inst_606 ( .Q(net_6592), .D(net_6592), .SE(net_3830), .SI(net_3806), .CK(net_9343) );
CLKBUF_X2 inst_12350 ( .A(net_12311), .Z(net_12312) );
NAND2_X2 inst_2942 ( .ZN(net_5504), .A1(net_4968), .A2(net_4967) );
CLKBUF_X2 inst_9929 ( .A(net_9109), .Z(net_9891) );
CLKBUF_X2 inst_13875 ( .A(net_13164), .Z(net_13837) );
CLKBUF_X2 inst_10138 ( .A(net_10099), .Z(net_10100) );
INV_X4 inst_5654 ( .A(net_6058), .ZN(net_416) );
INV_X4 inst_5089 ( .A(net_3243), .ZN(net_626) );
NAND2_X2 inst_3761 ( .A1(net_6775), .A2(net_1635), .ZN(net_1584) );
INV_X2 inst_5864 ( .A(net_831), .ZN(net_580) );
SDFF_X2 inst_853 ( .SI(net_7028), .Q(net_7028), .D(net_3792), .SE(net_3777), .CK(net_9024) );
CLKBUF_X2 inst_10287 ( .A(net_10248), .Z(net_10249) );
CLKBUF_X2 inst_8167 ( .A(net_8128), .Z(net_8129) );
SDFF_X2 inst_139 ( .QN(net_6239), .SI(net_6238), .SE(net_392), .D(net_145), .CK(net_13627) );
CLKBUF_X2 inst_13767 ( .A(net_13728), .Z(net_13729) );
SDFF_X2 inst_657 ( .Q(net_6714), .D(net_6714), .SE(net_3871), .SI(net_3805), .CK(net_10932) );
CLKBUF_X2 inst_10856 ( .A(net_10817), .Z(net_10818) );
CLKBUF_X2 inst_8903 ( .A(net_8864), .Z(net_8865) );
INV_X8 inst_4550 ( .ZN(net_1833), .A(net_704) );
CLKBUF_X2 inst_12803 ( .A(net_12764), .Z(net_12765) );
CLKBUF_X2 inst_12548 ( .A(net_11597), .Z(net_12510) );
SDFF_X2 inst_1316 ( .D(net_6382), .SE(net_5799), .SI(net_367), .Q(net_367), .CK(net_14293) );
OAI21_X2 inst_2098 ( .B2(net_4405), .ZN(net_4318), .B1(net_4030), .A(net_3518) );
CLKBUF_X2 inst_12465 ( .A(net_12426), .Z(net_12427) );
CLKBUF_X2 inst_8400 ( .A(net_8361), .Z(net_8362) );
NAND2_X2 inst_3551 ( .ZN(net_2516), .A2(net_2076), .A1(net_1767) );
INV_X4 inst_5528 ( .A(net_6132), .ZN(net_3629) );
OAI21_X2 inst_1921 ( .B1(net_5341), .ZN(net_5142), .A(net_4744), .B2(net_3941) );
CLKBUF_X2 inst_13890 ( .A(net_13634), .Z(net_13852) );
CLKBUF_X2 inst_12890 ( .A(net_12851), .Z(net_12852) );
DFF_X1 inst_6521 ( .QN(net_7437), .D(net_5430), .CK(net_12114) );
DFFR_X2 inst_6977 ( .QN(net_7784), .D(net_3991), .CK(net_10245), .RN(x1822) );
NAND2_X1 inst_4293 ( .ZN(net_4574), .A2(net_3867), .A1(net_1842) );
CLKBUF_X2 inst_13996 ( .A(net_13957), .Z(net_13958) );
SDFF_X2 inst_191 ( .Q(net_6263), .SI(net_6262), .D(net_3487), .SE(net_392), .CK(net_13468) );
CLKBUF_X2 inst_14285 ( .A(net_9102), .Z(net_14247) );
CLKBUF_X2 inst_10357 ( .A(net_10318), .Z(net_10319) );
NAND3_X2 inst_2638 ( .ZN(net_5691), .A1(net_5668), .A2(net_5296), .A3(net_4242) );
CLKBUF_X2 inst_8676 ( .A(net_8301), .Z(net_8638) );
CLKBUF_X2 inst_8908 ( .A(net_8869), .Z(net_8870) );
CLKBUF_X2 inst_9328 ( .A(net_9289), .Z(net_9290) );
CLKBUF_X2 inst_13485 ( .A(net_7849), .Z(net_13447) );
INV_X8 inst_4538 ( .ZN(net_2772), .A(net_1864) );
INV_X4 inst_5212 ( .ZN(net_485), .A(net_484) );
NAND2_X2 inst_3235 ( .ZN(net_4281), .A1(net_4280), .A2(net_1639) );
CLKBUF_X2 inst_14019 ( .A(net_13980), .Z(net_13981) );
CLKBUF_X2 inst_13988 ( .A(net_11284), .Z(net_13950) );
CLKBUF_X2 inst_8672 ( .A(net_8633), .Z(net_8634) );
CLKBUF_X2 inst_12786 ( .A(net_12747), .Z(net_12748) );
CLKBUF_X2 inst_9421 ( .A(net_9382), .Z(net_9383) );
DFF_X1 inst_6892 ( .D(net_2524), .Q(net_234), .CK(net_13140) );
CLKBUF_X2 inst_8711 ( .A(net_8672), .Z(net_8673) );
NAND2_X2 inst_3879 ( .A1(net_6575), .A2(net_1705), .ZN(net_1441) );
INV_X4 inst_5269 ( .A(net_1226), .ZN(net_422) );
DFF_X1 inst_6544 ( .QN(net_7321), .D(net_5340), .CK(net_12281) );
CLKBUF_X2 inst_12201 ( .A(net_9247), .Z(net_12163) );
CLKBUF_X2 inst_8125 ( .A(net_8086), .Z(net_8087) );
NOR4_X2 inst_2184 ( .ZN(net_1206), .A4(net_1040), .A1(x1209), .A3(x1203), .A2(x1193) );
CLKBUF_X2 inst_13296 ( .A(net_13257), .Z(net_13258) );
SDFF_X2 inst_892 ( .Q(net_7123), .D(net_7123), .SE(net_3888), .SI(net_3791), .CK(net_8722) );
NAND3_X2 inst_2665 ( .ZN(net_3967), .A2(net_3878), .A3(net_3740), .A1(net_2236) );
SDFF_X2 inst_1132 ( .SI(net_6684), .Q(net_6684), .D(net_3821), .SE(net_3471), .CK(net_9066) );
CLKBUF_X2 inst_14415 ( .A(net_14088), .Z(net_14377) );
NAND2_X2 inst_4100 ( .A1(net_6931), .A2(net_1654), .ZN(net_952) );
SDFF_X2 inst_968 ( .Q(net_6447), .D(net_6447), .SE(net_3820), .SI(net_3782), .CK(net_8072) );
INV_X4 inst_4700 ( .A(net_5980), .ZN(net_3363) );
CLKBUF_X2 inst_13531 ( .A(net_13492), .Z(net_13493) );
NAND2_X1 inst_4441 ( .A2(net_2131), .ZN(net_1345), .A1(net_1344) );
DFFR_X2 inst_6987 ( .D(net_3397), .QN(net_277), .CK(net_12804), .RN(x1822) );
OAI21_X2 inst_1803 ( .ZN(net_5387), .A(net_4714), .B2(net_3986), .B1(net_1108) );
NAND2_X2 inst_3153 ( .ZN(net_4810), .A2(net_4153), .A1(net_2111) );
NAND3_X2 inst_2814 ( .ZN(net_2284), .A3(net_1528), .A1(net_1317), .A2(net_943) );
INV_X2 inst_6076 ( .A(net_7468), .ZN(net_2124) );
CLKBUF_X2 inst_9819 ( .A(net_9780), .Z(net_9781) );
SDFF_X2 inst_936 ( .SI(net_7178), .Q(net_7178), .SE(net_3817), .D(net_3787), .CK(net_7848) );
NAND2_X2 inst_3809 ( .A1(net_6507), .A2(net_1642), .ZN(net_1536) );
CLKBUF_X2 inst_14357 ( .A(net_14318), .Z(net_14319) );
CLKBUF_X2 inst_11990 ( .A(net_11951), .Z(net_11952) );
NAND2_X2 inst_4004 ( .ZN(net_1280), .A1(net_664), .A2(net_632) );
CLKBUF_X2 inst_12708 ( .A(net_8500), .Z(net_12670) );
CLKBUF_X2 inst_11368 ( .A(net_11329), .Z(net_11330) );
CLKBUF_X2 inst_11838 ( .A(net_11799), .Z(net_11800) );
CLKBUF_X2 inst_10315 ( .A(net_10276), .Z(net_10277) );
HA_X1 inst_6171 ( .B(net_7785), .S(net_890), .CO(net_889), .A(net_888) );
CLKBUF_X2 inst_8887 ( .A(net_8848), .Z(net_8849) );
CLKBUF_X2 inst_14236 ( .A(net_14197), .Z(net_14198) );
NAND2_X2 inst_3798 ( .A1(net_6902), .A2(net_1639), .ZN(net_1547) );
DFF_X1 inst_6865 ( .D(net_2539), .Q(net_206), .CK(net_12463) );
INV_X4 inst_5232 ( .A(net_514), .ZN(net_458) );
NAND2_X2 inst_4109 ( .A1(net_6673), .A2(net_1655), .ZN(net_943) );
NAND2_X2 inst_4192 ( .A1(net_7691), .A2(net_916), .ZN(net_653) );
CLKBUF_X2 inst_12948 ( .A(net_12909), .Z(net_12910) );
CLKBUF_X2 inst_10048 ( .A(net_10009), .Z(net_10010) );
NAND2_X2 inst_3004 ( .A1(net_6884), .ZN(net_5007), .A2(net_5006) );
NAND2_X2 inst_3780 ( .A1(net_6905), .A2(net_1639), .ZN(net_1565) );
CLKBUF_X2 inst_12396 ( .A(net_12357), .Z(net_12358) );
CLKBUF_X2 inst_11305 ( .A(net_11266), .Z(net_11267) );
NAND3_X2 inst_2647 ( .ZN(net_5953), .A3(net_3959), .A2(net_1400), .A1(net_777) );
INV_X4 inst_4672 ( .ZN(net_4154), .A(net_3470) );
DFF_X1 inst_6576 ( .QN(net_7630), .D(net_5228), .CK(net_13091) );
CLKBUF_X2 inst_14438 ( .A(net_10724), .Z(net_14400) );
CLKBUF_X2 inst_12363 ( .A(net_12324), .Z(net_12325) );
NOR2_X2 inst_2456 ( .ZN(net_2814), .A2(net_2691), .A1(net_1162) );
CLKBUF_X2 inst_11959 ( .A(net_11832), .Z(net_11921) );
INV_X4 inst_5629 ( .A(net_6048), .ZN(net_2607) );
NAND3_X2 inst_2710 ( .ZN(net_2467), .A2(net_1813), .A3(net_1617), .A1(net_1355) );
SDFF_X2 inst_1058 ( .SI(net_7049), .Q(net_7049), .D(net_3836), .SE(net_3818), .CK(net_9007) );
NAND2_X4 inst_2887 ( .ZN(net_4132), .A2(net_3332), .A1(net_2968) );
CLKBUF_X2 inst_12162 ( .A(net_9975), .Z(net_12124) );
CLKBUF_X2 inst_12639 ( .A(net_9378), .Z(net_12601) );
CLKBUF_X2 inst_11120 ( .A(net_11081), .Z(net_11082) );
NAND2_X2 inst_3360 ( .ZN(net_3526), .A1(net_3525), .A2(net_3225) );
DFF_X1 inst_6821 ( .QN(net_5968), .D(net_3017), .CK(net_11418) );
INV_X4 inst_4984 ( .A(net_1144), .ZN(net_875) );
CLKBUF_X2 inst_8805 ( .A(net_8766), .Z(net_8767) );
OAI22_X2 inst_1473 ( .B1(net_4855), .A1(net_4228), .ZN(net_4224), .A2(net_4223), .B2(net_4222) );
INV_X4 inst_5334 ( .A(net_6114), .ZN(net_3701) );
CLKBUF_X2 inst_12793 ( .A(net_12754), .Z(net_12755) );
CLKBUF_X2 inst_14098 ( .A(net_10441), .Z(net_14060) );
OAI21_X2 inst_1788 ( .B1(net_5436), .ZN(net_5403), .A(net_4677), .B2(net_3988) );
CLKBUF_X2 inst_9306 ( .A(net_8355), .Z(net_9268) );
SDFF_X2 inst_1272 ( .Q(net_5858), .SE(net_3066), .SI(net_3065), .D(net_604), .CK(net_7981) );
NAND2_X2 inst_4182 ( .A1(net_7093), .ZN(net_704), .A2(net_683) );
SDFF_X2 inst_632 ( .SI(net_6643), .Q(net_6643), .SE(net_3851), .D(net_3783), .CK(net_9115) );
XOR2_X2 inst_0 ( .A(net_2565), .Z(net_1254), .B(net_1253) );
NAND2_X4 inst_2852 ( .ZN(net_5471), .A1(net_4911), .A2(net_4910) );
CLKBUF_X2 inst_13934 ( .A(net_13895), .Z(net_13896) );
DFF_X1 inst_6751 ( .QN(net_7635), .D(net_4845), .CK(net_13414) );
CLKBUF_X2 inst_11405 ( .A(net_11366), .Z(net_11367) );
CLKBUF_X2 inst_11199 ( .A(net_11160), .Z(net_11161) );
NAND2_X2 inst_3973 ( .ZN(net_1297), .A1(net_885), .A2(net_315) );
CLKBUF_X2 inst_12266 ( .A(net_12227), .Z(net_12228) );
AOI222_X2 inst_7584 ( .A1(net_7241), .ZN(net_5339), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_335), .C2(net_333) );
CLKBUF_X2 inst_8994 ( .A(net_8955), .Z(net_8956) );
SDFF_X2 inst_433 ( .Q(net_7398), .D(net_7398), .SE(net_3994), .SI(net_363), .CK(net_9642) );
CLKBUF_X2 inst_13520 ( .A(net_12049), .Z(net_13482) );
OAI21_X2 inst_1983 ( .B1(net_4853), .ZN(net_4846), .A(net_4583), .B2(net_3867) );
CLKBUF_X2 inst_13771 ( .A(net_13732), .Z(net_13733) );
CLKBUF_X2 inst_13249 ( .A(net_13210), .Z(net_13211) );
CLKBUF_X2 inst_11817 ( .A(net_11778), .Z(net_11779) );
INV_X4 inst_4939 ( .ZN(net_753), .A(net_752) );
CLKBUF_X2 inst_13748 ( .A(net_11588), .Z(net_13710) );
CLKBUF_X2 inst_13772 ( .A(net_13733), .Z(net_13734) );
CLKBUF_X2 inst_11312 ( .A(net_11273), .Z(net_11274) );
DFF_X1 inst_6417 ( .QN(net_6152), .D(net_5753), .CK(net_9049) );
CLKBUF_X2 inst_8984 ( .A(net_7847), .Z(net_8946) );
AOI22_X2 inst_7323 ( .ZN(net_3433), .A2(net_3432), .B2(net_3431), .A1(net_1307), .B1(net_908) );
OAI21_X2 inst_1948 ( .B1(net_5225), .ZN(net_5072), .A(net_4729), .B2(net_3986) );
CLKBUF_X2 inst_11955 ( .A(net_11916), .Z(net_11917) );
CLKBUF_X2 inst_8409 ( .A(net_8370), .Z(net_8371) );
CLKBUF_X2 inst_8638 ( .A(net_8599), .Z(net_8600) );
CLKBUF_X2 inst_9269 ( .A(net_9230), .Z(net_9231) );
CLKBUF_X2 inst_8266 ( .A(net_8227), .Z(net_8228) );
INV_X2 inst_5781 ( .ZN(net_2450), .A(net_2449) );
CLKBUF_X2 inst_13476 ( .A(net_10846), .Z(net_13438) );
SDFF_X2 inst_422 ( .D(net_6391), .SE(net_5799), .SI(net_376), .Q(net_376), .CK(net_14212) );
NOR2_X4 inst_2243 ( .ZN(net_5643), .A1(net_5489), .A2(net_4455) );
OAI22_X2 inst_1475 ( .B1(net_4855), .A1(net_4228), .B2(net_4223), .ZN(net_4219), .A2(net_4218) );
OR2_X2 inst_1426 ( .A2(net_6419), .A1(net_6418), .ZN(net_807) );
CLKBUF_X2 inst_9021 ( .A(net_8417), .Z(net_8983) );
INV_X4 inst_4812 ( .ZN(net_5107), .A(net_1166) );
NAND2_X2 inst_3090 ( .A1(net_6485), .A2(net_4927), .ZN(net_4913) );
OAI222_X2 inst_1637 ( .ZN(net_4302), .B2(net_4301), .C2(net_4300), .A2(net_4168), .A1(net_2451), .B1(net_1653), .C1(net_583) );
SDFFR_X2 inst_1352 ( .D(net_3782), .SE(net_3297), .SI(net_296), .Q(net_296), .CK(net_13184), .RN(x1822) );
CLKBUF_X2 inst_12338 ( .A(net_12299), .Z(net_12300) );
CLKBUF_X2 inst_10012 ( .A(net_9973), .Z(net_9974) );
CLKBUF_X2 inst_8355 ( .A(net_8316), .Z(net_8317) );
NOR2_X4 inst_2261 ( .ZN(net_5625), .A1(net_5470), .A2(net_4428) );
CLKBUF_X2 inst_9955 ( .A(net_9916), .Z(net_9917) );
INV_X4 inst_4879 ( .ZN(net_1082), .A(net_632) );
INV_X4 inst_4695 ( .A(net_5960), .ZN(net_3368) );
NAND2_X2 inst_4142 ( .A1(net_1151), .ZN(net_913), .A2(net_883) );
NAND2_X2 inst_3390 ( .ZN(net_3769), .A2(net_3367), .A1(net_2891) );
CLKBUF_X2 inst_12125 ( .A(net_10039), .Z(net_12087) );
CLKBUF_X2 inst_9076 ( .A(net_8888), .Z(net_9038) );
CLKBUF_X2 inst_8513 ( .A(net_8474), .Z(net_8475) );
CLKBUF_X2 inst_11260 ( .A(net_11221), .Z(net_11222) );
CLKBUF_X2 inst_9097 ( .A(net_9058), .Z(net_9059) );
CLKBUF_X2 inst_8178 ( .A(net_8139), .Z(net_8140) );
AOI222_X1 inst_7609 ( .C1(net_5941), .B1(net_2970), .ZN(net_2874), .A1(net_2872), .B2(net_259), .C2(net_222), .A2(net_185) );
NAND2_X2 inst_2930 ( .ZN(net_5522), .A1(net_4995), .A2(net_4994) );
CLKBUF_X2 inst_12680 ( .A(net_12641), .Z(net_12642) );
INV_X4 inst_5683 ( .A(net_6173), .ZN(net_3525) );
CLKBUF_X2 inst_12206 ( .A(net_8000), .Z(net_12168) );
INV_X4 inst_4790 ( .A(net_3052), .ZN(net_1721) );
CLKBUF_X2 inst_9851 ( .A(net_9812), .Z(net_9813) );
NAND2_X1 inst_4307 ( .ZN(net_4559), .A2(net_3866), .A1(net_2147) );
NAND2_X4 inst_2859 ( .A1(net_5887), .ZN(net_5054), .A2(net_4140) );
SDFF_X2 inst_397 ( .SI(net_7338), .Q(net_7338), .D(net_4780), .SE(net_3856), .CK(net_9404) );
SDFF_X2 inst_504 ( .SI(net_7031), .Q(net_7031), .D(net_3892), .SE(net_3818), .CK(net_11966) );
CLKBUF_X2 inst_8601 ( .A(net_8562), .Z(net_8563) );
NAND2_X2 inst_3192 ( .ZN(net_4734), .A2(net_3986), .A1(net_1906) );
INV_X4 inst_5006 ( .A(net_7808), .ZN(net_3787) );
CLKBUF_X2 inst_14240 ( .A(net_14201), .Z(net_14202) );
CLKBUF_X2 inst_9026 ( .A(net_7937), .Z(net_8988) );
CLKBUF_X2 inst_9780 ( .A(net_9741), .Z(net_9742) );
SDFF_X2 inst_1297 ( .D(net_6387), .SE(net_6052), .SI(net_312), .Q(net_312), .CK(net_13805) );
NAND2_X2 inst_3194 ( .ZN(net_4732), .A2(net_3986), .A1(net_1894) );
CLKBUF_X2 inst_13585 ( .A(net_13546), .Z(net_13547) );
CLKBUF_X2 inst_11129 ( .A(net_11090), .Z(net_11091) );
NAND2_X2 inst_3884 ( .A1(net_6967), .A2(net_1833), .ZN(net_1435) );
CLKBUF_X2 inst_13831 ( .A(net_8482), .Z(net_13793) );
CLKBUF_X2 inst_9146 ( .A(net_9107), .Z(net_9108) );
DFF_X2 inst_6296 ( .QN(net_5981), .D(net_1658), .CK(net_12526) );
NAND2_X1 inst_4246 ( .ZN(net_4681), .A2(net_3988), .A1(net_2201) );
SDFF_X2 inst_1173 ( .SI(net_6926), .Q(net_6926), .D(net_3806), .SE(net_3734), .CK(net_8912) );
NAND2_X2 inst_3904 ( .A1(net_7113), .A2(net_1675), .ZN(net_1406) );
CLKBUF_X2 inst_9708 ( .A(net_9669), .Z(net_9670) );
CLKBUF_X2 inst_10634 ( .A(net_10595), .Z(net_10596) );
NAND2_X2 inst_2908 ( .ZN(net_5789), .A2(net_5773), .A1(net_413) );
DFF_X2 inst_6333 ( .QN(net_7810), .CK(net_11274), .D(x1459) );
INV_X4 inst_5019 ( .A(net_770), .ZN(net_732) );
INV_X4 inst_5649 ( .A(net_7098), .ZN(net_2569) );
OR2_X4 inst_1393 ( .A2(net_7379), .A1(net_891), .ZN(net_778) );
DFF_X2 inst_6276 ( .D(net_2615), .QN(net_229), .CK(net_9503) );
NAND2_X2 inst_3519 ( .ZN(net_2548), .A2(net_2171), .A1(net_1432) );
NAND2_X2 inst_4075 ( .A1(net_6802), .A2(net_1651), .ZN(net_977) );
CLKBUF_X2 inst_13402 ( .A(net_9678), .Z(net_13364) );
CLKBUF_X2 inst_9507 ( .A(net_9468), .Z(net_9469) );
INV_X4 inst_4893 ( .A(net_3799), .ZN(net_3282) );
INV_X2 inst_5875 ( .A(net_7452), .ZN(net_1376) );
INV_X4 inst_5153 ( .ZN(net_620), .A(net_563) );
INV_X2 inst_5731 ( .ZN(net_3962), .A(net_3961) );
CLKBUF_X2 inst_11318 ( .A(net_10362), .Z(net_11280) );
CLKBUF_X2 inst_14264 ( .A(net_14225), .Z(net_14226) );
CLKBUF_X2 inst_8514 ( .A(net_8475), .Z(net_8476) );
DFF_X1 inst_6717 ( .QN(net_7318), .D(net_5346), .CK(net_10147) );
CLKBUF_X2 inst_8631 ( .A(net_7909), .Z(net_8593) );
CLKBUF_X2 inst_13118 ( .A(net_13079), .Z(net_13080) );
CLKBUF_X2 inst_9807 ( .A(net_9768), .Z(net_9769) );
CLKBUF_X2 inst_14446 ( .A(net_14407), .Z(net_14408) );
CLKBUF_X2 inst_9089 ( .A(net_9050), .Z(net_9051) );
CLKBUF_X2 inst_13684 ( .A(net_13645), .Z(net_13646) );
DFF_X1 inst_6459 ( .QN(net_6128), .D(net_5600), .CK(net_10961) );
INV_X4 inst_4791 ( .ZN(net_1271), .A(net_1270) );
CLKBUF_X2 inst_8007 ( .A(net_7968), .Z(net_7969) );
CLKBUF_X2 inst_9302 ( .A(net_9263), .Z(net_9264) );
AOI22_X2 inst_7244 ( .B1(net_6812), .A1(net_6780), .ZN(net_5318), .A2(net_5316), .B2(net_5315) );
NAND2_X2 inst_2937 ( .ZN(net_5509), .A1(net_4980), .A2(net_4978) );
CLKBUF_X2 inst_12995 ( .A(net_12304), .Z(net_12957) );
DFF_X2 inst_6283 ( .QN(net_7688), .D(net_2487), .CK(net_9497) );
AOI22_X2 inst_7380 ( .B1(net_7744), .A1(net_7715), .A2(net_5916), .B2(net_2957), .ZN(net_2941) );
CLKBUF_X2 inst_7864 ( .A(net_7825), .Z(net_7826) );
SDFF_X2 inst_687 ( .Q(net_6753), .D(net_6753), .SE(net_3815), .SI(net_3789), .CK(net_11333) );
AOI22_X2 inst_7387 ( .A2(net_5916), .B2(net_2957), .ZN(net_2933), .B1(net_2664), .A1(net_709) );
INV_X2 inst_5857 ( .ZN(net_636), .A(net_635) );
CLKBUF_X2 inst_9463 ( .A(net_9424), .Z(net_9425) );
OAI21_X2 inst_1774 ( .B1(net_5440), .ZN(net_5420), .A(net_4699), .B2(net_3989) );
NOR2_X2 inst_2319 ( .A2(net_6259), .A1(net_5840), .ZN(net_5822) );
DFFR_X2 inst_7091 ( .QN(net_6422), .D(net_2697), .CK(net_10239), .RN(x1822) );
CLKBUF_X2 inst_8032 ( .A(net_7993), .Z(net_7994) );
CLKBUF_X2 inst_12596 ( .A(net_12557), .Z(net_12558) );
INV_X4 inst_5519 ( .A(net_7579), .ZN(net_1881) );
SDFF_X2 inst_985 ( .Q(net_6471), .D(net_6471), .SE(net_3904), .SI(net_3810), .CK(net_11664) );
CLKBUF_X2 inst_7927 ( .A(net_7888), .Z(net_7889) );
NOR2_X4 inst_2225 ( .ZN(net_5673), .A1(net_5541), .A2(net_4510) );
CLKBUF_X2 inst_12473 ( .A(net_12434), .Z(net_12435) );
CLKBUF_X2 inst_13805 ( .A(net_13766), .Z(net_13767) );
DFF_X1 inst_6943 ( .QN(net_6050), .D(net_2223), .CK(net_14358) );
NOR2_X2 inst_2513 ( .A1(net_3046), .ZN(net_1160), .A2(net_1159) );
NAND2_X2 inst_4061 ( .A1(net_7211), .A2(net_1648), .ZN(net_991) );
NOR2_X4 inst_2254 ( .ZN(net_5632), .A1(net_5477), .A2(net_4435) );
AOI21_X2 inst_7775 ( .B1(net_6602), .ZN(net_4029), .B2(net_2583), .A(net_2329) );
DFF_X2 inst_6255 ( .Q(net_6388), .D(net_6387), .CK(net_13844) );
CLKBUF_X2 inst_10111 ( .A(net_10072), .Z(net_10073) );
CLKBUF_X2 inst_12985 ( .A(net_12077), .Z(net_12947) );
CLKBUF_X2 inst_10627 ( .A(net_10502), .Z(net_10589) );
CLKBUF_X2 inst_14208 ( .A(net_14169), .Z(net_14170) );
CLKBUF_X2 inst_12563 ( .A(net_12524), .Z(net_12525) );
INV_X2 inst_5918 ( .A(net_7316), .ZN(net_1795) );
CLKBUF_X2 inst_12969 ( .A(net_12930), .Z(net_12931) );
CLKBUF_X2 inst_9255 ( .A(net_9216), .Z(net_9217) );
OAI21_X2 inst_2007 ( .B1(net_5895), .B2(net_4518), .ZN(net_4504), .A(net_3674) );
CLKBUF_X2 inst_10922 ( .A(net_10883), .Z(net_10884) );
CLKBUF_X2 inst_12519 ( .A(net_12480), .Z(net_12481) );
NAND2_X2 inst_3644 ( .ZN(net_2226), .A2(net_1917), .A1(net_1693) );
CLKBUF_X2 inst_10965 ( .A(net_10926), .Z(net_10927) );
SDFF_X2 inst_805 ( .SI(net_7807), .Q(net_6978), .D(net_6978), .SE(net_3891), .CK(net_10870) );
CLKBUF_X2 inst_11755 ( .A(net_11716), .Z(net_11717) );
SDFF_X2 inst_354 ( .SI(net_7641), .Q(net_7641), .D(net_4797), .SE(net_3867), .CK(net_13260) );
CLKBUF_X2 inst_13794 ( .A(net_13755), .Z(net_13756) );
CLKBUF_X2 inst_9991 ( .A(net_9633), .Z(net_9953) );
INV_X2 inst_6005 ( .A(net_7633), .ZN(net_1846) );
SDFF_X2 inst_1145 ( .SI(net_6805), .Q(net_6805), .D(net_3810), .SE(net_3729), .CK(net_8491) );
CLKBUF_X2 inst_12859 ( .A(net_10038), .Z(net_12821) );
DFF_X2 inst_6235 ( .Q(net_7771), .D(net_5928), .CK(net_12378) );
CLKBUF_X2 inst_12387 ( .A(net_9950), .Z(net_12349) );
CLKBUF_X2 inst_12664 ( .A(net_12625), .Z(net_12626) );
CLKBUF_X2 inst_13735 ( .A(net_13696), .Z(net_13697) );
INV_X4 inst_5603 ( .A(net_6410), .ZN(net_1824) );
CLKBUF_X2 inst_14257 ( .A(net_14218), .Z(net_14219) );
DFF_X1 inst_6569 ( .QN(net_7505), .D(net_5093), .CK(net_12088) );
SDFF_X2 inst_373 ( .SI(net_7646), .Q(net_7646), .D(net_4785), .SE(net_3867), .CK(net_10271) );
AOI21_X2 inst_7731 ( .B1(net_6744), .ZN(net_4116), .B2(net_2581), .A(net_2366) );
OAI21_X2 inst_1868 ( .ZN(net_5246), .B1(net_5198), .A(net_4531), .B2(net_3870) );
CLKBUF_X2 inst_13672 ( .A(net_13633), .Z(net_13634) );
CLKBUF_X2 inst_11428 ( .A(net_11389), .Z(net_11390) );
CLKBUF_X2 inst_9537 ( .A(net_8764), .Z(net_9499) );
CLKBUF_X2 inst_8414 ( .A(net_8375), .Z(net_8376) );
XNOR2_X2 inst_22 ( .ZN(net_2577), .A(net_2273), .B(net_1928) );
CLKBUF_X2 inst_13914 ( .A(net_13875), .Z(net_13876) );
OAI21_X2 inst_1717 ( .ZN(net_5577), .B1(net_5545), .A(net_4687), .B2(net_3989) );
NAND2_X2 inst_3099 ( .A1(net_6445), .A2(net_4925), .ZN(net_4904) );
CLKBUF_X2 inst_13289 ( .A(net_13250), .Z(net_13251) );
DFFR_X2 inst_7034 ( .QN(net_6009), .D(net_3195), .CK(net_11431), .RN(x1822) );
NAND2_X4 inst_2901 ( .A1(net_5893), .ZN(net_3399), .A2(net_551) );
SDFF_X2 inst_767 ( .Q(net_6863), .D(net_6863), .SE(net_3901), .SI(net_3802), .CK(net_8933) );
AOI21_X2 inst_7657 ( .B2(net_3439), .ZN(net_3388), .A(net_3210), .B1(net_752) );
CLKBUF_X2 inst_14065 ( .A(net_14026), .Z(net_14027) );
INV_X2 inst_6080 ( .A(net_7648), .ZN(net_2128) );
NAND2_X2 inst_3356 ( .ZN(net_3533), .A1(net_3532), .A2(net_3225) );
SDFF_X2 inst_718 ( .SI(net_6762), .Q(net_6762), .SE(net_3872), .D(net_3799), .CK(net_11093) );
CLKBUF_X2 inst_10405 ( .A(net_9025), .Z(net_10367) );
NAND2_X2 inst_4024 ( .A1(net_6800), .A2(net_1651), .ZN(net_1028) );
CLKBUF_X2 inst_7914 ( .A(net_7875), .Z(net_7876) );
AOI22_X2 inst_7362 ( .A2(net_2994), .B2(net_2993), .ZN(net_2976), .A1(net_1205), .B1(net_1204) );
CLKBUF_X2 inst_8100 ( .A(net_8061), .Z(net_8062) );
CLKBUF_X2 inst_9166 ( .A(net_8310), .Z(net_9128) );
INV_X4 inst_5585 ( .A(net_7416), .ZN(net_2178) );
CLKBUF_X2 inst_8350 ( .A(net_8209), .Z(net_8312) );
NAND2_X1 inst_4310 ( .ZN(net_4556), .A2(net_3866), .A1(net_1986) );
CLKBUF_X2 inst_8943 ( .A(net_8904), .Z(net_8905) );
SDFF_X2 inst_526 ( .SI(net_6641), .Q(net_6641), .SE(net_3850), .D(net_3831), .CK(net_12044) );
OAI21_X2 inst_2147 ( .B1(net_5778), .ZN(net_2797), .A(net_2668), .B2(net_2666) );
CLKBUF_X2 inst_13171 ( .A(net_8053), .Z(net_13133) );
SDFF_X2 inst_1178 ( .SI(net_6950), .Q(net_6950), .D(net_3898), .SE(net_3741), .CK(net_8123) );
OAI21_X2 inst_2091 ( .B2(net_4506), .ZN(net_4325), .B1(net_4132), .A(net_3686) );
NAND2_X2 inst_3104 ( .A1(net_6582), .ZN(net_4898), .A2(net_4897) );
CLKBUF_X2 inst_9174 ( .A(net_8323), .Z(net_9136) );
OAI22_X2 inst_1450 ( .B1(net_4855), .ZN(net_4623), .A2(net_4622), .B2(net_4621), .A1(net_4218) );
CLKBUF_X2 inst_8423 ( .A(net_8384), .Z(net_8385) );
DFF_X1 inst_6689 ( .QN(net_7278), .D(net_5115), .CK(net_9452) );
CLKBUF_X2 inst_12247 ( .A(net_12208), .Z(net_12209) );
CLKBUF_X2 inst_10733 ( .A(net_10694), .Z(net_10695) );
INV_X4 inst_5511 ( .A(net_7570), .ZN(net_1861) );
NAND2_X2 inst_3123 ( .A1(net_6612), .A2(net_4899), .ZN(net_4878) );
CLKBUF_X2 inst_8066 ( .A(net_7892), .Z(net_8028) );
CLKBUF_X2 inst_11592 ( .A(net_9085), .Z(net_11554) );
CLKBUF_X2 inst_11149 ( .A(net_11110), .Z(net_11111) );
INV_X2 inst_5863 ( .A(net_835), .ZN(net_583) );
CLKBUF_X2 inst_10645 ( .A(net_10397), .Z(net_10607) );
NAND2_X2 inst_3725 ( .A1(net_6762), .A2(net_1635), .ZN(net_1620) );
INV_X4 inst_5400 ( .A(net_7267), .ZN(net_2051) );
SDFF_X2 inst_500 ( .Q(net_6974), .D(net_6974), .SI(net_3894), .SE(net_3891), .CK(net_8228) );
OAI22_X2 inst_1592 ( .A1(net_3273), .B2(net_3200), .A2(net_3196), .ZN(net_3161), .B1(net_470) );
INV_X4 inst_5348 ( .A(net_7746), .ZN(net_2938) );
OAI21_X2 inst_1770 ( .B1(net_5448), .ZN(net_5424), .A(net_4703), .B2(net_3989) );
CLKBUF_X2 inst_14403 ( .A(net_14364), .Z(net_14365) );
SDFF_X2 inst_550 ( .Q(net_6431), .D(net_6431), .SI(net_3883), .SE(net_3820), .CK(net_11671) );
NAND2_X2 inst_3413 ( .A2(net_5976), .ZN(net_3380), .A1(net_2880) );
INV_X2 inst_6095 ( .A(net_7294), .ZN(net_2077) );
DFF_X1 inst_6758 ( .QN(net_7301), .D(net_4871), .CK(net_9870) );
INV_X8 inst_4483 ( .ZN(net_4274), .A(net_3925) );
CLKBUF_X2 inst_12857 ( .A(net_12818), .Z(net_12819) );
INV_X2 inst_5913 ( .A(net_7662), .ZN(net_1850) );
CLKBUF_X2 inst_11972 ( .A(net_11933), .Z(net_11934) );
CLKBUF_X2 inst_13610 ( .A(net_13571), .Z(net_13572) );
CLKBUF_X2 inst_8311 ( .A(net_8272), .Z(net_8273) );
CLKBUF_X2 inst_8702 ( .A(net_8663), .Z(net_8664) );
CLKBUF_X2 inst_11109 ( .A(net_11070), .Z(net_11071) );
CLKBUF_X2 inst_14132 ( .A(net_14093), .Z(net_14094) );
INV_X4 inst_5471 ( .A(net_7726), .ZN(net_2647) );
OR2_X2 inst_1419 ( .ZN(net_3761), .A2(net_785), .A1(net_504) );
NAND3_X2 inst_2661 ( .ZN(net_3935), .A3(net_3396), .A2(net_2958), .A1(net_2840) );
CLKBUF_X2 inst_8237 ( .A(net_8133), .Z(net_8199) );
INV_X2 inst_6034 ( .A(net_7351), .ZN(net_2004) );
NOR2_X2 inst_2501 ( .ZN(net_2585), .A1(net_2489), .A2(net_689) );
NAND2_X2 inst_3548 ( .ZN(net_2519), .A2(net_2016), .A1(net_1755) );
SDFF_X2 inst_594 ( .Q(net_6564), .D(net_6564), .SE(net_3823), .SI(net_3798), .CK(net_12923) );
CLKBUF_X2 inst_13848 ( .A(net_8952), .Z(net_13810) );
NAND2_X1 inst_4435 ( .A2(net_2131), .ZN(net_1390), .A1(net_1389) );
CLKBUF_X2 inst_14164 ( .A(net_12964), .Z(net_14126) );
OAI222_X2 inst_1632 ( .A1(net_5866), .C2(net_5087), .ZN(net_5086), .A2(net_5085), .B2(net_5084), .B1(net_2450), .C1(net_599) );
NOR4_X2 inst_2175 ( .ZN(net_3246), .A4(net_3119), .A1(net_2640), .A3(net_2476), .A2(net_834) );
NAND2_X1 inst_4241 ( .ZN(net_4686), .A2(net_3989), .A1(net_2106) );
SDFF_X2 inst_925 ( .Q(net_7162), .D(net_7162), .SE(net_3903), .SI(net_3800), .CK(net_10640) );
CLKBUF_X2 inst_13314 ( .A(net_11356), .Z(net_13276) );
NOR3_X2 inst_2193 ( .ZN(net_3884), .A1(net_3387), .A3(net_1741), .A2(net_809) );
NOR2_X2 inst_2378 ( .ZN(net_5129), .A2(net_4607), .A1(net_4406) );
CLKBUF_X2 inst_10302 ( .A(net_10263), .Z(net_10264) );
DFF_X2 inst_6302 ( .D(net_1691), .QN(net_265), .CK(net_10780) );
CLKBUF_X2 inst_14137 ( .A(net_14098), .Z(net_14099) );
CLKBUF_X2 inst_9996 ( .A(net_9895), .Z(net_9958) );
CLKBUF_X2 inst_8734 ( .A(net_8695), .Z(net_8696) );
CLKBUF_X2 inst_9793 ( .A(net_8869), .Z(net_9755) );
CLKBUF_X2 inst_8999 ( .A(net_8960), .Z(net_8961) );
INV_X16 inst_6147 ( .A(net_5943), .ZN(net_5941) );
CLKBUF_X2 inst_14392 ( .A(net_12863), .Z(net_14354) );
OAI22_X2 inst_1536 ( .B1(net_4637), .A1(net_4030), .B2(net_4026), .ZN(net_4023), .A2(net_4022) );
SDFF_X2 inst_881 ( .Q(net_7111), .D(net_7111), .SE(net_3888), .SI(net_3812), .CK(net_12162) );
CLKBUF_X2 inst_13874 ( .A(net_13835), .Z(net_13836) );
CLKBUF_X2 inst_11300 ( .A(net_11261), .Z(net_11262) );
NAND2_X2 inst_3876 ( .A1(net_6837), .A2(net_1521), .ZN(net_1444) );
NAND2_X2 inst_3848 ( .A2(net_1696), .ZN(net_1489), .A1(net_1488) );
CLKBUF_X2 inst_13164 ( .A(net_13125), .Z(net_13126) );
DFFR_X2 inst_7001 ( .QN(net_7718), .D(net_3351), .CK(net_8603), .RN(x1822) );
CLKBUF_X2 inst_12175 ( .A(net_12136), .Z(net_12137) );
CLKBUF_X2 inst_12079 ( .A(net_12040), .Z(net_12041) );
NAND2_X2 inst_3706 ( .A1(net_7039), .A2(net_1975), .ZN(net_1644) );
CLKBUF_X2 inst_10072 ( .A(net_10033), .Z(net_10034) );
CLKBUF_X2 inst_13979 ( .A(net_8225), .Z(net_13941) );
CLKBUF_X2 inst_11153 ( .A(net_11114), .Z(net_11115) );
CLKBUF_X2 inst_9219 ( .A(net_9180), .Z(net_9181) );
SDFF_X2 inst_247 ( .Q(net_6347), .SI(net_6346), .D(net_3581), .SE(net_392), .CK(net_14130) );
DFFR_X2 inst_7066 ( .QN(net_6045), .D(net_3086), .CK(net_10005), .RN(x1822) );
INV_X2 inst_6089 ( .A(net_7290), .ZN(net_1991) );
SDFF_X2 inst_403 ( .SI(net_7366), .Q(net_7366), .D(net_4783), .SE(net_3853), .CK(net_9907) );
CLKBUF_X2 inst_12031 ( .A(net_11992), .Z(net_11993) );
DFF_X1 inst_6740 ( .QN(net_7332), .D(net_4865), .CK(net_12690) );
CLKBUF_X2 inst_10501 ( .A(net_10462), .Z(net_10463) );
NAND2_X2 inst_3446 ( .A1(net_7763), .ZN(net_3070), .A2(net_3057) );
NAND3_X2 inst_2728 ( .ZN(net_2373), .A3(net_1632), .A1(net_1461), .A2(net_1028) );
CLKBUF_X2 inst_10796 ( .A(net_10757), .Z(net_10758) );
CLKBUF_X2 inst_8847 ( .A(net_8808), .Z(net_8809) );
OAI22_X2 inst_1588 ( .A1(net_3268), .B2(net_3200), .A2(net_3196), .ZN(net_3185), .B1(net_575) );
NAND2_X2 inst_3801 ( .A1(net_6623), .A2(net_1624), .ZN(net_1544) );
NAND2_X2 inst_4177 ( .A2(net_6553), .ZN(net_774), .A1(net_581) );
CLKBUF_X2 inst_9350 ( .A(net_8506), .Z(net_9312) );
CLKBUF_X2 inst_8002 ( .A(net_7963), .Z(net_7964) );
CLKBUF_X2 inst_10996 ( .A(net_10957), .Z(net_10958) );
DFF_X1 inst_6491 ( .QN(net_7403), .D(net_5558), .CK(net_12126) );
NOR2_X2 inst_2516 ( .A1(net_5934), .ZN(net_2916), .A2(net_537) );
CLKBUF_X2 inst_13133 ( .A(net_13094), .Z(net_13095) );
CLKBUF_X2 inst_9193 ( .A(net_8249), .Z(net_9155) );
CLKBUF_X2 inst_13901 ( .A(net_13862), .Z(net_13863) );
OAI21_X2 inst_2155 ( .ZN(net_2690), .B2(net_2687), .A(net_2618), .B1(net_693) );
CLKBUF_X2 inst_12927 ( .A(net_12888), .Z(net_12889) );
CLKBUF_X2 inst_9567 ( .A(net_9528), .Z(net_9529) );
DFF_X1 inst_6352 ( .QN(net_6206), .D(net_5832), .CK(net_13709) );
OAI22_X2 inst_1506 ( .B1(net_4660), .B2(net_4500), .A2(net_4109), .A1(net_4105), .ZN(net_4086) );
CLKBUF_X2 inst_9494 ( .A(net_9455), .Z(net_9456) );
SDFF_X2 inst_464 ( .Q(net_6886), .D(net_6886), .SI(net_3902), .SE(net_3901), .CK(net_11517) );
CLKBUF_X2 inst_13428 ( .A(net_13389), .Z(net_13390) );
INV_X4 inst_5360 ( .A(net_7561), .ZN(net_1868) );
CLKBUF_X2 inst_13392 ( .A(net_13353), .Z(net_13354) );
CLKBUF_X2 inst_10455 ( .A(net_8679), .Z(net_10417) );
AOI222_X2 inst_7541 ( .C1(net_7676), .A1(net_7644), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1880), .B1(net_1879) );
INV_X2 inst_6058 ( .A(net_7624), .ZN(net_1842) );
SDFF_X2 inst_341 ( .SI(net_7374), .Q(net_7374), .D(net_4784), .SE(net_3853), .CK(net_12767) );
NAND2_X2 inst_3785 ( .A1(net_6501), .A2(net_1642), .ZN(net_1560) );
CLKBUF_X2 inst_12313 ( .A(net_11324), .Z(net_12275) );
CLKBUF_X2 inst_13090 ( .A(net_13051), .Z(net_13052) );
INV_X4 inst_5678 ( .A(net_6151), .ZN(net_3581) );
CLKBUF_X2 inst_14006 ( .A(net_13967), .Z(net_13968) );
CLKBUF_X2 inst_11095 ( .A(net_11056), .Z(net_11057) );
NOR2_X2 inst_2359 ( .ZN(net_5305), .A2(net_4635), .A1(net_4507) );
NAND2_X2 inst_3702 ( .A1(net_6441), .ZN(net_1678), .A2(net_1677) );
CLKBUF_X2 inst_11229 ( .A(net_11190), .Z(net_11191) );
CLKBUF_X2 inst_8526 ( .A(net_8487), .Z(net_8488) );
CLKBUF_X2 inst_13913 ( .A(net_13874), .Z(net_13875) );
CLKBUF_X2 inst_13031 ( .A(net_12426), .Z(net_12993) );
CLKBUF_X2 inst_8505 ( .A(net_8466), .Z(net_8467) );
AOI22_X2 inst_7454 ( .B2(net_7740), .A2(net_7739), .B1(net_7711), .A1(net_7710), .ZN(net_660) );
INV_X4 inst_5556 ( .A(net_7279), .ZN(net_2023) );
DFF_X1 inst_6826 ( .D(net_3005), .CK(net_13404), .Q(x179) );
SDFFR_X2 inst_1361 ( .SI(net_7741), .Q(net_7741), .D(net_4596), .SE(net_2604), .CK(net_13180), .RN(x1822) );
CLKBUF_X2 inst_10226 ( .A(net_10187), .Z(net_10188) );
NAND2_X2 inst_3401 ( .ZN(net_3461), .A2(net_3323), .A1(net_3233) );
CLKBUF_X2 inst_13105 ( .A(net_13066), .Z(net_13067) );
CLKBUF_X2 inst_12949 ( .A(net_8817), .Z(net_12911) );
CLKBUF_X2 inst_12688 ( .A(net_12649), .Z(net_12650) );
CLKBUF_X2 inst_12439 ( .A(net_12400), .Z(net_12401) );
CLKBUF_X2 inst_11916 ( .A(net_11877), .Z(net_11878) );
AOI222_X2 inst_7525 ( .C1(net_7518), .B1(net_7486), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_1990), .A1(net_1989) );
CLKBUF_X2 inst_8840 ( .A(net_8432), .Z(net_8802) );
INV_X4 inst_4968 ( .ZN(net_2249), .A(net_702) );
INV_X8 inst_4463 ( .ZN(net_5297), .A(net_4288) );
NOR3_X2 inst_2208 ( .ZN(net_2617), .A3(net_2616), .A1(net_2489), .A2(net_765) );
CLKBUF_X2 inst_14319 ( .A(net_14280), .Z(net_14281) );
INV_X4 inst_5598 ( .A(net_5985), .ZN(net_652) );
CLKBUF_X2 inst_8789 ( .A(net_8750), .Z(net_8751) );
CLKBUF_X2 inst_10698 ( .A(net_10659), .Z(net_10660) );
CLKBUF_X2 inst_10122 ( .A(net_10083), .Z(net_10084) );
NAND2_X2 inst_4162 ( .ZN(net_933), .A2(net_534), .A1(net_530) );
CLKBUF_X2 inst_8975 ( .A(net_8936), .Z(net_8937) );
CLKBUF_X2 inst_7873 ( .A(net_7829), .Z(net_7835) );
INV_X4 inst_5171 ( .A(net_1657), .ZN(net_537) );
CLKBUF_X2 inst_12936 ( .A(net_12897), .Z(net_12898) );
NOR4_X2 inst_2174 ( .ZN(net_3247), .A4(net_3123), .A1(net_2638), .A3(net_2484), .A2(net_830) );
DFF_X1 inst_6721 ( .QN(net_7323), .D(net_5336), .CK(net_10138) );
CLKBUF_X2 inst_14363 ( .A(net_14324), .Z(net_14325) );
NAND2_X2 inst_3201 ( .ZN(net_4725), .A2(net_3986), .A1(net_1884) );
CLKBUF_X2 inst_10779 ( .A(net_10537), .Z(net_10741) );
CLKBUF_X2 inst_13089 ( .A(net_13050), .Z(net_13051) );
AOI21_X2 inst_7702 ( .B1(net_6461), .ZN(net_5911), .B2(net_2580), .A(net_2305) );
XNOR2_X2 inst_14 ( .ZN(net_2641), .B(net_2640), .A(net_2477) );
CLKBUF_X2 inst_9366 ( .A(net_8196), .Z(net_9328) );
CLKBUF_X2 inst_7886 ( .A(net_7847), .Z(net_7848) );
CLKBUF_X2 inst_12068 ( .A(net_9644), .Z(net_12030) );
NOR2_X2 inst_2325 ( .A2(net_6293), .A1(net_5840), .ZN(net_5816) );
CLKBUF_X2 inst_12354 ( .A(net_12315), .Z(net_12316) );
SDFF_X2 inst_251 ( .Q(net_6343), .SI(net_6342), .D(net_3589), .SE(net_392), .CK(net_13499) );
CLKBUF_X2 inst_10651 ( .A(net_10612), .Z(net_10613) );
CLKBUF_X2 inst_7983 ( .A(net_7944), .Z(net_7945) );
SDFF_X2 inst_1074 ( .SI(net_7199), .Q(net_7199), .D(net_3799), .SE(net_3751), .CK(net_13315) );
AOI22_X2 inst_7375 ( .A2(net_5916), .B2(net_2957), .ZN(net_2946), .B1(net_2673), .A1(net_847) );
CLKBUF_X2 inst_10149 ( .A(net_10110), .Z(net_10111) );
OAI22_X2 inst_1552 ( .B2(net_3405), .A2(net_3360), .ZN(net_3353), .A1(net_3188), .B1(net_511) );
OAI22_X2 inst_1524 ( .B1(net_4644), .A1(net_4057), .B2(net_4051), .ZN(net_4048), .A2(net_4047) );
CLKBUF_X2 inst_13983 ( .A(net_11093), .Z(net_13945) );
CLKBUF_X2 inst_9369 ( .A(net_9330), .Z(net_9331) );
INV_X4 inst_4789 ( .A(net_2804), .ZN(net_1715) );
INV_X4 inst_4977 ( .A(net_3002), .ZN(net_879) );
CLKBUF_X2 inst_11100 ( .A(net_11061), .Z(net_11062) );
CLKBUF_X2 inst_9892 ( .A(net_9777), .Z(net_9854) );
CLKBUF_X2 inst_9883 ( .A(net_9844), .Z(net_9845) );
AOI21_X2 inst_7781 ( .B1(net_6608), .ZN(net_4016), .B2(net_2583), .A(net_2287) );
OAI22_X2 inst_1602 ( .B2(net_3200), .A2(net_3144), .ZN(net_3134), .A1(net_3133), .B1(net_767) );
SDFF_X2 inst_969 ( .Q(net_6448), .D(net_6448), .SE(net_3820), .SI(net_3796), .CK(net_10849) );
CLKBUF_X2 inst_8567 ( .A(net_8528), .Z(net_8529) );
DFF_X1 inst_6463 ( .QN(net_6148), .D(net_5596), .CK(net_11989) );
CLKBUF_X2 inst_13081 ( .A(net_13042), .Z(net_13043) );
CLKBUF_X2 inst_12487 ( .A(net_12448), .Z(net_12449) );
NOR2_X2 inst_2528 ( .ZN(net_2708), .A2(net_295), .A1(net_289) );
CLKBUF_X2 inst_9749 ( .A(net_9710), .Z(net_9711) );
INV_X4 inst_4917 ( .A(net_3813), .ZN(net_3268) );
CLKBUF_X2 inst_13628 ( .A(net_13589), .Z(net_13590) );
SDFF_X2 inst_898 ( .Q(net_7129), .D(net_7129), .SE(net_3888), .SI(net_3801), .CK(net_10644) );
DFFR_X2 inst_7049 ( .QN(net_6018), .D(net_3189), .CK(net_10436), .RN(x1822) );
OAI21_X2 inst_1977 ( .B1(net_4868), .ZN(net_4859), .A(net_4376), .B2(net_3853) );
OAI21_X2 inst_1793 ( .B1(net_5412), .ZN(net_5397), .A(net_4672), .B2(net_3988) );
NAND2_X1 inst_4227 ( .ZN(net_4700), .A2(net_3989), .A1(net_2193) );
CLKBUF_X2 inst_8012 ( .A(net_7973), .Z(net_7974) );
DFF_X1 inst_6840 ( .Q(net_389), .D(net_386), .CK(net_12239) );
CLKBUF_X2 inst_9800 ( .A(net_9761), .Z(net_9762) );
CLKBUF_X2 inst_9223 ( .A(net_9184), .Z(net_9185) );
CLKBUF_X2 inst_9747 ( .A(net_8930), .Z(net_9709) );
CLKBUF_X2 inst_11804 ( .A(net_11765), .Z(net_11766) );
INV_X4 inst_5299 ( .A(net_7233), .ZN(net_2567) );
CLKBUF_X2 inst_10824 ( .A(net_9371), .Z(net_10786) );
CLKBUF_X2 inst_10805 ( .A(net_10766), .Z(net_10767) );
INV_X4 inst_5697 ( .A(net_5916), .ZN(net_5915) );
CLKBUF_X2 inst_12290 ( .A(net_8724), .Z(net_12252) );
NOR2_X4 inst_2291 ( .A2(net_7791), .ZN(net_2865), .A1(net_416) );
NOR2_X2 inst_2343 ( .A2(net_5992), .A1(net_5778), .ZN(net_5710) );
CLKBUF_X2 inst_8230 ( .A(net_8191), .Z(net_8192) );
CLKBUF_X2 inst_11500 ( .A(net_11461), .Z(net_11462) );
NOR2_X2 inst_2538 ( .A2(net_7760), .A1(net_3208), .ZN(net_656) );
INV_X2 inst_5708 ( .ZN(net_4310), .A(net_4217) );
INV_X4 inst_4822 ( .ZN(net_1091), .A(net_1090) );
NAND2_X2 inst_3132 ( .ZN(net_4831), .A2(net_4153), .A1(net_2166) );
CLKBUF_X2 inst_13835 ( .A(net_13796), .Z(net_13797) );
AOI22_X2 inst_7395 ( .A2(net_3105), .B1(net_2970), .ZN(net_2846), .A1(net_645), .B2(net_255) );
INV_X4 inst_4999 ( .A(net_6823), .ZN(net_1150) );
INV_X2 inst_6071 ( .A(net_7365), .ZN(net_2042) );
INV_X2 inst_5819 ( .A(net_1308), .ZN(net_1051) );
NAND2_X2 inst_3910 ( .A1(net_6712), .A2(net_1497), .ZN(net_1397) );
CLKBUF_X2 inst_12303 ( .A(net_7846), .Z(net_12265) );
SDFFR_X2 inst_1332 ( .SE(net_4147), .D(net_4146), .SI(net_155), .Q(net_155), .CK(net_12363), .RN(x1822) );
CLKBUF_X2 inst_12427 ( .A(net_10551), .Z(net_12389) );
OAI21_X2 inst_1841 ( .B1(net_5359), .ZN(net_5331), .A(net_4371), .B2(net_3853) );
CLKBUF_X2 inst_11929 ( .A(net_11890), .Z(net_11891) );
NAND2_X2 inst_3345 ( .ZN(net_3557), .A1(net_3556), .A2(net_3225) );
NAND2_X2 inst_3264 ( .A2(net_3858), .ZN(net_3853), .A1(net_1646) );
CLKBUF_X2 inst_12584 ( .A(net_12545), .Z(net_12546) );
INV_X4 inst_5169 ( .ZN(net_540), .A(net_539) );
INV_X4 inst_4945 ( .ZN(net_743), .A(net_742) );
CLKBUF_X2 inst_8782 ( .A(net_8231), .Z(net_8744) );
NOR2_X2 inst_2332 ( .A2(net_6286), .A1(net_5840), .ZN(net_5809) );
CLKBUF_X2 inst_9982 ( .A(net_8293), .Z(net_9944) );
CLKBUF_X2 inst_13415 ( .A(net_13376), .Z(net_13377) );
CLKBUF_X2 inst_9082 ( .A(net_9043), .Z(net_9044) );
CLKBUF_X2 inst_13431 ( .A(net_13392), .Z(net_13393) );
CLKBUF_X2 inst_13908 ( .A(net_12809), .Z(net_13870) );
CLKBUF_X2 inst_10970 ( .A(net_10931), .Z(net_10932) );
INV_X2 inst_5946 ( .A(net_7471), .ZN(net_2110) );
NOR2_X2 inst_2310 ( .A2(net_6204), .A1(net_5840), .ZN(net_5831) );
CLKBUF_X2 inst_9720 ( .A(net_9681), .Z(net_9682) );
SDFF_X2 inst_1089 ( .SI(net_7075), .Q(net_7075), .D(net_3810), .SE(net_3742), .CK(net_11860) );
CLKBUF_X2 inst_10251 ( .A(net_7833), .Z(net_10213) );
DFF_X1 inst_6537 ( .QN(net_7469), .D(net_5579), .CK(net_12108) );
CLKBUF_X2 inst_14327 ( .A(net_10159), .Z(net_14289) );
DFF_X1 inst_6430 ( .QN(net_6173), .D(net_5740), .CK(net_11607) );
INV_X4 inst_5017 ( .A(net_7793), .ZN(net_3792) );
DFF_X1 inst_6932 ( .D(net_2400), .Q(net_246), .CK(net_8021) );
SDFF_X2 inst_1290 ( .D(net_3814), .SE(net_3256), .SI(net_138), .Q(net_138), .CK(net_8462) );
CLKBUF_X2 inst_7939 ( .A(net_7858), .Z(net_7901) );
CLKBUF_X2 inst_11451 ( .A(net_10239), .Z(net_11413) );
DFF_X1 inst_6342 ( .QN(net_6189), .D(net_5844), .CK(net_13647) );
INV_X4 inst_5367 ( .A(net_7229), .ZN(net_415) );
CLKBUF_X2 inst_9092 ( .A(net_9053), .Z(net_9054) );
INV_X2 inst_5845 ( .ZN(net_1951), .A(net_736) );
INV_X4 inst_5038 ( .A(net_7824), .ZN(net_3800) );
CLKBUF_X2 inst_13399 ( .A(net_13360), .Z(net_13361) );
INV_X4 inst_5142 ( .ZN(net_1144), .A(net_574) );
INV_X2 inst_5757 ( .A(net_3399), .ZN(net_3322) );
CLKBUF_X2 inst_12614 ( .A(net_12575), .Z(net_12576) );
INV_X4 inst_4899 ( .ZN(net_870), .A(net_869) );
OAI21_X2 inst_2046 ( .B2(net_4457), .ZN(net_4454), .B1(net_4083), .A(net_3522) );
CLKBUF_X2 inst_12021 ( .A(net_11982), .Z(net_11983) );
INV_X2 inst_6041 ( .A(net_7511), .ZN(net_2184) );
CLKBUF_X2 inst_12604 ( .A(net_12565), .Z(net_12566) );
INV_X4 inst_5079 ( .A(net_7793), .ZN(net_3797) );
NAND2_X2 inst_4129 ( .A2(net_1228), .ZN(net_1163), .A1(net_379) );
CLKBUF_X2 inst_11632 ( .A(net_11593), .Z(net_11594) );
AOI222_X2 inst_7505 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2052), .A1(net_2051), .B1(net_2050), .C1(net_2049) );
DFF_X1 inst_6340 ( .Q(net_6195), .D(net_5846), .CK(net_13773) );
DFF_X1 inst_6429 ( .QN(net_6172), .D(net_5741), .CK(net_11611) );
NAND2_X2 inst_3861 ( .A2(net_1696), .ZN(net_1472), .A1(net_1471) );
NAND2_X1 inst_4399 ( .A2(net_3297), .ZN(net_3081), .A1(net_3080) );
CLKBUF_X2 inst_14176 ( .A(net_14039), .Z(net_14138) );
CLKBUF_X2 inst_11547 ( .A(net_11508), .Z(net_11509) );
CLKBUF_X2 inst_9847 ( .A(net_9808), .Z(net_9809) );
CLKBUF_X2 inst_9840 ( .A(net_9801), .Z(net_9802) );
CLKBUF_X2 inst_14224 ( .A(net_14185), .Z(net_14186) );
CLKBUF_X2 inst_13783 ( .A(net_13744), .Z(net_13745) );
DFF_X1 inst_6533 ( .QN(net_7480), .D(net_5418), .CK(net_12478) );
NAND2_X2 inst_4196 ( .A1(net_2839), .ZN(net_1211), .A2(net_304) );
NAND2_X2 inst_3524 ( .ZN(net_2543), .A2(net_2098), .A1(net_1328) );
CLKBUF_X2 inst_12333 ( .A(net_12294), .Z(net_12295) );
CLKBUF_X2 inst_10672 ( .A(net_10633), .Z(net_10634) );
INV_X8 inst_4479 ( .ZN(net_4899), .A(net_4261) );
SDFF_X2 inst_1014 ( .SI(net_6489), .Q(net_6489), .SE(net_3886), .D(net_3806), .CK(net_8762) );
NOR2_X2 inst_2531 ( .ZN(net_3861), .A2(net_886), .A1(net_770) );
CLKBUF_X2 inst_10009 ( .A(net_9970), .Z(net_9971) );
DFF_X1 inst_6781 ( .QN(net_6165), .D(net_4321), .CK(net_7941) );
CLKBUF_X2 inst_11879 ( .A(net_11840), .Z(net_11841) );
CLKBUF_X2 inst_10882 ( .A(net_10275), .Z(net_10844) );
AOI21_X2 inst_7719 ( .B1(net_6870), .ZN(net_4103), .B2(net_2579), .A(net_2337) );
INV_X4 inst_4782 ( .ZN(net_2636), .A(net_1661) );
SDFFR_X2 inst_1347 ( .SE(net_3256), .D(net_718), .SI(net_146), .Q(net_146), .CK(net_10705), .RN(x1822) );
CLKBUF_X2 inst_11073 ( .A(net_11034), .Z(net_11035) );
SDFF_X2 inst_509 ( .SI(net_6761), .Q(net_6761), .D(net_3892), .SE(net_3872), .CK(net_8308) );
CLKBUF_X2 inst_12299 ( .A(net_12260), .Z(net_12261) );
NAND3_X2 inst_2687 ( .ZN(net_3176), .A2(net_3167), .A3(net_3047), .A1(net_3003) );
OAI221_X2 inst_1680 ( .ZN(net_3369), .A(net_3180), .B2(net_2983), .C2(net_2901), .C1(net_2858), .B1(net_1966) );
CLKBUF_X2 inst_11775 ( .A(net_10992), .Z(net_11737) );
CLKBUF_X2 inst_11473 ( .A(net_11434), .Z(net_11435) );
OAI22_X2 inst_1626 ( .B1(net_6420), .A2(net_2820), .B2(net_2718), .ZN(net_2717), .A1(net_1039) );
NAND3_X2 inst_2622 ( .ZN(net_5717), .A1(net_5612), .A2(net_5125), .A3(net_4176) );
SDFF_X2 inst_153 ( .Q(net_6225), .SI(net_6224), .SE(net_392), .D(net_131), .CK(net_14089) );
CLKBUF_X2 inst_12834 ( .A(net_11741), .Z(net_12796) );
INV_X4 inst_4856 ( .ZN(net_1057), .A(net_1045) );
CLKBUF_X2 inst_9751 ( .A(net_8988), .Z(net_9713) );
CLKBUF_X2 inst_12271 ( .A(net_12232), .Z(net_12233) );
OAI22_X2 inst_1459 ( .B2(net_5910), .B1(net_4644), .A2(net_4610), .ZN(net_4608), .A1(net_4041) );
NAND2_X2 inst_4094 ( .A1(net_6529), .A2(net_1645), .ZN(net_958) );
CLKBUF_X2 inst_10483 ( .A(net_10444), .Z(net_10445) );
DFF_X1 inst_6528 ( .QN(net_7475), .D(net_5423), .CK(net_10085) );
CLKBUF_X2 inst_9789 ( .A(net_9750), .Z(net_9751) );
CLKBUF_X2 inst_9117 ( .A(net_9078), .Z(net_9079) );
SDFF_X2 inst_209 ( .Q(net_6305), .SI(net_6304), .D(net_3677), .SE(net_392), .CK(net_13556) );
NAND2_X2 inst_3894 ( .A2(net_1696), .ZN(net_1422), .A1(net_1421) );
INV_X2 inst_6068 ( .A(net_7501), .ZN(net_2119) );
CLKBUF_X2 inst_8037 ( .A(net_7998), .Z(net_7999) );
CLKBUF_X2 inst_10132 ( .A(net_10093), .Z(net_10094) );
INV_X4 inst_5385 ( .A(net_6022), .ZN(net_472) );
SDFF_X2 inst_1087 ( .SI(net_7079), .Q(net_7079), .D(net_3784), .SE(net_3747), .CK(net_8998) );
DFF_X1 inst_6365 ( .QN(net_6297), .D(net_5819), .CK(net_13795) );
OAI21_X2 inst_1781 ( .ZN(net_5411), .B1(net_5410), .A(net_4691), .B2(net_3989) );
CLKBUF_X2 inst_13701 ( .A(net_13662), .Z(net_13663) );
NAND3_X2 inst_2769 ( .ZN(net_2331), .A3(net_1603), .A1(net_1393), .A2(net_951) );
CLKBUF_X2 inst_14453 ( .A(net_14414), .Z(net_14415) );
CLKBUF_X2 inst_10061 ( .A(net_9340), .Z(net_10023) );
OR2_X4 inst_1375 ( .ZN(net_3446), .A2(net_3250), .A1(net_2612) );
CLKBUF_X2 inst_11353 ( .A(net_10805), .Z(net_11315) );
DFF_X2 inst_6230 ( .QN(net_7233), .D(net_3717), .CK(net_12540) );
CLKBUF_X2 inst_12199 ( .A(net_12160), .Z(net_12161) );
CLKBUF_X2 inst_7966 ( .A(net_7927), .Z(net_7928) );
NAND2_X2 inst_3982 ( .ZN(net_1288), .A1(net_885), .A2(net_321) );
INV_X8 inst_4564 ( .ZN(net_1648), .A(net_487) );
DFF_X1 inst_6482 ( .QN(net_7413), .D(net_5570), .CK(net_9312) );
CLKBUF_X2 inst_14273 ( .A(net_14234), .Z(net_14235) );
CLKBUF_X2 inst_9290 ( .A(net_9251), .Z(net_9252) );
INV_X4 inst_5258 ( .ZN(net_1143), .A(net_433) );
NAND2_X2 inst_3215 ( .ZN(net_4711), .A2(net_3986), .A1(net_1858) );
CLKBUF_X2 inst_12235 ( .A(net_12196), .Z(net_12197) );
INV_X2 inst_5810 ( .ZN(net_1207), .A(net_1206) );
CLKBUF_X2 inst_11209 ( .A(net_8183), .Z(net_11171) );
NAND4_X2 inst_2564 ( .ZN(net_1673), .A1(net_854), .A4(net_840), .A2(net_714), .A3(net_711) );
CLKBUF_X2 inst_8462 ( .A(net_8337), .Z(net_8424) );
SDFF_X2 inst_1082 ( .SI(net_7068), .Q(net_7068), .D(net_3814), .SE(net_3742), .CK(net_9003) );
NAND2_X2 inst_4167 ( .A2(net_7228), .ZN(net_821), .A1(net_415) );
CLKBUF_X2 inst_9204 ( .A(net_9047), .Z(net_9166) );
NAND3_X2 inst_2677 ( .ZN(net_3459), .A3(net_3305), .A1(net_2964), .A2(net_2954) );
NAND2_X1 inst_4374 ( .ZN(net_4353), .A2(net_3856), .A1(net_1788) );
OAI21_X2 inst_1995 ( .ZN(net_4520), .B1(net_4519), .B2(net_4518), .A(net_3700) );
CLKBUF_X2 inst_10068 ( .A(net_9923), .Z(net_10030) );
XNOR2_X2 inst_105 ( .B(net_3004), .ZN(net_1659), .A(net_1148) );
CLKBUF_X2 inst_9145 ( .A(net_9106), .Z(net_9107) );
NAND2_X2 inst_3518 ( .ZN(net_2549), .A2(net_1982), .A1(net_1470) );
OAI21_X2 inst_2161 ( .ZN(net_2850), .A(net_303), .B2(net_302), .B1(net_268) );
CLKBUF_X2 inst_8294 ( .A(net_8255), .Z(net_8256) );
SDFF_X2 inst_625 ( .SI(net_6635), .Q(net_6635), .SE(net_3851), .D(net_3812), .CK(net_9159) );
AOI22_X2 inst_7405 ( .B1(net_5939), .A2(net_2838), .ZN(net_2832), .A1(net_496), .B2(net_195) );
CLKBUF_X2 inst_12736 ( .A(net_12697), .Z(net_12698) );
NAND2_X2 inst_3367 ( .ZN(net_3512), .A1(net_3511), .A2(net_3223) );
DFF_X1 inst_6747 ( .QN(net_7586), .D(net_4848), .CK(net_10292) );
CLKBUF_X2 inst_14041 ( .A(net_14002), .Z(net_14003) );
SDFF_X2 inst_568 ( .SI(net_6776), .Q(net_6776), .SE(net_3872), .D(net_3831), .CK(net_8531) );
OAI22_X2 inst_1483 ( .A2(net_4162), .B2(net_4161), .ZN(net_4160), .B1(net_1695), .A1(net_1694) );
SDFF_X2 inst_523 ( .D(net_7807), .SI(net_6637), .Q(net_6637), .SE(net_3851), .CK(net_9365) );
CLKBUF_X2 inst_8119 ( .A(net_8049), .Z(net_8081) );
CLKBUF_X2 inst_10202 ( .A(net_8123), .Z(net_10164) );
OAI22_X2 inst_1492 ( .B1(net_4666), .A1(net_4132), .B2(net_4120), .ZN(net_4117), .A2(net_4116) );
SDFF_X2 inst_181 ( .Q(net_6273), .SI(net_6272), .D(net_3509), .SE(net_392), .CK(net_13926) );
CLKBUF_X2 inst_13212 ( .A(net_13173), .Z(net_13174) );
CLKBUF_X2 inst_8964 ( .A(net_8925), .Z(net_8926) );
CLKBUF_X2 inst_8329 ( .A(net_8290), .Z(net_8291) );
INV_X4 inst_5215 ( .ZN(net_1730), .A(net_894) );
NAND2_X1 inst_4234 ( .ZN(net_4693), .A2(net_3989), .A1(net_2141) );
DFF_X1 inst_6722 ( .QN(net_7346), .D(net_5334), .CK(net_12702) );
CLKBUF_X2 inst_11982 ( .A(net_11943), .Z(net_11944) );
CLKBUF_X2 inst_10885 ( .A(net_10846), .Z(net_10847) );
CLKBUF_X2 inst_9738 ( .A(net_8955), .Z(net_9700) );
SDFF_X2 inst_713 ( .SI(net_6786), .Q(net_6786), .SE(net_3872), .D(net_3788), .CK(net_11137) );
CLKBUF_X2 inst_10125 ( .A(net_9172), .Z(net_10087) );
NAND2_X4 inst_2898 ( .A1(net_5892), .ZN(net_3401), .A2(net_589) );
DFF_X1 inst_6918 ( .D(net_2409), .Q(net_253), .CK(net_13271) );
CLKBUF_X2 inst_10280 ( .A(net_10241), .Z(net_10242) );
CLKBUF_X2 inst_8875 ( .A(net_8836), .Z(net_8837) );
CLKBUF_X2 inst_11508 ( .A(net_11469), .Z(net_11470) );
OR2_X4 inst_1368 ( .ZN(net_3977), .A2(net_3739), .A1(net_682) );
CLKBUF_X2 inst_13708 ( .A(net_13669), .Z(net_13670) );
AOI22_X2 inst_7282 ( .B1(net_7219), .A1(net_7187), .A2(net_5244), .B2(net_5243), .ZN(net_5239) );
DFF_X1 inst_6775 ( .QN(net_6064), .D(net_4320), .CK(net_8736) );
OAI21_X2 inst_2088 ( .B1(net_5912), .B2(net_4415), .ZN(net_4400), .A(net_3480) );
AOI21_X2 inst_7768 ( .B1(net_7149), .ZN(net_4035), .B2(net_2582), .A(net_2319) );
CLKBUF_X2 inst_14062 ( .A(net_14023), .Z(net_14024) );
NAND2_X2 inst_3208 ( .ZN(net_4718), .A2(net_3986), .A1(net_1887) );
AOI22_X2 inst_7410 ( .B1(net_5939), .A2(net_2838), .ZN(net_2825), .A1(net_750), .B2(net_205) );
DFF_X1 inst_6673 ( .QN(net_7269), .D(net_5156), .CK(net_9889) );
NAND2_X2 inst_4134 ( .A2(net_1228), .ZN(net_1165), .A1(net_380) );
NAND2_X2 inst_3507 ( .ZN(net_2560), .A2(net_2206), .A1(net_1495) );
OR2_X4 inst_1379 ( .ZN(net_4008), .A2(net_3442), .A1(net_3255) );
SDFF_X2 inst_271 ( .Q(net_6367), .SI(net_6366), .D(net_3554), .SE(net_392), .CK(net_13613) );
CLKBUF_X2 inst_11918 ( .A(net_7891), .Z(net_11880) );
CLKBUF_X2 inst_12326 ( .A(net_9312), .Z(net_12288) );
CLKBUF_X2 inst_9582 ( .A(net_9543), .Z(net_9544) );
DFF_X1 inst_6705 ( .QN(net_7288), .D(net_5370), .CK(net_12990) );
SDFF_X2 inst_1230 ( .SI(net_7197), .Q(net_7197), .D(net_3802), .SE(net_3750), .CK(net_10477) );
CLKBUF_X2 inst_10844 ( .A(net_10805), .Z(net_10806) );
AOI21_X2 inst_7691 ( .B1(net_6736), .ZN(net_4135), .B2(net_2581), .A(net_2373) );
AOI22_X2 inst_7262 ( .B1(net_6953), .A1(net_6921), .A2(net_5298), .B2(net_5297), .ZN(net_5292) );
NAND2_X2 inst_3535 ( .ZN(net_2532), .A2(net_2191), .A1(net_1359) );
CLKBUF_X2 inst_12217 ( .A(net_12178), .Z(net_12179) );
CLKBUF_X2 inst_9344 ( .A(net_9305), .Z(net_9306) );
CLKBUF_X2 inst_9221 ( .A(net_9028), .Z(net_9183) );
NAND2_X2 inst_3497 ( .ZN(net_3937), .A2(net_2644), .A1(net_1702) );
INV_X16 inst_6131 ( .ZN(net_4415), .A(net_3838) );
SDFF_X2 inst_1064 ( .Q(net_6736), .D(net_6736), .SI(net_3894), .SE(net_3815), .CK(net_11085) );
INV_X4 inst_5416 ( .ZN(net_517), .A(net_276) );
CLKBUF_X2 inst_13643 ( .A(net_13604), .Z(net_13605) );
CLKBUF_X2 inst_14229 ( .A(net_14190), .Z(net_14191) );
CLKBUF_X2 inst_11110 ( .A(net_11071), .Z(net_11072) );
INV_X2 inst_5796 ( .ZN(net_2229), .A(net_2228) );
NAND2_X2 inst_3599 ( .ZN(net_2401), .A2(net_1874), .A1(net_1321) );
CLKBUF_X2 inst_14335 ( .A(net_8490), .Z(net_14297) );
CLKBUF_X2 inst_9571 ( .A(net_9532), .Z(net_9533) );
CLKBUF_X2 inst_13727 ( .A(net_13688), .Z(net_13689) );
SDFF_X2 inst_583 ( .Q(net_6581), .D(net_6581), .SE(net_3823), .SI(net_3804), .CK(net_9186) );
CLKBUF_X2 inst_12124 ( .A(net_12085), .Z(net_12086) );
OAI21_X2 inst_1904 ( .B1(net_5361), .ZN(net_5165), .A(net_4765), .B2(net_3941) );
CLKBUF_X2 inst_13970 ( .A(net_13931), .Z(net_13932) );
INV_X4 inst_5208 ( .ZN(net_3167), .A(net_558) );
NAND2_X2 inst_3581 ( .ZN(net_2430), .A2(net_2429), .A1(net_880) );
CLKBUF_X2 inst_10732 ( .A(net_10693), .Z(net_10694) );
CLKBUF_X2 inst_9930 ( .A(net_9891), .Z(net_9892) );
CLKBUF_X2 inst_14146 ( .A(net_14107), .Z(net_14108) );
CLKBUF_X2 inst_10932 ( .A(net_10893), .Z(net_10894) );
NAND2_X1 inst_4325 ( .ZN(net_4539), .A2(net_3870), .A1(net_1413) );
CLKBUF_X2 inst_10441 ( .A(net_10402), .Z(net_10403) );
INV_X4 inst_4833 ( .ZN(net_3053), .A(net_1076) );
OAI21_X2 inst_2065 ( .B2(net_4436), .ZN(net_4430), .B1(net_4051), .A(net_3545) );
CLKBUF_X2 inst_10765 ( .A(net_10726), .Z(net_10727) );
NOR2_X4 inst_2251 ( .ZN(net_5635), .A1(net_5481), .A2(net_4441) );
NAND2_X2 inst_3987 ( .ZN(net_1283), .A1(net_885), .A2(net_316) );
DFF_X1 inst_6913 ( .Q(net_6055), .D(net_2385), .CK(net_14373) );
CLKBUF_X2 inst_12825 ( .A(net_12786), .Z(net_12787) );
CLKBUF_X2 inst_13720 ( .A(net_13681), .Z(net_13682) );
DFF_X1 inst_6788 ( .D(net_3946), .CK(net_9571), .Q(x744) );
INV_X4 inst_5124 ( .ZN(net_593), .A(net_592) );
CLKBUF_X2 inst_14346 ( .A(net_11756), .Z(net_14308) );
AOI21_X2 inst_7709 ( .B1(net_6868), .ZN(net_4498), .B2(net_2579), .A(net_2354) );
CLKBUF_X2 inst_13226 ( .A(net_13187), .Z(net_13188) );
INV_X4 inst_4863 ( .A(net_3046), .ZN(net_1076) );
CLKBUF_X2 inst_12513 ( .A(net_10145), .Z(net_12475) );
INV_X4 inst_4910 ( .ZN(net_864), .A(net_863) );
OAI21_X2 inst_1899 ( .B1(net_5200), .ZN(net_5177), .A(net_4554), .B2(net_3866) );
CLKBUF_X2 inst_9349 ( .A(net_8920), .Z(net_9311) );
CLKBUF_X2 inst_12113 ( .A(net_12074), .Z(net_12075) );
NAND3_X4 inst_2569 ( .ZN(net_4596), .A3(net_1664), .A1(net_1229), .A2(net_1050) );
CLKBUF_X2 inst_10573 ( .A(net_10534), .Z(net_10535) );
CLKBUF_X2 inst_9811 ( .A(net_9772), .Z(net_9773) );
CLKBUF_X2 inst_10197 ( .A(net_10158), .Z(net_10159) );
CLKBUF_X2 inst_9048 ( .A(net_9009), .Z(net_9010) );
NAND3_X2 inst_2716 ( .ZN(net_2460), .A2(net_1816), .A3(net_1583), .A1(net_1481) );
CLKBUF_X2 inst_8693 ( .A(net_8444), .Z(net_8655) );
INV_X2 inst_6025 ( .A(net_7286), .ZN(net_2214) );
NAND2_X2 inst_3228 ( .ZN(net_4527), .A2(net_4294), .A1(net_1735) );
CLKBUF_X2 inst_9212 ( .A(net_9173), .Z(net_9174) );
OAI21_X2 inst_2124 ( .B1(net_3265), .B2(net_3087), .ZN(net_3063), .A(net_2914) );
CLKBUF_X2 inst_13268 ( .A(net_13229), .Z(net_13230) );
NOR2_X4 inst_2289 ( .A2(net_7791), .ZN(net_2870), .A1(net_800) );
OAI22_X2 inst_1435 ( .B1(net_5854), .ZN(net_5794), .A2(net_5784), .B2(net_5783), .A1(net_5770) );
CLKBUF_X2 inst_11582 ( .A(net_11543), .Z(net_11544) );
NAND2_X2 inst_3746 ( .A1(net_6491), .A2(net_1642), .ZN(net_1599) );
CLKBUF_X2 inst_12288 ( .A(net_12249), .Z(net_12250) );
NAND3_X2 inst_2750 ( .ZN(net_2351), .A3(net_1542), .A1(net_1329), .A2(net_1006) );
CLKBUF_X2 inst_10810 ( .A(net_10771), .Z(net_10772) );
NAND2_X2 inst_4121 ( .A2(net_1228), .ZN(net_1174), .A1(net_382) );
INV_X2 inst_5800 ( .ZN(net_1924), .A(net_228) );
OAI22_X2 inst_1467 ( .B2(net_5057), .ZN(net_4395), .A1(net_4139), .A2(net_3826), .B1(net_1172) );
NAND3_X2 inst_2640 ( .ZN(net_5689), .A1(net_5666), .A2(net_5294), .A3(net_4240) );
CLKBUF_X2 inst_14313 ( .A(net_14274), .Z(net_14275) );
CLKBUF_X2 inst_10258 ( .A(net_10219), .Z(net_10220) );
INV_X2 inst_5772 ( .ZN(net_2981), .A(net_2980) );
CLKBUF_X2 inst_12732 ( .A(net_12693), .Z(net_12694) );
CLKBUF_X2 inst_8162 ( .A(net_8014), .Z(net_8124) );
CLKBUF_X2 inst_7908 ( .A(net_7869), .Z(net_7870) );
CLKBUF_X2 inst_10803 ( .A(net_10764), .Z(net_10765) );
NAND2_X1 inst_4448 ( .A2(net_1256), .ZN(net_1134), .A1(net_1133) );
CLKBUF_X2 inst_14102 ( .A(net_14063), .Z(net_14064) );
CLKBUF_X2 inst_13227 ( .A(net_13188), .Z(net_13189) );
DFF_X2 inst_6317 ( .QN(net_7797), .CK(net_10945), .D(x1564) );
NAND2_X4 inst_2834 ( .ZN(net_5559), .A1(net_5030), .A2(net_5029) );
INV_X4 inst_4784 ( .ZN(net_2638), .A(net_1659) );
CLKBUF_X2 inst_8130 ( .A(net_8091), .Z(net_8092) );
CLKBUF_X2 inst_12256 ( .A(net_12217), .Z(net_12218) );
OAI22_X2 inst_1513 ( .B1(net_4650), .A1(net_4080), .B2(net_4074), .ZN(net_4071), .A2(net_4070) );
CLKBUF_X2 inst_9864 ( .A(net_9825), .Z(net_9826) );
CLKBUF_X2 inst_11756 ( .A(net_11717), .Z(net_11718) );
CLKBUF_X2 inst_10916 ( .A(net_10877), .Z(net_10878) );
NAND2_X2 inst_3321 ( .ZN(net_3604), .A1(net_3603), .A2(net_3228) );
NAND2_X2 inst_4080 ( .A1(net_6526), .A2(net_1645), .ZN(net_972) );
CLKBUF_X2 inst_10846 ( .A(net_10807), .Z(net_10808) );
AOI21_X2 inst_7667 ( .ZN(net_3010), .B1(net_2857), .B2(net_2742), .A(net_933) );
CLKBUF_X2 inst_12750 ( .A(net_12711), .Z(net_12712) );
OAI22_X2 inst_1545 ( .B2(net_3405), .ZN(net_3361), .A2(net_3360), .A1(net_3268), .B1(net_456) );
SDFF_X2 inst_333 ( .D(net_6393), .SE(net_5799), .SI(net_378), .Q(net_378), .CK(net_13899) );
NAND2_X2 inst_3338 ( .ZN(net_3570), .A2(net_3225), .A1(net_2700) );
AOI21_X2 inst_7684 ( .B1(net_7010), .ZN(net_4225), .A(net_2465), .B2(net_1100) );
INV_X2 inst_5988 ( .ZN(net_1133), .A(net_114) );
CLKBUF_X2 inst_8368 ( .A(net_8329), .Z(net_8330) );
INV_X4 inst_5279 ( .A(net_7261), .ZN(net_2015) );
SDFF_X2 inst_406 ( .SI(net_7370), .Q(net_7370), .D(net_4780), .SE(net_3853), .CK(net_9398) );
CLKBUF_X2 inst_11934 ( .A(net_8704), .Z(net_11896) );
INV_X2 inst_5933 ( .A(net_7332), .ZN(net_1781) );
INV_X4 inst_4579 ( .ZN(net_5494), .A(net_5493) );
CLKBUF_X2 inst_13818 ( .A(net_13779), .Z(net_13780) );
SDFF_X2 inst_328 ( .SI(net_7493), .Q(net_7493), .D(net_5100), .SE(net_3989), .CK(net_12442) );
CLKBUF_X2 inst_11394 ( .A(net_8612), .Z(net_11356) );
CLKBUF_X2 inst_9335 ( .A(net_8280), .Z(net_9297) );
CLKBUF_X2 inst_10953 ( .A(net_9249), .Z(net_10915) );
CLKBUF_X2 inst_10897 ( .A(net_10858), .Z(net_10859) );
NAND2_X1 inst_4217 ( .ZN(net_4743), .A2(net_3988), .A1(net_2069) );
NAND3_X2 inst_2764 ( .ZN(net_2337), .A3(net_1547), .A1(net_1515), .A2(net_1003) );
CLKBUF_X2 inst_8496 ( .A(net_8457), .Z(net_8458) );
SDFF_X2 inst_818 ( .Q(net_6993), .D(net_6993), .SE(net_3891), .SI(net_3821), .CK(net_11014) );
CLKBUF_X2 inst_12373 ( .A(net_12334), .Z(net_12335) );
DFF_X2 inst_6246 ( .QN(net_7749), .D(net_3029), .CK(net_7931) );
CLKBUF_X2 inst_13755 ( .A(net_9829), .Z(net_13717) );
CLKBUF_X2 inst_11065 ( .A(net_11026), .Z(net_11027) );
INV_X1 inst_6155 ( .A(net_5852), .ZN(x84) );
INV_X2 inst_5774 ( .ZN(net_2917), .A(net_2852) );
CLKBUF_X2 inst_9664 ( .A(net_9625), .Z(net_9626) );
CLKBUF_X2 inst_8719 ( .A(net_7840), .Z(net_8681) );
CLKBUF_X2 inst_9902 ( .A(net_9725), .Z(net_9864) );
CLKBUF_X2 inst_11610 ( .A(net_8849), .Z(net_11572) );
CLKBUF_X2 inst_9825 ( .A(net_8821), .Z(net_9787) );
AOI222_X2 inst_7561 ( .ZN(net_5432), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_365), .C2(net_363), .A1(net_351) );
CLKBUF_X2 inst_10172 ( .A(net_8820), .Z(net_10134) );
NAND2_X2 inst_3178 ( .ZN(net_4755), .A2(net_3941), .A1(net_2087) );
NAND2_X2 inst_3274 ( .ZN(net_3698), .A1(net_3697), .A2(net_3231) );
CLKBUF_X2 inst_13920 ( .A(net_13881), .Z(net_13882) );
NAND2_X2 inst_4203 ( .A2(net_5988), .ZN(net_1737), .A1(net_573) );
CLKBUF_X2 inst_11776 ( .A(net_11737), .Z(net_11738) );
CLKBUF_X2 inst_12643 ( .A(net_11659), .Z(net_12605) );
CLKBUF_X2 inst_9972 ( .A(net_9933), .Z(net_9934) );
NAND2_X4 inst_2840 ( .ZN(net_5544), .A1(net_5018), .A2(net_5017) );
CLKBUF_X2 inst_12521 ( .A(net_12482), .Z(net_12483) );
CLKBUF_X2 inst_10939 ( .A(net_10900), .Z(net_10901) );
CLKBUF_X2 inst_9178 ( .A(net_9139), .Z(net_9140) );
CLKBUF_X2 inst_10066 ( .A(net_10027), .Z(net_10028) );
CLKBUF_X2 inst_14214 ( .A(net_12658), .Z(net_14176) );
CLKBUF_X2 inst_8360 ( .A(net_8309), .Z(net_8322) );
NAND3_X2 inst_2781 ( .ZN(net_2319), .A3(net_1610), .A1(net_1447), .A2(net_962) );
CLKBUF_X2 inst_9544 ( .A(net_9505), .Z(net_9506) );
DFF_X1 inst_6442 ( .QN(net_6073), .D(net_5728), .CK(net_10889) );
CLKBUF_X2 inst_13190 ( .A(net_12125), .Z(net_13152) );
SDFF_X2 inst_906 ( .Q(net_7142), .D(net_7142), .SE(net_3903), .SI(net_3813), .CK(net_7863) );
NAND2_X1 inst_4276 ( .ZN(net_4592), .A2(net_3867), .A1(net_1907) );
INV_X4 inst_5222 ( .ZN(net_470), .A(net_469) );
CLKBUF_X2 inst_13600 ( .A(net_13561), .Z(net_13562) );
INV_X4 inst_5098 ( .ZN(net_748), .A(net_620) );
CLKBUF_X2 inst_11043 ( .A(net_8412), .Z(net_11005) );
SDFF_X2 inst_1248 ( .SI(net_6544), .Q(net_6544), .D(net_3796), .SE(net_3755), .CK(net_11625) );
NAND3_X2 inst_2598 ( .ZN(net_5741), .A1(net_5636), .A2(net_5211), .A3(net_4200) );
CLKBUF_X2 inst_12780 ( .A(net_9591), .Z(net_12742) );
NOR2_X2 inst_2402 ( .ZN(net_3768), .A1(net_3767), .A2(net_3766) );
CLKBUF_X2 inst_8877 ( .A(net_8838), .Z(net_8839) );
NAND3_X2 inst_2616 ( .ZN(net_5723), .A1(net_5618), .A2(net_5135), .A3(net_4182) );
CLKBUF_X2 inst_8095 ( .A(net_8056), .Z(net_8057) );
NAND2_X2 inst_3998 ( .A2(net_1910), .ZN(net_1187), .A1(net_1186) );
CLKBUF_X2 inst_9035 ( .A(net_8996), .Z(net_8997) );
NAND2_X1 inst_4300 ( .ZN(net_4566), .A2(net_3866), .A1(net_1850) );
OAI21_X2 inst_2113 ( .ZN(net_3397), .B1(net_3321), .B2(net_2749), .A(net_543) );
CLKBUF_X2 inst_12000 ( .A(net_9371), .Z(net_11962) );
AOI21_X2 inst_7645 ( .B1(net_5891), .ZN(net_3906), .B2(net_3905), .A(net_2607) );
INV_X4 inst_5249 ( .ZN(net_443), .A(net_442) );
OAI21_X2 inst_1820 ( .ZN(net_5368), .B1(net_5337), .A(net_4335), .B2(net_3859) );
SDFF_X2 inst_183 ( .Q(net_6271), .SI(net_6270), .D(net_3513), .SE(net_392), .CK(net_13920) );
CLKBUF_X2 inst_8253 ( .A(net_8087), .Z(net_8215) );
DFFR_X2 inst_6998 ( .QN(net_7692), .D(net_3354), .CK(net_10358), .RN(x1822) );
AOI21_X2 inst_7748 ( .B1(net_6592), .ZN(net_4403), .B2(net_2583), .A(net_2282) );
DFF_X1 inst_6703 ( .QN(net_7286), .D(net_5372), .CK(net_10168) );
CLKBUF_X2 inst_8471 ( .A(net_8425), .Z(net_8433) );
INV_X2 inst_6065 ( .ZN(net_3082), .A(net_284) );
INV_X4 inst_4729 ( .A(net_3200), .ZN(net_3193) );
NOR2_X4 inst_2271 ( .ZN(net_5615), .A1(net_5460), .A2(net_4409) );
DFF_X2 inst_6209 ( .QN(net_7382), .D(net_4299), .CK(net_9522) );
AND4_X2 inst_7793 ( .ZN(net_2487), .A4(net_2486), .A2(net_1219), .A1(x1126), .A3(x1101) );
CLKBUF_X2 inst_10314 ( .A(net_10275), .Z(net_10276) );
CLKBUF_X2 inst_8081 ( .A(net_8042), .Z(net_8043) );
NAND2_X2 inst_3779 ( .A1(net_6910), .A2(net_1639), .ZN(net_1566) );
OAI21_X2 inst_1848 ( .B1(net_5345), .ZN(net_5324), .A(net_4384), .B2(net_3853) );
CLKBUF_X2 inst_12694 ( .A(net_12655), .Z(net_12656) );
NAND2_X1 inst_4451 ( .A2(net_1256), .ZN(net_1128), .A1(net_1127) );
CLKBUF_X2 inst_11644 ( .A(net_11605), .Z(net_11606) );
SDFF_X2 inst_697 ( .SI(net_7802), .Q(net_6735), .D(net_6735), .SE(net_3815), .CK(net_11096) );
CLKBUF_X2 inst_11150 ( .A(net_11111), .Z(net_11112) );
CLKBUF_X2 inst_14035 ( .A(net_13996), .Z(net_13997) );
SDFF_X2 inst_487 ( .D(net_7807), .SI(net_6502), .Q(net_6502), .SE(net_3889), .CK(net_8669) );
INV_X4 inst_5159 ( .A(net_713), .ZN(net_554) );
CLKBUF_X2 inst_11338 ( .A(net_11299), .Z(net_11300) );
CLKBUF_X2 inst_10350 ( .A(net_10311), .Z(net_10312) );
AOI222_X2 inst_7527 ( .C1(net_7524), .B1(net_7492), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_1984), .A1(net_1983) );
CLKBUF_X2 inst_13941 ( .A(net_13902), .Z(net_13903) );
INV_X4 inst_5315 ( .A(net_7504), .ZN(net_2105) );
CLKBUF_X2 inst_11512 ( .A(net_11473), .Z(net_11474) );
CLKBUF_X2 inst_13696 ( .A(net_13657), .Z(net_13658) );
OAI21_X2 inst_2133 ( .A(net_5920), .ZN(net_2900), .B1(net_2899), .B2(net_2898) );
OAI211_X2 inst_2163 ( .ZN(net_3376), .C1(net_3341), .C2(net_3089), .B(net_2842), .A(net_2775) );
CLKBUF_X2 inst_12307 ( .A(net_12268), .Z(net_12269) );
CLKBUF_X2 inst_9947 ( .A(net_9653), .Z(net_9909) );
INV_X2 inst_6051 ( .A(net_7301), .ZN(net_2041) );
INV_X4 inst_4668 ( .ZN(net_4007), .A(net_3732) );
CLKBUF_X2 inst_8758 ( .A(net_8719), .Z(net_8720) );
CLKBUF_X2 inst_12975 ( .A(net_12936), .Z(net_12937) );
INV_X4 inst_5497 ( .A(net_5984), .ZN(net_589) );
CLKBUF_X2 inst_13972 ( .A(net_11525), .Z(net_13934) );
OAI21_X2 inst_1861 ( .ZN(net_5256), .B1(net_5222), .A(net_4542), .B2(net_3870) );
NAND2_X2 inst_3570 ( .ZN(net_2497), .A2(net_1994), .A1(net_1789) );
CLKBUF_X2 inst_9133 ( .A(net_9094), .Z(net_9095) );
CLKBUF_X2 inst_14198 ( .A(net_14159), .Z(net_14160) );
AOI222_X2 inst_7598 ( .A1(net_7538), .ZN(net_4847), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_370), .C2(net_368) );
INV_X4 inst_4835 ( .ZN(net_4790), .A(net_1075) );
OAI21_X2 inst_2004 ( .B2(net_4518), .ZN(net_4509), .B1(net_4508), .A(net_3680) );
CLKBUF_X2 inst_8667 ( .A(net_8628), .Z(net_8629) );
NAND2_X4 inst_2857 ( .A1(net_5888), .ZN(net_5084), .A2(net_4149) );
SDFF_X2 inst_220 ( .Q(net_6334), .SI(net_6333), .D(net_3657), .SE(net_392), .CK(net_14051) );
OAI22_X2 inst_1585 ( .B2(net_3200), .A2(net_3193), .ZN(net_3191), .A1(net_3190), .B1(net_553) );
CLKBUF_X2 inst_11412 ( .A(net_11373), .Z(net_11374) );
CLKBUF_X2 inst_10754 ( .A(net_10715), .Z(net_10716) );
SDFF_X2 inst_245 ( .Q(net_6349), .SI(net_6348), .D(net_3579), .SE(net_392), .CK(net_14133) );
DFFR_X2 inst_6991 ( .QN(net_7706), .D(net_3356), .CK(net_13227), .RN(x1822) );
CLKBUF_X2 inst_11965 ( .A(net_11926), .Z(net_11927) );
CLKBUF_X2 inst_9779 ( .A(net_9740), .Z(net_9741) );
OAI21_X2 inst_1873 ( .ZN(net_5233), .B1(net_5232), .A(net_4589), .B2(net_3867) );
NAND2_X2 inst_4111 ( .A1(net_6657), .A2(net_1655), .ZN(net_941) );
CLKBUF_X2 inst_8388 ( .A(net_8163), .Z(net_8350) );
CLKBUF_X2 inst_8768 ( .A(net_8303), .Z(net_8730) );
AND2_X2 inst_7854 ( .ZN(net_3038), .A1(net_2936), .A2(net_2827) );
SDFF_X2 inst_147 ( .Q(net_6231), .SI(net_6230), .SE(net_392), .D(net_137), .CK(net_14110) );
INV_X16 inst_6135 ( .ZN(net_2957), .A(net_2625) );
SDFF_X2 inst_313 ( .SI(net_7455), .Q(net_7455), .D(net_5105), .SE(net_3993), .CK(net_12585) );
OAI221_X2 inst_1676 ( .C1(net_5940), .ZN(net_3939), .B2(net_3937), .A(net_3731), .B1(net_3055), .C2(net_201) );
NAND2_X2 inst_4170 ( .A2(net_6688), .ZN(net_813), .A1(net_471) );
CLKBUF_X2 inst_11765 ( .A(net_8030), .Z(net_11727) );
CLKBUF_X2 inst_8480 ( .A(net_8441), .Z(net_8442) );
SDFF_X2 inst_1041 ( .Q(net_7545), .D(net_7545), .SE(net_3896), .SI(net_379), .CK(net_13101) );
INV_X4 inst_5263 ( .ZN(net_662), .A(net_427) );
OAI21_X2 inst_2086 ( .B1(net_5902), .B2(net_4415), .ZN(net_4402), .A(net_3482) );
NAND2_X2 inst_3114 ( .A1(net_6587), .A2(net_4897), .ZN(net_4887) );
NAND2_X2 inst_3577 ( .ZN(net_2458), .A2(net_1974), .A1(net_1356) );
CLKBUF_X2 inst_9451 ( .A(net_9412), .Z(net_9413) );
CLKBUF_X2 inst_12918 ( .A(net_12151), .Z(net_12880) );
CLKBUF_X2 inst_8743 ( .A(net_7903), .Z(net_8705) );
CLKBUF_X2 inst_8570 ( .A(net_8201), .Z(net_8532) );
CLKBUF_X2 inst_8195 ( .A(net_8156), .Z(net_8157) );
CLKBUF_X2 inst_12789 ( .A(net_8793), .Z(net_12751) );
INV_X4 inst_4754 ( .ZN(net_2724), .A(x38) );
SDFF_X2 inst_553 ( .Q(net_6449), .D(net_6449), .SI(net_3898), .SE(net_3820), .CK(net_8423) );
CLKBUF_X2 inst_9271 ( .A(net_7991), .Z(net_9233) );
CLKBUF_X2 inst_10216 ( .A(net_10177), .Z(net_10178) );
NAND2_X2 inst_3331 ( .ZN(net_3584), .A1(net_3583), .A2(net_3228) );
CLKBUF_X2 inst_11554 ( .A(net_11515), .Z(net_11516) );
SDFF_X2 inst_242 ( .Q(net_6352), .SI(net_6351), .D(net_3609), .SE(net_392), .CK(net_13503) );
DFF_X1 inst_6589 ( .QN(net_7559), .D(net_5061), .CK(net_13451) );
INV_X4 inst_4680 ( .ZN(net_3383), .A(net_3382) );
CLKBUF_X2 inst_8950 ( .A(net_8911), .Z(net_8912) );
SDFF_X2 inst_1186 ( .D(net_7799), .SI(net_6931), .Q(net_6931), .SE(net_3734), .CK(net_11772) );
OAI21_X2 inst_1753 ( .ZN(net_5480), .A(net_4806), .B2(net_4805), .B1(net_4304) );
OAI21_X2 inst_1727 ( .ZN(net_5567), .B1(net_5436), .A(net_4832), .B2(net_4153) );
CLKBUF_X2 inst_9513 ( .A(net_9474), .Z(net_9475) );
CLKBUF_X2 inst_10542 ( .A(net_9362), .Z(net_10504) );
SDFF_X2 inst_1166 ( .SI(net_6935), .Q(net_6935), .D(net_3894), .SE(net_3734), .CK(net_11777) );
OAI21_X2 inst_1739 ( .ZN(net_5540), .B1(net_5539), .A(net_4808), .B2(net_4153) );
XNOR2_X2 inst_116 ( .A(net_2569), .ZN(net_817), .B(net_816) );
CLKBUF_X2 inst_13712 ( .A(net_7881), .Z(net_13674) );
DFF_X1 inst_6559 ( .QN(net_7452), .D(net_5047), .CK(net_9664) );
INV_X4 inst_5498 ( .A(net_7693), .ZN(net_710) );
CLKBUF_X2 inst_10142 ( .A(net_10103), .Z(net_10104) );
CLKBUF_X2 inst_12430 ( .A(net_10251), .Z(net_12392) );
SDFF_X2 inst_471 ( .Q(net_7014), .D(net_7014), .SE(net_3899), .SI(net_3897), .CK(net_11970) );
NAND2_X2 inst_4087 ( .A1(net_7214), .A2(net_1648), .ZN(net_965) );
CLKBUF_X2 inst_10680 ( .A(net_10641), .Z(net_10642) );
INV_X4 inst_5446 ( .A(net_6030), .ZN(net_496) );
CLKBUF_X2 inst_12104 ( .A(net_12065), .Z(net_12066) );
DFF_X1 inst_6557 ( .QN(net_7655), .D(net_5177), .CK(net_10604) );
INV_X4 inst_4956 ( .A(net_1216), .ZN(net_725) );
CLKBUF_X2 inst_11081 ( .A(net_10203), .Z(net_11043) );
NAND2_X2 inst_3609 ( .ZN(net_2387), .A2(net_1863), .A1(net_1345) );
SDFF_X2 inst_896 ( .Q(net_7128), .D(net_7128), .SE(net_3888), .SI(net_3821), .CK(net_8714) );
CLKBUF_X2 inst_8619 ( .A(net_8501), .Z(net_8581) );
CLKBUF_X2 inst_12315 ( .A(net_12276), .Z(net_12277) );
DFF_X1 inst_6649 ( .QN(net_7624), .D(net_5199), .CK(net_13151) );
CLKBUF_X2 inst_13338 ( .A(net_13299), .Z(net_13300) );
CLKBUF_X2 inst_9276 ( .A(net_9237), .Z(net_9238) );
CLKBUF_X2 inst_8221 ( .A(net_7849), .Z(net_8183) );
NAND3_X2 inst_2608 ( .ZN(net_5731), .A1(net_5626), .A2(net_5169), .A3(net_4191) );
INV_X2 inst_6008 ( .A(net_7656), .ZN(net_1840) );
CLKBUF_X2 inst_9317 ( .A(net_8268), .Z(net_9279) );
CLKBUF_X2 inst_11840 ( .A(net_11801), .Z(net_11802) );
AOI22_X2 inst_7445 ( .A2(net_2667), .B2(net_2650), .ZN(net_857), .A1(net_856), .B1(net_855) );
CLKBUF_X2 inst_12659 ( .A(net_12620), .Z(net_12621) );
CLKBUF_X2 inst_8577 ( .A(net_8538), .Z(net_8539) );
AOI22_X2 inst_7438 ( .ZN(net_4853), .A2(net_1228), .B1(net_1226), .B2(net_384), .A1(net_372) );
NAND4_X2 inst_2557 ( .ZN(net_3301), .A4(net_2977), .A2(net_2780), .A1(net_2756), .A3(net_2755) );
NOR2_X2 inst_2521 ( .ZN(net_1698), .A2(net_899), .A1(net_641) );
SDFF_X2 inst_385 ( .SI(net_7304), .Q(net_7304), .D(net_4782), .SE(net_3859), .CK(net_9927) );
NAND2_X2 inst_3319 ( .ZN(net_3608), .A1(net_3607), .A2(net_3226) );
CLKBUF_X2 inst_14110 ( .A(net_14071), .Z(net_14072) );
NAND3_X2 inst_2653 ( .ZN(net_3947), .A3(net_3398), .A2(net_2956), .A1(net_2837) );
CLKBUF_X2 inst_11062 ( .A(net_11023), .Z(net_11024) );
INV_X4 inst_4621 ( .ZN(net_4201), .A(net_4063) );
CLKBUF_X2 inst_11519 ( .A(net_11480), .Z(net_11481) );
CLKBUF_X2 inst_11324 ( .A(net_11285), .Z(net_11286) );
NOR2_X2 inst_2550 ( .A2(net_6413), .ZN(net_614), .A1(net_403) );
CLKBUF_X2 inst_10696 ( .A(net_8000), .Z(net_10658) );
CLKBUF_X2 inst_13150 ( .A(net_7855), .Z(net_13112) );
AOI222_X2 inst_7559 ( .A1(net_7391), .ZN(net_5545), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_354), .C2(net_352) );
NAND2_X1 inst_4281 ( .ZN(net_4586), .A2(net_3867), .A1(net_1899) );
SDFF_X2 inst_596 ( .Q(net_6567), .D(net_6567), .SE(net_3823), .SI(net_3814), .CK(net_12915) );
NAND3_X2 inst_2771 ( .ZN(net_2329), .A3(net_1537), .A1(net_1332), .A2(net_948) );
CLKBUF_X2 inst_8835 ( .A(net_8486), .Z(net_8797) );
INV_X4 inst_4687 ( .ZN(net_3736), .A(net_3364) );
OAI21_X2 inst_2142 ( .B1(net_5778), .ZN(net_2802), .A(net_2683), .B2(net_2681) );
CLKBUF_X2 inst_9245 ( .A(net_9206), .Z(net_9207) );
CLKBUF_X2 inst_12810 ( .A(net_12771), .Z(net_12772) );
OAI21_X2 inst_1705 ( .ZN(net_5589), .A(net_5212), .B2(net_4458), .B1(net_4080) );
CLKBUF_X2 inst_11286 ( .A(net_11247), .Z(net_11248) );
INV_X4 inst_5110 ( .A(net_848), .ZN(net_610) );
INV_X4 inst_4664 ( .A(net_4168), .ZN(net_3868) );
DFF_X1 inst_6817 ( .D(net_3157), .CK(net_10818), .Q(x234) );
INV_X4 inst_5003 ( .A(net_7817), .ZN(net_3779) );
NAND2_X1 inst_4458 ( .A2(net_1256), .ZN(net_1114), .A1(net_1113) );
CLKBUF_X2 inst_12215 ( .A(net_12176), .Z(net_12177) );
CLKBUF_X2 inst_9407 ( .A(net_9368), .Z(net_9369) );
INV_X2 inst_5798 ( .ZN(net_2225), .A(net_2224) );
NAND2_X2 inst_3253 ( .ZN(net_3929), .A2(net_3472), .A1(net_1727) );
INV_X4 inst_5321 ( .A(net_5999), .ZN(net_601) );
CLKBUF_X2 inst_14250 ( .A(net_14211), .Z(net_14212) );
CLKBUF_X2 inst_14055 ( .A(net_12742), .Z(net_14017) );
CLKBUF_X2 inst_10518 ( .A(net_9370), .Z(net_10480) );
INV_X4 inst_5184 ( .ZN(net_634), .A(net_523) );
INV_X4 inst_4596 ( .ZN(net_5075), .A(net_4293) );
CLKBUF_X2 inst_9013 ( .A(net_8974), .Z(net_8975) );
CLKBUF_X2 inst_8427 ( .A(net_8388), .Z(net_8389) );
SDFF_X2 inst_637 ( .SI(net_6650), .Q(net_6650), .SE(net_3850), .D(net_3794), .CK(net_12013) );
SDFF_X2 inst_547 ( .SI(net_6509), .Q(net_6509), .SE(net_3886), .D(net_3836), .CK(net_11673) );
CLKBUF_X2 inst_9107 ( .A(net_9068), .Z(net_9069) );
CLKBUF_X2 inst_13572 ( .A(net_13533), .Z(net_13534) );
OAI22_X2 inst_1607 ( .B2(net_3200), .A2(net_3193), .ZN(net_3126), .B1(net_1718), .A1(net_873) );
CLKBUF_X2 inst_13148 ( .A(net_12363), .Z(net_13110) );
CLKBUF_X2 inst_11847 ( .A(net_8016), .Z(net_11809) );
DFFR_X2 inst_7033 ( .QN(net_6019), .D(net_3191), .CK(net_8595), .RN(x1822) );
CLKBUF_X2 inst_8152 ( .A(net_8004), .Z(net_8114) );
CLKBUF_X2 inst_10159 ( .A(net_10120), .Z(net_10121) );
CLKBUF_X2 inst_10367 ( .A(net_7831), .Z(net_10329) );
INV_X4 inst_4762 ( .ZN(net_2784), .A(net_2772) );
SDFF_X2 inst_164 ( .Q(net_6250), .SI(net_6249), .D(net_3607), .SE(net_392), .CK(net_13983) );
CLKBUF_X2 inst_11623 ( .A(net_11584), .Z(net_11585) );
CLKBUF_X2 inst_8534 ( .A(net_8495), .Z(net_8496) );
CLKBUF_X2 inst_9002 ( .A(net_8963), .Z(net_8964) );
OAI21_X2 inst_1854 ( .ZN(net_5264), .B1(net_5240), .A(net_4549), .B2(net_3870) );
CLKBUF_X2 inst_12676 ( .A(net_12637), .Z(net_12638) );
INV_X2 inst_5922 ( .A(net_7353), .ZN(net_1996) );
OAI21_X2 inst_1710 ( .B2(net_5912), .ZN(net_5584), .A(net_5129), .B1(net_4030) );
AOI22_X2 inst_7295 ( .B1(net_6545), .A1(net_6513), .A2(net_5184), .B2(net_5183), .ZN(net_5176) );
NOR2_X2 inst_2407 ( .ZN(net_3865), .A2(net_3743), .A1(net_2805) );
CLKBUF_X2 inst_13814 ( .A(net_9790), .Z(net_13776) );
CLKBUF_X2 inst_8467 ( .A(net_8428), .Z(net_8429) );
INV_X4 inst_4884 ( .A(net_3807), .ZN(net_3194) );
AOI222_X2 inst_7516 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2022), .A1(net_2021), .B1(net_2020), .C1(net_2019) );
NAND2_X2 inst_3142 ( .ZN(net_4821), .A2(net_4153), .A1(net_2144) );
NOR2_X2 inst_2305 ( .A2(net_6209), .A1(net_5843), .ZN(net_5836) );
SDFF_X2 inst_753 ( .SI(net_7807), .Q(net_6875), .D(net_6875), .SE(net_3901), .CK(net_11482) );
CLKBUF_X2 inst_10079 ( .A(net_10040), .Z(net_10041) );
CLKBUF_X2 inst_9647 ( .A(net_9608), .Z(net_9609) );
OAI21_X2 inst_2150 ( .B1(net_5778), .ZN(net_2794), .A(net_2648), .B2(net_2646) );
INV_X4 inst_5486 ( .A(net_6145), .ZN(net_3593) );
NAND2_X2 inst_3427 ( .ZN(net_3221), .A2(net_3097), .A1(net_2770) );
CLKBUF_X2 inst_10930 ( .A(net_9115), .Z(net_10892) );
DFF_X2 inst_6262 ( .QN(net_5975), .D(net_2731), .CK(net_8559) );
INV_X2 inst_5768 ( .A(net_3256), .ZN(net_3008) );
CLKBUF_X2 inst_9770 ( .A(net_9731), .Z(net_9732) );
DFF_X1 inst_6946 ( .Q(net_6403), .D(net_688), .CK(net_12971) );
SDFF_X2 inst_946 ( .SI(net_7189), .Q(net_7189), .SE(net_3819), .D(net_3795), .CK(net_10637) );
OAI21_X2 inst_1954 ( .ZN(net_5066), .B1(net_4847), .A(net_4713), .B2(net_3986) );
NOR2_X4 inst_2260 ( .ZN(net_5626), .A1(net_5471), .A2(net_4429) );
CLKBUF_X2 inst_8141 ( .A(net_8003), .Z(net_8103) );
CLKBUF_X2 inst_13276 ( .A(net_13237), .Z(net_13238) );
NAND2_X2 inst_3941 ( .A1(net_6429), .A2(net_1677), .ZN(net_1350) );
CLKBUF_X2 inst_13543 ( .A(net_10445), .Z(net_13505) );
AND2_X4 inst_7815 ( .ZN(net_3822), .A2(net_3240), .A1(net_691) );
CLKBUF_X2 inst_12746 ( .A(net_12707), .Z(net_12708) );
CLKBUF_X2 inst_10588 ( .A(net_10549), .Z(net_10550) );
DFFR_X2 inst_7014 ( .D(net_3300), .QN(net_284), .CK(net_12864), .RN(x1822) );
NAND2_X2 inst_3858 ( .A1(net_6834), .A2(net_1521), .ZN(net_1475) );
CLKBUF_X2 inst_13129 ( .A(net_13090), .Z(net_13091) );
CLKBUF_X2 inst_11700 ( .A(net_11661), .Z(net_11662) );
INV_X4 inst_4625 ( .ZN(net_4197), .A(net_4054) );
DFFS_X2 inst_6951 ( .QN(net_6406), .D(net_2723), .CK(net_14405), .SN(x1822) );
NAND2_X2 inst_3922 ( .A1(net_7111), .A2(net_1675), .ZN(net_1380) );
OAI21_X2 inst_2053 ( .B2(net_4457), .ZN(net_4446), .B1(net_4445), .A(net_3572) );
CLKBUF_X2 inst_13949 ( .A(net_13763), .Z(net_13911) );
CLKBUF_X2 inst_10539 ( .A(net_10500), .Z(net_10501) );
CLKBUF_X2 inst_10038 ( .A(net_9393), .Z(net_10000) );
SDFF_X2 inst_1325 ( .D(net_6384), .SE(net_5800), .SI(net_349), .Q(net_349), .CK(net_13656) );
CLKBUF_X2 inst_8859 ( .A(net_8820), .Z(net_8821) );
CLKBUF_X2 inst_13503 ( .A(net_13464), .Z(net_13465) );
CLKBUF_X2 inst_13008 ( .A(net_12969), .Z(net_12970) );
DFF_X1 inst_6873 ( .D(net_2532), .Q(net_202), .CK(net_10059) );
CLKBUF_X2 inst_14087 ( .A(net_14048), .Z(net_14049) );
AOI22_X2 inst_7342 ( .ZN(net_3181), .A2(net_2986), .B2(net_2904), .A1(net_1746), .B1(net_1049) );
CLKBUF_X2 inst_8818 ( .A(net_8779), .Z(net_8780) );
INV_X4 inst_5105 ( .A(net_7812), .ZN(net_3807) );
NAND2_X2 inst_3312 ( .ZN(net_3622), .A1(net_3621), .A2(net_3226) );
CLKBUF_X2 inst_9207 ( .A(net_9168), .Z(net_9169) );
CLKBUF_X2 inst_12725 ( .A(net_12686), .Z(net_12687) );
CLKBUF_X2 inst_12143 ( .A(net_12104), .Z(net_12105) );
SDFF_X2 inst_1235 ( .SI(net_7203), .Q(net_7203), .D(net_3814), .SE(net_3750), .CK(net_10473) );
NAND2_X2 inst_3561 ( .ZN(net_2506), .A2(net_2026), .A1(net_1790) );
CLKBUF_X2 inst_14107 ( .A(net_14068), .Z(net_14069) );
CLKBUF_X2 inst_14286 ( .A(net_8496), .Z(net_14248) );
CLKBUF_X2 inst_13143 ( .A(net_13104), .Z(net_13105) );
NAND2_X2 inst_3046 ( .A1(net_6995), .A2(net_4977), .ZN(net_4961) );
CLKBUF_X2 inst_8751 ( .A(net_7994), .Z(net_8713) );
NAND2_X2 inst_3626 ( .ZN(net_1957), .A1(net_1286), .A2(net_1124) );
NAND2_X2 inst_4036 ( .A1(net_6534), .A2(net_1645), .ZN(net_1016) );
INV_X4 inst_4644 ( .ZN(net_4178), .A(net_4015) );
INV_X4 inst_5244 ( .A(net_495), .ZN(net_446) );
INV_X4 inst_4844 ( .ZN(net_4779), .A(net_1066) );
NAND2_X2 inst_3757 ( .A1(net_6492), .A2(net_1642), .ZN(net_1588) );
SDFF_X2 inst_917 ( .Q(net_7154), .D(net_7154), .SE(net_3903), .SI(net_3782), .CK(net_11571) );
NAND2_X2 inst_3712 ( .A1(net_6764), .A2(net_1635), .ZN(net_1634) );
CLKBUF_X2 inst_13457 ( .A(net_8139), .Z(net_13419) );
OAI21_X2 inst_1743 ( .ZN(net_5530), .A(net_4824), .B2(net_4153), .B1(net_1255) );
CLKBUF_X2 inst_11713 ( .A(net_11674), .Z(net_11675) );
CLKBUF_X2 inst_13403 ( .A(net_13364), .Z(net_13365) );
OAI22_X2 inst_1600 ( .A1(net_3280), .B2(net_3200), .A2(net_3193), .ZN(net_3136), .B1(net_695) );
INV_X4 inst_5022 ( .A(net_1147), .ZN(net_747) );
SDFF_X2 inst_215 ( .Q(net_6339), .SI(net_6338), .D(net_3645), .SE(net_392), .CK(net_14065) );
NAND2_X4 inst_2850 ( .ZN(net_5473), .A1(net_4915), .A2(net_4914) );
CLKBUF_X2 inst_14268 ( .A(net_14229), .Z(net_14230) );
INV_X4 inst_5163 ( .ZN(net_548), .A(net_547) );
NAND3_X2 inst_2624 ( .ZN(net_5705), .A1(net_5682), .A2(net_5318), .A3(net_4256) );
CLKBUF_X2 inst_9590 ( .A(net_9551), .Z(net_9552) );
AOI21_X2 inst_7677 ( .B1(net_7013), .ZN(net_4218), .A(net_2456), .B2(net_1100) );
SDFF_X2 inst_849 ( .Q(net_7001), .D(net_7001), .SE(net_3899), .SI(net_3798), .CK(net_11945) );
AOI22_X2 inst_7393 ( .A2(net_2925), .B2(net_2924), .ZN(net_2875), .A1(net_1156), .B1(net_1142) );
DFF_X2 inst_6258 ( .QN(net_5967), .D(net_2737), .CK(net_9708) );
AOI222_X2 inst_7550 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1853), .A1(net_1852), .B1(net_1851), .C1(net_1850) );
XOR2_X2 inst_3 ( .A(net_2567), .Z(net_1248), .B(net_1247) );
CLKBUF_X2 inst_11293 ( .A(net_11254), .Z(net_11255) );
NAND2_X2 inst_3060 ( .A1(net_7157), .A2(net_4954), .ZN(net_4945) );
INV_X2 inst_5812 ( .ZN(net_1104), .A(net_1103) );
CLKBUF_X2 inst_10041 ( .A(net_10002), .Z(net_10003) );
SDFF_X2 inst_566 ( .SI(net_7807), .Q(net_6573), .D(net_6573), .SE(net_3823), .CK(net_9699) );
OR2_X4 inst_1399 ( .A2(net_6959), .A1(net_6958), .ZN(net_478) );
CLKBUF_X2 inst_8912 ( .A(net_8483), .Z(net_8874) );
CLKBUF_X2 inst_12301 ( .A(net_12262), .Z(net_12263) );
CLKBUF_X2 inst_10613 ( .A(net_10574), .Z(net_10575) );
NAND2_X1 inst_4357 ( .ZN(net_4370), .A2(net_3853), .A1(net_2062) );
INV_X4 inst_4819 ( .ZN(net_4785), .A(net_1094) );
NAND2_X1 inst_4327 ( .ZN(net_4537), .A2(net_3870), .A1(net_2146) );
CLKBUF_X2 inst_12997 ( .A(net_12958), .Z(net_12959) );
CLKBUF_X2 inst_11375 ( .A(net_11336), .Z(net_11337) );
INV_X4 inst_4774 ( .ZN(net_1720), .A(net_1719) );
CLKBUF_X2 inst_8622 ( .A(net_8262), .Z(net_8584) );
CLKBUF_X2 inst_10419 ( .A(net_10380), .Z(net_10381) );
NOR2_X2 inst_2333 ( .A2(net_6285), .A1(net_5840), .ZN(net_5808) );
CLKBUF_X2 inst_12401 ( .A(net_12362), .Z(net_12363) );
DFFR_X2 inst_7047 ( .QN(net_6011), .D(net_3140), .CK(net_10438), .RN(x1822) );
CLKBUF_X2 inst_11345 ( .A(net_11306), .Z(net_11307) );
INV_X2 inst_5928 ( .A(net_7322), .ZN(net_1788) );
INV_X4 inst_5056 ( .ZN(net_750), .A(net_643) );
NAND2_X2 inst_4016 ( .A1(net_6933), .A2(net_1654), .ZN(net_1036) );
INV_X4 inst_5370 ( .A(net_7783), .ZN(net_510) );
OAI21_X2 inst_1732 ( .ZN(net_5560), .B1(net_5412), .A(net_4827), .B2(net_4153) );
NAND2_X2 inst_2914 ( .ZN(net_5713), .A2(net_5712), .A1(net_2949) );
AOI21_X2 inst_7648 ( .ZN(net_3440), .B2(net_3439), .A(net_3211), .B1(net_728) );
NAND2_X2 inst_3294 ( .ZN(net_3658), .A1(net_3657), .A2(net_3229) );
AOI22_X2 inst_7256 ( .B1(net_6947), .A1(net_6915), .ZN(net_5300), .A2(net_5298), .B2(net_5297) );
NAND3_X2 inst_2741 ( .ZN(net_2360), .A3(net_1619), .A1(net_1479), .A2(net_1012) );
CLKBUF_X2 inst_11825 ( .A(net_11786), .Z(net_11787) );
CLKBUF_X2 inst_11966 ( .A(net_11927), .Z(net_11928) );
INV_X2 inst_6119 ( .ZN(net_5936), .A(x1286) );
CLKBUF_X2 inst_14380 ( .A(net_8818), .Z(net_14342) );
OAI22_X2 inst_1522 ( .B1(net_4644), .A1(net_4057), .B2(net_4056), .ZN(net_4052), .A2(net_4051) );
CLKBUF_X2 inst_12135 ( .A(net_11701), .Z(net_12097) );
CLKBUF_X2 inst_11455 ( .A(net_11416), .Z(net_11417) );
DFF_X2 inst_6269 ( .QN(net_5970), .D(net_2635), .CK(net_11409) );
CLKBUF_X2 inst_13955 ( .A(net_12769), .Z(net_13917) );
CLKBUF_X2 inst_13247 ( .A(net_13208), .Z(net_13209) );
CLKBUF_X2 inst_9481 ( .A(net_9442), .Z(net_9443) );
INV_X2 inst_5858 ( .A(net_796), .ZN(net_623) );
NAND2_X2 inst_3069 ( .A1(net_7162), .A2(net_4954), .ZN(net_4936) );
CLKBUF_X2 inst_8645 ( .A(net_8606), .Z(net_8607) );
NAND2_X2 inst_3631 ( .ZN(net_1952), .A1(net_1287), .A2(net_1128) );
INV_X2 inst_5761 ( .ZN(net_3034), .A(net_2976) );
DFFR_X2 inst_6964 ( .QN(net_7782), .D(net_4163), .CK(net_10254), .RN(x1822) );
CLKBUF_X2 inst_12809 ( .A(net_12770), .Z(net_12771) );
CLKBUF_X2 inst_12520 ( .A(net_12481), .Z(net_12482) );
SDFF_X2 inst_1101 ( .SI(net_6820), .Q(net_6820), .D(net_3801), .SE(net_3722), .CK(net_8349) );
CLKBUF_X2 inst_8596 ( .A(net_8557), .Z(net_8558) );
CLKBUF_X2 inst_9528 ( .A(net_8757), .Z(net_9490) );
DFF_X1 inst_6652 ( .QN(net_7659), .D(net_5193), .CK(net_10555) );
NAND2_X2 inst_2950 ( .ZN(net_5490), .A1(net_4949), .A2(net_4948) );
CLKBUF_X2 inst_11889 ( .A(net_11850), .Z(net_11851) );
CLKBUF_X2 inst_8584 ( .A(net_8545), .Z(net_8546) );
CLKBUF_X2 inst_7902 ( .A(net_7858), .Z(net_7864) );
INV_X4 inst_5691 ( .A(net_7382), .ZN(net_892) );
CLKBUF_X2 inst_8392 ( .A(net_7898), .Z(net_8354) );
SDFF_X2 inst_861 ( .SI(net_7047), .Q(net_7047), .D(net_3784), .SE(net_3777), .CK(net_11876) );
CLKBUF_X2 inst_11549 ( .A(net_11510), .Z(net_11511) );
AOI22_X2 inst_7431 ( .A1(net_2970), .B1(net_2772), .ZN(net_2761), .A2(net_233), .B2(net_159) );
CLKBUF_X2 inst_12013 ( .A(net_11974), .Z(net_11975) );
NAND2_X2 inst_2990 ( .A1(net_6722), .A2(net_5031), .ZN(net_5021) );
AOI222_X2 inst_7495 ( .B1(net_7367), .C1(net_7303), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2088), .A1(net_2087) );
SDFF_X2 inst_1283 ( .D(net_7807), .SE(net_3256), .SI(net_144), .Q(net_144), .CK(net_10690) );
NOR2_X2 inst_2451 ( .ZN(net_2819), .A2(net_2696), .A1(net_1182) );
CLKBUF_X2 inst_11225 ( .A(net_11186), .Z(net_11187) );
CLKBUF_X2 inst_10625 ( .A(net_10586), .Z(net_10587) );
SDFF_X2 inst_1202 ( .SI(net_7085), .Q(net_7085), .D(net_3898), .SE(net_3747), .CK(net_10979) );
NAND2_X1 inst_4290 ( .ZN(net_4577), .A2(net_3867), .A1(net_1184) );
DFFR_X2 inst_7020 ( .D(net_3295), .QN(net_295), .CK(net_11435), .RN(x1822) );
NOR2_X4 inst_2227 ( .ZN(net_5671), .A1(net_5535), .A2(net_4502) );
CLKBUF_X2 inst_12594 ( .A(net_12555), .Z(net_12556) );
SDFF_X2 inst_660 ( .Q(net_6718), .D(net_6718), .SE(net_3871), .SI(net_3791), .CK(net_8154) );
NOR2_X2 inst_2490 ( .ZN(net_2394), .A1(net_2393), .A2(net_2230) );
CLKBUF_X2 inst_11027 ( .A(net_10988), .Z(net_10989) );
CLKBUF_X2 inst_10238 ( .A(net_10199), .Z(net_10200) );
CLKBUF_X2 inst_10150 ( .A(net_10111), .Z(net_10112) );
INV_X4 inst_5195 ( .ZN(net_506), .A(net_505) );
OAI22_X2 inst_1576 ( .A2(net_3297), .B2(net_3286), .ZN(net_3269), .A1(net_3268), .B1(net_463) );
CLKBUF_X2 inst_11532 ( .A(net_11493), .Z(net_11494) );
NAND2_X2 inst_3462 ( .A2(net_5982), .ZN(net_2888), .A1(net_2887) );
CLKBUF_X2 inst_8288 ( .A(net_8135), .Z(net_8250) );
NAND2_X1 inst_4254 ( .ZN(net_4672), .A2(net_3988), .A1(net_2180) );
INV_X4 inst_5642 ( .ZN(net_1224), .A(net_280) );
NAND2_X1 inst_4330 ( .ZN(net_4534), .A2(net_3870), .A1(net_1985) );
AOI222_X2 inst_7459 ( .ZN(net_2221), .A1(net_2220), .B1(net_2219), .C1(net_2218), .A2(net_2204), .B2(net_2202), .C2(net_2200) );
CLKBUF_X2 inst_11898 ( .A(net_11859), .Z(net_11860) );
CLKBUF_X2 inst_10031 ( .A(net_9992), .Z(net_9993) );
CLKBUF_X2 inst_8390 ( .A(net_8351), .Z(net_8352) );
CLKBUF_X2 inst_14220 ( .A(net_14181), .Z(net_14182) );
CLKBUF_X2 inst_11925 ( .A(net_11886), .Z(net_11887) );
DFF_X1 inst_6659 ( .QN(net_7651), .D(net_5182), .CK(net_12263) );
AND2_X4 inst_7828 ( .ZN(net_3017), .A2(net_2819), .A1(net_2258) );
NAND2_X1 inst_4368 ( .ZN(net_4359), .A2(net_3856), .A1(net_1759) );
CLKBUF_X2 inst_10331 ( .A(net_8312), .Z(net_10293) );
CLKBUF_X2 inst_12204 ( .A(net_12165), .Z(net_12166) );
CLKBUF_X2 inst_11137 ( .A(net_8832), .Z(net_11099) );
CLKBUF_X2 inst_9388 ( .A(net_9349), .Z(net_9350) );
SDFF_X2 inst_794 ( .SI(net_6923), .Q(net_6923), .SE(net_3887), .D(net_3801), .CK(net_8131) );
NAND3_X2 inst_2754 ( .ZN(net_2347), .A3(net_1599), .A1(net_1434), .A2(net_970) );
AOI22_X2 inst_7354 ( .B2(net_3105), .ZN(net_3096), .A2(net_2712), .A1(net_1127), .B1(net_652) );
CLKBUF_X2 inst_12049 ( .A(net_12010), .Z(net_12011) );
NAND3_X2 inst_2759 ( .ZN(net_2342), .A3(net_1640), .A1(net_1509), .A2(net_990) );
CLKBUF_X2 inst_12092 ( .A(net_12053), .Z(net_12054) );
SDFF_X2 inst_1147 ( .SI(net_6808), .Q(net_6808), .D(net_3897), .SE(net_3722), .CK(net_11697) );
OAI21_X2 inst_1768 ( .B1(net_5539), .ZN(net_5426), .A(net_4640), .B2(net_3993) );
DFF_X1 inst_6410 ( .QN(net_6157), .D(net_5760), .CK(net_11054) );
CLKBUF_X2 inst_12865 ( .A(net_12826), .Z(net_12827) );
CLKBUF_X2 inst_11165 ( .A(net_11126), .Z(net_11127) );
CLKBUF_X2 inst_8256 ( .A(net_8217), .Z(net_8218) );
NAND2_X2 inst_2917 ( .ZN(net_5707), .A2(net_5706), .A1(net_2757) );
NOR2_X2 inst_2423 ( .A2(net_5892), .ZN(net_3226), .A1(net_687) );
OR2_X2 inst_1408 ( .A1(net_4152), .ZN(net_1690), .A2(net_1689) );
SDFF_X2 inst_996 ( .Q(net_6484), .D(net_6484), .SE(net_3904), .SI(net_3788), .CK(net_10835) );
CLKBUF_X2 inst_10963 ( .A(net_8283), .Z(net_10925) );
INV_X2 inst_5889 ( .A(net_7328), .ZN(net_1768) );
CLKBUF_X2 inst_12074 ( .A(net_11086), .Z(net_12036) );
CLKBUF_X2 inst_13563 ( .A(net_13524), .Z(net_13525) );
OAI21_X2 inst_1889 ( .B1(net_5232), .ZN(net_5192), .A(net_4568), .B2(net_3866) );
OAI22_X2 inst_1527 ( .B1(net_4644), .A1(net_4057), .B2(net_4045), .ZN(net_4042), .A2(net_4041) );
INV_X16 inst_6142 ( .ZN(net_1975), .A(net_915) );
OAI21_X2 inst_2011 ( .ZN(net_4499), .B1(net_4498), .B2(net_4497), .A(net_3664) );
CLKBUF_X2 inst_13495 ( .A(net_13456), .Z(net_13457) );
OAI21_X2 inst_1761 ( .ZN(net_5435), .B1(net_5434), .A(net_4658), .B2(net_3993) );
SDFF_X2 inst_740 ( .Q(net_6858), .D(net_6858), .SE(net_3893), .SI(net_3821), .CK(net_11499) );
DFF_X1 inst_6582 ( .QN(net_7571), .D(net_5068), .CK(net_13453) );
CLKBUF_X2 inst_9418 ( .A(net_8767), .Z(net_9380) );
AND3_X2 inst_7803 ( .A1(net_2616), .ZN(net_2563), .A3(net_1206), .A2(x1155) );
INV_X4 inst_5474 ( .A(net_5990), .ZN(net_606) );
NAND2_X2 inst_4189 ( .A2(net_6032), .ZN(net_1159), .A1(net_467) );
XNOR2_X2 inst_84 ( .B(net_2256), .ZN(net_1307), .A(net_1306) );
DFF_X1 inst_6803 ( .D(net_3864), .CK(net_9564), .Q(x765) );
INV_X2 inst_5974 ( .A(net_7506), .ZN(net_2188) );
OAI21_X2 inst_1937 ( .B1(net_5548), .ZN(net_5108), .A(net_4740), .B2(net_3988) );
SDFF_X2 inst_173 ( .Q(net_6241), .SI(net_6240), .D(net_3536), .SE(net_392), .CK(net_13519) );
AOI21_X2 inst_7660 ( .B2(net_5927), .ZN(net_3320), .A(net_3319), .B1(net_1829) );
INV_X4 inst_5568 ( .A(net_7409), .ZN(net_2097) );
NAND2_X1 inst_4405 ( .A2(net_3087), .ZN(net_2913), .A1(net_2839) );
SDFF_X2 inst_611 ( .Q(net_6617), .D(net_6617), .SE(net_3830), .SI(net_3795), .CK(net_12029) );
CLKBUF_X2 inst_10550 ( .A(net_8549), .Z(net_10512) );
NOR2_X2 inst_2487 ( .A2(net_5778), .ZN(net_2593), .A1(net_917) );
CLKBUF_X2 inst_12417 ( .A(net_11398), .Z(net_12379) );
INV_X2 inst_5821 ( .ZN(net_1047), .A(net_1046) );
INV_X2 inst_5713 ( .ZN(net_4253), .A(net_4127) );
CLKBUF_X2 inst_12462 ( .A(net_9783), .Z(net_12424) );
CLKBUF_X2 inst_10493 ( .A(net_10454), .Z(net_10455) );
CLKBUF_X2 inst_12549 ( .A(net_12510), .Z(net_12511) );
CLKBUF_X2 inst_8723 ( .A(net_8684), .Z(net_8685) );
CLKBUF_X2 inst_13047 ( .A(net_10508), .Z(net_13009) );
AND3_X2 inst_7802 ( .A1(net_2590), .ZN(net_2586), .A2(net_2585), .A3(net_2584) );
OAI21_X2 inst_1943 ( .B1(net_5237), .ZN(net_5082), .A(net_4734), .B2(net_3986) );
AND2_X4 inst_7847 ( .ZN(net_1960), .A2(net_796), .A1(net_677) );
SDFF_X2 inst_490 ( .Q(net_6854), .D(net_6854), .SI(net_3898), .SE(net_3893), .CK(net_11512) );
INV_X4 inst_5573 ( .A(net_6075), .ZN(net_3558) );
AOI22_X2 inst_7305 ( .B1(net_6678), .A1(net_6646), .ZN(net_5140), .A2(net_5139), .B2(net_5138) );
CLKBUF_X2 inst_13378 ( .A(net_10733), .Z(net_13340) );
CLKBUF_X2 inst_8375 ( .A(net_7907), .Z(net_8337) );
NOR2_X4 inst_2218 ( .ZN(net_5680), .A1(net_5559), .A2(net_4517) );
SDFF_X2 inst_1309 ( .D(net_6386), .SE(net_5801), .SI(net_331), .Q(net_331), .CK(net_14299) );
OAI22_X2 inst_1531 ( .B1(net_4650), .A1(net_4080), .B2(net_4068), .ZN(net_4036), .A2(net_4035) );
AOI21_X2 inst_7640 ( .B1(net_5892), .ZN(net_3916), .B2(net_3915), .A(net_2594) );
DFFR_X2 inst_7083 ( .QN(net_7727), .D(net_2793), .CK(net_9989), .RN(x1822) );
CLKBUF_X2 inst_11706 ( .A(net_10987), .Z(net_11668) );
INV_X4 inst_4938 ( .ZN(net_902), .A(net_754) );
NAND2_X2 inst_2922 ( .A2(net_7776), .ZN(net_5770), .A1(net_5606) );
NAND2_X2 inst_3803 ( .A1(net_6906), .A2(net_1639), .ZN(net_1542) );
CLKBUF_X2 inst_13234 ( .A(net_9945), .Z(net_13196) );
CLKBUF_X2 inst_11831 ( .A(net_11792), .Z(net_11793) );
CLKBUF_X2 inst_11649 ( .A(net_11610), .Z(net_11611) );
CLKBUF_X2 inst_10242 ( .A(net_9439), .Z(net_10204) );
NAND2_X2 inst_3183 ( .ZN(net_4750), .A2(net_3941), .A1(net_2017) );
CLKBUF_X2 inst_10410 ( .A(net_9530), .Z(net_10372) );
CLKBUF_X2 inst_10860 ( .A(net_10821), .Z(net_10822) );
CLKBUF_X2 inst_13301 ( .A(net_13262), .Z(net_13263) );
CLKBUF_X2 inst_11256 ( .A(net_9145), .Z(net_11218) );
NAND2_X1 inst_4312 ( .ZN(net_4554), .A2(net_3866), .A1(net_1871) );
CLKBUF_X2 inst_12950 ( .A(net_12911), .Z(net_12912) );
INV_X4 inst_5328 ( .ZN(net_500), .A(net_154) );
CLKBUF_X2 inst_8410 ( .A(net_8007), .Z(net_8372) );
CLKBUF_X2 inst_13161 ( .A(net_13122), .Z(net_13123) );
DFF_X2 inst_6226 ( .QN(net_6693), .D(net_3721), .CK(net_9713) );
SDFF_X2 inst_1037 ( .Q(net_7539), .D(net_7539), .SE(net_3896), .SI(net_373), .CK(net_10264) );
AOI21_X2 inst_7777 ( .B1(net_6597), .ZN(net_4418), .B2(net_2583), .A(net_2302) );
CLKBUF_X2 inst_8652 ( .A(net_8321), .Z(net_8614) );
SDFF_X2 inst_300 ( .SI(net_7518), .Q(net_7518), .D(net_5107), .SE(net_3988), .CK(net_9800) );
NAND2_X2 inst_3596 ( .ZN(net_2404), .A2(net_1876), .A1(net_1439) );
SDFF_X2 inst_1250 ( .SI(net_6546), .Q(net_6546), .D(net_3795), .SE(net_3756), .CK(net_11222) );
SDFF_X2 inst_1226 ( .SI(net_7219), .Q(net_7219), .D(net_3796), .SE(net_3751), .CK(net_8686) );
DFFR_X2 inst_7071 ( .QN(net_6034), .D(net_3062), .CK(net_12639), .RN(x1822) );
CLKBUF_X2 inst_10240 ( .A(net_9504), .Z(net_10202) );
INV_X2 inst_5964 ( .A(net_7667), .ZN(net_1883) );
CLKBUF_X2 inst_8802 ( .A(net_8763), .Z(net_8764) );
SDFF_X2 inst_446 ( .Q(net_7399), .D(net_7399), .SE(net_3994), .SI(net_364), .CK(net_9621) );
OAI21_X2 inst_1979 ( .ZN(net_4854), .B1(net_4853), .A(net_4540), .B2(net_3870) );
SDFF_X2 inst_364 ( .SI(net_7614), .Q(net_7614), .D(net_4785), .SE(net_3870), .CK(net_10274) );
CLKBUF_X2 inst_11586 ( .A(net_10009), .Z(net_11548) );
CLKBUF_X2 inst_9253 ( .A(net_9214), .Z(net_9215) );
INV_X4 inst_4923 ( .A(net_3804), .ZN(net_3142) );
CLKBUF_X2 inst_9283 ( .A(net_9244), .Z(net_9245) );
SDFF_X2 inst_824 ( .SI(net_7799), .Q(net_6970), .D(net_6970), .SE(net_3891), .CK(net_11956) );
NAND2_X2 inst_2997 ( .A1(net_6746), .A2(net_5033), .ZN(net_5014) );
NAND2_X2 inst_3533 ( .ZN(net_2534), .A2(net_2139), .A1(net_1438) );
AND2_X4 inst_7839 ( .ZN(net_1967), .A2(net_784), .A1(net_662) );
INV_X4 inst_4712 ( .ZN(net_3120), .A(net_3051) );
SDFF_X2 inst_411 ( .SI(net_7376), .Q(net_7376), .D(net_4777), .SE(net_3853), .CK(net_12207) );
CLKBUF_X2 inst_12897 ( .A(net_12858), .Z(net_12859) );
CLKBUF_X2 inst_9055 ( .A(net_7876), .Z(net_9017) );
CLKBUF_X2 inst_10393 ( .A(net_10354), .Z(net_10355) );
CLKBUF_X2 inst_10380 ( .A(net_10341), .Z(net_10342) );
DFF_X1 inst_6600 ( .QN(net_7507), .D(net_5408), .CK(net_10071) );
CLKBUF_X2 inst_13691 ( .A(net_13652), .Z(net_13653) );
CLKBUF_X2 inst_9007 ( .A(net_8968), .Z(net_8969) );
NAND2_X2 inst_3750 ( .A1(net_6497), .A2(net_1642), .ZN(net_1595) );
NAND2_X2 inst_4026 ( .A1(net_6662), .A2(net_1655), .ZN(net_1026) );
CLKBUF_X2 inst_11173 ( .A(net_11134), .Z(net_11135) );
CLKBUF_X2 inst_9395 ( .A(net_9356), .Z(net_9357) );
CLKBUF_X2 inst_11333 ( .A(net_11294), .Z(net_11295) );
CLKBUF_X2 inst_10668 ( .A(net_10417), .Z(net_10630) );
NAND2_X2 inst_4056 ( .A1(net_6801), .A2(net_1651), .ZN(net_996) );
CLKBUF_X2 inst_11010 ( .A(net_10971), .Z(net_10972) );
NAND2_X1 inst_4382 ( .ZN(net_4345), .A2(net_3859), .A1(net_2073) );
CLKBUF_X2 inst_10908 ( .A(net_7837), .Z(net_10870) );
NAND2_X1 inst_4401 ( .A2(net_3297), .ZN(net_3078), .A1(net_3077) );
CLKBUF_X2 inst_14426 ( .A(net_14387), .Z(net_14388) );
CLKBUF_X2 inst_10388 ( .A(net_10349), .Z(net_10350) );
NAND2_X2 inst_3430 ( .ZN(net_3218), .A2(net_3107), .A1(net_2768) );
CLKBUF_X2 inst_13480 ( .A(net_13441), .Z(net_13442) );
CLKBUF_X2 inst_8708 ( .A(net_8454), .Z(net_8670) );
CLKBUF_X2 inst_13297 ( .A(net_10150), .Z(net_13259) );
CLKBUF_X2 inst_14020 ( .A(net_13981), .Z(net_13982) );
CLKBUF_X2 inst_13368 ( .A(net_13329), .Z(net_13330) );
CLKBUF_X2 inst_9874 ( .A(net_9835), .Z(net_9836) );
INV_X4 inst_5538 ( .ZN(net_563), .A(net_282) );
INV_X4 inst_5462 ( .A(net_7281), .ZN(net_2011) );
NAND2_X2 inst_3439 ( .ZN(net_3209), .A2(net_3032), .A1(net_2767) );
CLKBUF_X2 inst_13968 ( .A(net_13929), .Z(net_13930) );
CLKBUF_X2 inst_8308 ( .A(net_8083), .Z(net_8270) );
INV_X4 inst_5412 ( .A(net_6423), .ZN(net_2453) );
XNOR2_X2 inst_61 ( .A(net_6403), .B(net_6402), .ZN(net_1837) );
SDFF_X2 inst_203 ( .Q(net_6311), .SI(net_6310), .D(net_3699), .SE(net_392), .CK(net_13570) );
INV_X2 inst_5834 ( .A(net_1304), .ZN(net_900) );
CLKBUF_X2 inst_10901 ( .A(net_10282), .Z(net_10863) );
CLKBUF_X2 inst_14077 ( .A(net_14038), .Z(net_14039) );
CLKBUF_X2 inst_10014 ( .A(net_9975), .Z(net_9976) );
SDFF_X2 inst_1139 ( .SI(net_6663), .Q(net_6663), .D(net_3814), .SE(net_3465), .CK(net_12886) );
CLKBUF_X2 inst_10597 ( .A(net_10558), .Z(net_10559) );
CLKBUF_X2 inst_12459 ( .A(net_12420), .Z(net_12421) );
CLKBUF_X2 inst_8852 ( .A(net_8813), .Z(net_8814) );
CLKBUF_X2 inst_8520 ( .A(net_8322), .Z(net_8482) );
DFF_X1 inst_6601 ( .QN(net_7508), .D(net_5407), .CK(net_10070) );
INV_X8 inst_4507 ( .ZN(net_3819), .A(net_3260) );
CLKBUF_X2 inst_9968 ( .A(net_9929), .Z(net_9930) );
OAI22_X2 inst_1571 ( .A2(net_3297), .B2(net_3286), .ZN(net_3278), .A1(net_3277), .B1(net_1714) );
AOI21_X2 inst_7631 ( .ZN(net_4298), .B2(net_3451), .B1(net_3179), .A(x889) );
CLKBUF_X2 inst_12009 ( .A(net_11009), .Z(net_11971) );
DFF_X1 inst_6607 ( .QN(net_7514), .D(net_5401), .CK(net_9651) );
SDFF_X2 inst_456 ( .Q(net_6057), .SI(net_3918), .SE(net_3312), .D(net_3311), .CK(net_10322) );
SDFF_X2 inst_832 ( .Q(net_7011), .D(net_7011), .SE(net_3899), .SI(net_3787), .CK(net_8081) );
CLKBUF_X2 inst_8214 ( .A(net_8175), .Z(net_8176) );
CLKBUF_X2 inst_11246 ( .A(net_8931), .Z(net_11208) );
DFF_X1 inst_6511 ( .QN(net_7433), .D(net_5449), .CK(net_9814) );
OR2_X2 inst_1402 ( .ZN(net_4161), .A2(net_3895), .A1(net_3452) );
CLKBUF_X2 inst_8102 ( .A(net_8063), .Z(net_8064) );
SDFF_X2 inst_275 ( .D(net_6399), .SE(net_6052), .SI(net_324), .Q(net_324), .CK(net_13832) );
CLKBUF_X2 inst_11492 ( .A(net_11453), .Z(net_11454) );
NAND2_X2 inst_3106 ( .A1(net_6583), .A2(net_4897), .ZN(net_4895) );
DFF_X1 inst_6810 ( .D(net_3458), .CK(net_10820), .Q(x379) );
NAND2_X2 inst_3728 ( .A1(net_7040), .A2(net_1975), .ZN(net_1617) );
CLKBUF_X2 inst_11576 ( .A(net_11537), .Z(net_11538) );
CLKBUF_X2 inst_13379 ( .A(net_13340), .Z(net_13341) );
DFF_X1 inst_6843 ( .D(net_2557), .Q(net_208), .CK(net_9745) );
NOR2_X2 inst_2416 ( .A1(net_5997), .ZN(net_3407), .A2(net_3399) );
DFF_X2 inst_6270 ( .QN(net_6415), .D(net_2688), .CK(net_10208) );
INV_X4 inst_5453 ( .ZN(net_486), .A(x1215) );
NAND2_X2 inst_3812 ( .A1(net_6637), .A2(net_1624), .ZN(net_1533) );
INV_X4 inst_5405 ( .A(net_7273), .ZN(net_2158) );
CLKBUF_X2 inst_8810 ( .A(net_8771), .Z(net_8772) );
CLKBUF_X2 inst_13317 ( .A(net_9506), .Z(net_13279) );
CLKBUF_X2 inst_7879 ( .A(net_7840), .Z(net_7841) );
NAND2_X2 inst_3959 ( .A1(net_6843), .A2(net_1521), .ZN(net_1325) );
NOR2_X2 inst_2503 ( .ZN(net_1242), .A2(net_671), .A1(net_630) );
CLKBUF_X2 inst_9839 ( .A(net_8962), .Z(net_9801) );
INV_X4 inst_5420 ( .A(net_6104), .ZN(net_3703) );
INV_X4 inst_4877 ( .ZN(net_1084), .A(net_905) );
INV_X8 inst_4518 ( .ZN(net_3465), .A(net_3118) );
CLKBUF_X2 inst_11185 ( .A(net_11146), .Z(net_11147) );
CLKBUF_X2 inst_9994 ( .A(net_9955), .Z(net_9956) );
CLKBUF_X2 inst_10348 ( .A(net_10309), .Z(net_10310) );
XNOR2_X2 inst_94 ( .B(net_2999), .ZN(net_1660), .A(net_1151) );
CLKBUF_X2 inst_9726 ( .A(net_9687), .Z(net_9688) );
CLKBUF_X2 inst_10946 ( .A(net_10907), .Z(net_10908) );
DFF_X1 inst_6832 ( .D(net_2592), .QN(net_227), .CK(net_12300) );
CLKBUF_X2 inst_14234 ( .A(net_14195), .Z(net_14196) );
CLKBUF_X2 inst_7958 ( .A(net_7919), .Z(net_7920) );
CLKBUF_X2 inst_11858 ( .A(net_11819), .Z(net_11820) );
CLKBUF_X2 inst_13060 ( .A(net_13021), .Z(net_13022) );
CLKBUF_X2 inst_11237 ( .A(net_11198), .Z(net_11199) );
NAND2_X1 inst_4345 ( .ZN(net_4382), .A2(net_3856), .A1(net_1754) );
SDFF_X2 inst_424 ( .D(net_6391), .SE(net_6051), .SI(net_308), .Q(net_308), .CK(net_13734) );
SDFF_X2 inst_591 ( .Q(net_6589), .D(net_6589), .SE(net_3823), .SI(net_3801), .CK(net_12030) );
NAND2_X2 inst_3166 ( .ZN(net_4767), .A2(net_3941), .A1(net_2162) );
CLKBUF_X2 inst_14218 ( .A(net_14179), .Z(net_14180) );
AOI22_X2 inst_7452 ( .B2(net_2931), .A2(net_2647), .ZN(net_714), .A1(net_713), .B1(net_712) );
CLKBUF_X2 inst_13807 ( .A(net_9277), .Z(net_13769) );
CLKBUF_X2 inst_10428 ( .A(net_10389), .Z(net_10390) );
NAND2_X2 inst_3656 ( .A1(net_7062), .ZN(net_1807), .A2(net_791) );
CLKBUF_X2 inst_12497 ( .A(net_11848), .Z(net_12459) );
NOR2_X4 inst_2237 ( .ZN(net_5661), .A1(net_5516), .A2(net_4489) );
NAND2_X1 inst_4417 ( .ZN(net_2740), .A2(net_266), .A1(net_265) );
CLKBUF_X2 inst_10784 ( .A(net_10745), .Z(net_10746) );
CLKBUF_X2 inst_9155 ( .A(net_9116), .Z(net_9117) );
CLKBUF_X2 inst_8320 ( .A(net_8281), .Z(net_8282) );
DFF_X1 inst_6834 ( .D(net_2621), .CK(net_9560), .Q(x149) );
INV_X2 inst_5727 ( .ZN(net_3999), .A(net_3906) );
CLKBUF_X2 inst_14012 ( .A(net_10823), .Z(net_13974) );
CLKBUF_X2 inst_11861 ( .A(net_11347), .Z(net_11823) );
DFF_X1 inst_6853 ( .D(net_2552), .Q(net_218), .CK(net_9537) );
NAND3_X2 inst_2706 ( .ZN(net_2471), .A2(net_1815), .A3(net_1545), .A1(net_1416) );
CLKBUF_X2 inst_8640 ( .A(net_8601), .Z(net_8602) );
SDFF_X2 inst_476 ( .Q(net_6985), .D(net_6985), .SI(net_3900), .SE(net_3891), .CK(net_9042) );
CLKBUF_X2 inst_10249 ( .A(net_10210), .Z(net_10211) );
DFF_X1 inst_6684 ( .QN(net_7272), .D(net_5120), .CK(net_9964) );
NAND2_X2 inst_3742 ( .A1(net_6908), .A2(net_1639), .ZN(net_1603) );
CLKBUF_X2 inst_10701 ( .A(net_10662), .Z(net_10663) );
NOR2_X2 inst_2499 ( .A1(net_3044), .ZN(net_1740), .A2(net_1739) );
NAND3_X2 inst_2827 ( .ZN(net_1217), .A2(net_1216), .A3(net_1215), .A1(net_680) );
CLKBUF_X2 inst_11542 ( .A(net_11503), .Z(net_11504) );
CLKBUF_X2 inst_9062 ( .A(net_9023), .Z(net_9024) );
XNOR2_X2 inst_20 ( .ZN(net_2614), .A(net_2248), .B(net_1208) );
NOR2_X2 inst_2448 ( .A2(net_5922), .ZN(net_2973), .A1(net_549) );
CLKBUF_X2 inst_10007 ( .A(net_9168), .Z(net_9969) );
CLKBUF_X2 inst_13421 ( .A(net_13382), .Z(net_13383) );
INV_X4 inst_5549 ( .A(net_6180), .ZN(net_3564) );
INV_X4 inst_4994 ( .A(net_781), .ZN(net_752) );
NOR2_X2 inst_2541 ( .ZN(net_5889), .A1(net_486), .A2(x1286) );
CLKBUF_X2 inst_13590 ( .A(net_8014), .Z(net_13552) );
SDFF_X2 inst_576 ( .Q(net_6572), .D(net_6572), .SE(net_3823), .SI(net_3811), .CK(net_9355) );
OAI21_X2 inst_1693 ( .ZN(net_5601), .A(net_5303), .B2(net_4519), .B1(net_4132) );
CLKBUF_X2 inst_14398 ( .A(net_14359), .Z(net_14360) );
CLKBUF_X2 inst_10182 ( .A(net_10143), .Z(net_10144) );
CLKBUF_X2 inst_10131 ( .A(net_9423), .Z(net_10093) );
NAND2_X2 inst_3306 ( .ZN(net_3634), .A1(net_3633), .A2(net_3229) );
SDFF_X2 inst_1020 ( .SI(net_6516), .Q(net_6516), .SE(net_3886), .D(net_3788), .CK(net_11239) );
CLKBUF_X2 inst_11007 ( .A(net_10968), .Z(net_10969) );
CLKBUF_X2 inst_10376 ( .A(net_10337), .Z(net_10338) );
AOI21_X2 inst_7721 ( .B1(net_6866), .ZN(net_5907), .B2(net_2579), .A(net_2341) );
NAND2_X4 inst_2876 ( .A1(net_5883), .ZN(net_4263), .A2(net_2580) );
NAND2_X2 inst_3055 ( .A1(net_7122), .ZN(net_4951), .A2(net_4950) );
CLKBUF_X2 inst_11057 ( .A(net_8603), .Z(net_11019) );
CLKBUF_X2 inst_13886 ( .A(net_13847), .Z(net_13848) );
SDFF_X2 inst_976 ( .Q(net_6428), .D(net_6428), .SE(net_3820), .SI(net_3799), .CK(net_8853) );
NAND2_X2 inst_3952 ( .A1(net_6437), .A2(net_1677), .ZN(net_1333) );
CLKBUF_X2 inst_9919 ( .A(net_9880), .Z(net_9881) );
CLKBUF_X2 inst_12084 ( .A(net_12045), .Z(net_12046) );
SDFF_X2 inst_1279 ( .D(net_3792), .SE(net_3256), .SI(net_130), .Q(net_130), .CK(net_8479) );
NAND2_X2 inst_3588 ( .ZN(net_2412), .A2(net_1900), .A1(net_1456) );
DFFR_X2 inst_7027 ( .D(net_3283), .QN(net_271), .CK(net_12332), .RN(x1822) );
DFF_X1 inst_6562 ( .QN(net_7435), .D(net_5045), .CK(net_12097) );
INV_X4 inst_5559 ( .A(net_7419), .ZN(net_2170) );
SDFF_X2 inst_1096 ( .SI(net_6940), .Q(net_6940), .D(net_3787), .SE(net_3734), .CK(net_8842) );
CLKBUF_X2 inst_13011 ( .A(net_12972), .Z(net_12973) );
AOI222_X2 inst_7474 ( .C1(net_7519), .B1(net_7487), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2157), .A1(net_2156) );
CLKBUF_X2 inst_13280 ( .A(net_13241), .Z(net_13242) );
CLKBUF_X2 inst_13287 ( .A(net_13248), .Z(net_13249) );
INV_X8 inst_4552 ( .ZN(net_1256), .A(net_885) );
CLKBUF_X2 inst_11036 ( .A(net_10997), .Z(net_10998) );
CLKBUF_X2 inst_8025 ( .A(net_7986), .Z(net_7987) );
CLKBUF_X2 inst_9260 ( .A(net_7990), .Z(net_9222) );
INV_X4 inst_5637 ( .A(net_7735), .ZN(net_2676) );
OAI21_X2 inst_1839 ( .B1(net_5363), .ZN(net_5333), .A(net_4373), .B2(net_3853) );
CLKBUF_X2 inst_8041 ( .A(net_8002), .Z(net_8003) );
AOI21_X2 inst_7723 ( .B1(net_6729), .ZN(net_5895), .B2(net_2581), .A(net_2363) );
NAND2_X2 inst_3399 ( .ZN(net_3468), .A2(net_3329), .A1(net_3242) );
NAND2_X2 inst_3414 ( .ZN(net_3259), .A1(net_3258), .A2(net_499) );
CLKBUF_X2 inst_13095 ( .A(net_13056), .Z(net_13057) );
INV_X8 inst_4495 ( .ZN(net_3899), .A(net_3148) );
OAI22_X2 inst_1432 ( .B1(net_5857), .ZN(net_5797), .A2(net_5790), .B2(net_5789), .A1(net_5773) );
SDFF_X2 inst_725 ( .Q(net_6841), .D(net_6841), .SE(net_3893), .SI(net_3812), .CK(net_8654) );
INV_X4 inst_5667 ( .A(net_7574), .ZN(net_1891) );
CLKBUF_X2 inst_12840 ( .A(net_12801), .Z(net_12802) );
CLKBUF_X2 inst_12159 ( .A(net_12120), .Z(net_12121) );
DFF_X2 inst_6326 ( .QN(net_7803), .CK(net_11528), .D(x1519) );
NAND2_X2 inst_3084 ( .A1(net_6482), .A2(net_4927), .ZN(net_4919) );
CLKBUF_X2 inst_11739 ( .A(net_11700), .Z(net_11701) );
SDFFR_X2 inst_1337 ( .Q(net_7691), .D(net_7691), .SI(net_3797), .SE(net_3405), .CK(net_13195), .RN(x1822) );
CLKBUF_X2 inst_9790 ( .A(net_9394), .Z(net_9752) );
INV_X4 inst_5375 ( .A(net_6166), .ZN(net_3530) );
NOR2_X2 inst_2464 ( .ZN(net_2734), .A2(net_2733), .A1(net_2730) );
NAND2_X2 inst_3096 ( .A1(net_6476), .A2(net_4927), .ZN(net_4907) );
CLKBUF_X2 inst_8776 ( .A(net_8677), .Z(net_8738) );
NAND2_X2 inst_3015 ( .A1(net_6857), .A2(net_5004), .ZN(net_4994) );
CLKBUF_X2 inst_11197 ( .A(net_11158), .Z(net_11159) );
CLKBUF_X2 inst_9433 ( .A(net_9394), .Z(net_9395) );
CLKBUF_X2 inst_14432 ( .A(net_11849), .Z(net_14394) );
NAND2_X2 inst_4010 ( .ZN(net_1260), .A2(net_1225), .A1(net_358) );
CLKBUF_X2 inst_13254 ( .A(net_9668), .Z(net_13216) );
CLKBUF_X2 inst_9677 ( .A(net_9638), .Z(net_9639) );
NAND2_X2 inst_3328 ( .ZN(net_3590), .A1(net_3589), .A2(net_3228) );
CLKBUF_X2 inst_11618 ( .A(net_11579), .Z(net_11580) );
NOR2_X2 inst_2441 ( .A2(net_5971), .ZN(net_3166), .A1(net_3003) );
CLKBUF_X2 inst_8399 ( .A(net_8360), .Z(net_8361) );
SDFF_X2 inst_1111 ( .SI(net_6656), .Q(net_6656), .D(net_3806), .SE(net_3465), .CK(net_9329) );
CLKBUF_X2 inst_11945 ( .A(net_11906), .Z(net_11907) );
CLKBUF_X2 inst_9122 ( .A(net_7829), .Z(net_9084) );
NAND3_X2 inst_2658 ( .ZN(net_3942), .A3(net_3388), .A2(net_2932), .A1(net_2824) );
CLKBUF_X2 inst_9714 ( .A(net_9675), .Z(net_9676) );
AOI22_X2 inst_7427 ( .A1(net_2970), .B1(net_2772), .ZN(net_2765), .A2(net_243), .B2(net_169) );
SDFF_X2 inst_878 ( .D(net_7802), .SI(net_7037), .Q(net_7037), .SE(net_3777), .CK(net_8201) );
CLKBUF_X2 inst_11496 ( .A(net_11457), .Z(net_11458) );
INV_X4 inst_4959 ( .ZN(net_1170), .A(net_722) );
CLKBUF_X2 inst_13442 ( .A(net_13403), .Z(net_13404) );
DFF_X1 inst_6782 ( .QN(net_6084), .D(net_4318), .CK(net_12946) );
SDFF_X2 inst_480 ( .SI(net_6506), .Q(net_6506), .SE(net_3886), .D(net_3831), .CK(net_8805) );
OAI21_X2 inst_1926 ( .ZN(net_5119), .A(net_4754), .B2(net_3941), .B1(net_1177) );
INV_X4 inst_4631 ( .ZN(net_4191), .A(net_4042) );
NAND2_X1 inst_4351 ( .ZN(net_4376), .A2(net_3853), .A1(net_2038) );
DFF_X2 inst_6211 ( .QN(net_7686), .D(net_4009), .CK(net_8321) );
CLKBUF_X2 inst_12761 ( .A(net_12722), .Z(net_12723) );
DFF_X1 inst_6383 ( .QN(net_6114), .D(net_5705), .CK(net_11207) );
SDFF_X2 inst_564 ( .Q(net_6569), .D(net_6569), .SI(net_3894), .SE(net_3823), .CK(net_9193) );
NAND2_X2 inst_2986 ( .A1(net_6720), .A2(net_5031), .ZN(net_5025) );
CLKBUF_X2 inst_8074 ( .A(net_8035), .Z(net_8036) );
NOR3_X2 inst_2206 ( .A3(net_5922), .ZN(net_3039), .A2(net_2851), .A1(net_2850) );
CLKBUF_X2 inst_13597 ( .A(net_13558), .Z(net_13559) );
NAND3_X2 inst_2792 ( .ZN(net_2308), .A3(net_1549), .A1(net_1275), .A2(net_971) );
CLKBUF_X2 inst_12795 ( .A(net_12052), .Z(net_12757) );
CLKBUF_X2 inst_10262 ( .A(net_9403), .Z(net_10224) );
SDFF_X2 inst_739 ( .Q(net_6857), .D(net_6857), .SE(net_3893), .SI(net_3788), .CK(net_11501) );
CLKBUF_X2 inst_11210 ( .A(net_11171), .Z(net_11172) );
DFF_X1 inst_6637 ( .QN(net_7593), .D(net_5242), .CK(net_10568) );
DFF_X1 inst_6500 ( .QN(net_7422), .D(net_5532), .CK(net_12627) );
XNOR2_X2 inst_46 ( .B(net_7230), .ZN(net_2440), .A(net_1062) );
SDFF_X2 inst_934 ( .SI(net_7176), .Q(net_7176), .SE(net_3817), .D(net_3811), .CK(net_7849) );
NOR2_X2 inst_2537 ( .A2(net_7750), .A1(net_3208), .ZN(net_657) );
SDFF_X2 inst_1000 ( .Q(net_6487), .D(net_6487), .SE(net_3904), .SI(net_3800), .CK(net_8057) );
CLKBUF_X2 inst_12361 ( .A(net_12322), .Z(net_12323) );
SDFF_X2 inst_1126 ( .SI(net_6676), .Q(net_6676), .D(net_3836), .SE(net_3471), .CK(net_9080) );
CLKBUF_X2 inst_13065 ( .A(net_13026), .Z(net_13027) );
NAND2_X2 inst_3470 ( .ZN(net_2745), .A1(net_2709), .A2(net_229) );
SDFF_X2 inst_796 ( .SI(net_6897), .Q(net_6897), .SE(net_3887), .D(net_3799), .CK(net_11795) );
NAND3_X2 inst_2585 ( .ZN(net_5754), .A1(net_5649), .A2(net_5271), .A3(net_4309) );
CLKBUF_X2 inst_12044 ( .A(net_11020), .Z(net_12006) );
NOR2_X2 inst_2364 ( .ZN(net_5286), .A2(net_4628), .A1(net_4484) );
CLKBUF_X2 inst_14135 ( .A(net_14096), .Z(net_14097) );
CLKBUF_X2 inst_11727 ( .A(net_11688), .Z(net_11689) );
NAND2_X1 inst_4299 ( .ZN(net_4567), .A2(net_3866), .A1(net_1901) );
CLKBUF_X2 inst_11281 ( .A(net_11242), .Z(net_11243) );
OAI21_X2 inst_1882 ( .ZN(net_5203), .B1(net_5202), .A(net_4576), .B2(net_3867) );
CLKBUF_X2 inst_13787 ( .A(net_13748), .Z(net_13749) );
AND2_X4 inst_7812 ( .A1(net_7791), .A2(net_7771), .ZN(net_4145) );
AOI21_X2 inst_7628 ( .B2(net_5951), .B1(net_5950), .ZN(net_5607), .A(x977) );
DFF_X1 inst_6699 ( .QN(net_7297), .D(net_5376), .CK(net_12251) );
CLKBUF_X2 inst_8441 ( .A(net_8402), .Z(net_8403) );
CLKBUF_X2 inst_8218 ( .A(net_8179), .Z(net_8180) );
DFF_X1 inst_6578 ( .QN(net_7567), .D(net_5072), .CK(net_13461) );
OAI22_X2 inst_1499 ( .B1(net_4660), .A1(net_4105), .B2(net_4104), .ZN(net_4100), .A2(net_4099) );
NAND2_X2 inst_2972 ( .ZN(net_5497), .A2(net_5258), .A1(net_406) );
CLKBUF_X2 inst_12849 ( .A(net_12810), .Z(net_12811) );
CLKBUF_X2 inst_9470 ( .A(net_9374), .Z(net_9432) );
INV_X4 inst_5531 ( .A(net_7701), .ZN(net_845) );
INV_X4 inst_5397 ( .A(net_6139), .ZN(net_3655) );
SDFF_X2 inst_727 ( .SI(net_7807), .Q(net_6843), .D(net_6843), .SE(net_3893), .CK(net_11506) );
CLKBUF_X2 inst_11795 ( .A(net_9550), .Z(net_11757) );
INV_X4 inst_4804 ( .ZN(net_5094), .A(net_1178) );
CLKBUF_X2 inst_11686 ( .A(net_11647), .Z(net_11648) );
CLKBUF_X2 inst_9293 ( .A(net_9254), .Z(net_9255) );
NAND2_X4 inst_2874 ( .A1(net_4278), .ZN(net_4265), .A2(net_1833) );
CLKBUF_X2 inst_12345 ( .A(net_12306), .Z(net_12307) );
DFF_X1 inst_6485 ( .QN(net_7416), .D(net_5567), .CK(net_12509) );
INV_X4 inst_4607 ( .ZN(net_4237), .A(net_4092) );
NOR2_X2 inst_2431 ( .ZN(net_3423), .A2(net_3119), .A1(net_3042) );
NAND2_X2 inst_3297 ( .ZN(net_3652), .A1(net_3651), .A2(net_3229) );
CLKBUF_X2 inst_8861 ( .A(net_8011), .Z(net_8823) );
INV_X2 inst_5931 ( .A(net_7651), .ZN(net_2134) );
INV_X4 inst_5429 ( .A(net_6140), .ZN(net_3653) );
CLKBUF_X2 inst_12556 ( .A(net_10955), .Z(net_12518) );
CLKBUF_X2 inst_12052 ( .A(net_9717), .Z(net_12014) );
NAND2_X1 inst_4423 ( .A1(net_7611), .A2(net_2131), .ZN(net_1478) );
CLKBUF_X2 inst_10438 ( .A(net_10399), .Z(net_10400) );
CLKBUF_X2 inst_13384 ( .A(net_8286), .Z(net_13346) );
CLKBUF_X2 inst_11880 ( .A(net_10609), .Z(net_11842) );
CLKBUF_X2 inst_8274 ( .A(net_8235), .Z(net_8236) );
AOI222_X2 inst_7607 ( .A1(net_7398), .ZN(net_5440), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_361), .C2(net_359) );
SDFF_X2 inst_953 ( .SI(net_7168), .Q(net_7168), .SE(net_3817), .D(net_3798), .CK(net_13332) );
CLKBUF_X2 inst_13674 ( .A(net_10916), .Z(net_13636) );
CLKBUF_X2 inst_11524 ( .A(net_7942), .Z(net_11486) );
NAND2_X1 inst_4342 ( .ZN(net_4385), .A2(net_3856), .A1(net_1785) );
INV_X4 inst_5483 ( .A(net_7583), .ZN(net_1858) );
CLKBUF_X2 inst_8664 ( .A(net_8625), .Z(net_8626) );
CLKBUF_X2 inst_12887 ( .A(net_12848), .Z(net_12849) );
CLKBUF_X2 inst_10398 ( .A(net_10359), .Z(net_10360) );
INV_X4 inst_5060 ( .ZN(net_736), .A(net_637) );
NAND2_X1 inst_4339 ( .ZN(net_4388), .A2(net_3856), .A1(net_1778) );
CLKBUF_X2 inst_14187 ( .A(net_14148), .Z(net_14149) );
OR2_X2 inst_1421 ( .A2(net_6409), .A1(net_6408), .ZN(net_1920) );
DFF_X1 inst_6694 ( .QN(net_7292), .D(net_5381), .CK(net_12995) );
NAND2_X2 inst_3373 ( .ZN(net_3500), .A1(net_3499), .A2(net_3223) );
CLKBUF_X2 inst_8919 ( .A(net_8744), .Z(net_8881) );
CLKBUF_X2 inst_12819 ( .A(net_12780), .Z(net_12781) );
INV_X4 inst_4902 ( .ZN(net_1240), .A(net_867) );
NAND2_X1 inst_4262 ( .ZN(net_4658), .A2(net_3993), .A1(net_1476) );
CLKBUF_X2 inst_12607 ( .A(net_10931), .Z(net_12569) );
CLKBUF_X2 inst_8298 ( .A(net_7993), .Z(net_8260) );
CLKBUF_X2 inst_10406 ( .A(net_9891), .Z(net_10368) );
CLKBUF_X2 inst_13882 ( .A(net_13843), .Z(net_13844) );
CLKBUF_X2 inst_9688 ( .A(net_9649), .Z(net_9650) );
NAND2_X2 inst_3664 ( .A1(net_7345), .A2(net_1798), .ZN(net_1797) );
CLKBUF_X2 inst_9961 ( .A(net_9922), .Z(net_9923) );
AOI221_X2 inst_7613 ( .C2(net_3105), .B1(net_2970), .ZN(net_2967), .A(net_2789), .C1(net_465), .B2(net_248) );
CLKBUF_X2 inst_11464 ( .A(net_11425), .Z(net_11426) );
CLKBUF_X2 inst_10536 ( .A(net_10497), .Z(net_10498) );
INV_X2 inst_6011 ( .A(net_7296), .ZN(net_2057) );
DFFR_X2 inst_6956 ( .QN(net_7731), .D(net_5780), .CK(net_7979), .RN(x1822) );
INV_X4 inst_4720 ( .ZN(net_3022), .A(net_2865) );
NAND2_X2 inst_3486 ( .ZN(net_2662), .A1(net_2661), .A2(net_2660) );
CLKBUF_X2 inst_13246 ( .A(net_13207), .Z(net_13208) );
CLKBUF_X2 inst_11488 ( .A(net_11449), .Z(net_11450) );
CLKBUF_X2 inst_8833 ( .A(net_8794), .Z(net_8795) );
CLKBUF_X2 inst_13961 ( .A(net_13922), .Z(net_13923) );
INV_X4 inst_4986 ( .A(net_7817), .ZN(net_3791) );
CLKBUF_X2 inst_9636 ( .A(net_9597), .Z(net_9598) );
DFF_X1 inst_6378 ( .QN(net_6284), .D(net_5806), .CK(net_13695) );
SDFF_X2 inst_294 ( .D(net_6395), .SE(net_6052), .SI(net_320), .Q(net_320), .CK(net_13824) );
CLKBUF_X2 inst_13510 ( .A(net_8592), .Z(net_13472) );
CLKBUF_X2 inst_8970 ( .A(net_8931), .Z(net_8932) );
CLKBUF_X2 inst_13358 ( .A(net_11458), .Z(net_13320) );
CLKBUF_X2 inst_12099 ( .A(net_8907), .Z(net_12061) );
CLKBUF_X2 inst_8275 ( .A(net_8236), .Z(net_8237) );
AND2_X4 inst_7842 ( .ZN(net_1484), .A2(net_792), .A1(net_643) );
CLKBUF_X2 inst_13769 ( .A(net_8433), .Z(net_13731) );
NAND2_X2 inst_3384 ( .ZN(net_3478), .A1(net_3477), .A2(net_3226) );
CLKBUF_X2 inst_11202 ( .A(net_10766), .Z(net_11164) );
DFF_X1 inst_6628 ( .QN(net_7599), .D(net_5257), .CK(net_10575) );
CLKBUF_X2 inst_10029 ( .A(net_9990), .Z(net_9991) );
AOI21_X4 inst_7621 ( .B2(net_5953), .B1(net_5952), .ZN(net_5606), .A(x940) );
SDFF_X2 inst_810 ( .Q(net_6965), .D(net_6965), .SE(net_3891), .SI(net_3778), .CK(net_10648) );
CLKBUF_X2 inst_13877 ( .A(net_13838), .Z(net_13839) );
CLKBUF_X2 inst_8982 ( .A(net_8943), .Z(net_8944) );
SDFF_X2 inst_230 ( .Q(net_6324), .SI(net_6323), .D(net_3637), .SE(net_392), .CK(net_14019) );
INV_X2 inst_5903 ( .A(net_7347), .ZN(net_2038) );
CLKBUF_X2 inst_9511 ( .A(net_9472), .Z(net_9473) );
CLKBUF_X2 inst_9767 ( .A(net_9728), .Z(net_9729) );
NAND2_X2 inst_3035 ( .A1(net_7022), .A2(net_4979), .ZN(net_4972) );
CLKBUF_X2 inst_10089 ( .A(net_10050), .Z(net_10051) );
OAI21_X2 inst_1893 ( .B1(net_5222), .ZN(net_5188), .A(net_4564), .B2(net_3866) );
CLKBUF_X2 inst_12063 ( .A(net_12024), .Z(net_12025) );
INV_X4 inst_4728 ( .A(net_5983), .ZN(net_3041) );
INV_X4 inst_5101 ( .ZN(net_2384), .A(net_1068) );
CLKBUF_X2 inst_8325 ( .A(net_7973), .Z(net_8287) );
DFF_X1 inst_6480 ( .QN(net_7411), .D(net_5572), .CK(net_10104) );
NAND2_X1 inst_4385 ( .ZN(net_4342), .A2(net_3859), .A1(net_2041) );
AND2_X4 inst_7836 ( .A1(net_6417), .A2(net_3452), .ZN(net_2714) );
CLKBUF_X2 inst_10010 ( .A(net_9971), .Z(net_9972) );
CLKBUF_X2 inst_11984 ( .A(net_10645), .Z(net_11946) );
SDFF_X2 inst_481 ( .Q(net_7006), .D(net_7006), .SE(net_3899), .SI(net_3894), .CK(net_8232) );
INV_X2 inst_5992 ( .A(net_7482), .ZN(net_2219) );
INV_X4 inst_4606 ( .ZN(net_4238), .A(net_4094) );
CLKBUF_X2 inst_8633 ( .A(net_8594), .Z(net_8595) );
CLKBUF_X2 inst_14375 ( .A(net_11188), .Z(net_14337) );
SDFF_X2 inst_452 ( .Q(net_6061), .SI(net_3922), .SE(net_3320), .D(net_3319), .CK(net_10328) );
CLKBUF_X2 inst_10338 ( .A(net_10299), .Z(net_10300) );
CLKBUF_X2 inst_9392 ( .A(net_9353), .Z(net_9354) );
CLKBUF_X2 inst_13699 ( .A(net_13660), .Z(net_13661) );
CLKBUF_X2 inst_8397 ( .A(net_7875), .Z(net_8359) );
NAND2_X2 inst_3061 ( .A1(net_7125), .A2(net_4950), .ZN(net_4944) );
DFF_X2 inst_6208 ( .QN(net_7684), .D(net_4171), .CK(net_10797) );
CLKBUF_X2 inst_13146 ( .A(net_13107), .Z(net_13108) );
CLKBUF_X2 inst_14000 ( .A(net_13386), .Z(net_13962) );
NAND2_X2 inst_4144 ( .A1(net_1148), .ZN(net_911), .A2(net_716) );
CLKBUF_X2 inst_10254 ( .A(net_10215), .Z(net_10216) );
CLKBUF_X2 inst_14308 ( .A(net_14269), .Z(net_14270) );
CLKBUF_X2 inst_11180 ( .A(net_11141), .Z(net_11142) );
SDFF_X2 inst_728 ( .Q(net_6844), .D(net_6844), .SE(net_3893), .SI(net_3787), .CK(net_8884) );
CLKBUF_X2 inst_13056 ( .A(net_13017), .Z(net_13018) );
CLKBUF_X2 inst_10372 ( .A(net_8410), .Z(net_10334) );
NAND3_X2 inst_2780 ( .ZN(net_2320), .A3(net_1560), .A1(net_1333), .A2(net_1001) );
NAND2_X2 inst_3121 ( .A1(net_6611), .A2(net_4899), .ZN(net_4880) );
NOR2_X2 inst_2485 ( .A2(net_5778), .ZN(net_2649), .A1(net_431) );
CLKBUF_X2 inst_9087 ( .A(net_9048), .Z(net_9049) );
CLKBUF_X2 inst_10584 ( .A(net_10545), .Z(net_10546) );
DFF_X1 inst_6655 ( .QN(net_7662), .D(net_5190), .CK(net_13061) );
CLKBUF_X2 inst_13353 ( .A(net_13314), .Z(net_13315) );
NAND2_X2 inst_4152 ( .A2(net_1225), .ZN(net_1065), .A1(net_361) );
NOR2_X4 inst_2217 ( .ZN(net_5681), .A1(net_5561), .A2(net_4520) );
CLKBUF_X2 inst_13707 ( .A(net_13668), .Z(net_13669) );
CLKBUF_X2 inst_11031 ( .A(net_10992), .Z(net_10993) );
SDFF_X2 inst_850 ( .SI(net_7799), .Q(net_7002), .D(net_7002), .SE(net_3899), .CK(net_11942) );
NAND2_X4 inst_2844 ( .ZN(net_5479), .A1(net_4930), .A2(net_4929) );
AOI221_X2 inst_7612 ( .C2(net_3105), .B1(net_2970), .ZN(net_2969), .C1(net_2968), .A(net_2785), .B2(net_249) );
NOR2_X2 inst_2492 ( .ZN(net_2591), .A2(net_2489), .A1(net_1277) );
CLKBUF_X2 inst_11175 ( .A(net_7919), .Z(net_11137) );
NAND2_X2 inst_3582 ( .ZN(net_2428), .A2(net_2427), .A1(net_799) );
NAND2_X2 inst_3480 ( .ZN(net_2680), .A1(net_2679), .A2(net_2678) );
CLKBUF_X2 inst_14125 ( .A(net_13246), .Z(net_14087) );
CLKBUF_X2 inst_12642 ( .A(net_12603), .Z(net_12604) );
CLKBUF_X2 inst_11721 ( .A(net_11682), .Z(net_11683) );
NOR2_X2 inst_2438 ( .ZN(net_3428), .A1(net_3044), .A2(net_3043) );
INV_X32 inst_5705 ( .ZN(net_5778), .A(net_4596) );
CLKBUF_X2 inst_10879 ( .A(net_10840), .Z(net_10841) );
CLKBUF_X2 inst_10391 ( .A(net_10352), .Z(net_10353) );
INV_X4 inst_5479 ( .A(net_6090), .ZN(net_3481) );
SDFF_X2 inst_237 ( .Q(net_6357), .SI(net_6356), .D(net_3599), .SE(net_392), .CK(net_13959) );
NOR2_X2 inst_2543 ( .A2(net_1699), .ZN(net_651), .A1(net_546) );
NAND3_X2 inst_2772 ( .ZN(net_2328), .A3(net_1608), .A1(net_1446), .A2(net_1008) );
CLKBUF_X2 inst_11449 ( .A(net_10970), .Z(net_11411) );
CLKBUF_X2 inst_8836 ( .A(net_8000), .Z(net_8798) );
CLKBUF_X2 inst_13178 ( .A(net_13139), .Z(net_13140) );
AOI21_X2 inst_7638 ( .ZN(net_3952), .B2(net_3760), .B1(net_2886), .A(net_929) );
CLKBUF_X2 inst_8056 ( .A(net_8017), .Z(net_8018) );
CLKBUF_X2 inst_11017 ( .A(net_10978), .Z(net_10979) );
DFFR_X2 inst_7093 ( .QN(net_6420), .D(net_2717), .CK(net_13018), .RN(x1822) );
INV_X4 inst_4818 ( .ZN(net_4802), .A(net_1108) );
XNOR2_X2 inst_51 ( .ZN(net_2254), .A(net_2253), .B(net_2252) );
SDFF_X2 inst_813 ( .Q(net_6987), .D(net_6987), .SE(net_3891), .SI(net_3803), .CK(net_11905) );
CLKBUF_X2 inst_10379 ( .A(net_10340), .Z(net_10341) );
DFF_X1 inst_6691 ( .QN(net_7280), .D(net_5113), .CK(net_12254) );
CLKBUF_X2 inst_13373 ( .A(net_13334), .Z(net_13335) );
CLKBUF_X2 inst_11195 ( .A(net_11156), .Z(net_11157) );
CLKBUF_X2 inst_10381 ( .A(net_8028), .Z(net_10343) );
OAI21_X2 inst_1837 ( .ZN(net_5336), .B1(net_5335), .A(net_4378), .B2(net_3856) );
SDFF_X2 inst_974 ( .Q(net_6454), .D(net_6454), .SE(net_3820), .SI(net_3801), .CK(net_8070) );
CLKBUF_X2 inst_13198 ( .A(net_13159), .Z(net_13160) );
CLKBUF_X2 inst_9100 ( .A(net_9061), .Z(net_9062) );
INV_X4 inst_5686 ( .A(net_6127), .ZN(net_3639) );
CLKBUF_X2 inst_10944 ( .A(net_10559), .Z(net_10906) );
NAND2_X2 inst_3291 ( .ZN(net_3664), .A1(net_3663), .A2(net_3229) );
XNOR2_X2 inst_64 ( .ZN(net_1727), .B(net_1726), .A(net_1270) );
SDFF_X2 inst_1001 ( .Q(net_6460), .D(net_6460), .SE(net_3904), .SI(net_3799), .CK(net_11655) );
CLKBUF_X2 inst_13964 ( .A(net_13925), .Z(net_13926) );
SDFF_X2 inst_743 ( .Q(net_6860), .D(net_6860), .SE(net_3893), .SI(net_3800), .CK(net_11746) );
OAI21_X2 inst_2106 ( .ZN(net_3972), .A(net_3971), .B2(net_3874), .B1(net_865) );
NAND2_X2 inst_4051 ( .A1(net_6533), .A2(net_1645), .ZN(net_1001) );
NAND3_X2 inst_2723 ( .ZN(net_2378), .A3(net_1631), .A1(net_1442), .A2(net_967) );
NAND2_X2 inst_3033 ( .A1(net_7021), .A2(net_4979), .ZN(net_4974) );
INV_X2 inst_5825 ( .ZN(net_930), .A(net_929) );
NAND2_X2 inst_2925 ( .ZN(net_5531), .A1(net_5007), .A2(net_5005) );
AND2_X4 inst_7843 ( .ZN(net_1969), .A2(net_788), .A1(net_638) );
CLKBUF_X2 inst_9141 ( .A(net_9102), .Z(net_9103) );
NAND2_X1 inst_4265 ( .ZN(net_4655), .A2(net_3993), .A1(net_1376) );
CLKBUF_X2 inst_10537 ( .A(net_10498), .Z(net_10499) );
CLKBUF_X2 inst_9510 ( .A(net_9463), .Z(net_9472) );
OAI21_X2 inst_1828 ( .ZN(net_5354), .B1(net_5353), .A(net_4390), .B2(net_3856) );
CLKBUF_X2 inst_8628 ( .A(net_8589), .Z(net_8590) );
OAI21_X2 inst_1809 ( .ZN(net_5379), .B1(net_5359), .A(net_4349), .B2(net_3859) );
NAND2_X2 inst_3388 ( .ZN(net_3895), .A1(net_936), .A2(net_113) );
NAND2_X2 inst_3735 ( .A1(net_7181), .A2(net_1637), .ZN(net_1610) );
DFF_X1 inst_6664 ( .QN(net_7657), .D(net_5174), .CK(net_10550) );
CLKBUF_X2 inst_11238 ( .A(net_9562), .Z(net_11200) );
NAND3_X2 inst_2675 ( .ZN(net_3748), .A3(net_3307), .A1(net_2967), .A2(net_2945) );
INV_X4 inst_5311 ( .A(net_6015), .ZN(net_2596) );
CLKBUF_X2 inst_8272 ( .A(net_8144), .Z(net_8234) );
CLKBUF_X2 inst_12172 ( .A(net_12133), .Z(net_12134) );
CLKBUF_X2 inst_11866 ( .A(net_10995), .Z(net_11828) );
SDFF_X2 inst_141 ( .Q(net_6237), .SI(net_6236), .SE(net_392), .D(net_143), .CK(net_13620) );
CLKBUF_X2 inst_10578 ( .A(net_10539), .Z(net_10540) );
NOR2_X2 inst_2520 ( .A1(net_7093), .ZN(net_1100), .A2(net_867) );
NAND2_X1 inst_4344 ( .ZN(net_4383), .A2(net_3856), .A1(net_1774) );
CLKBUF_X2 inst_8111 ( .A(net_8035), .Z(net_8073) );
CLKBUF_X2 inst_8541 ( .A(net_8502), .Z(net_8503) );
SDFF_X2 inst_571 ( .Q(net_6729), .D(net_6729), .SI(net_3892), .SE(net_3815), .CK(net_11118) );
NAND2_X2 inst_4011 ( .A1(net_6941), .A2(net_1654), .ZN(net_1044) );
OAI21_X2 inst_1974 ( .B1(net_4866), .ZN(net_4862), .A(net_4392), .B2(net_3856) );
INV_X2 inst_6007 ( .A(net_7500), .ZN(net_2123) );
CLKBUF_X2 inst_11478 ( .A(net_11439), .Z(net_11440) );
CLKBUF_X2 inst_10432 ( .A(net_10393), .Z(net_10394) );
OAI21_X2 inst_2017 ( .B2(net_4497), .ZN(net_4491), .B1(net_4099), .A(net_3652) );
SDFF_X2 inst_1154 ( .SI(net_6816), .Q(net_6816), .D(net_3790), .SE(net_3722), .CK(net_8336) );
AOI21_X2 inst_7728 ( .B1(net_6456), .ZN(net_4426), .B2(net_2580), .A(net_2332) );
CLKBUF_X2 inst_12413 ( .A(net_12374), .Z(net_12375) );
DFF_X1 inst_6445 ( .QN(net_6096), .D(net_5725), .CK(net_9221) );
CLKBUF_X2 inst_9584 ( .A(net_7907), .Z(net_9546) );
CLKBUF_X2 inst_8045 ( .A(net_8006), .Z(net_8007) );
AOI22_X2 inst_7436 ( .B1(net_7078), .A1(net_7046), .A2(net_1975), .ZN(net_1974), .B2(net_791) );
SDFF_X2 inst_469 ( .Q(net_7021), .D(net_7021), .SE(net_3899), .SI(net_3898), .CK(net_10878) );
CLKBUF_X2 inst_8598 ( .A(net_8437), .Z(net_8560) );
AOI222_X2 inst_7468 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2179), .A1(net_2178), .B1(net_2177), .C1(net_2176) );
CLKBUF_X2 inst_11689 ( .A(net_9809), .Z(net_11651) );
NAND2_X2 inst_2980 ( .A1(net_6717), .ZN(net_5032), .A2(net_5031) );
INV_X4 inst_5197 ( .ZN(net_643), .A(net_547) );
DFF_X1 inst_6837 ( .D(net_2502), .Q(net_159), .CK(net_9436) );
CLKBUF_X2 inst_10184 ( .A(net_10145), .Z(net_10146) );
SDFF_X2 inst_915 ( .Q(net_7151), .D(net_7151), .SE(net_3903), .SI(net_3805), .CK(net_11580) );
CLKBUF_X2 inst_9869 ( .A(net_9830), .Z(net_9831) );
CLKBUF_X2 inst_8866 ( .A(net_8455), .Z(net_8828) );
DFF_X1 inst_6507 ( .QN(net_7429), .D(net_5517), .CK(net_12498) );
DFF_X1 inst_6642 ( .QN(net_7631), .D(net_5226), .CK(net_10562) );
NAND2_X1 inst_4416 ( .ZN(net_2741), .A2(net_192), .A1(net_191) );
CLKBUF_X2 inst_10008 ( .A(net_9969), .Z(net_9970) );
NOR2_X2 inst_2339 ( .A2(net_6319), .A1(net_5840), .ZN(net_5802) );
CLKBUF_X2 inst_12300 ( .A(net_12261), .Z(net_12262) );
INV_X4 inst_5660 ( .A(net_7702), .ZN(net_851) );
CLKBUF_X2 inst_14017 ( .A(net_13978), .Z(net_13979) );
CLKBUF_X2 inst_11603 ( .A(net_11564), .Z(net_11565) );
SDFF_X2 inst_1216 ( .SI(net_7206), .Q(net_7206), .D(net_3813), .SE(net_3750), .CK(net_13313) );
CLKBUF_X2 inst_8260 ( .A(net_8080), .Z(net_8222) );
DFF_X1 inst_6697 ( .QN(net_7295), .D(net_5378), .CK(net_10172) );
CLKBUF_X2 inst_9552 ( .A(net_9367), .Z(net_9514) );
CLKBUF_X2 inst_12591 ( .A(net_8700), .Z(net_12553) );
SDFF_X2 inst_952 ( .SI(net_7167), .Q(net_7167), .SE(net_3817), .D(net_3799), .CK(net_13333) );
INV_X4 inst_4807 ( .ZN(net_4780), .A(net_1175) );
OAI221_X2 inst_1668 ( .C2(net_5902), .ZN(net_4641), .B1(net_4637), .B2(net_4405), .C1(net_4030), .A(net_3490) );
INV_X2 inst_5972 ( .A(net_7617), .ZN(net_1186) );
CLKBUF_X2 inst_11169 ( .A(net_11130), .Z(net_11131) );
CLKBUF_X2 inst_9987 ( .A(net_9063), .Z(net_9949) );
AOI22_X2 inst_7254 ( .B1(net_6810), .A1(net_6778), .A2(net_5316), .B2(net_5315), .ZN(net_5302) );
INV_X4 inst_4811 ( .ZN(net_4787), .A(net_1167) );
CLKBUF_X2 inst_11942 ( .A(net_11903), .Z(net_11904) );
DFFR_X2 inst_7068 ( .QN(net_6030), .D(net_3088), .CK(net_10000), .RN(x1822) );
SDFF_X2 inst_721 ( .SI(net_6766), .Q(net_6766), .SE(net_3816), .D(net_3814), .CK(net_8957) );
CLKBUF_X2 inst_11135 ( .A(net_11006), .Z(net_11097) );
CLKBUF_X2 inst_10838 ( .A(net_10799), .Z(net_10800) );
SDFF_X2 inst_293 ( .D(net_6395), .SE(net_5799), .SI(net_380), .Q(net_380), .CK(net_14325) );
INV_X4 inst_4741 ( .ZN(net_2749), .A(net_2748) );
CLKBUF_X2 inst_11078 ( .A(net_10758), .Z(net_11040) );
CLKBUF_X2 inst_13667 ( .A(net_13628), .Z(net_13629) );
OR2_X4 inst_1366 ( .ZN(net_4168), .A2(net_3746), .A1(net_3338) );
NAND2_X2 inst_3009 ( .A1(net_6854), .A2(net_5004), .ZN(net_5000) );
NAND2_X2 inst_3744 ( .A1(net_6505), .A2(net_1642), .ZN(net_1601) );
CLKBUF_X2 inst_13079 ( .A(net_13040), .Z(net_13041) );
OAI21_X2 inst_1915 ( .B1(net_5347), .ZN(net_5150), .A(net_4749), .B2(net_3941) );
NAND3_X2 inst_2794 ( .ZN(net_2306), .A3(net_1588), .A1(net_1418), .A2(net_969) );
INV_X4 inst_5402 ( .ZN(net_1223), .A(net_281) );
SDFF_X2 inst_1254 ( .SI(net_6551), .Q(net_6551), .D(net_3800), .SE(net_3755), .CK(net_11618) );
NAND2_X2 inst_2953 ( .ZN(net_5487), .A1(net_4943), .A2(net_4942) );
DFFR_X2 inst_7111 ( .D(net_1944), .QN(net_119), .CK(net_9576), .RN(x1822) );
CLKBUF_X2 inst_14412 ( .A(net_13282), .Z(net_14374) );
CLKBUF_X2 inst_14031 ( .A(net_13992), .Z(net_13993) );
NAND2_X2 inst_3553 ( .ZN(net_2514), .A2(net_2044), .A1(net_1750) );
CLKBUF_X2 inst_13000 ( .A(net_12961), .Z(net_12962) );
CLKBUF_X2 inst_8219 ( .A(net_8178), .Z(net_8181) );
XNOR2_X2 inst_98 ( .ZN(net_2245), .A(net_1153), .B(net_1146) );
OAI21_X2 inst_1811 ( .ZN(net_5377), .B1(net_5355), .A(net_4347), .B2(net_3859) );
INV_X8 inst_4544 ( .ZN(net_2580), .A(net_1278) );
CLKBUF_X2 inst_11147 ( .A(net_11108), .Z(net_11109) );
CLKBUF_X2 inst_11351 ( .A(net_11312), .Z(net_11313) );
NAND2_X2 inst_3087 ( .A1(net_6451), .A2(net_4925), .ZN(net_4916) );
SDFF_X2 inst_959 ( .Q(net_6436), .D(net_6436), .SE(net_3820), .SI(net_3812), .CK(net_8650) );
CLKBUF_X2 inst_10801 ( .A(net_10762), .Z(net_10763) );
CLKBUF_X2 inst_10102 ( .A(net_10063), .Z(net_10064) );
DFFR_X2 inst_7054 ( .QN(net_5987), .D(net_3146), .CK(net_10746), .RN(x1822) );
CLKBUF_X2 inst_8826 ( .A(net_8787), .Z(net_8788) );
CLKBUF_X2 inst_9156 ( .A(net_9117), .Z(net_9118) );
SDFF_X2 inst_163 ( .Q(net_6251), .SI(net_6250), .D(net_3558), .SE(net_392), .CK(net_13987) );
CLKBUF_X2 inst_8455 ( .A(net_8416), .Z(net_8417) );
SDFF_X2 inst_394 ( .SI(net_7335), .Q(net_7335), .D(net_4874), .SE(net_3856), .CK(net_9843) );
CLKBUF_X2 inst_13343 ( .A(net_8428), .Z(net_13305) );
CLKBUF_X2 inst_11619 ( .A(net_8117), .Z(net_11581) );
AOI21_X4 inst_7626 ( .B1(net_7001), .ZN(net_4617), .A(net_2459), .B2(net_1100) );
SDFF_X2 inst_605 ( .Q(net_6610), .D(net_6610), .SE(net_3830), .SI(net_3807), .CK(net_12169) );
CLKBUF_X2 inst_9998 ( .A(net_9959), .Z(net_9960) );
OAI21_X2 inst_1814 ( .ZN(net_5374), .B1(net_5349), .A(net_4344), .B2(net_3859) );
AOI222_X2 inst_7481 ( .C1(net_7523), .B1(net_7491), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2139), .A1(net_2138) );
NAND3_X2 inst_2799 ( .ZN(net_2301), .A3(net_1553), .A1(net_1419), .A2(net_979) );
INV_X8 inst_4470 ( .ZN(net_5280), .A(net_4279) );
CLKBUF_X2 inst_10988 ( .A(net_9530), .Z(net_10950) );
CLKBUF_X2 inst_10875 ( .A(net_10836), .Z(net_10837) );
OAI21_X2 inst_2048 ( .B2(net_4457), .ZN(net_4452), .B1(net_4076), .A(net_3565) );
SDFF_X2 inst_361 ( .SI(net_7610), .Q(net_7610), .D(net_4788), .SE(net_3870), .CK(net_13396) );
NAND2_X2 inst_2948 ( .ZN(net_5492), .A1(net_4955), .A2(net_4953) );
CLKBUF_X2 inst_7900 ( .A(net_7861), .Z(net_7862) );
CLKBUF_X2 inst_11358 ( .A(net_11319), .Z(net_11320) );
CLKBUF_X2 inst_10396 ( .A(net_8220), .Z(net_10358) );
NAND2_X2 inst_3400 ( .ZN(net_3466), .A2(net_3333), .A1(net_3244) );
CLKBUF_X2 inst_8127 ( .A(net_8005), .Z(net_8089) );
CLKBUF_X2 inst_11643 ( .A(net_8821), .Z(net_11605) );
CLKBUF_X2 inst_13850 ( .A(net_13811), .Z(net_13812) );
CLKBUF_X2 inst_12134 ( .A(net_12095), .Z(net_12096) );
OAI21_X2 inst_1931 ( .ZN(net_5114), .A(net_4751), .B2(net_3941), .B1(net_1137) );
CLKBUF_X2 inst_8082 ( .A(net_7862), .Z(net_8044) );
CLKBUF_X2 inst_11008 ( .A(net_9055), .Z(net_10970) );
INV_X4 inst_4735 ( .A(net_5978), .ZN(net_3874) );
DFF_X1 inst_6631 ( .QN(net_7587), .D(net_5252), .CK(net_10300) );
CLKBUF_X2 inst_11926 ( .A(net_10116), .Z(net_11888) );
CLKBUF_X2 inst_8402 ( .A(net_8363), .Z(net_8364) );
NAND2_X2 inst_3002 ( .A1(net_6883), .ZN(net_5009), .A2(net_5006) );
CLKBUF_X2 inst_13007 ( .A(net_12968), .Z(net_12969) );
NAND2_X1 inst_4389 ( .ZN(net_4338), .A2(net_3859), .A1(net_2003) );
SDFF_X2 inst_786 ( .SI(net_6915), .Q(net_6915), .D(net_3804), .SE(net_3781), .CK(net_8145) );
DFF_X1 inst_6828 ( .Q(net_390), .D(net_387), .CK(net_12784) );
NAND2_X2 inst_2940 ( .ZN(net_5506), .A1(net_4972), .A2(net_4971) );
CLKBUF_X2 inst_11855 ( .A(net_11816), .Z(net_11817) );
AOI222_X2 inst_7533 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1904), .A1(net_1903), .B1(net_1902), .C1(net_1901) );
CLKBUF_X2 inst_9383 ( .A(net_9344), .Z(net_9345) );
DFF_X1 inst_6606 ( .QN(net_7513), .D(net_5402), .CK(net_12084) );
XOR2_X2 inst_2 ( .A(net_2573), .Z(net_1250), .B(net_1249) );
CLKBUF_X2 inst_11267 ( .A(net_10225), .Z(net_11229) );
CLKBUF_X2 inst_11003 ( .A(net_10933), .Z(net_10965) );
DFFR_X2 inst_7022 ( .D(net_3266), .QN(net_270), .CK(net_12338), .RN(x1822) );
NAND2_X2 inst_3474 ( .ZN(net_2867), .A1(net_2709), .A2(net_2631) );
CLKBUF_X2 inst_12328 ( .A(net_12289), .Z(net_12290) );
SDFF_X2 inst_578 ( .Q(net_6575), .D(net_6575), .SE(net_3823), .SI(net_3809), .CK(net_7886) );
SDFF_X2 inst_888 ( .Q(net_7100), .D(net_7100), .SE(net_3888), .SI(net_3806), .CK(net_7915) );
CLKBUF_X2 inst_12306 ( .A(net_12267), .Z(net_12268) );
OAI21_X2 inst_1769 ( .B1(net_5537), .ZN(net_5425), .A(net_4639), .B2(net_3993) );
NAND2_X2 inst_3625 ( .ZN(net_1958), .A1(net_1291), .A2(net_1134) );
INV_X2 inst_5999 ( .A(net_6412), .ZN(net_403) );
CLKBUF_X2 inst_14197 ( .A(net_14158), .Z(net_14159) );
CLKBUF_X2 inst_13063 ( .A(net_9532), .Z(net_13025) );
DFF_X1 inst_6598 ( .QN(net_7467), .D(net_5411), .CK(net_12086) );
INV_X2 inst_5979 ( .A(net_7481), .ZN(net_2165) );
AOI22_X2 inst_7317 ( .ZN(net_4594), .B2(net_3978), .A2(net_3386), .A1(net_1742), .B1(net_924) );
AND2_X4 inst_7817 ( .ZN(net_3263), .A2(net_3162), .A1(net_539) );
NAND3_X2 inst_2581 ( .ZN(net_5758), .A1(net_5653), .A2(net_5275), .A3(net_4313) );
NAND2_X2 inst_4110 ( .A1(net_6656), .A2(net_1655), .ZN(net_942) );
OAI211_X2 inst_2164 ( .ZN(net_2725), .B(net_2724), .A(net_2599), .C2(net_2598), .C1(net_2384) );
OAI22_X2 inst_1498 ( .B1(net_4660), .B2(net_4110), .A1(net_4105), .ZN(net_4102), .A2(net_4101) );
SDFFR_X2 inst_1358 ( .Q(net_6024), .D(net_6024), .SI(net_3800), .SE(net_3200), .CK(net_10396), .RN(x1822) );
CLKBUF_X2 inst_13208 ( .A(net_10815), .Z(net_13170) );
CLKBUF_X2 inst_8343 ( .A(net_7983), .Z(net_8305) );
CLKBUF_X2 inst_11696 ( .A(net_11657), .Z(net_11658) );
NAND2_X1 inst_4392 ( .ZN(net_4335), .A2(net_3859), .A1(net_1991) );
CLKBUF_X2 inst_11093 ( .A(net_9292), .Z(net_11055) );
CLKBUF_X2 inst_8590 ( .A(net_8551), .Z(net_8552) );
INV_X4 inst_4915 ( .A(net_3801), .ZN(net_828) );
CLKBUF_X2 inst_14424 ( .A(net_12215), .Z(net_14386) );
CLKBUF_X2 inst_12456 ( .A(net_12417), .Z(net_12418) );
INV_X4 inst_4775 ( .ZN(net_1718), .A(net_1717) );
CLKBUF_X2 inst_8530 ( .A(net_8075), .Z(net_8492) );
CLKBUF_X2 inst_9655 ( .A(net_9130), .Z(net_9617) );
CLKBUF_X2 inst_11245 ( .A(net_7874), .Z(net_11207) );
CLKBUF_X2 inst_10831 ( .A(net_10792), .Z(net_10793) );
NAND2_X1 inst_4450 ( .A2(net_1256), .ZN(net_1130), .A1(net_1129) );
CLKBUF_X2 inst_12817 ( .A(net_12778), .Z(net_12779) );
CLKBUF_X2 inst_12460 ( .A(net_12421), .Z(net_12422) );
NAND2_X2 inst_3182 ( .ZN(net_4751), .A2(net_3941), .A1(net_2023) );
NAND2_X2 inst_3385 ( .ZN(net_3476), .A1(net_3475), .A2(net_3223) );
OAI22_X2 inst_1572 ( .A2(net_3297), .B2(net_3286), .ZN(net_3276), .A1(net_3275), .B1(net_1720) );
CLKBUF_X2 inst_11753 ( .A(net_11714), .Z(net_11715) );
NAND2_X4 inst_2866 ( .ZN(net_4285), .A1(net_4274), .A2(net_1645) );
DFF_X1 inst_6805 ( .D(net_3748), .CK(net_8322), .Q(x390) );
INV_X4 inst_4906 ( .A(net_3795), .ZN(net_3190) );
CLKBUF_X2 inst_11528 ( .A(net_11489), .Z(net_11490) );
CLKBUF_X2 inst_11546 ( .A(net_11507), .Z(net_11508) );
INV_X4 inst_5379 ( .A(net_6126), .ZN(net_3641) );
SDFF_X2 inst_838 ( .Q(net_7018), .D(net_7018), .SE(net_3899), .SI(net_3804), .CK(net_11004) );
CLKBUF_X2 inst_14026 ( .A(net_10979), .Z(net_13988) );
CLKBUF_X2 inst_10221 ( .A(net_10182), .Z(net_10183) );
CLKBUF_X2 inst_12905 ( .A(net_9326), .Z(net_12867) );
INV_X4 inst_4978 ( .A(net_787), .ZN(net_737) );
OR2_X2 inst_1405 ( .ZN(net_3040), .A2(net_3039), .A1(net_2917) );
CLKBUF_X2 inst_7875 ( .A(net_7834), .Z(net_7837) );
DFF_X1 inst_6811 ( .D(net_3376), .CK(net_13413), .Q(x172) );
NAND2_X2 inst_4058 ( .A1(net_6539), .A2(net_1645), .ZN(net_994) );
DFF_X1 inst_6786 ( .Q(net_7780), .D(net_4297), .CK(net_13058) );
CLKBUF_X2 inst_9172 ( .A(net_9133), .Z(net_9134) );
NAND3_X2 inst_2749 ( .ZN(net_2352), .A3(net_1565), .A1(net_1342), .A2(net_976) );
INV_X4 inst_5584 ( .A(net_7787), .ZN(net_1699) );
CLKBUF_X2 inst_9721 ( .A(net_9682), .Z(net_9683) );
DFFR_X2 inst_6963 ( .QN(net_7721), .D(net_4597), .CK(net_12424), .RN(x1822) );
CLKBUF_X2 inst_12048 ( .A(net_12009), .Z(net_12010) );
CLKBUF_X2 inst_8823 ( .A(net_8784), .Z(net_8785) );
CLKBUF_X2 inst_11118 ( .A(net_11079), .Z(net_11080) );
INV_X4 inst_5567 ( .A(net_7727), .ZN(net_2658) );
CLKBUF_X2 inst_10346 ( .A(net_8577), .Z(net_10308) );
NAND2_X1 inst_4367 ( .ZN(net_4360), .A2(net_3853), .A1(net_2210) );
OAI21_X2 inst_2013 ( .B2(net_4497), .ZN(net_4495), .B1(net_4103), .A(net_3660) );
INV_X8 inst_4506 ( .ZN(net_3817), .A(net_3260) );
NAND3_X2 inst_2756 ( .ZN(net_2345), .A3(net_1616), .A1(net_1468), .A2(net_1034) );
AOI21_X2 inst_7712 ( .B1(net_6877), .ZN(net_4093), .B2(net_2579), .A(net_2349) );
CLKBUF_X2 inst_10071 ( .A(net_9584), .Z(net_10033) );
SDFF_X2 inst_492 ( .Q(net_6839), .D(net_6839), .SI(net_3894), .SE(net_3893), .CK(net_11815) );
OAI21_X2 inst_1731 ( .ZN(net_5562), .B1(net_5414), .A(net_4828), .B2(net_4153) );
CLKBUF_X2 inst_8635 ( .A(net_8596), .Z(net_8597) );
INV_X4 inst_5414 ( .A(net_5860), .ZN(net_508) );
NAND2_X2 inst_2960 ( .ZN(net_5467), .A1(net_4902), .A2(net_4901) );
CLKBUF_X2 inst_7960 ( .A(net_7827), .Z(net_7922) );
OAI21_X2 inst_1909 ( .B1(net_5351), .ZN(net_5159), .A(net_4760), .B2(net_3941) );
CLKBUF_X2 inst_12589 ( .A(net_12550), .Z(net_12551) );
NAND2_X1 inst_4318 ( .ZN(net_4546), .A2(net_3870), .A1(net_1428) );
DFF_X1 inst_6616 ( .QN(net_7577), .D(net_5391), .CK(net_13283) );
CLKBUF_X2 inst_12292 ( .A(net_12253), .Z(net_12254) );
CLKBUF_X2 inst_11080 ( .A(net_11041), .Z(net_11042) );
XNOR2_X2 inst_82 ( .B(net_2252), .ZN(net_1335), .A(net_1334) );
NAND2_X1 inst_4335 ( .ZN(net_4392), .A2(net_3856), .A1(net_1795) );
NAND2_X2 inst_4187 ( .ZN(net_1743), .A1(net_586), .A2(net_293) );
NAND2_X1 inst_4239 ( .ZN(net_4688), .A2(net_3989), .A1(net_2114) );
CLKBUF_X2 inst_11669 ( .A(net_9070), .Z(net_11631) );
AOI22_X2 inst_7335 ( .B2(net_3439), .ZN(net_3307), .A2(net_2712), .B1(net_1227), .A1(net_148) );
CLKBUF_X2 inst_7991 ( .A(net_7951), .Z(net_7953) );
CLKBUF_X2 inst_9063 ( .A(net_8379), .Z(net_9025) );
CLKBUF_X2 inst_12171 ( .A(net_8386), .Z(net_12133) );
CLKBUF_X2 inst_8443 ( .A(net_8229), .Z(net_8405) );
SDFF_X2 inst_1121 ( .SI(net_6670), .Q(net_6670), .D(net_3787), .SE(net_3465), .CK(net_7840) );
AOI22_X2 inst_7455 ( .B2(net_7744), .A2(net_7742), .B1(net_7715), .A1(net_7713), .ZN(net_659) );
CLKBUF_X2 inst_12185 ( .A(net_12146), .Z(net_12147) );
CLKBUF_X2 inst_8932 ( .A(net_8893), .Z(net_8894) );
NAND2_X2 inst_3161 ( .ZN(net_4772), .A2(net_3941), .A1(net_2011) );
NAND2_X2 inst_3187 ( .ZN(net_4746), .A2(net_3941), .A1(net_1997) );
CLKBUF_X2 inst_11053 ( .A(net_10928), .Z(net_11015) );
SDFF_X2 inst_307 ( .SI(net_7528), .Q(net_7528), .D(net_5099), .SE(net_3988), .CK(net_9968) );
CLKBUF_X2 inst_8411 ( .A(net_8372), .Z(net_8373) );
CLKBUF_X2 inst_8292 ( .A(net_8253), .Z(net_8254) );
CLKBUF_X2 inst_10032 ( .A(net_8392), .Z(net_9994) );
CLKBUF_X2 inst_12663 ( .A(net_11394), .Z(net_12625) );
CLKBUF_X2 inst_11462 ( .A(net_11423), .Z(net_11424) );
NAND3_X2 inst_2816 ( .ZN(net_2282), .A3(net_1526), .A1(net_1437), .A2(net_942) );
OAI21_X2 inst_2034 ( .B2(net_4476), .ZN(net_4469), .B1(net_4225), .A(net_3598) );
SDFF_X2 inst_276 ( .D(net_6398), .SE(net_5801), .SI(net_343), .Q(net_343), .CK(net_14336) );
SDFF_X2 inst_717 ( .SI(net_6789), .Q(net_6789), .SE(net_3816), .D(net_3800), .CK(net_11320) );
OAI22_X2 inst_1505 ( .B1(net_4660), .A1(net_4105), .B2(net_4091), .ZN(net_4088), .A2(net_4087) );
CLKBUF_X2 inst_13380 ( .A(net_13341), .Z(net_13342) );
CLKBUF_X2 inst_10439 ( .A(net_10400), .Z(net_10401) );
NAND2_X2 inst_3339 ( .ZN(net_3569), .A1(net_3568), .A2(net_3225) );
CLKBUF_X2 inst_8460 ( .A(net_8171), .Z(net_8422) );
NAND2_X2 inst_3791 ( .A1(net_7172), .A2(net_1637), .ZN(net_1554) );
CLKBUF_X2 inst_11557 ( .A(net_11518), .Z(net_11519) );
INV_X4 inst_5297 ( .A(net_7096), .ZN(net_532) );
XNOR2_X2 inst_91 ( .ZN(net_1200), .B(net_1199), .A(net_779) );
OAI21_X2 inst_1762 ( .ZN(net_5433), .B1(net_5432), .A(net_4657), .B2(net_3993) );
OAI21_X2 inst_2023 ( .B1(net_5897), .B2(net_4497), .ZN(net_4483), .A(net_3632) );
NAND3_X2 inst_2779 ( .ZN(net_2321), .A3(net_1614), .A1(net_1406), .A2(net_1022) );
CLKBUF_X2 inst_7944 ( .A(net_7905), .Z(net_7906) );
NAND2_X2 inst_3686 ( .A2(net_1798), .ZN(net_1762), .A1(net_1761) );
NAND2_X2 inst_3842 ( .A1(net_7104), .A2(net_1675), .ZN(net_1496) );
DFF_X1 inst_6508 ( .QN(net_7430), .D(net_5515), .CK(net_12493) );
CLKBUF_X2 inst_12186 ( .A(net_12147), .Z(net_12148) );
OAI21_X2 inst_1703 ( .B2(net_5909), .ZN(net_5591), .A(net_5214), .B1(net_4080) );
INV_X4 inst_4919 ( .A(net_3814), .ZN(net_3275) );
CLKBUF_X2 inst_13250 ( .A(net_9940), .Z(net_13212) );
INV_X2 inst_5886 ( .A(net_7654), .ZN(net_2090) );
DFF_X1 inst_6566 ( .QN(net_7502), .D(net_5108), .CK(net_12091) );
INV_X4 inst_4715 ( .ZN(net_3123), .A(net_3043) );
AOI22_X2 inst_7424 ( .A1(net_2970), .B1(net_2772), .ZN(net_2768), .A2(net_241), .B2(net_167) );
CLKBUF_X2 inst_14139 ( .A(net_7950), .Z(net_14101) );
CLKBUF_X2 inst_13680 ( .A(net_13641), .Z(net_13642) );
AOI21_X2 inst_7788 ( .ZN(net_1942), .A(net_1941), .B1(net_1823), .B2(net_1233) );
CLKBUF_X2 inst_8934 ( .A(net_8895), .Z(net_8896) );
SDFF_X2 inst_614 ( .Q(net_6620), .D(net_6620), .SE(net_3830), .SI(net_3821), .CK(net_12019) );
CLKBUF_X2 inst_14079 ( .A(net_14040), .Z(net_14041) );
CLKBUF_X2 inst_11897 ( .A(net_11858), .Z(net_11859) );
DFF_X1 inst_6648 ( .QN(net_7622), .D(net_5203), .CK(net_10560) );
CLKBUF_X2 inst_9080 ( .A(net_9041), .Z(net_9042) );
CLKBUF_X2 inst_8851 ( .A(net_8812), .Z(net_8813) );
CLKBUF_X2 inst_12197 ( .A(net_10784), .Z(net_12159) );
OAI21_X2 inst_1896 ( .B1(net_5206), .ZN(net_5180), .A(net_4557), .B2(net_3866) );
SDFF_X2 inst_1031 ( .Q(net_7546), .D(net_7546), .SE(net_3896), .SI(net_380), .CK(net_13117) );
CLKBUF_X2 inst_8075 ( .A(net_8036), .Z(net_8037) );
SDFF_X2 inst_945 ( .Q(net_7235), .D(net_7235), .SE(net_3822), .SI(net_331), .CK(net_9834) );
CLKBUF_X2 inst_11187 ( .A(net_11148), .Z(net_11149) );
SDFF_X2 inst_369 ( .SI(net_7640), .Q(net_7640), .D(net_4789), .SE(net_3867), .CK(net_13247) );
DFF_X1 inst_6415 ( .QN(net_6162), .D(net_5755), .CK(net_11042) );
INV_X4 inst_5161 ( .ZN(net_682), .A(net_551) );
OAI21_X2 inst_1900 ( .B1(net_5198), .ZN(net_5175), .A(net_4553), .B2(net_3866) );
CLKBUF_X2 inst_12899 ( .A(net_12860), .Z(net_12861) );
CLKBUF_X2 inst_7984 ( .A(net_7878), .Z(net_7946) );
CLKBUF_X2 inst_12850 ( .A(net_11263), .Z(net_12812) );
DFF_X1 inst_6489 ( .QN(net_7420), .D(net_5562), .CK(net_9683) );
INV_X4 inst_5695 ( .A(net_6067), .ZN(net_3577) );
NAND2_X2 inst_2916 ( .ZN(net_5709), .A2(net_5708), .A1(net_2931) );
SDFF_X2 inst_266 ( .Q(net_6368), .SI(net_6367), .D(net_3552), .SE(net_392), .CK(net_14069) );
SDFF_X2 inst_1286 ( .D(net_3892), .SE(net_3256), .SI(net_133), .Q(net_133), .CK(net_8473) );
CLKBUF_X2 inst_9288 ( .A(net_9249), .Z(net_9250) );
OAI21_X2 inst_2051 ( .B2(net_4457), .ZN(net_4449), .B1(net_4070), .A(net_3533) );
CLKBUF_X2 inst_8382 ( .A(net_8343), .Z(net_8344) );
CLKBUF_X2 inst_8812 ( .A(net_8356), .Z(net_8774) );
SDFF_X2 inst_1198 ( .SI(net_7080), .Q(net_7080), .D(net_3783), .SE(net_3747), .CK(net_8990) );
SDFF_X2 inst_171 ( .Q(net_6243), .SI(net_6242), .D(net_3577), .SE(net_392), .CK(net_13523) );
XNOR2_X2 inst_77 ( .ZN(net_1933), .A(net_1240), .B(net_622) );
DFF_X1 inst_6399 ( .QN(net_6138), .D(net_5689), .CK(net_8172) );
CLKBUF_X2 inst_8224 ( .A(net_8185), .Z(net_8186) );
CLKBUF_X2 inst_10950 ( .A(net_10911), .Z(net_10912) );
SDFF_X2 inst_374 ( .SI(net_7647), .Q(net_7647), .D(net_4793), .SE(net_3867), .CK(net_13387) );
CLKBUF_X2 inst_12832 ( .A(net_7947), .Z(net_12794) );
XNOR2_X2 inst_103 ( .ZN(net_1919), .B(net_1142), .A(net_732) );
CLKBUF_X2 inst_13328 ( .A(net_13289), .Z(net_13290) );
NAND2_X2 inst_3690 ( .A2(net_1798), .ZN(net_1755), .A1(net_1754) );
CLKBUF_X2 inst_11710 ( .A(net_8388), .Z(net_11672) );
CLKBUF_X2 inst_10763 ( .A(net_10015), .Z(net_10725) );
DFFR_X2 inst_7086 ( .QN(net_7736), .D(net_2799), .CK(net_10522), .RN(x1822) );
CLKBUF_X2 inst_9642 ( .A(net_9603), .Z(net_9604) );
CLKBUF_X2 inst_11716 ( .A(net_9441), .Z(net_11678) );
INV_X2 inst_6061 ( .ZN(net_1119), .A(net_124) );
DFF_X1 inst_6353 ( .QN(net_6205), .D(net_5831), .CK(net_13705) );
CLKBUF_X2 inst_9905 ( .A(net_9866), .Z(net_9867) );
NAND2_X2 inst_3738 ( .A1(net_6899), .A2(net_1639), .ZN(net_1607) );
CLKBUF_X2 inst_11881 ( .A(net_11842), .Z(net_11843) );
NAND2_X4 inst_2855 ( .ZN(net_5468), .A1(net_4905), .A2(net_4904) );
CLKBUF_X2 inst_8247 ( .A(net_8208), .Z(net_8209) );
CLKBUF_X2 inst_10097 ( .A(net_9627), .Z(net_10059) );
DFF_X1 inst_6749 ( .QN(net_7634), .D(net_4846), .CK(net_13418) );
CLKBUF_X2 inst_13553 ( .A(net_13514), .Z(net_13515) );
SDFF_X2 inst_809 ( .Q(net_6983), .D(net_6983), .SE(net_3891), .SI(net_3807), .CK(net_9037) );
OAI21_X2 inst_2058 ( .ZN(net_4440), .B1(net_4439), .B2(net_4436), .A(net_3608) );
CLKBUF_X2 inst_9637 ( .A(net_9598), .Z(net_9599) );
NAND2_X2 inst_3675 ( .A2(net_1798), .ZN(net_1782), .A1(net_1781) );
AND2_X4 inst_7816 ( .ZN(net_3264), .A2(net_3154), .A1(net_587) );
SDFF_X2 inst_1234 ( .SI(net_7202), .Q(net_7202), .D(net_3883), .SE(net_3751), .CK(net_13304) );
NAND4_X2 inst_2562 ( .ZN(net_1822), .A1(net_1821), .A4(net_1820), .A2(net_1053), .A3(net_757) );
CLKBUF_X2 inst_10040 ( .A(net_10001), .Z(net_10002) );
CLKBUF_X2 inst_14245 ( .A(net_14206), .Z(net_14207) );
NOR2_X2 inst_2398 ( .A1(net_5778), .ZN(net_3930), .A2(net_286) );
CLKBUF_X2 inst_13925 ( .A(net_13886), .Z(net_13887) );
SDFF_X2 inst_1022 ( .SI(net_6490), .Q(net_6490), .SE(net_3889), .D(net_3802), .CK(net_11640) );
NAND3_X2 inst_2595 ( .ZN(net_5744), .A1(net_5639), .A2(net_5218), .A3(net_4203) );
INV_X4 inst_5614 ( .A(net_7559), .ZN(net_1872) );
CLKBUF_X2 inst_9248 ( .A(net_9209), .Z(net_9210) );
CLKBUF_X2 inst_11938 ( .A(net_11899), .Z(net_11900) );
CLKBUF_X2 inst_9400 ( .A(net_9361), .Z(net_9362) );
NOR2_X2 inst_2371 ( .ZN(net_5214), .A2(net_4615), .A1(net_4446) );
NAND2_X2 inst_2939 ( .ZN(net_5507), .A1(net_4974), .A2(net_4973) );
DFF_X1 inst_6818 ( .Q(net_5849), .D(net_3072), .CK(net_10230) );
CLKBUF_X2 inst_10416 ( .A(net_10377), .Z(net_10378) );
SDFF_X2 inst_1223 ( .SI(net_7215), .Q(net_7215), .D(net_3805), .SE(net_3751), .CK(net_11539) );
NAND3_X2 inst_2785 ( .ZN(net_2315), .A3(net_1568), .A1(net_1367), .A2(net_981) );
CLKBUF_X2 inst_13636 ( .A(net_11924), .Z(net_13598) );
NAND2_X2 inst_3906 ( .A1(net_6561), .A2(net_1705), .ZN(net_1404) );
DFF_X2 inst_6241 ( .QN(net_7380), .D(net_3033), .CK(net_9507) );
CLKBUF_X2 inst_8928 ( .A(net_8889), .Z(net_8890) );
DFF_X1 inst_6574 ( .QN(net_7564), .D(net_5080), .CK(net_13098) );
SDFF_X2 inst_681 ( .Q(net_6727), .D(net_6727), .SE(net_3815), .SI(net_3806), .CK(net_8284) );
CLKBUF_X2 inst_8657 ( .A(net_8618), .Z(net_8619) );
INV_X4 inst_5432 ( .A(net_6149), .ZN(net_3573) );
CLKBUF_X2 inst_13785 ( .A(net_12092), .Z(net_13747) );
AOI21_X2 inst_7665 ( .B2(net_5926), .ZN(net_3310), .A(net_3309), .B1(net_1212) );
INV_X4 inst_4886 ( .ZN(net_906), .A(net_882) );
CLKBUF_X2 inst_9322 ( .A(net_8008), .Z(net_9284) );
OAI21_X2 inst_2010 ( .ZN(net_4501), .B1(net_4500), .B2(net_4497), .A(net_3666) );
CLKBUF_X2 inst_13181 ( .A(net_11647), .Z(net_13143) );
CLKBUF_X2 inst_11575 ( .A(net_8074), .Z(net_11537) );
CLKBUF_X2 inst_10665 ( .A(net_10626), .Z(net_10627) );
INV_X4 inst_5547 ( .A(net_7534), .ZN(net_527) );
NAND2_X2 inst_2915 ( .ZN(net_5711), .A2(net_5710), .A1(net_2934) );
NAND2_X2 inst_3296 ( .ZN(net_3654), .A1(net_3653), .A2(net_3229) );
CLKBUF_X2 inst_9135 ( .A(net_9096), .Z(net_9097) );
SDFF_X2 inst_871 ( .SI(net_7030), .Q(net_7030), .D(net_3802), .SE(net_3777), .CK(net_11937) );
INV_X1 inst_6148 ( .A(net_3406), .ZN(net_3332) );
NAND3_X2 inst_2684 ( .ZN(net_3179), .A3(net_2980), .A2(net_1971), .A1(net_1102) );
DFF_X2 inst_6320 ( .QN(net_7822), .CK(net_8249), .D(x1358) );
DFF_X1 inst_6379 ( .QN(net_6283), .D(net_5805), .CK(net_13694) );
SDFF_X2 inst_532 ( .Q(net_6609), .D(net_6609), .SI(net_3897), .SE(net_3830), .CK(net_12041) );
DFF_X1 inst_6842 ( .D(net_2518), .Q(net_169), .CK(net_10107) );
SDFF_X2 inst_1171 ( .SI(net_6942), .Q(net_6942), .D(net_3776), .SE(net_3734), .CK(net_8837) );
NOR2_X2 inst_2382 ( .ZN(net_4804), .A2(net_4803), .A1(net_500) );
NAND2_X2 inst_2965 ( .ZN(net_5462), .A1(net_4890), .A2(net_4889) );
NAND2_X2 inst_3164 ( .ZN(net_4769), .A2(net_3941), .A1(net_2021) );
CLKBUF_X2 inst_12228 ( .A(net_12189), .Z(net_12190) );
NAND2_X2 inst_2969 ( .ZN(net_5458), .A1(net_4882), .A2(net_4881) );
INV_X4 inst_5274 ( .ZN(net_419), .A(net_418) );
INV_X4 inst_5493 ( .A(net_6017), .ZN(net_582) );
NAND2_X2 inst_3314 ( .ZN(net_3618), .A1(net_3617), .A2(net_3231) );
INV_X4 inst_5616 ( .A(net_7729), .ZN(net_2655) );
CLKBUF_X2 inst_8192 ( .A(net_8153), .Z(net_8154) );
INV_X2 inst_5766 ( .ZN(net_3021), .A(net_3020) );
NAND3_X2 inst_2594 ( .ZN(net_5745), .A1(net_5640), .A2(net_5219), .A3(net_4204) );
INV_X4 inst_5113 ( .A(net_2843), .ZN(net_605) );
CLKBUF_X2 inst_14052 ( .A(net_7906), .Z(net_14014) );
NAND2_X2 inst_4037 ( .A1(net_6658), .A2(net_1655), .ZN(net_1015) );
NAND2_X2 inst_3976 ( .ZN(net_1294), .A1(net_885), .A2(net_324) );
CLKBUF_X2 inst_13277 ( .A(net_12447), .Z(net_13239) );
CLKBUF_X2 inst_13566 ( .A(net_13111), .Z(net_13528) );
CLKBUF_X2 inst_12073 ( .A(net_12034), .Z(net_12035) );
SDFF_X2 inst_1327 ( .SE(net_6412), .Q(net_6412), .D(net_2715), .SI(net_2714), .CK(net_10197) );
CLKBUF_X2 inst_10598 ( .A(net_10559), .Z(net_10560) );
CLKBUF_X2 inst_11715 ( .A(net_11676), .Z(net_11677) );
CLKBUF_X2 inst_11773 ( .A(net_11734), .Z(net_11735) );
CLKBUF_X2 inst_9444 ( .A(net_9405), .Z(net_9406) );
SDFF_X2 inst_1119 ( .SI(net_6668), .Q(net_6668), .D(net_3811), .SE(net_3465), .CK(net_9320) );
NAND2_X2 inst_3699 ( .A1(net_6559), .ZN(net_1706), .A2(net_1705) );
INV_X4 inst_5082 ( .A(net_7794), .ZN(net_3806) );
CLKBUF_X2 inst_9684 ( .A(net_9645), .Z(net_9646) );
SDFF_X2 inst_1255 ( .SI(net_6523), .Q(net_6523), .D(net_3892), .SE(net_3756), .CK(net_8753) );
INV_X2 inst_6066 ( .A(net_7447), .ZN(net_1395) );
CLKBUF_X2 inst_9844 ( .A(net_8360), .Z(net_9806) );
INV_X4 inst_5050 ( .A(net_1145), .ZN(net_759) );
CLKBUF_X2 inst_10947 ( .A(net_10908), .Z(net_10909) );
CLKBUF_X2 inst_9279 ( .A(net_8548), .Z(net_9241) );
OAI21_X2 inst_1791 ( .ZN(net_5400), .B1(net_5399), .A(net_4674), .B2(net_3988) );
CLKBUF_X2 inst_9112 ( .A(net_9073), .Z(net_9074) );
NAND2_X2 inst_3420 ( .A2(net_5917), .ZN(net_3242), .A1(net_3241) );
INV_X4 inst_4925 ( .A(net_3793), .ZN(net_3131) );
CLKBUF_X2 inst_8834 ( .A(net_8795), .Z(net_8796) );
DFFR_X2 inst_7021 ( .D(net_3271), .QN(net_269), .CK(net_12340), .RN(x1822) );
NAND2_X1 inst_4457 ( .A2(net_1256), .ZN(net_1116), .A1(net_1115) );
INV_X16 inst_6133 ( .ZN(net_3200), .A(net_2743) );
CLKBUF_X2 inst_12341 ( .A(net_11223), .Z(net_12303) );
INV_X4 inst_5064 ( .ZN(net_715), .A(net_633) );
CLKBUF_X2 inst_11827 ( .A(net_11788), .Z(net_11789) );
SDFF_X2 inst_528 ( .Q(net_6598), .D(net_6598), .SI(net_3883), .SE(net_3830), .CK(net_12202) );
CLKBUF_X2 inst_9360 ( .A(net_9321), .Z(net_9322) );
SDFF_X2 inst_903 ( .Q(net_7107), .D(net_7107), .SE(net_3888), .SI(net_3814), .CK(net_10489) );
CLKBUF_X2 inst_13574 ( .A(net_9928), .Z(net_13536) );
CLKBUF_X2 inst_9782 ( .A(net_8881), .Z(net_9744) );
OAI21_X2 inst_1725 ( .ZN(net_5569), .B1(net_5440), .A(net_4834), .B2(net_4153) );
INV_X4 inst_5391 ( .A(net_7573), .ZN(net_1865) );
CLKBUF_X2 inst_13173 ( .A(net_11730), .Z(net_13135) );
INV_X4 inst_4957 ( .ZN(net_3048), .A(net_1216) );
CLKBUF_X2 inst_8607 ( .A(net_8568), .Z(net_8569) );
CLKBUF_X2 inst_11377 ( .A(net_10663), .Z(net_11339) );
CLKBUF_X2 inst_8602 ( .A(net_8563), .Z(net_8564) );
SDFF_X2 inst_846 ( .Q(net_7026), .D(net_7026), .SE(net_3899), .SI(net_3801), .CK(net_10989) );
INV_X2 inst_5925 ( .A(net_7315), .ZN(net_1764) );
CLKBUF_X2 inst_9700 ( .A(net_9661), .Z(net_9662) );
NAND2_X2 inst_3504 ( .A1(net_6417), .ZN(net_2687), .A2(net_2262) );
NAND2_X2 inst_3924 ( .A2(net_1696), .ZN(net_1377), .A1(net_1376) );
OAI21_X2 inst_1734 ( .ZN(net_5555), .B1(net_5554), .A(net_4813), .B2(net_4153) );
CLKBUF_X2 inst_14408 ( .A(net_14369), .Z(net_14370) );
INV_X8 inst_4510 ( .ZN(net_3871), .A(net_3168) );
DFFR_X2 inst_7036 ( .QN(net_5998), .D(net_3185), .CK(net_12561), .RN(x1822) );
INV_X4 inst_4646 ( .ZN(net_4176), .A(net_4011) );
CLKBUF_X2 inst_9548 ( .A(net_9061), .Z(net_9510) );
INV_X4 inst_4572 ( .ZN(net_5790), .A(net_5789) );
INV_X4 inst_5189 ( .ZN(net_677), .A(net_514) );
CLKBUF_X2 inst_13053 ( .A(net_13014), .Z(net_13015) );
CLKBUF_X2 inst_11203 ( .A(net_11164), .Z(net_11165) );
NAND2_X2 inst_3464 ( .A2(net_5970), .ZN(net_2884), .A1(net_2883) );
SDFF_X2 inst_1044 ( .Q(net_7244), .D(net_7244), .SE(net_3822), .SI(net_340), .CK(net_12669) );
CLKBUF_X2 inst_9233 ( .A(net_9194), .Z(net_9195) );
NAND2_X2 inst_3354 ( .ZN(net_3537), .A1(net_3536), .A2(net_3226) );
DFF_X2 inst_6187 ( .QN(net_6825), .D(net_5086), .CK(net_10800) );
CLKBUF_X2 inst_10309 ( .A(net_10270), .Z(net_10271) );
INV_X4 inst_4993 ( .A(net_788), .ZN(net_696) );
AOI222_X2 inst_7554 ( .C1(net_7668), .A1(net_7636), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1839), .B1(net_1838) );
CLKBUF_X2 inst_9509 ( .A(net_9470), .Z(net_9471) );
CLKBUF_X2 inst_14389 ( .A(net_14350), .Z(net_14351) );
CLKBUF_X2 inst_9500 ( .A(net_7850), .Z(net_9462) );
CLKBUF_X2 inst_8327 ( .A(net_8137), .Z(net_8289) );
NAND2_X2 inst_3014 ( .A1(net_6889), .A2(net_5006), .ZN(net_4995) );
CLKBUF_X2 inst_8199 ( .A(net_8115), .Z(net_8161) );
DFF_X2 inst_6256 ( .QN(net_6414), .D(net_2790), .CK(net_10212) );
SDFF_X2 inst_227 ( .Q(net_6327), .SI(net_6326), .D(net_3631), .SE(net_392), .CK(net_14027) );
OAI22_X2 inst_1532 ( .B1(net_4637), .ZN(net_4034), .A2(net_4033), .B2(net_4032), .A1(net_4030) );
NAND2_X1 inst_4303 ( .ZN(net_4563), .A2(net_3866), .A1(net_1844) );
INV_X2 inst_5861 ( .A(net_818), .ZN(net_599) );
OAI21_X2 inst_2136 ( .ZN(net_2821), .B1(net_2820), .A(net_2707), .B2(net_2454) );
NAND3_X2 inst_2718 ( .ZN(net_2457), .A2(net_1814), .A3(net_1594), .A1(net_1506) );
NAND2_X4 inst_2891 ( .ZN(net_4030), .A2(net_3322), .A1(net_3106) );
NAND2_X2 inst_3927 ( .A1(net_6846), .A2(net_1521), .ZN(net_1371) );
XNOR2_X2 inst_58 ( .B(net_4152), .ZN(net_1927), .A(net_1689) );
CLKBUF_X2 inst_11653 ( .A(net_11614), .Z(net_11615) );
CLKBUF_X2 inst_9574 ( .A(net_9535), .Z(net_9536) );
NAND2_X2 inst_3633 ( .ZN(net_1950), .A1(net_1298), .A2(net_1262) );
AOI222_X2 inst_7557 ( .A1(net_7394), .ZN(net_5537), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_357), .C2(net_355) );
CLKBUF_X2 inst_8642 ( .A(net_8598), .Z(net_8604) );
INV_X2 inst_6036 ( .A(net_7594), .ZN(net_1465) );
CLKBUF_X2 inst_9775 ( .A(net_9736), .Z(net_9737) );
CLKBUF_X2 inst_13792 ( .A(net_13753), .Z(net_13754) );
OAI22_X2 inst_1469 ( .B2(net_5043), .ZN(net_4393), .A1(net_4137), .A2(net_3824), .B1(net_1170) );
CLKBUF_X2 inst_12056 ( .A(net_12017), .Z(net_12018) );
CLKBUF_X2 inst_10295 ( .A(net_10256), .Z(net_10257) );
CLKBUF_X2 inst_9944 ( .A(net_9905), .Z(net_9906) );
INV_X4 inst_5029 ( .A(net_7823), .ZN(net_3801) );
CLKBUF_X2 inst_12878 ( .A(net_9058), .Z(net_12840) );
INV_X4 inst_5690 ( .A(net_7731), .ZN(net_2952) );
CLKBUF_X2 inst_10200 ( .A(net_10161), .Z(net_10162) );
CLKBUF_X2 inst_9592 ( .A(net_9553), .Z(net_9554) );
SDFF_X2 inst_581 ( .Q(net_6560), .D(net_6560), .SE(net_3823), .SI(net_3806), .CK(net_9351) );
NOR2_X2 inst_2551 ( .A1(net_6001), .A2(net_5995), .ZN(net_2891) );
INV_X4 inst_5288 ( .A(net_6692), .ZN(net_587) );
XNOR2_X2 inst_28 ( .ZN(net_2566), .B(net_2565), .A(net_2445) );
NAND2_X1 inst_4407 ( .A2(net_3087), .ZN(net_2910), .A1(net_2828) );
NOR2_X2 inst_2424 ( .A2(net_5891), .ZN(net_3225), .A1(net_3224) );
INV_X8 inst_4517 ( .ZN(net_3471), .A(net_3118) );
CLKBUF_X2 inst_9410 ( .A(net_8541), .Z(net_9372) );
CLKBUF_X2 inst_12656 ( .A(net_12617), .Z(net_12618) );
CLKBUF_X2 inst_9434 ( .A(net_9395), .Z(net_9396) );
CLKBUF_X2 inst_13719 ( .A(net_8034), .Z(net_13681) );
CLKBUF_X2 inst_9401 ( .A(net_9362), .Z(net_9363) );
AOI22_X2 inst_7440 ( .ZN(net_4851), .A2(net_1228), .B1(net_1226), .B2(net_385), .A1(net_373) );
NAND2_X2 inst_3144 ( .ZN(net_4819), .A2(net_4153), .A1(net_1983) );
CLKBUF_X2 inst_13386 ( .A(net_13347), .Z(net_13348) );
SDFF_X2 inst_592 ( .Q(net_6590), .D(net_6590), .SE(net_3823), .SI(net_3800), .CK(net_9182) );
INV_X16 inst_6124 ( .ZN(net_4925), .A(net_4262) );
AOI22_X2 inst_7289 ( .B1(net_7226), .A1(net_7194), .A2(net_5244), .B2(net_5243), .ZN(net_5216) );
CLKBUF_X2 inst_13841 ( .A(net_8549), .Z(net_13803) );
CLKBUF_X2 inst_11530 ( .A(net_11491), .Z(net_11492) );
SDFF_X2 inst_993 ( .Q(net_6480), .D(net_6480), .SE(net_3904), .SI(net_3796), .CK(net_10838) );
NAND2_X2 inst_3666 ( .A2(net_1798), .ZN(net_1794), .A1(net_1793) );
INV_X4 inst_5143 ( .ZN(net_784), .A(net_573) );
INV_X4 inst_5177 ( .ZN(net_618), .A(net_529) );
DFF_X1 inst_6407 ( .QN(net_6154), .D(net_5763), .CK(net_8256) );
AOI22_X2 inst_7264 ( .B1(net_6955), .A1(net_6923), .A2(net_5298), .B2(net_5297), .ZN(net_5290) );
CLKBUF_X2 inst_13855 ( .A(net_13816), .Z(net_13817) );
CLKBUF_X2 inst_13504 ( .A(net_10406), .Z(net_13466) );
AND2_X2 inst_7858 ( .ZN(net_2273), .A1(net_2272), .A2(net_2271) );
CLKBUF_X2 inst_12876 ( .A(net_12837), .Z(net_12838) );
INV_X4 inst_5096 ( .A(net_7811), .ZN(net_3897) );
SDFF_X2 inst_630 ( .SI(net_6642), .Q(net_6642), .SE(net_3851), .D(net_3784), .CK(net_9154) );
NAND2_X2 inst_3948 ( .A1(net_6431), .A2(net_1677), .ZN(net_1340) );
INV_X4 inst_5535 ( .ZN(net_1219), .A(x1155) );
CLKBUF_X2 inst_11413 ( .A(net_11374), .Z(net_11375) );
INV_X4 inst_5227 ( .ZN(net_3227), .A(net_462) );
CLKBUF_X2 inst_14157 ( .A(net_14118), .Z(net_14119) );
INV_X4 inst_5268 ( .ZN(net_3147), .A(net_539) );
CLKBUF_X2 inst_11796 ( .A(net_11757), .Z(net_11758) );
CLKBUF_X2 inst_9662 ( .A(net_8531), .Z(net_9624) );
SDFF_X2 inst_1273 ( .D(net_6388), .SE(net_5799), .SI(net_373), .Q(net_373), .CK(net_14205) );
CLKBUF_X2 inst_12791 ( .A(net_12752), .Z(net_12753) );
CLKBUF_X2 inst_11337 ( .A(net_11298), .Z(net_11299) );
SDFF_X2 inst_512 ( .SI(net_6779), .Q(net_6779), .SE(net_3872), .D(net_3836), .CK(net_8382) );
CLKBUF_X2 inst_11808 ( .A(net_9108), .Z(net_11770) );
INV_X4 inst_4966 ( .ZN(net_2489), .A(net_708) );
SDFF_X2 inst_1301 ( .SE(net_7529), .Q(net_7529), .D(net_2994), .SI(net_2993), .CK(net_12578) );
CLKBUF_X2 inst_14307 ( .A(net_14268), .Z(net_14269) );
CLKBUF_X2 inst_12278 ( .A(net_11262), .Z(net_12240) );
OAI21_X2 inst_2151 ( .B1(net_5778), .ZN(net_2793), .A(net_2659), .B2(net_2657) );
CLKBUF_X2 inst_14109 ( .A(net_14070), .Z(net_14071) );
SDFF_X2 inst_647 ( .D(net_7802), .SI(net_6632), .Q(net_6632), .SE(net_3851), .CK(net_9149) );
NAND3_X2 inst_2830 ( .A1(net_2382), .A2(net_2299), .ZN(net_1154), .A3(net_460) );
NAND2_X2 inst_3054 ( .A1(net_7154), .A2(net_4954), .ZN(net_4952) );
CLKBUF_X2 inst_12871 ( .A(net_9155), .Z(net_12833) );
CLKBUF_X2 inst_11744 ( .A(net_11705), .Z(net_11706) );
INV_X4 inst_4764 ( .ZN(net_2425), .A(net_1940) );
INV_X4 inst_5137 ( .ZN(net_792), .A(net_578) );
CLKBUF_X2 inst_13271 ( .A(net_10897), .Z(net_13233) );
NAND2_X2 inst_2985 ( .A1(net_6752), .A2(net_5033), .ZN(net_5026) );
CLKBUF_X2 inst_9821 ( .A(net_9782), .Z(net_9783) );
CLKBUF_X2 inst_8156 ( .A(net_8117), .Z(net_8118) );
SDFF_X2 inst_833 ( .Q(net_7012), .D(net_7012), .SE(net_3899), .SI(net_3809), .CK(net_11902) );
NAND2_X2 inst_3772 ( .A1(net_6898), .A2(net_1639), .ZN(net_1573) );
NAND2_X2 inst_4210 ( .A2(net_6009), .A1(net_6008), .ZN(net_3241) );
CLKBUF_X2 inst_11968 ( .A(net_11929), .Z(net_11930) );
SDFF_X2 inst_960 ( .Q(net_6437), .D(net_6437), .SE(net_3820), .SI(net_3811), .CK(net_8646) );
OAI21_X2 inst_2043 ( .ZN(net_4459), .B1(net_4458), .B2(net_4457), .A(net_3712) );
XNOR2_X2 inst_118 ( .ZN(net_5864), .B(net_1655), .A(net_823) );
INV_X4 inst_4924 ( .A(net_3812), .ZN(net_3289) );
NOR2_X2 inst_2411 ( .A1(net_6008), .ZN(net_3412), .A2(net_3406) );
CLKBUF_X2 inst_12709 ( .A(net_10494), .Z(net_12671) );
CLKBUF_X2 inst_14433 ( .A(net_14394), .Z(net_14395) );
CLKBUF_X2 inst_10781 ( .A(net_10742), .Z(net_10743) );
XNOR2_X2 inst_38 ( .ZN(net_2444), .A(net_1686), .B(net_535) );
DFF_X1 inst_6591 ( .QN(net_7561), .D(net_5059), .CK(net_10584) );
SDFF_X2 inst_381 ( .SI(net_7676), .Q(net_7676), .D(net_4786), .SE(net_3866), .CK(net_7983) );
OAI21_X2 inst_2037 ( .B1(net_4598), .B2(net_4476), .ZN(net_4466), .A(net_3574) );
NAND3_X2 inst_2601 ( .ZN(net_5738), .A1(net_5633), .A2(net_5185), .A3(net_4198) );
CLKBUF_X2 inst_8578 ( .A(net_7886), .Z(net_8540) );
CLKBUF_X2 inst_13532 ( .A(net_13493), .Z(net_13494) );
CLKBUF_X2 inst_9448 ( .A(net_9409), .Z(net_9410) );
DFF_X1 inst_6930 ( .D(net_2402), .Q(net_247), .CK(net_10414) );
CLKBUF_X2 inst_9102 ( .A(net_8555), .Z(net_9064) );
NAND2_X2 inst_3837 ( .A1(net_6426), .A2(net_1677), .ZN(net_1502) );
CLKBUF_X2 inst_12276 ( .A(net_12237), .Z(net_12238) );
SDFF_X2 inst_883 ( .SI(net_7807), .Q(net_7113), .D(net_7113), .SE(net_3888), .CK(net_12155) );
DFF_X1 inst_6876 ( .D(net_2497), .Q(net_164), .CK(net_12233) );
AOI222_X2 inst_7577 ( .A1(net_7542), .ZN(net_5202), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_374), .C2(net_372) );
CLKBUF_X2 inst_12536 ( .A(net_12497), .Z(net_12498) );
CLKBUF_X2 inst_13108 ( .A(net_9536), .Z(net_13070) );
CLKBUF_X2 inst_12710 ( .A(net_10578), .Z(net_12672) );
CLKBUF_X2 inst_10355 ( .A(net_10316), .Z(net_10317) );
SDFF_X2 inst_756 ( .Q(net_6878), .D(net_6878), .SE(net_3901), .SI(net_3808), .CK(net_11736) );
CLKBUF_X2 inst_8068 ( .A(net_8029), .Z(net_8030) );
INV_X4 inst_5496 ( .A(net_7277), .ZN(net_2027) );
CLKBUF_X2 inst_13880 ( .A(net_13841), .Z(net_13842) );
INV_X2 inst_6002 ( .A(net_7435), .ZN(net_1452) );
CLKBUF_X2 inst_13423 ( .A(net_13384), .Z(net_13385) );
CLKBUF_X2 inst_10228 ( .A(net_10189), .Z(net_10190) );
CLKBUF_X2 inst_9270 ( .A(net_9231), .Z(net_9232) );
SDFF_X2 inst_1188 ( .D(net_7802), .SI(net_6934), .Q(net_6934), .SE(net_3734), .CK(net_11769) );
INV_X4 inst_4597 ( .ZN(net_5050), .A(net_4292) );
INV_X4 inst_5503 ( .A(net_7275), .ZN(net_2029) );
CLKBUF_X2 inst_9873 ( .A(net_7877), .Z(net_9835) );
CLKBUF_X2 inst_9685 ( .A(net_9108), .Z(net_9647) );
SDFF_X2 inst_1165 ( .SI(net_6925), .Q(net_6925), .D(net_3792), .SE(net_3734), .CK(net_8914) );
INV_X4 inst_5439 ( .A(net_7420), .ZN(net_2142) );
CLKBUF_X2 inst_11029 ( .A(net_10990), .Z(net_10991) );
CLKBUF_X2 inst_8891 ( .A(net_7834), .Z(net_8853) );
NAND3_X2 inst_2644 ( .ZN(net_5947), .A3(net_3965), .A2(net_1969), .A1(net_810) );
DFF_X1 inst_6922 ( .D(net_2405), .Q(net_259), .CK(net_12394) );
NAND3_X2 inst_2626 ( .ZN(net_5703), .A1(net_5680), .A2(net_5314), .A3(net_4254) );
CLKBUF_X2 inst_13462 ( .A(net_13423), .Z(net_13424) );
CLKBUF_X2 inst_9960 ( .A(net_9921), .Z(net_9922) );
CLKBUF_X2 inst_9314 ( .A(net_8790), .Z(net_9276) );
INV_X4 inst_4629 ( .ZN(net_4193), .A(net_4046) );
DFFR_X2 inst_6957 ( .QN(net_7734), .D(net_5779), .CK(net_10536), .RN(x1822) );
CLKBUF_X2 inst_8966 ( .A(net_8927), .Z(net_8928) );
CLKBUF_X2 inst_14140 ( .A(net_14101), .Z(net_14102) );
INV_X2 inst_5983 ( .A(net_7469), .ZN(net_2120) );
CLKBUF_X2 inst_9056 ( .A(net_9017), .Z(net_9018) );
CLKBUF_X2 inst_8363 ( .A(net_8324), .Z(net_8325) );
NAND2_X2 inst_3873 ( .A2(net_1696), .ZN(net_1449), .A1(net_1448) );
DFF_X1 inst_6883 ( .Q(net_6416), .D(net_2491), .CK(net_14385) );
SDFF_X2 inst_992 ( .Q(net_6479), .D(net_6479), .SE(net_3904), .SI(net_3803), .CK(net_8065) );
SDFF_X2 inst_488 ( .Q(net_7102), .D(net_7102), .SI(net_3892), .SE(net_3888), .CK(net_10507) );
CLKBUF_X2 inst_14085 ( .A(net_8049), .Z(net_14047) );
AND2_X4 inst_7809 ( .ZN(net_3842), .A2(net_3841), .A1(net_1143) );
SDFF_X2 inst_387 ( .SI(net_7306), .Q(net_7306), .D(net_4780), .SE(net_3859), .CK(net_9407) );
INV_X4 inst_5196 ( .A(net_572), .ZN(net_504) );
CLKBUF_X2 inst_8666 ( .A(net_8268), .Z(net_8628) );
AOI22_X2 inst_7308 ( .B1(net_6681), .A1(net_6649), .A2(net_5139), .B2(net_5138), .ZN(net_5135) );
SDFF_X2 inst_254 ( .SI(net_6379), .Q(net_6340), .D(net_3615), .SE(net_392), .CK(net_13502) );
INV_X2 inst_6053 ( .A(net_7498), .ZN(net_2180) );
INV_X4 inst_4601 ( .ZN(net_4243), .A(net_4106) );
CLKBUF_X2 inst_9543 ( .A(net_8042), .Z(net_9505) );
CLKBUF_X2 inst_12784 ( .A(net_12745), .Z(net_12746) );
CLKBUF_X2 inst_8801 ( .A(net_8085), .Z(net_8763) );
OAI21_X2 inst_2129 ( .B2(net_5915), .ZN(net_2960), .B1(net_2959), .A(net_2758) );
OR2_X2 inst_1412 ( .A1(net_6420), .ZN(net_1071), .A2(net_807) );
INV_X2 inst_5750 ( .ZN(net_3913), .A(net_3739) );
CLKBUF_X2 inst_11273 ( .A(net_9907), .Z(net_11235) );
CLKBUF_X2 inst_9862 ( .A(net_9753), .Z(net_9824) );
SDFF_X2 inst_1181 ( .SI(net_6954), .Q(net_6954), .D(net_3821), .SE(net_3741), .CK(net_11685) );
CLKBUF_X2 inst_10957 ( .A(net_9714), .Z(net_10919) );
CLKBUF_X2 inst_8986 ( .A(net_8947), .Z(net_8948) );
HA_X1 inst_6165 ( .S(net_1710), .CO(net_1709), .B(net_1222), .A(net_906) );
CLKBUF_X2 inst_13364 ( .A(net_13325), .Z(net_13326) );
CLKBUF_X2 inst_12774 ( .A(net_11484), .Z(net_12736) );
INV_X4 inst_5045 ( .A(net_3241), .ZN(net_648) );
SDFF_X2 inst_661 ( .Q(net_6720), .D(net_6720), .SE(net_3871), .SI(net_3790), .CK(net_10924) );
DFF_X2 inst_6265 ( .QN(net_5982), .D(net_2641), .CK(net_12532) );
AOI22_X2 inst_7416 ( .B1(net_5939), .ZN(net_2778), .A1(net_2777), .B2(net_219), .A2(net_182) );
OAI22_X2 inst_1548 ( .B2(net_3405), .A2(net_3360), .ZN(net_3357), .A1(net_3299), .B1(net_434) );
CLKBUF_X2 inst_10817 ( .A(net_7985), .Z(net_10779) );
OAI21_X2 inst_2073 ( .B1(net_5911), .B2(net_4436), .ZN(net_4420), .A(net_3529) );
AOI22_X2 inst_7346 ( .B1(net_3857), .B2(net_3105), .ZN(net_3104), .A2(net_2712), .A1(net_1115) );
CLKBUF_X2 inst_9913 ( .A(net_9874), .Z(net_9875) );
CLKBUF_X2 inst_8661 ( .A(net_7864), .Z(net_8623) );
CLKBUF_X2 inst_11418 ( .A(net_8656), .Z(net_11380) );
CLKBUF_X2 inst_14255 ( .A(net_10074), .Z(net_14217) );
CLKBUF_X2 inst_9457 ( .A(net_9418), .Z(net_9419) );
NAND2_X2 inst_3984 ( .ZN(net_1286), .A1(net_885), .A2(net_313) );
INV_X4 inst_4682 ( .ZN(net_3378), .A(net_3377) );
DFFR_X2 inst_7013 ( .D(net_3288), .QN(net_283), .CK(net_12866), .RN(x1822) );
CLKBUF_X2 inst_11310 ( .A(net_11271), .Z(net_11272) );
SDFF_X2 inst_419 ( .D(net_6391), .SE(net_5800), .SI(net_356), .Q(net_356), .CK(net_14149) );
CLKBUF_X2 inst_10899 ( .A(net_10860), .Z(net_10861) );
AOI222_X2 inst_7488 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2112), .A1(net_2111), .B1(net_2110), .C1(net_2109) );
CLKBUF_X2 inst_12546 ( .A(net_12507), .Z(net_12508) );
CLKBUF_X2 inst_12098 ( .A(net_12059), .Z(net_12060) );
INV_X2 inst_5715 ( .ZN(net_4251), .A(net_4123) );
DFF_X1 inst_6495 ( .QN(net_7407), .D(net_5546), .CK(net_9304) );
CLKBUF_X2 inst_8470 ( .A(net_8431), .Z(net_8432) );
DFF_X1 inst_6941 ( .Q(net_7792), .D(net_7790), .CK(net_12388) );
CLKBUF_X2 inst_10462 ( .A(net_10423), .Z(net_10424) );
AND3_X4 inst_7799 ( .A3(net_2590), .ZN(net_1229), .A1(net_708), .A2(net_624) );
CLKBUF_X2 inst_10629 ( .A(net_10590), .Z(net_10591) );
CLKBUF_X2 inst_14298 ( .A(net_11630), .Z(net_14260) );
CLKBUF_X2 inst_14283 ( .A(net_14244), .Z(net_14245) );
CLKBUF_X2 inst_12018 ( .A(net_11979), .Z(net_11980) );
CLKBUF_X2 inst_12377 ( .A(net_9860), .Z(net_12339) );
CLKBUF_X2 inst_7898 ( .A(net_7859), .Z(net_7860) );
INV_X4 inst_5130 ( .A(net_1657), .ZN(net_689) );
CLKBUF_X2 inst_12749 ( .A(net_9591), .Z(net_12711) );
CLKBUF_X2 inst_11160 ( .A(net_11121), .Z(net_11122) );
XNOR2_X2 inst_34 ( .ZN(net_2475), .A(net_2474), .B(net_914) );
NAND2_X2 inst_3717 ( .A1(net_7166), .A2(net_1637), .ZN(net_1629) );
CLKBUF_X2 inst_9120 ( .A(net_9081), .Z(net_9082) );
XNOR2_X2 inst_12 ( .A(net_4138), .ZN(net_3824), .B(net_722) );
CLKBUF_X2 inst_12690 ( .A(net_12651), .Z(net_12652) );
CLKBUF_X2 inst_9823 ( .A(net_9784), .Z(net_9785) );
INV_X4 inst_5489 ( .A(net_7253), .ZN(net_2009) );
CLKBUF_X2 inst_13946 ( .A(net_12341), .Z(net_13908) );
AOI21_X2 inst_7765 ( .B1(net_7133), .ZN(net_5898), .B2(net_2582), .A(net_2317) );
CLKBUF_X2 inst_9856 ( .A(net_9561), .Z(net_9818) );
CLKBUF_X2 inst_9760 ( .A(net_9721), .Z(net_9722) );
CLKBUF_X2 inst_8682 ( .A(net_8643), .Z(net_8644) );
OR2_X2 inst_1424 ( .A2(net_7093), .A1(net_7092), .ZN(net_621) );
INV_X4 inst_5290 ( .A(net_6962), .ZN(net_525) );
CLKBUF_X2 inst_10239 ( .A(net_10200), .Z(net_10201) );
OR2_X2 inst_1425 ( .A2(net_6958), .A1(net_6957), .ZN(net_675) );
CLKBUF_X2 inst_8585 ( .A(net_8546), .Z(net_8547) );
NOR2_X2 inst_2307 ( .A2(net_6207), .A1(net_5840), .ZN(net_5834) );
NOR3_X2 inst_2198 ( .ZN(net_3451), .A3(net_3156), .A2(net_3009), .A1(net_2862) );
CLKBUF_X2 inst_11611 ( .A(net_11572), .Z(net_11573) );
SDFF_X2 inst_258 ( .Q(net_6376), .SI(net_6375), .D(net_3564), .SE(net_392), .CK(net_13961) );
NAND3_X2 inst_2611 ( .ZN(net_5728), .A1(net_5623), .A2(net_5145), .A3(net_4188) );
CLKBUF_X2 inst_13469 ( .A(net_13430), .Z(net_13431) );
INV_X4 inst_5004 ( .A(net_7813), .ZN(net_3805) );
CLKBUF_X2 inst_9926 ( .A(net_7944), .Z(net_9888) );
NOR2_X2 inst_2405 ( .ZN(net_3759), .A1(net_3758), .A2(net_3757) );
CLKBUF_X2 inst_13126 ( .A(net_13087), .Z(net_13088) );
NAND2_X2 inst_2994 ( .A1(net_6724), .A2(net_5031), .ZN(net_5017) );
NAND2_X2 inst_3023 ( .A1(net_6849), .A2(net_5004), .ZN(net_4986) );
SDFF_X2 inst_1243 ( .SI(net_6538), .Q(net_6538), .D(net_3897), .SE(net_3756), .CK(net_8827) );
CLKBUF_X2 inst_13155 ( .A(net_13116), .Z(net_13117) );
CLKBUF_X2 inst_13074 ( .A(net_13035), .Z(net_13036) );
CLKBUF_X2 inst_9512 ( .A(net_9473), .Z(net_9474) );
NAND2_X2 inst_3076 ( .A1(net_6446), .ZN(net_4929), .A2(net_4925) );
CLKBUF_X2 inst_10964 ( .A(net_10925), .Z(net_10926) );
SDFF_X2 inst_482 ( .Q(net_6971), .D(net_6971), .SE(net_3891), .SI(net_3890), .CK(net_8101) );
CLKBUF_X2 inst_10514 ( .A(net_10475), .Z(net_10476) );
CLKBUF_X2 inst_9804 ( .A(net_9732), .Z(net_9766) );
NAND2_X2 inst_3534 ( .ZN(net_2533), .A2(net_2082), .A1(net_1520) );
NAND2_X2 inst_3276 ( .ZN(net_3694), .A1(net_3693), .A2(net_3231) );
INV_X2 inst_5958 ( .A(net_7324), .ZN(net_1774) );
CLKBUF_X2 inst_10230 ( .A(net_10191), .Z(net_10192) );
SDFF_X2 inst_1093 ( .SI(net_6927), .Q(net_6927), .D(net_3802), .SE(net_3741), .CK(net_11780) );
NAND2_X2 inst_3996 ( .A2(net_1910), .ZN(net_1192), .A1(net_1191) );
DFFR_X2 inst_7059 ( .QN(net_6040), .D(net_3090), .CK(net_12853), .RN(x1822) );
SDFF_X2 inst_539 ( .Q(net_6580), .D(net_6580), .SI(net_3900), .SE(net_3823), .CK(net_12195) );
AOI21_X2 inst_7646 ( .B2(net_5849), .ZN(net_3753), .A(net_1930), .B1(x38) );
CLKBUF_X2 inst_12915 ( .A(net_8775), .Z(net_12877) );
CLKBUF_X2 inst_11066 ( .A(net_10681), .Z(net_11028) );
SDFF_X2 inst_895 ( .Q(net_7127), .D(net_7127), .SE(net_3888), .SI(net_3793), .CK(net_11864) );
CLKBUF_X2 inst_11042 ( .A(net_11003), .Z(net_11004) );
CLKBUF_X2 inst_10054 ( .A(net_10015), .Z(net_10016) );
CLKBUF_X2 inst_10707 ( .A(net_9559), .Z(net_10669) );
OR2_X2 inst_1430 ( .A2(net_6405), .A1(net_6404), .ZN(net_938) );
NAND2_X2 inst_3271 ( .ZN(net_3704), .A1(net_3703), .A2(net_3231) );
NAND2_X2 inst_3257 ( .A2(net_3869), .ZN(net_3866), .A1(net_1649) );
CLKBUF_X2 inst_10759 ( .A(net_10720), .Z(net_10721) );
DFF_X1 inst_6583 ( .QN(net_7553), .D(net_5067), .CK(net_10315) );
CLKBUF_X2 inst_14081 ( .A(net_14042), .Z(net_14043) );
CLKBUF_X2 inst_11498 ( .A(net_8077), .Z(net_11460) );
CLKBUF_X2 inst_10034 ( .A(net_9995), .Z(net_9996) );
NOR2_X2 inst_2341 ( .A2(net_6036), .A1(net_5778), .ZN(net_5712) );
INV_X4 inst_5526 ( .A(net_6158), .ZN(net_3603) );
CLKBUF_X2 inst_10685 ( .A(net_10646), .Z(net_10647) );
CLKBUF_X2 inst_10616 ( .A(net_10577), .Z(net_10578) );
CLKBUF_X2 inst_9979 ( .A(net_9639), .Z(net_9941) );
NAND2_X2 inst_4122 ( .A2(net_1222), .ZN(net_1169), .A1(net_342) );
CLKBUF_X2 inst_12557 ( .A(net_11154), .Z(net_12519) );
SDFF_X2 inst_763 ( .Q(net_6887), .D(net_6887), .SE(net_3901), .SI(net_3795), .CK(net_11481) );
NOR2_X2 inst_2330 ( .A2(net_6288), .A1(net_5840), .ZN(net_5811) );
AOI22_X2 inst_7377 ( .B1(net_7740), .A1(net_7711), .A2(net_5916), .B2(net_2957), .ZN(net_2944) );
NAND2_X2 inst_3636 ( .ZN(net_1947), .A1(net_1284), .A2(net_1258) );
CLKBUF_X2 inst_13184 ( .A(net_13145), .Z(net_13146) );
CLKBUF_X2 inst_11069 ( .A(net_11030), .Z(net_11031) );
CLKBUF_X2 inst_14018 ( .A(net_13979), .Z(net_13980) );
CLKBUF_X2 inst_9901 ( .A(net_9862), .Z(net_9863) );
CLKBUF_X2 inst_10324 ( .A(net_10057), .Z(net_10286) );
CLKBUF_X2 inst_13754 ( .A(net_13715), .Z(net_13716) );
CLKBUF_X2 inst_9189 ( .A(net_9150), .Z(net_9151) );
SDFF_X2 inst_537 ( .Q(net_6562), .D(net_6562), .SI(net_3892), .SE(net_3823), .CK(net_10058) );
INV_X4 inst_4797 ( .ZN(net_5103), .A(net_1260) );
INV_X2 inst_6082 ( .A(net_7650), .ZN(net_2147) );
CLKBUF_X2 inst_8482 ( .A(net_8443), .Z(net_8444) );
SDFF_X2 inst_826 ( .SI(net_7802), .Q(net_6973), .D(net_6973), .SE(net_3891), .CK(net_11950) );
CLKBUF_X2 inst_9343 ( .A(net_9094), .Z(net_9305) );
NAND2_X2 inst_4002 ( .ZN(net_1282), .A1(net_665), .A2(net_611) );
INV_X4 inst_5069 ( .A(net_3147), .ZN(net_699) );
CLKBUF_X2 inst_14009 ( .A(net_13970), .Z(net_13971) );
CLKBUF_X2 inst_10362 ( .A(net_10323), .Z(net_10324) );
SDFF_X2 inst_159 ( .Q(net_6255), .SI(net_6254), .D(net_3548), .SE(net_392), .CK(net_13538) );
DFFR_X2 inst_7042 ( .QN(net_6006), .D(net_3127), .CK(net_11427), .RN(x1822) );
CLKBUF_X2 inst_13220 ( .A(net_13181), .Z(net_13182) );
CLKBUF_X2 inst_9572 ( .A(net_9533), .Z(net_9534) );
CLKBUF_X2 inst_14341 ( .A(net_14302), .Z(net_14303) );
INV_X2 inst_5759 ( .ZN(net_3036), .A(net_2995) );
CLKBUF_X2 inst_13657 ( .A(net_13618), .Z(net_13619) );
CLKBUF_X2 inst_11005 ( .A(net_10966), .Z(net_10967) );
CLKBUF_X2 inst_10786 ( .A(net_9837), .Z(net_10748) );
CLKBUF_X2 inst_8431 ( .A(net_8344), .Z(net_8393) );
DFF_X2 inst_6318 ( .QN(net_7798), .CK(net_10942), .D(x1557) );
AOI22_X2 inst_7379 ( .B1(net_7742), .A1(net_7713), .A2(net_5916), .B2(net_2957), .ZN(net_2942) );
CLKBUF_X2 inst_8863 ( .A(net_8824), .Z(net_8825) );
NAND2_X2 inst_3950 ( .A1(net_6980), .A2(net_1833), .ZN(net_1338) );
NAND2_X1 inst_4288 ( .ZN(net_4579), .A2(net_3867), .A1(net_1188) );
SDFF_X2 inst_869 ( .SI(net_7056), .Q(net_7056), .SE(net_3818), .D(net_3788), .CK(net_8212) );
CLKBUF_X2 inst_10671 ( .A(net_10632), .Z(net_10633) );
CLKBUF_X2 inst_8339 ( .A(net_8300), .Z(net_8301) );
XNOR2_X2 inst_19 ( .ZN(net_2615), .A(net_2255), .B(net_1209) );
NAND3_X2 inst_2646 ( .ZN(net_5951), .A3(net_3961), .A2(net_1960), .A1(net_701) );
CLKBUF_X2 inst_13623 ( .A(net_13584), .Z(net_13585) );
CLKBUF_X2 inst_11509 ( .A(net_10414), .Z(net_11471) );
CLKBUF_X2 inst_10378 ( .A(net_10339), .Z(net_10340) );
CLKBUF_X2 inst_13599 ( .A(net_13560), .Z(net_13561) );
DFF_X1 inst_6543 ( .QN(net_7360), .D(net_5329), .CK(net_13016) );
CLKBUF_X2 inst_13229 ( .A(net_10259), .Z(net_13191) );
CLKBUF_X2 inst_9753 ( .A(net_8632), .Z(net_9715) );
NAND2_X1 inst_4268 ( .ZN(net_4649), .A2(net_3993), .A1(net_1471) );
CLKBUF_X2 inst_14170 ( .A(net_14131), .Z(net_14132) );
NAND2_X2 inst_3830 ( .A1(net_7114), .A2(net_1675), .ZN(net_1511) );
CLKBUF_X2 inst_13649 ( .A(net_11683), .Z(net_13611) );
CLKBUF_X2 inst_9849 ( .A(net_7908), .Z(net_9811) );
NAND2_X2 inst_3267 ( .ZN(net_3712), .A1(net_3711), .A2(net_3225) );
CLKBUF_X2 inst_12287 ( .A(net_9446), .Z(net_12249) );
OAI21_X2 inst_1686 ( .ZN(net_5779), .B1(net_5778), .A(net_5713), .B2(net_5712) );
NAND2_X2 inst_3205 ( .ZN(net_4721), .A2(net_3986), .A1(net_1909) );
CLKBUF_X2 inst_14315 ( .A(net_14276), .Z(net_14277) );
CLKBUF_X2 inst_10541 ( .A(net_10502), .Z(net_10503) );
INV_X2 inst_6048 ( .A(net_7664), .ZN(net_1854) );
CLKBUF_X2 inst_8945 ( .A(net_8906), .Z(net_8907) );
SDFF_X2 inst_612 ( .Q(net_6618), .D(net_6618), .SE(net_3830), .SI(net_3794), .CK(net_12027) );
CLKBUF_X2 inst_12505 ( .A(net_12466), .Z(net_12467) );
OAI21_X2 inst_1789 ( .B1(net_5434), .ZN(net_5402), .A(net_4676), .B2(net_3988) );
OAI21_X2 inst_1692 ( .ZN(net_5602), .A(net_5304), .B2(net_4521), .B1(net_4132) );
DFF_X2 inst_6185 ( .QN(net_6689), .D(net_5384), .CK(net_9726) );
NAND2_X2 inst_3986 ( .ZN(net_1284), .A1(net_885), .A2(net_325) );
AOI21_X4 inst_7627 ( .B1(net_7000), .ZN(net_4619), .A(net_2460), .B2(net_1100) );
CLKBUF_X2 inst_9437 ( .A(net_8099), .Z(net_9399) );
NAND2_X2 inst_3441 ( .ZN(net_3168), .A1(net_3167), .A2(net_3166) );
DFFS_X2 inst_6955 ( .QN(net_6410), .D(net_2689), .CK(net_14393), .SN(x1822) );
CLKBUF_X2 inst_13137 ( .A(net_13067), .Z(net_13099) );
CLKBUF_X2 inst_14328 ( .A(net_14289), .Z(net_14290) );
AOI22_X2 inst_7275 ( .B1(net_7089), .A1(net_7057), .A2(net_5280), .B2(net_5279), .ZN(net_5273) );
CLKBUF_X2 inst_10819 ( .A(net_9275), .Z(net_10781) );
CLKBUF_X2 inst_12332 ( .A(net_12293), .Z(net_12294) );
CLKBUF_X2 inst_9413 ( .A(net_8690), .Z(net_9375) );
NOR2_X2 inst_2455 ( .ZN(net_2815), .A2(net_2693), .A1(net_1180) );
CLKBUF_X2 inst_8000 ( .A(net_7961), .Z(net_7962) );
CLKBUF_X2 inst_12923 ( .A(net_12884), .Z(net_12885) );
CLKBUF_X2 inst_11535 ( .A(net_11496), .Z(net_11497) );
CLKBUF_X2 inst_10575 ( .A(net_9733), .Z(net_10537) );
DFF_X1 inst_6724 ( .QN(net_7357), .D(net_5332), .CK(net_10133) );
CLKBUF_X2 inst_11581 ( .A(net_11542), .Z(net_11543) );
INV_X4 inst_4828 ( .ZN(net_1083), .A(net_1082) );
INV_X4 inst_5218 ( .ZN(net_475), .A(net_474) );
INV_X4 inst_5389 ( .A(net_6021), .ZN(net_514) );
CLKBUF_X2 inst_12516 ( .A(net_12477), .Z(net_12478) );
INV_X4 inst_4860 ( .A(net_7807), .ZN(net_3299) );
CLKBUF_X2 inst_12226 ( .A(net_12187), .Z(net_12188) );
DFF_X1 inst_6770 ( .QN(net_6066), .D(net_4647), .CK(net_8737) );
SDFFR_X2 inst_1344 ( .Q(net_7712), .D(net_7712), .SI(net_3900), .SE(net_3405), .CK(net_13186), .RN(x1822) );
OAI22_X2 inst_1460 ( .B2(net_5902), .B1(net_4637), .ZN(net_4607), .A2(net_4605), .A1(net_4018) );
NOR2_X4 inst_2287 ( .ZN(net_5890), .A2(net_5872), .A1(net_3022) );
SDFF_X2 inst_885 ( .Q(net_7115), .D(net_7115), .SE(net_3888), .SI(net_3786), .CK(net_7918) );
CLKBUF_X2 inst_8968 ( .A(net_8929), .Z(net_8930) );
NAND3_X2 inst_2630 ( .ZN(net_5699), .A1(net_5676), .A2(net_5310), .A3(net_4250) );
INV_X2 inst_5803 ( .ZN(net_1725), .A(net_1100) );
CLKBUF_X2 inst_10748 ( .A(net_10709), .Z(net_10710) );
OAI22_X2 inst_1443 ( .B2(net_5905), .B1(net_4666), .A2(net_4634), .ZN(net_4632), .A1(net_4114) );
SDFF_X2 inst_1028 ( .D(net_7802), .SI(net_6497), .Q(net_6497), .SE(net_3889), .CK(net_11228) );
INV_X2 inst_5891 ( .A(net_7450), .ZN(net_1365) );
CLKBUF_X2 inst_10107 ( .A(net_8107), .Z(net_10069) );
NAND2_X2 inst_3935 ( .A2(net_1696), .ZN(net_1359), .A1(net_1358) );
NAND2_X2 inst_3610 ( .ZN(net_2386), .A2(net_1839), .A1(net_1378) );
CLKBUF_X2 inst_13097 ( .A(net_12156), .Z(net_13059) );
NAND2_X2 inst_2999 ( .A1(net_6747), .A2(net_5033), .ZN(net_5012) );
CLKBUF_X2 inst_9645 ( .A(net_9606), .Z(net_9607) );
SDFF_X2 inst_1271 ( .Q(net_5861), .SE(net_3040), .SI(net_3039), .D(net_550), .CK(net_12741) );
CLKBUF_X2 inst_12822 ( .A(net_12783), .Z(net_12784) );
CLKBUF_X2 inst_8351 ( .A(net_7863), .Z(net_8313) );
CLKBUF_X2 inst_12110 ( .A(net_12071), .Z(net_12072) );
NOR2_X2 inst_2321 ( .A2(net_6297), .A1(net_5840), .ZN(net_5820) );
CLKBUF_X2 inst_8188 ( .A(net_8149), .Z(net_8150) );
INV_X2 inst_5956 ( .A(net_7325), .ZN(net_1754) );
CLKBUF_X2 inst_13927 ( .A(net_13888), .Z(net_13889) );
NAND2_X2 inst_4156 ( .ZN(net_921), .A2(net_560), .A1(net_523) );
INV_X4 inst_5305 ( .A(net_6128), .ZN(net_3637) );
CLKBUF_X2 inst_9875 ( .A(net_9836), .Z(net_9837) );
CLKBUF_X2 inst_9928 ( .A(net_9393), .Z(net_9890) );
SDFF_X2 inst_200 ( .Q(net_6314), .SI(net_6313), .D(net_3473), .SE(net_392), .CK(net_13581) );
NAND2_X1 inst_4425 ( .A2(net_2131), .ZN(net_1456), .A1(net_1455) );
CLKBUF_X2 inst_11986 ( .A(net_11947), .Z(net_11948) );
CLKBUF_X2 inst_9727 ( .A(net_8342), .Z(net_9689) );
MUX2_X1 inst_4461 ( .S(net_7781), .Z(net_5862), .A(net_4162), .B(net_4161) );
DFF_X1 inst_6626 ( .QN(net_7596), .D(net_5261), .CK(net_13082) );
CLKBUF_X2 inst_14332 ( .A(net_13120), .Z(net_14294) );
NAND2_X1 inst_4373 ( .ZN(net_4354), .A2(net_3853), .A1(net_1992) );
CLKBUF_X2 inst_9939 ( .A(net_9900), .Z(net_9901) );
CLKBUF_X2 inst_9198 ( .A(net_7836), .Z(net_9160) );
AOI22_X2 inst_7407 ( .B1(net_5939), .A2(net_2838), .ZN(net_2829), .A1(net_2828), .B2(net_199) );
CLKBUF_X2 inst_12343 ( .A(net_12304), .Z(net_12305) );
OAI21_X2 inst_1750 ( .ZN(net_5515), .A(net_4817), .B2(net_4153), .B1(net_1070) );
CLKBUF_X2 inst_10807 ( .A(net_9643), .Z(net_10769) );
INV_X4 inst_5242 ( .ZN(net_3150), .A(net_525) );
NOR2_X4 inst_2236 ( .ZN(net_5662), .A1(net_5518), .A2(net_4490) );
NAND2_X2 inst_3368 ( .ZN(net_3510), .A1(net_3509), .A2(net_3223) );
AOI22_X2 inst_7307 ( .B1(net_6680), .A1(net_6648), .A2(net_5139), .B2(net_5138), .ZN(net_5136) );
OAI22_X2 inst_1553 ( .B2(net_3405), .A2(net_3360), .ZN(net_3352), .A1(net_3190), .B1(net_424) );
CLKBUF_X2 inst_13038 ( .A(net_12999), .Z(net_13000) );
CLKBUF_X2 inst_13937 ( .A(net_13898), .Z(net_13899) );
CLKBUF_X2 inst_10458 ( .A(net_10419), .Z(net_10420) );
CLKBUF_X2 inst_10155 ( .A(net_8954), .Z(net_10117) );
AOI21_X2 inst_7758 ( .B1(net_6475), .ZN(net_4039), .B2(net_2580), .A(net_2309) );
AOI222_X2 inst_7593 ( .A1(net_7392), .ZN(net_5542), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_355), .C2(net_353) );
OAI222_X2 inst_1635 ( .A1(net_5867), .C2(net_5052), .ZN(net_5051), .A2(net_5050), .B2(net_5049), .B1(net_2441), .C1(net_561) );
NAND2_X2 inst_4130 ( .ZN(net_939), .A2(net_938), .A1(net_679) );
CLKBUF_X2 inst_12121 ( .A(net_7930), .Z(net_12083) );
CLKBUF_X2 inst_9569 ( .A(net_9530), .Z(net_9531) );
CLKBUF_X2 inst_13102 ( .A(net_10664), .Z(net_13064) );
OAI22_X2 inst_1500 ( .B1(net_4660), .A1(net_4105), .B2(net_4101), .ZN(net_4098), .A2(net_4097) );
CLKBUF_X2 inst_11731 ( .A(net_9114), .Z(net_11693) );
CLKBUF_X2 inst_12294 ( .A(net_12255), .Z(net_12256) );
NAND3_X2 inst_2805 ( .ZN(net_2293), .A3(net_1541), .A1(net_1326), .A2(net_956) );
DFF_X1 inst_6438 ( .QN(net_6081), .D(net_5732), .CK(net_11280) );
NAND2_X2 inst_3499 ( .A2(net_2714), .ZN(net_2619), .A1(net_2421) );
NAND2_X2 inst_2932 ( .ZN(net_5518), .A1(net_4991), .A2(net_4990) );
SDFF_X2 inst_893 ( .Q(net_7125), .D(net_7125), .SE(net_3888), .SI(net_3795), .CK(net_8718) );
DFF_X1 inst_6917 ( .D(net_2395), .Q(net_251), .CK(net_8023) );
CLKBUF_X2 inst_9483 ( .A(net_9444), .Z(net_9445) );
NAND2_X2 inst_3048 ( .A1(net_6984), .A2(net_4977), .ZN(net_4959) );
CLKBUF_X2 inst_10911 ( .A(net_10872), .Z(net_10873) );
INV_X4 inst_4854 ( .ZN(net_1050), .A(net_689) );
CLKBUF_X2 inst_8128 ( .A(net_8089), .Z(net_8090) );
CLKBUF_X2 inst_13862 ( .A(net_13823), .Z(net_13824) );
SDFF_X2 inst_569 ( .Q(net_6733), .D(net_6733), .SI(net_3890), .SE(net_3815), .CK(net_11357) );
NAND2_X2 inst_3346 ( .ZN(net_3555), .A1(net_3554), .A2(net_3225) );
NAND2_X2 inst_2992 ( .A1(net_6723), .A2(net_5031), .ZN(net_5019) );
CLKBUF_X2 inst_9209 ( .A(net_8035), .Z(net_9171) );
CLKBUF_X2 inst_12763 ( .A(net_12724), .Z(net_12725) );
SDFF_X2 inst_1080 ( .Q(net_6362), .SI(net_6361), .D(net_3530), .SE(net_392), .CK(net_13600) );
DFF_X1 inst_6405 ( .QN(net_6132), .D(net_5765), .CK(net_10969) );
NOR2_X2 inst_2374 ( .ZN(net_5161), .A2(net_4611), .A1(net_4427) );
CLKBUF_X2 inst_14451 ( .A(net_11479), .Z(net_14413) );
AOI222_X2 inst_7473 ( .B1(net_7369), .C1(net_7305), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2159), .A1(net_2158) );
CLKBUF_X2 inst_12554 ( .A(net_12515), .Z(net_12516) );
SDFF_X2 inst_1103 ( .SI(net_6802), .Q(net_6802), .D(net_3812), .SE(net_3729), .CK(net_8266) );
DFF_X1 inst_6535 ( .QN(net_7482), .D(net_5416), .CK(net_9672) );
CLKBUF_X2 inst_8620 ( .A(net_8581), .Z(net_8582) );
CLKBUF_X2 inst_10678 ( .A(net_10639), .Z(net_10640) );
CLKBUF_X2 inst_9256 ( .A(net_9217), .Z(net_9218) );
AOI222_X2 inst_7494 ( .A2(net_2135), .B2(net_2133), .C2(net_2131), .ZN(net_2092), .A1(net_2091), .B1(net_2090), .C1(net_2089) );
SDFF_X2 inst_549 ( .Q(net_6466), .D(net_6466), .SE(net_3904), .SI(net_3894), .CK(net_11267) );
NAND2_X1 inst_4329 ( .ZN(net_4535), .A2(net_3870), .A1(net_1977) );
CLKBUF_X2 inst_12566 ( .A(net_12527), .Z(net_12528) );
NAND2_X1 inst_4220 ( .ZN(net_4740), .A2(net_3988), .A1(net_2113) );
INV_X4 inst_4708 ( .ZN(net_2989), .A(net_2988) );
SDFF_X2 inst_522 ( .SI(net_6630), .Q(net_6630), .D(net_3890), .SE(net_3851), .CK(net_7894) );
INV_X4 inst_5202 ( .A(net_541), .ZN(net_498) );
CLKBUF_X2 inst_13617 ( .A(net_13578), .Z(net_13579) );
INV_X4 inst_5040 ( .ZN(net_1218), .A(net_1040) );
CLKBUF_X2 inst_12408 ( .A(net_12369), .Z(net_12370) );
CLKBUF_X2 inst_9037 ( .A(net_8112), .Z(net_8999) );
CLKBUF_X2 inst_9842 ( .A(net_9803), .Z(net_9804) );
DFF_X2 inst_6231 ( .QN(net_6558), .D(net_3716), .CK(net_10733) );
NAND3_X2 inst_2809 ( .ZN(net_2289), .A3(net_1533), .A1(net_1512), .A2(net_1033) );
CLKBUF_X2 inst_14011 ( .A(net_10468), .Z(net_13973) );
CLKBUF_X2 inst_9654 ( .A(net_9615), .Z(net_9616) );
CLKBUF_X2 inst_13776 ( .A(net_13737), .Z(net_13738) );
CLKBUF_X2 inst_12478 ( .A(net_12439), .Z(net_12440) );
CLKBUF_X2 inst_13141 ( .A(net_13102), .Z(net_13103) );
DFF_X2 inst_6331 ( .QN(net_7796), .CK(net_11820), .D(x1572) );
CLKBUF_X2 inst_12797 ( .A(net_12758), .Z(net_12759) );
CLKBUF_X2 inst_9737 ( .A(net_9698), .Z(net_9699) );
NAND3_X2 inst_2673 ( .ZN(net_3752), .A3(net_3303), .A1(net_2963), .A2(net_2943) );
CLKBUF_X2 inst_13592 ( .A(net_13553), .Z(net_13554) );
OAI22_X2 inst_1618 ( .B1(net_5942), .ZN(net_2788), .A1(net_2786), .B2(net_209), .A2(net_172) );
INV_X4 inst_5062 ( .A(net_3159), .ZN(net_880) );
DFF_X1 inst_6936 ( .D(net_2403), .Q(net_261), .CK(net_8019) );
CLKBUF_X2 inst_14166 ( .A(net_14127), .Z(net_14128) );
OAI21_X2 inst_2126 ( .B2(net_3087), .B1(net_3071), .ZN(net_3061), .A(net_2908) );
CLKBUF_X2 inst_10484 ( .A(net_10445), .Z(net_10446) );
DFF_X1 inst_6911 ( .Q(net_6054), .D(net_2383), .CK(net_14380) );
CLKBUF_X2 inst_9144 ( .A(net_9105), .Z(net_9106) );
AOI21_X2 inst_7776 ( .B1(net_6603), .ZN(net_4026), .B2(net_2583), .A(net_2339) );
CLKBUF_X2 inst_11131 ( .A(net_11092), .Z(net_11093) );
CLKBUF_X2 inst_8997 ( .A(net_8958), .Z(net_8959) );
NAND3_X2 inst_2765 ( .ZN(net_2335), .A3(net_1550), .A1(net_1440), .A2(net_991) );
NAND2_X2 inst_3600 ( .ZN(net_2400), .A2(net_1857), .A1(net_1353) );
DFF_X1 inst_6493 ( .QN(net_7405), .D(net_5552), .CK(net_9306) );
SDFF_X2 inst_219 ( .Q(net_6335), .SI(net_6334), .D(net_3655), .SE(net_392), .CK(net_14054) );
SDFF_X2 inst_719 ( .SI(net_6763), .Q(net_6763), .SE(net_3872), .D(net_3798), .CK(net_11091) );
CLKBUF_X2 inst_10195 ( .A(net_10156), .Z(net_10157) );
NAND2_X2 inst_4166 ( .ZN(net_1682), .A2(net_825), .A1(net_485) );
INV_X4 inst_4881 ( .ZN(net_2704), .A(net_902) );
CLKBUF_X2 inst_8980 ( .A(net_8941), .Z(net_8942) );
CLKBUF_X2 inst_8695 ( .A(net_8656), .Z(net_8657) );
NAND2_X2 inst_3868 ( .A1(net_6704), .A2(net_1497), .ZN(net_1461) );
SDFF_X2 inst_1134 ( .SI(net_6686), .Q(net_6686), .D(net_3800), .SE(net_3465), .CK(net_11993) );
INV_X4 inst_5501 ( .A(net_6161), .ZN(net_3599) );
NOR3_X2 inst_2204 ( .A3(net_5920), .ZN(net_3183), .A2(net_2899), .A1(net_2898) );
OAI22_X2 inst_1609 ( .A1(net_3270), .ZN(net_3088), .A2(net_3087), .B2(net_3084), .B1(net_497) );
NAND2_X2 inst_4105 ( .A1(net_6668), .A2(net_1655), .ZN(net_947) );
NAND2_X2 inst_3546 ( .ZN(net_2521), .A2(net_2088), .A1(net_1787) );
SDFF_X2 inst_408 ( .SI(net_7372), .Q(net_7372), .D(net_4779), .SE(net_3853), .CK(net_9895) );
INV_X2 inst_5748 ( .ZN(net_3716), .A(net_3413) );
SDFF_X2 inst_1144 ( .D(net_7807), .SI(net_6804), .Q(net_6804), .SE(net_3729), .CK(net_10773) );
INV_X4 inst_4701 ( .ZN(net_3441), .A(net_3339) );
INV_X4 inst_5165 ( .A(net_645), .ZN(net_545) );
INV_X4 inst_5644 ( .A(net_6033), .ZN(net_467) );
CLKBUF_X2 inst_12419 ( .A(net_12380), .Z(net_12381) );
CLKBUF_X2 inst_11212 ( .A(net_7987), .Z(net_11174) );
INV_X4 inst_5366 ( .A(net_5998), .ZN(net_3106) );
DFF_X1 inst_6426 ( .QN(net_6181), .D(net_5744), .CK(net_10677) );
INV_X4 inst_5551 ( .A(net_6168), .ZN(net_3560) );
NAND3_X4 inst_2568 ( .A1(net_5943), .ZN(net_2488), .A2(net_1864), .A3(net_1819) );
INV_X4 inst_5596 ( .A(net_6008), .ZN(net_465) );
NOR2_X4 inst_2295 ( .ZN(net_2709), .A2(net_284), .A1(net_278) );
CLKBUF_X2 inst_13021 ( .A(net_8449), .Z(net_12983) );
CLKBUF_X2 inst_11591 ( .A(net_11552), .Z(net_11553) );
CLKBUF_X2 inst_10719 ( .A(net_10680), .Z(net_10681) );
NAND2_X2 inst_3814 ( .A1(net_6494), .A2(net_1642), .ZN(net_1531) );
CLKBUF_X2 inst_12968 ( .A(net_12929), .Z(net_12930) );
CLKBUF_X2 inst_8498 ( .A(net_8459), .Z(net_8460) );
NAND2_X2 inst_3028 ( .A1(net_6986), .ZN(net_4981), .A2(net_4977) );
NAND2_X2 inst_3532 ( .ZN(net_2535), .A2(net_2143), .A1(net_1377) );
CLKBUF_X2 inst_9190 ( .A(net_9151), .Z(net_9152) );
CLKBUF_X2 inst_9432 ( .A(net_8084), .Z(net_9394) );
NAND2_X2 inst_3854 ( .A1(net_6968), .A2(net_1833), .ZN(net_1481) );
CLKBUF_X2 inst_7871 ( .A(net_7832), .Z(net_7833) );
CLKBUF_X2 inst_10881 ( .A(net_10842), .Z(net_10843) );
NAND2_X2 inst_3514 ( .ZN(net_2553), .A2(net_2151), .A1(net_1385) );
CLKBUF_X2 inst_10826 ( .A(net_10787), .Z(net_10788) );
OAI22_X2 inst_1530 ( .B1(net_4644), .B2(net_4437), .A1(net_4057), .A2(net_4055), .ZN(net_4037) );
DFFR_X2 inst_7089 ( .QN(net_7729), .D(net_2792), .CK(net_13216), .RN(x1822) );
OAI22_X2 inst_1510 ( .B1(net_4650), .B2(net_4083), .A1(net_4080), .ZN(net_4077), .A2(net_4076) );
XNOR2_X2 inst_121 ( .ZN(net_5867), .B(net_1648), .A(net_833) );
INV_X4 inst_5421 ( .A(net_6084), .ZN(net_3517) );
CLKBUF_X2 inst_12449 ( .A(net_12410), .Z(net_12411) );
SDFF_X2 inst_1065 ( .SI(net_7038), .Q(net_7038), .D(net_3894), .SE(net_3777), .CK(net_8198) );
AOI21_X2 inst_7635 ( .ZN(net_3955), .B2(net_3769), .B1(net_2892), .A(net_923) );
CLKBUF_X2 inst_12002 ( .A(net_11963), .Z(net_11964) );
DFF_X2 inst_6308 ( .QN(net_7808), .CK(net_11279), .D(x1479) );
CLKBUF_X2 inst_11599 ( .A(net_11450), .Z(net_11561) );
NAND2_X2 inst_4119 ( .A2(net_1228), .ZN(net_1081), .A1(net_374) );
INV_X2 inst_5948 ( .ZN(net_1129), .A(net_126) );
NAND2_X1 inst_4332 ( .ZN(net_4532), .A2(net_3870), .A1(net_1320) );
CLKBUF_X2 inst_13766 ( .A(net_13727), .Z(net_13728) );
CLKBUF_X2 inst_9340 ( .A(net_9301), .Z(net_9302) );
CLKBUF_X2 inst_13318 ( .A(net_13279), .Z(net_13280) );
CLKBUF_X2 inst_10955 ( .A(net_10916), .Z(net_10917) );
CLKBUF_X2 inst_10076 ( .A(net_8323), .Z(net_10038) );
DFF_X2 inst_6282 ( .Q(net_6385), .D(net_6384), .CK(net_14172) );
CLKBUF_X2 inst_12111 ( .A(net_9168), .Z(net_12073) );
CLKBUF_X2 inst_14348 ( .A(net_10955), .Z(net_14310) );
CLKBUF_X2 inst_9495 ( .A(net_9037), .Z(net_9457) );
INV_X4 inst_5353 ( .A(net_6154), .ZN(net_3613) );
CLKBUF_X2 inst_14189 ( .A(net_14150), .Z(net_14151) );
CLKBUF_X2 inst_13876 ( .A(net_13837), .Z(net_13838) );
CLKBUF_X2 inst_9981 ( .A(net_9942), .Z(net_9943) );
CLKBUF_X2 inst_12586 ( .A(net_12547), .Z(net_12548) );
INV_X4 inst_4671 ( .A(net_4155), .ZN(net_3472) );
DFF_X2 inst_6244 ( .QN(net_7681), .D(net_2972), .CK(net_8320) );
CLKBUF_X2 inst_8753 ( .A(net_8217), .Z(net_8715) );
NAND2_X2 inst_4174 ( .A1(net_6823), .ZN(net_786), .A2(net_630) );
SDFF_X2 inst_530 ( .Q(net_6594), .D(net_6594), .SI(net_3892), .SE(net_3830), .CK(net_12935) );
CLKBUF_X2 inst_9009 ( .A(net_8970), .Z(net_8971) );
CLKBUF_X2 inst_8004 ( .A(net_7965), .Z(net_7966) );
SDFFR_X2 inst_1353 ( .D(net_3883), .SE(net_3297), .SI(net_274), .Q(net_274), .CK(net_12819), .RN(x1822) );
DFF_X1 inst_6369 ( .QN(net_6293), .D(net_5815), .CK(net_13786) );
AOI22_X2 inst_7370 ( .ZN(net_5957), .A2(net_5916), .B2(net_2957), .B1(net_2952), .A1(net_851) );
NOR2_X2 inst_2502 ( .A1(net_3042), .ZN(net_1264), .A2(net_1263) );
SDFF_X2 inst_769 ( .Q(net_6892), .D(net_6892), .SE(net_3901), .SI(net_3800), .CK(net_11724) );
CLKBUF_X2 inst_13334 ( .A(net_9886), .Z(net_13296) );
CLKBUF_X2 inst_12429 ( .A(net_12390), .Z(net_12391) );
SDFF_X2 inst_1200 ( .SI(net_7083), .Q(net_7083), .D(net_3780), .SE(net_3742), .CK(net_11841) );
CLKBUF_X2 inst_10888 ( .A(net_10038), .Z(net_10850) );
CLKBUF_X2 inst_10120 ( .A(net_10081), .Z(net_10082) );
CLKBUF_X2 inst_9114 ( .A(net_8302), .Z(net_9076) );
CLKBUF_X2 inst_11233 ( .A(net_9192), .Z(net_11195) );
CLKBUF_X2 inst_10918 ( .A(net_10879), .Z(net_10880) );
CLKBUF_X2 inst_8523 ( .A(net_8484), .Z(net_8485) );
NAND2_X2 inst_3021 ( .A1(net_6860), .A2(net_5004), .ZN(net_4988) );
NAND2_X2 inst_3974 ( .ZN(net_1296), .A1(net_885), .A2(net_319) );
DFF_X1 inst_6349 ( .QN(net_6209), .D(net_5835), .CK(net_14287) );
CLKBUF_X2 inst_13290 ( .A(net_13251), .Z(net_13252) );
AOI22_X2 inst_7365 ( .A2(net_5916), .ZN(net_2958), .B2(net_2957), .B1(net_2655), .A1(net_844) );
DFF_X1 inst_6474 ( .QN(net_6071), .D(net_5585), .CK(net_11675) );
CLKBUF_X2 inst_12601 ( .A(net_12562), .Z(net_12563) );
CLKBUF_X2 inst_12232 ( .A(net_12193), .Z(net_12194) );
CLKBUF_X2 inst_11664 ( .A(net_10610), .Z(net_11626) );
CLKBUF_X2 inst_11501 ( .A(net_11462), .Z(net_11463) );
SDFF_X2 inst_213 ( .Q(net_6301), .SI(net_6300), .D(net_3685), .SE(net_392), .CK(net_13545) );
CLKBUF_X2 inst_12618 ( .A(net_12579), .Z(net_12580) );
SDFF_X2 inst_205 ( .Q(net_6309), .SI(net_6308), .D(net_3669), .SE(net_392), .CK(net_13567) );
OAI221_X2 inst_1645 ( .ZN(net_5450), .B2(net_5043), .C2(net_5041), .A(net_4903), .C1(net_1153), .B1(net_723) );
CLKBUF_X2 inst_13045 ( .A(net_13006), .Z(net_13007) );
CLKBUF_X2 inst_7904 ( .A(net_7828), .Z(net_7866) );
NAND2_X2 inst_3722 ( .A1(net_6759), .A2(net_1635), .ZN(net_1623) );
INV_X4 inst_5410 ( .A(net_6159), .ZN(net_3601) );
CLKBUF_X2 inst_8043 ( .A(net_8004), .Z(net_8005) );
NAND2_X1 inst_4311 ( .ZN(net_4555), .A2(net_3866), .A1(net_2090) );
CLKBUF_X2 inst_11922 ( .A(net_10298), .Z(net_11884) );
NAND2_X2 inst_3911 ( .A2(net_1696), .ZN(net_1396), .A1(net_1395) );
OAI22_X2 inst_1515 ( .B1(net_4650), .A1(net_4080), .B2(net_4070), .ZN(net_4067), .A2(net_4066) );
DFF_X1 inst_6777 ( .QN(net_6124), .D(net_4324), .CK(net_10950) );
CLKBUF_X2 inst_9743 ( .A(net_9704), .Z(net_9705) );
AOI222_X2 inst_7546 ( .C1(net_7669), .A1(net_7637), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1866), .B1(net_1865) );
CLKBUF_X2 inst_13088 ( .A(net_8279), .Z(net_13050) );
CLKBUF_X2 inst_14117 ( .A(net_11422), .Z(net_14079) );
OAI21_X2 inst_1782 ( .B1(net_5448), .ZN(net_5409), .A(net_4683), .B2(net_3988) );
INV_X4 inst_5173 ( .A(net_586), .ZN(net_534) );
NAND2_X2 inst_2951 ( .ZN(net_5489), .A1(net_4947), .A2(net_4946) );
DFF_X1 inst_6464 ( .QN(net_6149), .D(net_5595), .CK(net_11985) );
CLKBUF_X2 inst_9176 ( .A(net_9137), .Z(net_9138) );
NAND2_X2 inst_3890 ( .A1(net_6571), .A2(net_1705), .ZN(net_1426) );
INV_X8 inst_4472 ( .ZN(net_5184), .A(net_4275) );
AOI222_X2 inst_7513 ( .B1(net_7373), .C1(net_7309), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2028), .A1(net_2027) );
SDFF_X2 inst_1015 ( .SI(net_6508), .Q(net_6508), .SE(net_3889), .D(net_3783), .CK(net_8404) );
DFFR_X2 inst_7003 ( .QN(net_7693), .D(net_3349), .CK(net_12878), .RN(x1822) );
CLKBUF_X2 inst_14390 ( .A(net_14351), .Z(net_14352) );
NAND2_X2 inst_3899 ( .A1(net_6973), .A2(net_1833), .ZN(net_1415) );
CLKBUF_X2 inst_13526 ( .A(net_13487), .Z(net_13488) );
CLKBUF_X2 inst_14226 ( .A(net_14187), .Z(net_14188) );
NAND2_X2 inst_3213 ( .ZN(net_4713), .A2(net_3986), .A1(net_2148) );
CLKBUF_X2 inst_10209 ( .A(net_10170), .Z(net_10171) );
NOR2_X2 inst_2535 ( .A2(net_7097), .ZN(net_1245), .A1(net_532) );
INV_X8 inst_4569 ( .A(net_7791), .ZN(net_5925) );
OAI221_X2 inst_1661 ( .C2(net_5895), .ZN(net_4667), .B1(net_4666), .B2(net_4506), .C1(net_4132), .A(net_3684) );
CLKBUF_X2 inst_12393 ( .A(net_12354), .Z(net_12355) );
INV_X8 inst_4480 ( .ZN(net_4282), .A(net_3928) );
CLKBUF_X2 inst_13583 ( .A(net_13544), .Z(net_13545) );
SDFF_X2 inst_283 ( .D(net_6397), .SE(net_5799), .SI(net_382), .Q(net_382), .CK(net_13904) );
CLKBUF_X2 inst_10723 ( .A(net_10684), .Z(net_10685) );
DFF_X1 inst_6676 ( .QN(net_7254), .D(net_5148), .CK(net_10183) );
NOR2_X2 inst_2519 ( .ZN(net_917), .A1(net_916), .A2(net_885) );
NAND2_X2 inst_3406 ( .A2(net_5968), .ZN(net_3384), .A1(net_2877) );
CLKBUF_X2 inst_9378 ( .A(net_8659), .Z(net_9340) );
OAI22_X2 inst_1597 ( .B2(net_3200), .A2(net_3196), .ZN(net_3140), .A1(net_3139), .B1(net_864) );
INV_X4 inst_5639 ( .A(net_6089), .ZN(net_3483) );
NAND2_X2 inst_3502 ( .ZN(net_2599), .A2(net_2598), .A1(net_429) );
AOI222_X2 inst_7574 ( .A1(net_7537), .ZN(net_4849), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_369), .C2(net_367) );
NAND2_X2 inst_3473 ( .ZN(net_2710), .A2(net_2706), .A1(net_396) );
INV_X2 inst_6018 ( .ZN(net_1123), .A(net_117) );
CLKBUF_X2 inst_9942 ( .A(net_9903), .Z(net_9904) );
CLKBUF_X2 inst_8502 ( .A(net_8463), .Z(net_8464) );
AOI21_X2 inst_7705 ( .B1(net_6467), .ZN(net_4056), .B2(net_2580), .A(net_2324) );
INV_X2 inst_5822 ( .ZN(net_937), .A(net_936) );
SDFF_X2 inst_431 ( .Q(net_7385), .D(net_7385), .SE(net_3994), .SI(net_350), .CK(net_9754) );
INV_X2 inst_6063 ( .A(net_7753), .ZN(net_5870) );
DFF_X1 inst_6448 ( .QN(net_6099), .D(net_5722), .CK(net_12058) );
SDFF_X2 inst_348 ( .SI(net_7679), .Q(net_7679), .D(net_4793), .SE(net_3866), .CK(net_13399) );
CLKBUF_X2 inst_11331 ( .A(net_11292), .Z(net_11293) );
AOI21_X2 inst_7676 ( .B1(net_7012), .ZN(net_4220), .A(net_2473), .B2(net_1100) );
DFF_X1 inst_6906 ( .D(net_2503), .Q(net_186), .CK(net_12402) );
AOI22_X2 inst_7429 ( .A1(net_2970), .B1(net_2772), .ZN(net_2763), .A2(net_245), .B2(net_171) );
CLKBUF_X2 inst_8737 ( .A(net_8210), .Z(net_8699) );
NAND3_X2 inst_2686 ( .ZN(net_3177), .A3(net_2982), .A2(net_1964), .A1(net_1104) );
INV_X4 inst_5123 ( .A(net_629), .ZN(net_594) );
CLKBUF_X2 inst_10774 ( .A(net_10735), .Z(net_10736) );
NAND2_X2 inst_3740 ( .A1(net_6900), .A2(net_1639), .ZN(net_1605) );
CLKBUF_X2 inst_9600 ( .A(net_9561), .Z(net_9562) );
NOR2_X4 inst_2293 ( .A2(net_7791), .ZN(net_2863), .A1(net_802) );
SDFFR_X2 inst_1364 ( .SI(net_7739), .Q(net_7739), .D(net_4596), .SE(net_2606), .CK(net_10330), .RN(x1822) );
CLKBUF_X2 inst_11299 ( .A(net_11260), .Z(net_11261) );
CLKBUF_X2 inst_11514 ( .A(net_11475), .Z(net_11476) );
SDFF_X2 inst_645 ( .D(net_7799), .SI(net_6629), .Q(net_6629), .SE(net_3850), .CK(net_12899) );
CLKBUF_X2 inst_13299 ( .A(net_10001), .Z(net_13261) );
NAND2_X2 inst_3041 ( .A1(net_7025), .A2(net_4979), .ZN(net_4966) );
NOR2_X2 inst_2352 ( .ZN(net_5652), .A1(net_5504), .A2(net_4471) );
NAND3_X2 inst_2719 ( .ZN(net_2456), .A2(net_1804), .A3(net_1591), .A1(net_1360) );
SDFF_X2 inst_269 ( .D(net_6400), .SE(net_5799), .SI(net_385), .Q(net_385), .CK(net_13910) );
DFF_X1 inst_6847 ( .D(net_2538), .QN(net_210), .CK(net_12614) );
DFF_X1 inst_6864 ( .D(net_2543), .QN(net_201), .CK(net_12465) );
CLKBUF_X2 inst_12534 ( .A(net_12495), .Z(net_12496) );
CLKBUF_X2 inst_14278 ( .A(net_12002), .Z(net_14240) );
CLKBUF_X2 inst_11278 ( .A(net_8187), .Z(net_11240) );
CLKBUF_X2 inst_9560 ( .A(net_9521), .Z(net_9522) );
NOR2_X2 inst_2544 ( .A1(net_3374), .A2(net_3372), .ZN(net_647) );
CLKBUF_X2 inst_9796 ( .A(net_8683), .Z(net_9758) );
SDFF_X2 inst_514 ( .Q(net_6697), .D(net_6697), .SI(net_3892), .SE(net_3871), .CK(net_8304) );
CLKBUF_X2 inst_14364 ( .A(net_8752), .Z(net_14326) );
CLKBUF_X2 inst_12707 ( .A(net_12668), .Z(net_12669) );
OAI22_X2 inst_1541 ( .B1(net_4637), .A1(net_4030), .B2(net_4016), .ZN(net_4013), .A2(net_4012) );
NAND2_X1 inst_4236 ( .ZN(net_4691), .A2(net_3989), .A1(net_2070) );
SDFF_X2 inst_685 ( .Q(net_6750), .D(net_6750), .SE(net_3815), .SI(net_3791), .CK(net_8371) );
CLKBUF_X2 inst_13281 ( .A(net_13242), .Z(net_13243) );
CLKBUF_X2 inst_9586 ( .A(net_9547), .Z(net_9548) );
CLKBUF_X2 inst_12952 ( .A(net_12913), .Z(net_12914) );
CLKBUF_X2 inst_13829 ( .A(net_13790), .Z(net_13791) );
CLKBUF_X2 inst_14061 ( .A(net_14022), .Z(net_14023) );
INV_X4 inst_4656 ( .ZN(net_5878), .A(net_4143) );
CLKBUF_X2 inst_10658 ( .A(net_10619), .Z(net_10620) );
CLKBUF_X2 inst_9150 ( .A(net_9111), .Z(net_9112) );
DFF_X2 inst_6338 ( .QN(net_7801), .CK(net_8159), .D(x1534) );
CLKBUF_X2 inst_14358 ( .A(net_14319), .Z(net_14320) );
INV_X4 inst_5621 ( .A(net_6098), .ZN(net_3507) );
CLKBUF_X2 inst_11585 ( .A(net_11546), .Z(net_11547) );
CLKBUF_X2 inst_10636 ( .A(net_10597), .Z(net_10598) );
NAND2_X2 inst_3432 ( .ZN(net_3216), .A2(net_3100), .A1(net_2765) );
CLKBUF_X2 inst_14047 ( .A(net_12339), .Z(net_14009) );
AOI21_X2 inst_7693 ( .B1(net_6735), .ZN(net_4130), .B2(net_2581), .A(net_2371) );
DFF_X1 inst_6561 ( .QN(net_7434), .D(net_5046), .CK(net_12552) );
CLKBUF_X2 inst_12700 ( .A(net_11125), .Z(net_12662) );
CLKBUF_X2 inst_12678 ( .A(net_8659), .Z(net_12640) );
CLKBUF_X2 inst_13984 ( .A(net_13945), .Z(net_13946) );
DFF_X1 inst_6886 ( .D(net_2519), .Q(net_167), .CK(net_12230) );
CLKBUF_X2 inst_8959 ( .A(net_8920), .Z(net_8921) );
SDFF_X2 inst_427 ( .SI(net_7752), .Q(net_7752), .SE(net_5925), .D(net_3913), .CK(net_12517) );
NAND2_X2 inst_3840 ( .A1(net_6442), .A2(net_1677), .ZN(net_1499) );
DFF_X1 inst_6881 ( .D(net_2515), .QN(net_174), .CK(net_9858) );
CLKBUF_X2 inst_13113 ( .A(net_13074), .Z(net_13075) );
CLKBUF_X2 inst_8905 ( .A(net_8866), .Z(net_8867) );
CLKBUF_X2 inst_13852 ( .A(net_13813), .Z(net_13814) );
CLKBUF_X2 inst_9477 ( .A(net_8629), .Z(net_9439) );
CLKBUF_X2 inst_11952 ( .A(net_11913), .Z(net_11914) );
OAI21_X2 inst_2144 ( .B1(net_5778), .ZN(net_2800), .A(net_2677), .B2(net_2675) );
INV_X2 inst_5721 ( .ZN(net_4245), .A(net_4112) );
INV_X16 inst_6121 ( .ZN(net_5004), .A(net_4267) );
SDFF_X2 inst_138 ( .Q(net_6212), .SI(net_6211), .SE(net_392), .D(net_146), .CK(net_14224) );
DFF_X1 inst_6793 ( .D(net_3948), .CK(net_12839), .Q(x718) );
DFFR_X2 inst_6973 ( .QN(net_7789), .D(net_3987), .CK(net_10247), .RN(x1822) );
NAND3_X2 inst_2810 ( .ZN(net_2288), .A3(net_1625), .A1(net_1348), .A2(net_953) );
INV_X4 inst_5333 ( .A(net_6122), .ZN(net_3689) );
CLKBUF_X2 inst_13971 ( .A(net_13932), .Z(net_13933) );
SDFF_X2 inst_899 ( .Q(net_7130), .D(net_7130), .SE(net_3888), .SI(net_3800), .CK(net_10642) );
INV_X4 inst_4944 ( .ZN(net_1306), .A(net_744) );
CLKBUF_X2 inst_10975 ( .A(net_10936), .Z(net_10937) );
CLKBUF_X2 inst_10259 ( .A(net_10220), .Z(net_10221) );
CLKBUF_X2 inst_12304 ( .A(net_12265), .Z(net_12266) );
SDFF_X2 inst_312 ( .SI(net_7454), .Q(net_7454), .D(net_5107), .SE(net_3993), .CK(net_12589) );
CLKBUF_X2 inst_13346 ( .A(net_13307), .Z(net_13308) );
CLKBUF_X2 inst_13256 ( .A(net_13217), .Z(net_13218) );
CLKBUF_X2 inst_13429 ( .A(net_13390), .Z(net_13391) );
CLKBUF_X2 inst_9554 ( .A(net_9515), .Z(net_9516) );
SDFF_X2 inst_309 ( .D(net_6393), .SE(net_6050), .SI(net_302), .Q(net_302), .CK(net_14216) );
CLKBUF_X2 inst_9889 ( .A(net_9850), .Z(net_9851) );
NAND2_X2 inst_3416 ( .ZN(net_3245), .A1(net_3240), .A2(net_602) );
OAI21_X2 inst_2149 ( .B1(net_5778), .ZN(net_2795), .A(net_2662), .B2(net_2660) );
CLKBUF_X2 inst_13765 ( .A(net_9964), .Z(net_13727) );
CLKBUF_X2 inst_8356 ( .A(net_8317), .Z(net_8318) );
DFFR_X2 inst_6980 ( .QN(net_5994), .D(net_3448), .CK(net_10760), .RN(x1822) );
INV_X4 inst_5001 ( .ZN(net_755), .A(net_707) );
CLKBUF_X2 inst_9365 ( .A(net_8146), .Z(net_9327) );
CLKBUF_X2 inst_11875 ( .A(net_11836), .Z(net_11837) );
AOI22_X2 inst_7265 ( .B1(net_6956), .A1(net_6924), .A2(net_5298), .B2(net_5297), .ZN(net_5289) );
CLKBUF_X2 inst_9833 ( .A(net_9794), .Z(net_9795) );
NAND3_X2 inst_2694 ( .ZN(net_2982), .A3(net_2896), .A2(net_2752), .A1(net_1923) );
AOI22_X2 inst_7386 ( .ZN(net_5959), .A2(net_5916), .B2(net_2957), .B1(net_2661), .A1(net_839) );
CLKBUF_X2 inst_8038 ( .A(net_7999), .Z(net_8000) );
CLKBUF_X2 inst_9950 ( .A(net_9911), .Z(net_9912) );
CLKBUF_X2 inst_9319 ( .A(net_9280), .Z(net_9281) );
CLKBUF_X2 inst_8172 ( .A(net_8133), .Z(net_8134) );
CLKBUF_X2 inst_13899 ( .A(net_8494), .Z(net_13861) );
CLKBUF_X2 inst_8876 ( .A(net_8032), .Z(net_8838) );
OAI21_X2 inst_1968 ( .ZN(net_4871), .B1(net_4870), .A(net_4342), .B2(net_3859) );
CLKBUF_X2 inst_12983 ( .A(net_12944), .Z(net_12945) );
NAND2_X2 inst_4078 ( .A1(net_6536), .A2(net_1645), .ZN(net_974) );
CLKBUF_X2 inst_12168 ( .A(net_12129), .Z(net_12130) );
NAND2_X2 inst_4067 ( .A1(net_7204), .A2(net_1648), .ZN(net_985) );
CLKBUF_X2 inst_12038 ( .A(net_11999), .Z(net_12000) );
SDFFR_X2 inst_1330 ( .Q(net_7770), .D(net_7770), .SE(net_4303), .SI(net_4165), .CK(net_12372), .RN(x1822) );
CLKBUF_X2 inst_13963 ( .A(net_13924), .Z(net_13925) );
CLKBUF_X2 inst_13728 ( .A(net_13689), .Z(net_13690) );
CLKBUF_X2 inst_12410 ( .A(net_12371), .Z(net_12372) );
CLKBUF_X2 inst_9109 ( .A(net_9070), .Z(net_9071) );
CLKBUF_X2 inst_8894 ( .A(net_8488), .Z(net_8856) );
OAI21_X2 inst_1898 ( .B1(net_5202), .ZN(net_5178), .A(net_4555), .B2(net_3866) );
CLKBUF_X2 inst_10175 ( .A(net_10136), .Z(net_10137) );
CLKBUF_X2 inst_14180 ( .A(net_14141), .Z(net_14142) );
CLKBUF_X2 inst_8885 ( .A(net_8846), .Z(net_8847) );
NAND2_X2 inst_3883 ( .A1(net_6424), .A2(net_1677), .ZN(net_1436) );
CLKBUF_X2 inst_10020 ( .A(net_9981), .Z(net_9982) );
CLKBUF_X2 inst_8551 ( .A(net_8459), .Z(net_8513) );
OAI21_X2 inst_1714 ( .ZN(net_5580), .B1(net_5554), .A(net_4690), .B2(net_3989) );
DFF_X2 inst_6275 ( .QN(net_5922), .D(net_389), .CK(net_12214) );
CLKBUF_X2 inst_11811 ( .A(net_8125), .Z(net_11773) );
CLKBUF_X2 inst_13451 ( .A(net_13412), .Z(net_13413) );
CLKBUF_X2 inst_9164 ( .A(net_8778), .Z(net_9126) );
CLKBUF_X2 inst_9096 ( .A(net_9057), .Z(net_9058) );
CLKBUF_X2 inst_9428 ( .A(net_9389), .Z(net_9390) );
INV_X4 inst_4777 ( .A(net_1965), .ZN(net_1714) );
CLKBUF_X2 inst_10851 ( .A(net_10812), .Z(net_10813) );
CLKBUF_X2 inst_10762 ( .A(net_10723), .Z(net_10724) );
INV_X2 inst_5818 ( .A(net_1637), .ZN(net_1095) );
CLKBUF_X2 inst_11292 ( .A(net_11253), .Z(net_11254) );
OAI22_X2 inst_1496 ( .B1(net_4660), .ZN(net_4111), .A2(net_4110), .B2(net_4109), .A1(net_4105) );
INV_X4 inst_5510 ( .A(net_7566), .ZN(net_1851) );
CLKBUF_X2 inst_9091 ( .A(net_9052), .Z(net_9053) );
DFFR_X2 inst_7041 ( .QN(net_6001), .D(net_3172), .CK(net_12861), .RN(x1822) );
CLKBUF_X2 inst_13005 ( .A(net_12966), .Z(net_12967) );
CLKBUF_X2 inst_9381 ( .A(net_9342), .Z(net_9343) );
NAND2_X1 inst_4297 ( .ZN(net_4569), .A2(net_3866), .A1(net_1912) );
SDFF_X2 inst_924 ( .Q(net_7161), .D(net_7161), .SE(net_3903), .SI(net_3801), .CK(net_8076) );
OAI22_X2 inst_1565 ( .A2(net_3297), .ZN(net_3288), .A1(net_3287), .B2(net_3286), .B1(net_756) );
CLKBUF_X2 inst_8415 ( .A(net_7856), .Z(net_8377) );
CLKBUF_X2 inst_12632 ( .A(net_12593), .Z(net_12594) );
CLKBUF_X2 inst_10308 ( .A(net_9624), .Z(net_10270) );
SDFF_X2 inst_287 ( .D(net_6396), .SE(net_5799), .SI(net_381), .Q(net_381), .CK(net_14329) );
CLKBUF_X2 inst_10614 ( .A(net_10237), .Z(net_10576) );
NAND3_X2 inst_2577 ( .ZN(net_5762), .A1(net_5657), .A2(net_5281), .A3(net_4306) );
CLKBUF_X2 inst_7929 ( .A(net_7890), .Z(net_7891) );
CLKBUF_X2 inst_12030 ( .A(net_11991), .Z(net_11992) );
AOI222_X2 inst_7565 ( .A1(net_7388), .ZN(net_5554), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_351), .C2(net_349) );
NAND2_X2 inst_3094 ( .A1(net_6487), .A2(net_4927), .ZN(net_4909) );
CLKBUF_X2 inst_13267 ( .A(net_13228), .Z(net_13229) );
CLKBUF_X2 inst_13830 ( .A(net_10840), .Z(net_13792) );
NAND2_X4 inst_2903 ( .ZN(net_3256), .A1(net_2916), .A2(net_2915) );
NAND2_X2 inst_4045 ( .A1(net_6935), .A2(net_1654), .ZN(net_1007) );
DFF_X1 inst_6431 ( .QN(net_6074), .D(net_5739), .CK(net_8450) );
CLKBUF_X2 inst_12623 ( .A(net_12584), .Z(net_12585) );
INV_X4 inst_4890 ( .ZN(net_877), .A(net_876) );
SDFF_X2 inst_984 ( .Q(net_6469), .D(net_6469), .SE(net_3904), .SI(net_3811), .CK(net_11667) );
NAND2_X2 inst_3804 ( .A1(net_6631), .A2(net_1624), .ZN(net_1541) );
DFF_X1 inst_6734 ( .QN(net_7353), .D(net_5321), .CK(net_10116) );
OAI21_X2 inst_2064 ( .B2(net_4436), .ZN(net_4431), .B1(net_4053), .A(net_3547) );
NOR2_X4 inst_2266 ( .ZN(net_5620), .A1(net_5465), .A2(net_4414) );
CLKBUF_X2 inst_14331 ( .A(net_14292), .Z(net_14293) );
SDFF_X2 inst_1292 ( .D(net_3806), .SE(net_3256), .SI(net_131), .Q(net_131), .CK(net_8455) );
CLKBUF_X2 inst_13206 ( .A(net_13167), .Z(net_13168) );
INV_X4 inst_5014 ( .A(net_1146), .ZN(net_722) );
OAI21_X2 inst_1963 ( .B1(net_5414), .ZN(net_5047), .A(net_4655), .B2(net_3993) );
SDFF_X2 inst_1056 ( .Q(net_6747), .D(net_6747), .SI(net_3900), .SE(net_3815), .CK(net_8353) );
CLKBUF_X2 inst_11818 ( .A(net_11779), .Z(net_11780) );
CLKBUF_X2 inst_13440 ( .A(net_13401), .Z(net_13402) );
NAND2_X2 inst_3648 ( .A1(net_7066), .ZN(net_1815), .A2(net_791) );
NAND2_X1 inst_4247 ( .ZN(net_4680), .A2(net_3988), .A1(net_2192) );
CLKBUF_X2 inst_14434 ( .A(net_14395), .Z(net_14396) );
CLKBUF_X2 inst_8744 ( .A(net_8705), .Z(net_8706) );
CLKBUF_X2 inst_12023 ( .A(net_11984), .Z(net_11985) );
CLKBUF_X2 inst_13437 ( .A(net_13398), .Z(net_13399) );
NOR2_X2 inst_2514 ( .A1(net_3048), .ZN(net_1158), .A2(net_1157) );
CLKBUF_X2 inst_7869 ( .A(net_7830), .Z(net_7831) );
CLKBUF_X2 inst_14359 ( .A(net_14320), .Z(net_14321) );
SDFF_X2 inst_1128 ( .SI(net_6679), .Q(net_6679), .D(net_3779), .SE(net_3465), .CK(net_9075) );
INV_X4 inst_4988 ( .ZN(net_867), .A(net_683) );
DFF_X1 inst_6524 ( .QN(net_7440), .D(net_5427), .CK(net_10089) );
CLKBUF_X2 inst_8009 ( .A(net_7970), .Z(net_7971) );
CLKBUF_X2 inst_11325 ( .A(net_9111), .Z(net_11287) );
NAND2_X2 inst_3222 ( .ZN(net_4704), .A2(net_3986), .A1(net_1868) );
NAND2_X2 inst_3759 ( .A1(net_6776), .A2(net_1635), .ZN(net_1586) );
CLKBUF_X2 inst_10928 ( .A(net_8856), .Z(net_10890) );
AOI22_X2 inst_7422 ( .A1(net_2970), .B1(net_2772), .ZN(net_2770), .A2(net_240), .B2(net_166) );
CLKBUF_X2 inst_14216 ( .A(net_14177), .Z(net_14178) );
CLKBUF_X2 inst_11677 ( .A(net_9144), .Z(net_11639) );
CLKBUF_X2 inst_11559 ( .A(net_10597), .Z(net_11521) );
CLKBUF_X2 inst_10064 ( .A(net_10025), .Z(net_10026) );
CLKBUF_X2 inst_10999 ( .A(net_10960), .Z(net_10961) );
NAND2_X2 inst_4070 ( .A1(net_7203), .A2(net_1648), .ZN(net_982) );
CLKBUF_X2 inst_9077 ( .A(net_8955), .Z(net_9039) );
OAI21_X2 inst_1924 ( .ZN(net_5121), .A(net_4755), .B2(net_3941), .B1(net_1073) );
CLKBUF_X2 inst_9023 ( .A(net_8984), .Z(net_8985) );
CLKBUF_X2 inst_12714 ( .A(net_12675), .Z(net_12676) );
CLKBUF_X2 inst_10502 ( .A(net_10463), .Z(net_10464) );
CLKBUF_X2 inst_10244 ( .A(net_7996), .Z(net_10206) );
AOI21_X2 inst_7650 ( .B2(net_3439), .ZN(net_3396), .A(net_3219), .B1(net_3073) );
INV_X4 inst_4748 ( .ZN(net_2752), .A(net_2629) );
NAND2_X2 inst_4160 ( .A1(net_7529), .ZN(net_919), .A2(net_635) );
INV_X4 inst_5685 ( .A(net_6081), .ZN(net_3544) );
CLKBUF_X2 inst_8296 ( .A(net_8257), .Z(net_8258) );
CLKBUF_X2 inst_12160 ( .A(net_12121), .Z(net_12122) );
SDFF_X2 inst_961 ( .Q(net_6439), .D(net_6439), .SE(net_3820), .SI(net_3810), .CK(net_8862) );
NAND2_X2 inst_3255 ( .ZN(net_3870), .A2(net_3869), .A1(net_3862) );
CLKBUF_X2 inst_12246 ( .A(net_10499), .Z(net_12208) );
CLKBUF_X2 inst_13119 ( .A(net_13080), .Z(net_13081) );
OAI22_X2 inst_1590 ( .A1(net_3299), .B2(net_3200), .A2(net_3187), .ZN(net_3172), .B1(net_453) );
CLKBUF_X2 inst_11082 ( .A(net_11043), .Z(net_11044) );
AOI222_X2 inst_7591 ( .A1(net_7387), .ZN(net_5410), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_350), .C2(net_348) );
CLKBUF_X2 inst_12800 ( .A(net_9097), .Z(net_12762) );
CLKBUF_X2 inst_8077 ( .A(net_8038), .Z(net_8039) );
CLKBUF_X2 inst_10931 ( .A(net_10892), .Z(net_10893) );
CLKBUF_X2 inst_10648 ( .A(net_10609), .Z(net_10610) );
CLKBUF_X2 inst_8332 ( .A(net_8253), .Z(net_8294) );
DFF_X2 inst_6229 ( .QN(net_7098), .D(net_3718), .CK(net_9712) );
SDFF_X2 inst_399 ( .SI(net_7341), .Q(net_7341), .D(net_4778), .SE(net_3856), .CK(net_9908) );
NOR2_X2 inst_2318 ( .A2(net_6220), .A1(net_5840), .ZN(net_5823) );
INV_X4 inst_5347 ( .A(net_6138), .ZN(net_3657) );
CLKBUF_X2 inst_12433 ( .A(net_11325), .Z(net_12395) );
INV_X4 inst_5103 ( .ZN(net_708), .A(net_615) );
NAND2_X2 inst_3957 ( .A2(net_1696), .ZN(net_1328), .A1(net_1327) );
CLKBUF_X2 inst_11364 ( .A(net_8662), .Z(net_11326) );
CLKBUF_X2 inst_9953 ( .A(net_8145), .Z(net_9915) );
NAND2_X2 inst_4020 ( .A1(net_6527), .A2(net_1645), .ZN(net_1032) );
CLKBUF_X2 inst_13404 ( .A(net_13365), .Z(net_13366) );
CLKBUF_X2 inst_8489 ( .A(net_7976), .Z(net_8451) );
NOR2_X2 inst_2316 ( .A2(net_6222), .A1(net_5840), .ZN(net_5825) );
NAND3_X2 inst_2737 ( .ZN(net_2364), .A3(net_1563), .A1(net_1427), .A2(net_999) );
DFF_X1 inst_6654 ( .QN(net_7661), .D(net_5191), .CK(net_13063) );
CLKBUF_X2 inst_14266 ( .A(net_7899), .Z(net_14228) );
SDFF_X2 inst_499 ( .Q(net_7117), .D(net_7117), .SI(net_3897), .SE(net_3888), .CK(net_7921) );
SDFF_X2 inst_1299 ( .Q(net_6361), .SI(net_6360), .D(net_3125), .SE(net_392), .CK(net_13597) );
CLKBUF_X2 inst_8404 ( .A(net_8365), .Z(net_8366) );
DFF_X1 inst_6450 ( .QN(net_6101), .D(net_5720), .CK(net_12054) );
CLKBUF_X2 inst_13487 ( .A(net_13448), .Z(net_13449) );
CLKBUF_X2 inst_10404 ( .A(net_9396), .Z(net_10366) );
DFF_X2 inst_6175 ( .Q(net_6399), .D(net_6398), .CK(net_14194) );
CLKBUF_X2 inst_9468 ( .A(net_9429), .Z(net_9430) );
SDFF_X2 inst_674 ( .Q(net_6738), .D(net_6738), .SE(net_3815), .SI(net_3812), .CK(net_11161) );
NOR2_X2 inst_2400 ( .ZN(net_3774), .A1(net_3773), .A2(net_3772) );
INV_X4 inst_5259 ( .ZN(net_861), .A(net_484) );
OAI22_X2 inst_1451 ( .B1(net_4855), .A2(net_4622), .ZN(net_4620), .B2(net_4619), .A1(net_4216) );
NAND2_X2 inst_4082 ( .A1(net_6523), .A2(net_1645), .ZN(net_970) );
INV_X4 inst_4781 ( .ZN(net_2632), .A(net_1662) );
INV_X4 inst_5518 ( .A(net_6160), .ZN(net_3523) );
CLKBUF_X2 inst_14151 ( .A(net_13627), .Z(net_14113) );
CLKBUF_X2 inst_14207 ( .A(net_11427), .Z(net_14169) );
CLKBUF_X2 inst_10859 ( .A(net_8646), .Z(net_10821) );
NOR2_X4 inst_2253 ( .ZN(net_5633), .A1(net_5478), .A2(net_4438) );
CLKBUF_X2 inst_13670 ( .A(net_10827), .Z(net_13632) );
OAI21_X2 inst_2009 ( .B1(net_5905), .B2(net_4518), .ZN(net_4502), .A(net_3670) );
CLKBUF_X2 inst_10115 ( .A(net_10076), .Z(net_10077) );
CLKBUF_X2 inst_9674 ( .A(net_9635), .Z(net_9636) );
SDFF_X2 inst_501 ( .Q(net_6481), .D(net_6481), .SE(net_3904), .SI(net_3898), .CK(net_8429) );
NAND2_X4 inst_2868 ( .A1(net_5885), .ZN(net_4271), .A2(net_2581) );
CLKBUF_X2 inst_12254 ( .A(net_12215), .Z(net_12216) );
OAI21_X2 inst_2093 ( .B2(net_4485), .ZN(net_4323), .B1(net_4105), .A(net_3644) );
DFF_X1 inst_6522 ( .QN(net_7438), .D(net_5429), .CK(net_9283) );
SDFF_X2 inst_1081 ( .SI(net_7208), .Q(net_7208), .D(net_3811), .SE(net_3750), .CK(net_12145) );
NAND2_X2 inst_3195 ( .ZN(net_4731), .A2(net_3986), .A1(net_1902) );
CLKBUF_X2 inst_8873 ( .A(net_8834), .Z(net_8835) );
CLKBUF_X2 inst_10731 ( .A(net_10692), .Z(net_10693) );
CLKBUF_X2 inst_12261 ( .A(net_12222), .Z(net_12223) );
OAI21_X2 inst_1832 ( .ZN(net_5346), .B1(net_5345), .A(net_4359), .B2(net_3856) );
NAND2_X4 inst_2905 ( .A2(net_5876), .ZN(net_2627), .A1(net_2626) );
CLKBUF_X2 inst_13241 ( .A(net_13202), .Z(net_13203) );
NAND3_X2 inst_2819 ( .ZN(net_2279), .A3(net_1606), .A1(net_1314), .A2(net_1015) );
CLKBUF_X2 inst_12263 ( .A(net_12224), .Z(net_12225) );
SDFF_X2 inst_640 ( .SI(net_6625), .Q(net_6625), .SE(net_3851), .D(net_3802), .CK(net_10052) );
INV_X8 inst_4562 ( .A(net_3222), .ZN(net_1222) );
CLKBUF_X2 inst_9893 ( .A(net_9854), .Z(net_9855) );
AOI222_X2 inst_7500 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2072), .A1(net_2071), .B1(net_2070), .C1(net_2069) );
DFF_X2 inst_6293 ( .Q(net_6383), .D(net_6382), .CK(net_14166) );
OAI22_X2 inst_1478 ( .B1(net_4855), .B2(net_4479), .A2(net_4230), .A1(net_4228), .ZN(net_4213) );
INV_X2 inst_6098 ( .A(net_7320), .ZN(net_1772) );
CLKBUF_X2 inst_9963 ( .A(net_9924), .Z(net_9925) );
SDFF_X2 inst_1114 ( .Q(net_6826), .D(net_3432), .SI(net_3431), .SE(net_2256), .CK(net_11382) );
CLKBUF_X2 inst_7982 ( .A(net_7943), .Z(net_7944) );
CLKBUF_X2 inst_9327 ( .A(net_9288), .Z(net_9289) );
CLKBUF_X2 inst_9535 ( .A(net_9496), .Z(net_9497) );
NAND2_X2 inst_4163 ( .ZN(net_927), .A1(net_547), .A2(net_477) );
CLKBUF_X2 inst_9020 ( .A(net_8610), .Z(net_8982) );
CLKBUF_X2 inst_12957 ( .A(net_12918), .Z(net_12919) );
CLKBUF_X2 inst_9085 ( .A(net_9041), .Z(net_9047) );
CLKBUF_X2 inst_13739 ( .A(net_11390), .Z(net_13701) );
OAI21_X2 inst_1982 ( .ZN(net_4848), .B1(net_4847), .A(net_4537), .B2(net_3870) );
INV_X2 inst_6075 ( .A(net_7467), .ZN(net_2070) );
OAI21_X2 inst_2089 ( .B1(net_5913), .B2(net_4415), .ZN(net_4399), .A(net_3476) );
CLKBUF_X2 inst_11805 ( .A(net_11766), .Z(net_11767) );
CLKBUF_X2 inst_11378 ( .A(net_11339), .Z(net_11340) );
OAI21_X2 inst_1849 ( .B1(net_5343), .ZN(net_5323), .A(net_4363), .B2(net_3853) );
OAI221_X2 inst_1679 ( .ZN(net_3370), .A(net_3181), .B2(net_2985), .C2(net_2903), .C1(net_2868), .B1(net_1963) );
INV_X4 inst_5540 ( .A(net_6133), .ZN(net_3627) );
CLKBUF_X2 inst_11123 ( .A(net_8589), .Z(net_11085) );
OAI21_X2 inst_1976 ( .B1(net_4870), .ZN(net_4860), .A(net_4365), .B2(net_3853) );
INV_X4 inst_4932 ( .ZN(net_764), .A(net_763) );
NAND3_X2 inst_2744 ( .ZN(net_2357), .A3(net_1607), .A1(net_1319), .A2(net_952) );
NAND2_X2 inst_3681 ( .A2(net_1798), .ZN(net_1771), .A1(net_1770) );
DFF_X1 inst_6909 ( .D(net_2530), .Q(net_156), .CK(net_9420) );
CLKBUF_X2 inst_13238 ( .A(net_8178), .Z(net_13200) );
NOR3_X2 inst_2215 ( .A3(net_2222), .ZN(net_1835), .A1(net_861), .A2(net_437) );
SDFF_X2 inst_337 ( .SI(net_7462), .Q(net_7462), .D(net_5095), .SE(net_3993), .CK(net_12521) );
OAI21_X2 inst_1855 ( .ZN(net_5263), .B1(net_5237), .A(net_4548), .B2(net_3870) );
INV_X4 inst_5277 ( .ZN(net_3919), .A(net_416) );
NOR2_X2 inst_2384 ( .ZN(net_4295), .A1(net_4151), .A2(net_4150) );
INV_X4 inst_4614 ( .ZN(net_4208), .A(net_4077) );
CLKBUF_X2 inst_11564 ( .A(net_11525), .Z(net_11526) );
CLKBUF_X2 inst_9606 ( .A(net_8296), .Z(net_9568) );
SDFF_X2 inst_1212 ( .D(net_7802), .SI(net_7069), .Q(net_7069), .SE(net_3742), .CK(net_8985) );
CLKBUF_X2 inst_11193 ( .A(net_11154), .Z(net_11155) );
SDFF_X2 inst_670 ( .Q(net_6702), .D(net_6702), .SE(net_3871), .SI(net_3814), .CK(net_8967) );
DFF_X2 inst_6220 ( .QN(net_6692), .D(net_3728), .CK(net_9716) );
CLKBUF_X2 inst_13355 ( .A(net_13316), .Z(net_13317) );
NAND2_X2 inst_4180 ( .A1(net_5935), .ZN(net_2730), .A2(net_769) );
INV_X2 inst_5789 ( .A(net_5973), .ZN(net_2239) );
CLKBUF_X2 inst_11105 ( .A(net_11066), .Z(net_11067) );
CLKBUF_X2 inst_13775 ( .A(net_13736), .Z(net_13737) );
CLKBUF_X2 inst_9612 ( .A(net_9573), .Z(net_9574) );
NAND2_X2 inst_3901 ( .A2(net_1696), .ZN(net_1410), .A1(net_1409) );
CLKBUF_X2 inst_9262 ( .A(net_9223), .Z(net_9224) );
DFF_X1 inst_6679 ( .QN(net_7257), .D(net_5146), .CK(net_12258) );
AOI21_X2 inst_7738 ( .B1(net_7138), .ZN(net_4458), .B2(net_2582), .A(net_2296) );
NOR2_X2 inst_2396 ( .A2(net_3996), .ZN(net_3987), .A1(net_2577) );
CLKBUF_X2 inst_10232 ( .A(net_9694), .Z(net_10194) );
CLKBUF_X2 inst_10281 ( .A(net_10242), .Z(net_10243) );
CLKBUF_X2 inst_14295 ( .A(net_14256), .Z(net_14257) );
CLKBUF_X2 inst_14093 ( .A(net_8326), .Z(net_14055) );
INV_X2 inst_5898 ( .A(net_7355), .ZN(net_2210) );
CLKBUF_X2 inst_8647 ( .A(net_8608), .Z(net_8609) );
CLKBUF_X2 inst_10845 ( .A(net_10480), .Z(net_10807) );
SDFF_X2 inst_246 ( .Q(net_6348), .SI(net_6347), .D(net_3619), .SE(net_392), .CK(net_14132) );
INV_X2 inst_5908 ( .A(net_7354), .ZN(net_1992) );
CLKBUF_X2 inst_12384 ( .A(net_12345), .Z(net_12346) );
SDFF_X2 inst_635 ( .SI(net_6647), .Q(net_6647), .SE(net_3851), .D(net_3796), .CK(net_10652) );
NAND2_X1 inst_4443 ( .A2(net_2131), .ZN(net_1321), .A1(net_1320) );
CLKBUF_X2 inst_9814 ( .A(net_9775), .Z(net_9776) );
INV_X2 inst_5787 ( .A(net_3452), .ZN(net_2262) );
SDFF_X2 inst_807 ( .Q(net_6980), .D(net_6980), .SE(net_3891), .SI(net_3786), .CK(net_11907) );
SDFF_X2 inst_705 ( .SI(net_6777), .Q(net_6777), .SE(net_3816), .D(net_3784), .CK(net_11327) );
CLKBUF_X2 inst_10569 ( .A(net_10530), .Z(net_10531) );
CLKBUF_X2 inst_8510 ( .A(net_8374), .Z(net_8472) );
SDFF_X2 inst_911 ( .Q(net_7148), .D(net_7148), .SE(net_3903), .SI(net_3808), .CK(net_7852) );
SDFF_X2 inst_519 ( .SI(net_6626), .Q(net_6626), .D(net_3892), .SE(net_3850), .CK(net_12938) );
CLKBUF_X2 inst_10921 ( .A(net_10106), .Z(net_10883) );
AOI21_X2 inst_7641 ( .B1(net_5893), .ZN(net_3914), .B2(net_3913), .A(net_2600) );
NAND2_X2 inst_3796 ( .A1(net_6489), .A2(net_1642), .ZN(net_1549) );
CLKBUF_X2 inst_9359 ( .A(net_9145), .Z(net_9321) );
SDFF_X2 inst_1003 ( .SI(net_7799), .Q(net_6462), .D(net_6462), .SE(net_3904), .CK(net_11252) );
CLKBUF_X2 inst_13804 ( .A(net_13765), .Z(net_13766) );
CLKBUF_X2 inst_12758 ( .A(net_12719), .Z(net_12720) );
CLKBUF_X2 inst_12174 ( .A(net_9826), .Z(net_12136) );
SDFF_X2 inst_1053 ( .Q(net_7242), .D(net_7242), .SE(net_3822), .SI(net_338), .CK(net_12654) );
INV_X4 inst_5158 ( .A(net_1227), .ZN(net_555) );
CLKBUF_X2 inst_10284 ( .A(net_9025), .Z(net_10246) );
NAND2_X2 inst_3469 ( .A1(net_6013), .A2(net_3105), .ZN(net_2755) );
NAND3_X2 inst_2774 ( .ZN(net_2326), .A3(net_1641), .A1(net_1392), .A2(net_955) );
INV_X2 inst_6026 ( .A(net_7626), .ZN(net_1907) );
DFF_X1 inst_6871 ( .D(net_2559), .Q(net_205), .CK(net_10062) );
CLKBUF_X2 inst_12202 ( .A(net_9564), .Z(net_12164) );
INV_X4 inst_5456 ( .A(net_7530), .ZN(net_600) );
SDFF_X2 inst_239 ( .Q(net_6355), .SI(net_6354), .D(net_3601), .SE(net_392), .CK(net_13953) );
INV_X4 inst_4577 ( .ZN(net_5498), .A(net_5497) );
SDFF_X2 inst_1193 ( .D(net_7807), .SI(net_7074), .Q(net_7074), .SE(net_3742), .CK(net_8051) );
OAI21_X2 inst_2080 ( .B2(net_4415), .ZN(net_4410), .B1(net_4026), .A(net_3504) );
OAI22_X2 inst_1625 ( .B2(net_2820), .ZN(net_2719), .A2(net_2718), .B1(net_896), .A1(net_515) );
AOI21_X2 inst_7710 ( .B1(net_6872), .ZN(net_4104), .B2(net_2579), .A(net_2353) );
SDFF_X2 inst_593 ( .Q(net_6563), .D(net_6563), .SE(net_3823), .SI(net_3799), .CK(net_10055) );
INV_X2 inst_5707 ( .ZN(net_4311), .A(net_4219) );
NOR2_X4 inst_2223 ( .ZN(net_5675), .A1(net_5547), .A2(net_4512) );
CLKBUF_X2 inst_10582 ( .A(net_8415), .Z(net_10544) );
INV_X8 inst_4522 ( .ZN(net_3734), .A(net_3116) );
INV_X16 inst_6137 ( .ZN(net_1635), .A(net_771) );
CLKBUF_X2 inst_12426 ( .A(net_12387), .Z(net_12388) );
CLKBUF_X2 inst_10099 ( .A(net_10060), .Z(net_10061) );
CLKBUF_X2 inst_12395 ( .A(net_12356), .Z(net_12357) );
SDFF_X2 inst_601 ( .Q(net_6604), .D(net_6604), .SE(net_3830), .SI(net_3811), .CK(net_9346) );
INV_X2 inst_5738 ( .ZN(net_3727), .A(net_3433) );
INV_X2 inst_6091 ( .A(net_7291), .ZN(net_2208) );
CLKBUF_X2 inst_13709 ( .A(net_8714), .Z(net_13671) );
AOI22_X2 inst_7391 ( .A2(net_3439), .B1(net_2970), .ZN(net_2928), .A1(net_2927), .B2(net_231) );
CLKBUF_X2 inst_7952 ( .A(net_7913), .Z(net_7914) );
AND2_X4 inst_7845 ( .A2(net_6410), .ZN(net_1668), .A1(net_618) );
CLKBUF_X2 inst_8097 ( .A(net_8058), .Z(net_8059) );
CLKBUF_X2 inst_9065 ( .A(net_9026), .Z(net_9027) );
CLKBUF_X2 inst_10045 ( .A(net_10006), .Z(net_10007) );
SDFF_X2 inst_479 ( .Q(net_6836), .D(net_6836), .SE(net_3893), .SI(net_3890), .CK(net_8900) );
OAI21_X2 inst_1773 ( .B1(net_5442), .ZN(net_5421), .A(net_4700), .B2(net_3989) );
CLKBUF_X2 inst_10448 ( .A(net_10409), .Z(net_10410) );
NOR2_X2 inst_2344 ( .A2(net_6003), .A1(net_5778), .ZN(net_5708) );
CLKBUF_X2 inst_10278 ( .A(net_8049), .Z(net_10240) );
CLKBUF_X2 inst_10133 ( .A(net_10054), .Z(net_10095) );
NAND2_X2 inst_3326 ( .ZN(net_3594), .A1(net_3593), .A2(net_3228) );
AOI22_X2 inst_7288 ( .B1(net_7225), .A1(net_7193), .A2(net_5244), .B2(net_5243), .ZN(net_5217) );
AOI21_X2 inst_7683 ( .B1(net_7002), .ZN(net_4479), .A(net_2471), .B2(net_1100) );
SDFF_X2 inst_771 ( .Q(net_6866), .D(net_6866), .SE(net_3901), .SI(net_3798), .CK(net_8932) );
OAI22_X2 inst_1583 ( .B2(net_3200), .ZN(net_3195), .A1(net_3194), .A2(net_3193), .B1(net_591) );
CLKBUF_X2 inst_12892 ( .A(net_11542), .Z(net_12854) );
NAND2_X1 inst_4387 ( .ZN(net_4340), .A2(net_3859), .A1(net_2007) );
CLKBUF_X2 inst_9420 ( .A(net_9381), .Z(net_9382) );
DFF_X2 inst_6325 ( .QN(net_7805), .CK(net_8679), .D(x1501) );
CLKBUF_X2 inst_11552 ( .A(net_11513), .Z(net_11514) );
DFFR_X1 inst_7113 ( .QN(net_5857), .D(net_5797), .CK(net_12428), .RN(x1822) );
INV_X2 inst_5780 ( .ZN(net_2699), .A(net_392) );
AOI22_X2 inst_7324 ( .ZN(net_3430), .A2(net_3429), .B2(net_3428), .A1(net_1303), .B1(net_904) );
CLKBUF_X2 inst_9334 ( .A(net_9295), .Z(net_9296) );
AOI22_X2 inst_7402 ( .B1(net_5939), .A1(net_2911), .A2(net_2838), .ZN(net_2836), .B2(net_204) );
CLKBUF_X2 inst_8169 ( .A(net_8130), .Z(net_8131) );
CLKBUF_X2 inst_12945 ( .A(net_11375), .Z(net_12907) );
CLKBUF_X2 inst_10523 ( .A(net_10484), .Z(net_10485) );
CLKBUF_X2 inst_13873 ( .A(net_13834), .Z(net_13835) );
INV_X2 inst_5782 ( .ZN(net_2448), .A(net_2447) );
CLKBUF_X2 inst_10520 ( .A(net_7922), .Z(net_10482) );
INV_X8 inst_4497 ( .ZN(net_3901), .A(net_3151) );
SDFF_X2 inst_1319 ( .D(net_6385), .SE(net_5801), .SI(net_330), .Q(net_330), .CK(net_13858) );
NAND3_X2 inst_2651 ( .A3(net_5957), .A2(net_5956), .ZN(net_3949), .A1(net_2836) );
INV_X4 inst_4756 ( .A(net_3252), .ZN(net_2777) );
NAND2_X2 inst_4201 ( .A2(net_769), .ZN(net_625), .A1(net_624) );
INV_X4 inst_5658 ( .A(net_7567), .ZN(net_1898) );
XNOR2_X2 inst_48 ( .ZN(net_2261), .A(net_2260), .B(net_2259) );
SDFF_X2 inst_358 ( .SI(net_7606), .Q(net_7606), .D(net_4791), .SE(net_3870), .CK(net_13256) );
INV_X8 inst_4462 ( .ZN(net_5315), .A(net_4289) );
OAI21_X2 inst_1756 ( .ZN(net_5445), .B1(net_5444), .A(net_4668), .B2(net_3993) );
NOR2_X4 inst_2246 ( .ZN(net_5640), .A1(net_5486), .A2(net_4452) );
AOI222_X2 inst_7507 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2044), .A1(net_2043), .B1(net_2042), .C1(net_2041) );
CLKBUF_X2 inst_14037 ( .A(net_13998), .Z(net_13999) );
CLKBUF_X2 inst_8794 ( .A(net_8755), .Z(net_8756) );
DFF_X1 inst_6766 ( .QN(net_6126), .D(net_4663), .CK(net_7827) );
CLKBUF_X2 inst_9309 ( .A(net_9005), .Z(net_9271) );
DFFR_X2 inst_7108 ( .D(net_1948), .QN(net_118), .CK(net_9580), .RN(x1822) );
SDFF_X2 inst_443 ( .Q(net_7397), .D(net_7397), .SE(net_3994), .SI(net_362), .CK(net_9628) );
CLKBUF_X2 inst_14177 ( .A(net_14138), .Z(net_14139) );
CLKBUF_X2 inst_11022 ( .A(net_10983), .Z(net_10984) );
CLKBUF_X2 inst_8766 ( .A(net_8727), .Z(net_8728) );
SDFF_X2 inst_655 ( .Q(net_6713), .D(net_6713), .SE(net_3871), .SI(net_3807), .CK(net_11355) );
NAND2_X1 inst_4259 ( .ZN(net_4664), .A2(net_3993), .A1(net_1361) );
INV_X2 inst_5914 ( .A(net_7361), .ZN(net_2054) );
CLKBUF_X2 inst_12152 ( .A(net_12113), .Z(net_12114) );
INV_X2 inst_5817 ( .A(net_1635), .ZN(net_1096) );
CLKBUF_X2 inst_9060 ( .A(net_7998), .Z(net_9022) );
CLKBUF_X2 inst_8422 ( .A(net_7960), .Z(net_8384) );
INV_X2 inst_5934 ( .A(net_7446), .ZN(net_1361) );
CLKBUF_X2 inst_9373 ( .A(net_9334), .Z(net_9335) );
OAI21_X2 inst_1700 ( .ZN(net_5594), .A(net_5268), .B2(net_4479), .B1(net_4228) );
CLKBUF_X2 inst_11316 ( .A(net_11277), .Z(net_11278) );
NAND3_X2 inst_2571 ( .ZN(net_5768), .A1(net_5663), .A2(net_5291), .A3(net_4237) );
NAND2_X1 inst_4438 ( .A2(net_2131), .ZN(net_1364), .A1(net_1363) );
CLKBUF_X2 inst_12481 ( .A(net_10310), .Z(net_12443) );
DFF_X1 inst_6662 ( .QN(net_7654), .D(net_5178), .CK(net_10553) );
CLKBUF_X2 inst_8800 ( .A(net_8761), .Z(net_8762) );
SDFF_X2 inst_730 ( .Q(net_6846), .D(net_6846), .SE(net_3893), .SI(net_3808), .CK(net_8880) );
CLKBUF_X2 inst_11430 ( .A(net_11391), .Z(net_11392) );
CLKBUF_X2 inst_10116 ( .A(net_10077), .Z(net_10078) );
DFF_X2 inst_6303 ( .Q(net_6382), .D(net_6381), .CK(net_14162) );
DFF_X1 inst_6754 ( .QN(net_6146), .D(net_4857), .CK(net_9140) );
SDFF_X2 inst_321 ( .SI(net_7485), .Q(net_7485), .D(net_5098), .SE(net_3989), .CK(net_12583) );
INV_X4 inst_5623 ( .A(net_6152), .ZN(net_3619) );
CLKBUF_X2 inst_10977 ( .A(net_7981), .Z(net_10939) );
CLKBUF_X2 inst_9669 ( .A(net_9630), .Z(net_9631) );
CLKBUF_X2 inst_11996 ( .A(net_11957), .Z(net_11958) );
CLKBUF_X2 inst_11516 ( .A(net_11477), .Z(net_11478) );
XNOR2_X2 inst_41 ( .ZN(net_2274), .B(net_1938), .A(net_1937) );
CLKBUF_X2 inst_12569 ( .A(net_9962), .Z(net_12531) );
CLKBUF_X2 inst_11743 ( .A(net_11704), .Z(net_11705) );
NAND2_X2 inst_3131 ( .ZN(net_4832), .A2(net_4153), .A1(net_2178) );
CLKBUF_X2 inst_12684 ( .A(net_12645), .Z(net_12646) );
CLKBUF_X2 inst_13308 ( .A(net_13269), .Z(net_13270) );
CLKBUF_X2 inst_11868 ( .A(net_11829), .Z(net_11830) );
OAI21_X2 inst_1989 ( .B1(net_4849), .ZN(net_4840), .A(net_4560), .B2(net_3866) );
CLKBUF_X2 inst_13260 ( .A(net_11246), .Z(net_13222) );
CLKBUF_X2 inst_9694 ( .A(net_9655), .Z(net_9656) );
SDFF_X2 inst_152 ( .Q(net_6226), .SI(net_6225), .SE(net_392), .D(net_132), .CK(net_14091) );
CLKBUF_X2 inst_8264 ( .A(net_8225), .Z(net_8226) );
INV_X4 inst_5609 ( .ZN(net_608), .A(net_283) );
CLKBUF_X2 inst_11111 ( .A(net_11072), .Z(net_11073) );
DFF_X1 inst_6944 ( .D(net_2233), .Q(net_386), .CK(net_14353) );
CLKBUF_X2 inst_12314 ( .A(net_12275), .Z(net_12276) );
SDFF_X2 inst_1152 ( .SI(net_6814), .Q(net_6814), .D(net_3779), .SE(net_3729), .CK(net_11291) );
DFF_X1 inst_6878 ( .D(net_2513), .Q(net_157), .CK(net_9555) );
DFF_X1 inst_6388 ( .QN(net_6119), .D(net_5700), .CK(net_11199) );
OR2_X4 inst_1400 ( .A2(net_6824), .A1(net_6823), .ZN(net_476) );
CLKBUF_X2 inst_14374 ( .A(net_14335), .Z(net_14336) );
DFF_X1 inst_6517 ( .QN(net_7448), .D(net_5437), .CK(net_9749) );
XNOR2_X2 inst_89 ( .ZN(net_1205), .B(net_1204), .A(net_790) );
INV_X4 inst_5233 ( .A(net_522), .ZN(net_457) );
OAI22_X2 inst_1520 ( .B1(net_4644), .ZN(net_4058), .A1(net_4057), .A2(net_4056), .B2(net_4055) );
DFF_X1 inst_6823 ( .QN(net_5976), .D(net_3015), .CK(net_9748) );
OAI22_X2 inst_1535 ( .B1(net_4637), .A1(net_4030), .B2(net_4029), .ZN(net_4025), .A2(net_4024) );
CLKBUF_X2 inst_14112 ( .A(net_9472), .Z(net_14074) );
CLKBUF_X2 inst_13609 ( .A(net_10519), .Z(net_13571) );
CLKBUF_X2 inst_8670 ( .A(net_8631), .Z(net_8632) );
SDFF_X2 inst_182 ( .Q(net_6272), .SI(net_6271), .D(net_3511), .SE(net_392), .CK(net_13923) );
SDFF_X2 inst_788 ( .SI(net_6917), .Q(net_6917), .SE(net_3781), .D(net_3779), .CK(net_8140) );
SDFF_X2 inst_931 ( .SI(net_7163), .Q(net_7163), .SE(net_3819), .D(net_3797), .CK(net_10488) );
CLKBUF_X2 inst_9205 ( .A(net_9166), .Z(net_9167) );
NAND2_X2 inst_3174 ( .ZN(net_4759), .A2(net_3941), .A1(net_2047) );
AOI222_X2 inst_7526 ( .A2(net_2135), .B2(net_2133), .C2(net_2131), .ZN(net_1988), .A1(net_1987), .B1(net_1986), .C1(net_1985) );
CLKBUF_X2 inst_13391 ( .A(net_11402), .Z(net_13353) );
OAI221_X2 inst_1674 ( .ZN(net_4158), .C2(net_4157), .B2(net_4155), .C1(net_3940), .A(net_3835), .B1(net_1925) );
NAND2_X2 inst_3824 ( .A1(net_7453), .A2(net_1696), .ZN(net_1520) );
INV_X2 inst_5990 ( .A(net_6045), .ZN(net_2834) );
DFF_X1 inst_6895 ( .D(net_2522), .Q(net_168), .CK(net_10221) );
CLKBUF_X2 inst_12807 ( .A(net_12768), .Z(net_12769) );
CLKBUF_X2 inst_8438 ( .A(net_8399), .Z(net_8400) );
OAI22_X2 inst_1579 ( .A1(net_3291), .ZN(net_3206), .B2(net_3200), .A2(net_3144), .B1(net_594) );
INV_X4 inst_5407 ( .A(net_6063), .ZN(net_3374) );
CLKBUF_X2 inst_13482 ( .A(net_13443), .Z(net_13444) );
CLKBUF_X2 inst_8315 ( .A(net_8276), .Z(net_8277) );
SDFF_X2 inst_193 ( .Q(net_6261), .SI(net_6260), .D(net_3493), .SE(net_392), .CK(net_13467) );
NAND2_X2 inst_4089 ( .A1(net_6932), .A2(net_1654), .ZN(net_963) );
CLKBUF_X2 inst_14320 ( .A(net_14281), .Z(net_14282) );
CLKBUF_X2 inst_11704 ( .A(net_11665), .Z(net_11666) );
OR2_X2 inst_1415 ( .ZN(net_3764), .A2(net_796), .A1(net_458) );
OAI21_X2 inst_1709 ( .ZN(net_5585), .A(net_5152), .B2(net_4437), .B1(net_4057) );
CLKBUF_X2 inst_12089 ( .A(net_12050), .Z(net_12051) );
CLKBUF_X2 inst_13631 ( .A(net_13592), .Z(net_13593) );
NAND2_X2 inst_3301 ( .ZN(net_3644), .A1(net_3643), .A2(net_3229) );
INV_X2 inst_5997 ( .A(net_7478), .ZN(net_2084) );
DFF_X1 inst_6469 ( .QN(net_6170), .D(net_5590), .CK(net_7962) );
NOR3_X2 inst_2202 ( .ZN(net_3156), .A1(net_2989), .A3(net_1747), .A2(net_1101) );
AOI222_X2 inst_7531 ( .C1(net_7671), .A1(net_7639), .B2(net_2135), .C2(net_2133), .ZN(net_1911), .A2(net_1910), .B1(net_1909) );
CLKBUF_X2 inst_11673 ( .A(net_11634), .Z(net_11635) );
NAND2_X2 inst_3180 ( .ZN(net_4753), .A2(net_3941), .A1(net_2029) );
CLKBUF_X2 inst_7969 ( .A(net_7930), .Z(net_7931) );
INV_X4 inst_4737 ( .A(net_5974), .ZN(net_3875) );
CLKBUF_X2 inst_9965 ( .A(net_9926), .Z(net_9927) );
CLKBUF_X2 inst_10618 ( .A(net_10579), .Z(net_10580) );
NAND2_X2 inst_2987 ( .A1(net_6753), .A2(net_5033), .ZN(net_5024) );
CLKBUF_X2 inst_12571 ( .A(net_12326), .Z(net_12533) );
CLKBUF_X2 inst_11645 ( .A(net_11606), .Z(net_11607) );
CLKBUF_X2 inst_13433 ( .A(net_13394), .Z(net_13395) );
INV_X4 inst_5578 ( .A(net_7698), .ZN(net_853) );
CLKBUF_X2 inst_11853 ( .A(net_11814), .Z(net_11815) );
INV_X2 inst_5884 ( .A(net_7616), .ZN(net_1193) );
CLKBUF_X2 inst_13396 ( .A(net_9623), .Z(net_13358) );
CLKBUF_X2 inst_11170 ( .A(net_11131), .Z(net_11132) );
CLKBUF_X2 inst_8655 ( .A(net_8616), .Z(net_8617) );
CLKBUF_X2 inst_11459 ( .A(net_10775), .Z(net_11421) );
INV_X4 inst_4599 ( .ZN(net_5041), .A(net_4290) );
CLKBUF_X2 inst_8147 ( .A(net_8108), .Z(net_8109) );
INV_X2 inst_5906 ( .A(net_7513), .ZN(net_2164) );
INV_X4 inst_4677 ( .ZN(net_3454), .A(net_3453) );
CLKBUF_X2 inst_12874 ( .A(net_12835), .Z(net_12836) );
NOR2_X2 inst_2473 ( .A2(net_5778), .ZN(net_2672), .A1(net_2609) );
INV_X4 inst_5516 ( .A(net_6824), .ZN(net_450) );
OAI21_X2 inst_1698 ( .ZN(net_5596), .A(net_5270), .B2(net_4619), .B1(net_4228) );
CLKBUF_X2 inst_11698 ( .A(net_10075), .Z(net_11660) );
SDFF_X2 inst_944 ( .SI(net_7187), .Q(net_7187), .SE(net_3819), .D(net_3796), .CK(net_8698) );
INV_X4 inst_5248 ( .A(net_838), .ZN(net_444) );
DFFR_X1 inst_7125 ( .Q(net_6003), .D(net_4799), .CK(net_10032), .RN(x1822) );
CLKBUF_X2 inst_12442 ( .A(net_12403), .Z(net_12404) );
INV_X8 inst_4516 ( .ZN(net_3904), .A(net_3203) );
CLKBUF_X2 inst_7992 ( .A(net_7953), .Z(net_7954) );
CLKBUF_X2 inst_13952 ( .A(net_13913), .Z(net_13914) );
SDFF_X2 inst_459 ( .SI(net_7807), .Q(net_7145), .D(net_7145), .SE(net_3903), .CK(net_7899) );
CLKBUF_X2 inst_8259 ( .A(net_7939), .Z(net_8221) );
CLKBUF_X2 inst_11737 ( .A(net_11698), .Z(net_11699) );
CLKBUF_X2 inst_8532 ( .A(net_8493), .Z(net_8494) );
NAND2_X4 inst_2864 ( .ZN(net_4287), .A1(net_4278), .A2(net_791) );
NAND2_X2 inst_3476 ( .ZN(net_2707), .A2(net_2706), .A1(net_2453) );
CLKBUF_X2 inst_10084 ( .A(net_10045), .Z(net_10046) );
AOI222_X2 inst_7461 ( .ZN(net_2213), .A1(net_2212), .A2(net_2211), .B1(net_2210), .B2(net_2209), .C1(net_2208), .C2(net_2207) );
CLKBUF_X2 inst_12861 ( .A(net_12822), .Z(net_12823) );
NAND2_X2 inst_3789 ( .A1(net_6901), .A2(net_1639), .ZN(net_1556) );
DFFR_X2 inst_7096 ( .D(net_1955), .QN(net_124), .CK(net_12329), .RN(x1822) );
CLKBUF_X2 inst_13723 ( .A(net_13684), .Z(net_13685) );
NAND2_X2 inst_3393 ( .ZN(net_3760), .A2(net_3364), .A1(net_2885) );
CLKBUF_X2 inst_8613 ( .A(net_8574), .Z(net_8575) );
SDFF_X2 inst_367 ( .SI(net_7638), .Q(net_7638), .D(net_4791), .SE(net_3867), .CK(net_13249) );
CLKBUF_X2 inst_8148 ( .A(net_7834), .Z(net_8110) );
CLKBUF_X2 inst_11589 ( .A(net_8029), .Z(net_11551) );
SDFF_X2 inst_957 ( .Q(net_6424), .D(net_6424), .SE(net_3820), .SI(net_3792), .CK(net_11556) );
INV_X4 inst_4976 ( .ZN(net_863), .A(net_795) );
CLKBUF_X2 inst_9657 ( .A(net_9618), .Z(net_9619) );
NAND2_X2 inst_3409 ( .ZN(net_4107), .A2(net_3337), .A1(net_2704) );
OAI21_X2 inst_1871 ( .ZN(net_5238), .B1(net_5237), .A(net_4592), .B2(net_3867) );
CLKBUF_X2 inst_13252 ( .A(net_13213), .Z(net_13214) );
NAND2_X2 inst_3591 ( .ZN(net_2409), .A2(net_1911), .A1(net_1346) );
NOR2_X2 inst_2300 ( .A2(net_6187), .A1(net_5843), .ZN(net_5842) );
INV_X2 inst_5970 ( .A(net_7657), .ZN(net_1867) );
DFF_X1 inst_6460 ( .QN(net_6129), .D(net_5599), .CK(net_10959) );
AOI222_X2 inst_7552 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1847), .A1(net_1846), .B1(net_1845), .C1(net_1844) );
CLKBUF_X2 inst_10800 ( .A(net_10761), .Z(net_10762) );
SDFF_X2 inst_450 ( .D(net_6390), .SE(net_6052), .SI(net_315), .Q(net_315), .CK(net_13730) );
CLKBUF_X2 inst_9723 ( .A(net_9684), .Z(net_9685) );
CLKBUF_X2 inst_11694 ( .A(net_9290), .Z(net_11656) );
SDFF_X2 inst_745 ( .Q(net_6834), .D(net_6834), .SE(net_3893), .SI(net_3798), .CK(net_8942) );
SDFF_X2 inst_520 ( .SI(net_7807), .Q(net_6708), .D(net_6708), .SE(net_3871), .CK(net_10778) );
INV_X2 inst_5717 ( .ZN(net_4249), .A(net_4119) );
NAND2_X2 inst_3658 ( .A1(net_7069), .ZN(net_1805), .A2(net_791) );
DFFR_X2 inst_7024 ( .D(net_3276), .QN(net_278), .CK(net_12643), .RN(x1822) );
CLKBUF_X2 inst_10019 ( .A(net_9980), .Z(net_9981) );
CLKBUF_X2 inst_11622 ( .A(net_9290), .Z(net_11584) );
CLKBUF_X2 inst_11667 ( .A(net_11470), .Z(net_11629) );
OAI21_X2 inst_2032 ( .B2(net_4476), .ZN(net_4471), .B1(net_4227), .A(net_3524) );
INV_X8 inst_4554 ( .ZN(net_2207), .A(net_811) );
INV_X2 inst_5977 ( .A(net_7358), .ZN(net_2078) );
NAND2_X2 inst_4113 ( .A2(net_1228), .ZN(net_1183), .A1(net_385) );
OAI21_X2 inst_2026 ( .ZN(net_4480), .B1(net_4479), .B2(net_4476), .A(net_3614) );
XNOR2_X2 inst_80 ( .ZN(net_1650), .A(net_1649), .B(net_820) );
NAND2_X2 inst_3623 ( .ZN(net_1961), .A2(net_1960), .A1(net_1717) );
SDFF_X2 inst_836 ( .Q(net_6997), .D(net_6997), .SE(net_3899), .SI(net_3778), .CK(net_10647) );
AOI21_X2 inst_7698 ( .B1(net_6745), .ZN(net_4114), .B2(net_2581), .A(net_2365) );
OAI22_X2 inst_1556 ( .B2(net_3405), .A2(net_3360), .ZN(net_3349), .A1(net_3270), .B1(net_577) );
CLKBUF_X2 inst_9228 ( .A(net_9189), .Z(net_9190) );
CLKBUF_X2 inst_9521 ( .A(net_9374), .Z(net_9483) );
CLKBUF_X2 inst_8821 ( .A(net_8782), .Z(net_8783) );
DFF_X1 inst_6796 ( .D(net_3942), .CK(net_12307), .Q(x681) );
CLKBUF_X2 inst_10771 ( .A(net_10732), .Z(net_10733) );
DFF_X1 inst_6564 ( .QN(net_7623), .D(net_5201), .CK(net_13465) );
CLKBUF_X2 inst_11243 ( .A(net_8839), .Z(net_11205) );
CLKBUF_X2 inst_9562 ( .A(net_9523), .Z(net_9524) );
CLKBUF_X2 inst_12075 ( .A(net_12036), .Z(net_12037) );
SDFF_X2 inst_241 ( .Q(net_6353), .SI(net_6352), .D(net_3605), .SE(net_392), .CK(net_13944) );
NAND2_X1 inst_4409 ( .A2(net_3087), .ZN(net_2908), .A1(net_2809) );
INV_X4 inst_5120 ( .ZN(net_3159), .A(net_597) );
INV_X4 inst_4934 ( .ZN(net_1161), .A(net_759) );
CLKBUF_X2 inst_14410 ( .A(net_14371), .Z(net_14372) );
SDFF_X2 inst_862 ( .SI(net_7029), .Q(net_7029), .SE(net_3818), .D(net_3806), .CK(net_11873) );
NAND2_X1 inst_4358 ( .ZN(net_4369), .A2(net_3853), .A1(net_2058) );
NAND2_X1 inst_4390 ( .ZN(net_4337), .A2(net_3859), .A1(net_1999) );
DFF_X1 inst_6690 ( .QN(net_7279), .D(net_5114), .CK(net_9449) );
CLKBUF_X2 inst_14142 ( .A(net_14103), .Z(net_14104) );
CLKBUF_X2 inst_13491 ( .A(net_13452), .Z(net_13453) );
NAND2_X2 inst_3918 ( .A1(net_7457), .A2(net_1696), .ZN(net_1385) );
NAND3_X2 inst_2758 ( .ZN(net_2343), .A3(net_1622), .A1(net_1430), .A2(net_1020) );
SDFF_X2 inst_1116 ( .SI(net_6655), .Q(net_6655), .D(net_3792), .SE(net_3465), .CK(net_9693) );
INV_X8 inst_4504 ( .ZN(net_3887), .A(net_3261) );
CLKBUF_X2 inst_7947 ( .A(net_7908), .Z(net_7909) );
CLKBUF_X2 inst_10620 ( .A(net_10581), .Z(net_10582) );
NAND2_X2 inst_3753 ( .A1(net_6630), .A2(net_1624), .ZN(net_1592) );
INV_X4 inst_5545 ( .ZN(net_523), .A(net_271) );
OAI21_X2 inst_1764 ( .B1(net_5551), .ZN(net_5430), .A(net_4648), .B2(net_3993) );
CLKBUF_X2 inst_14024 ( .A(net_13985), .Z(net_13986) );
INV_X4 inst_5271 ( .A(net_847), .ZN(net_420) );
CLKBUF_X2 inst_12050 ( .A(net_10555), .Z(net_12012) );
INV_X4 inst_5323 ( .A(net_6061), .ZN(net_801) );
AOI222_X2 inst_7472 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2163), .A1(net_2162), .B1(net_2161), .C1(net_2160) );
CLKBUF_X2 inst_11555 ( .A(net_11516), .Z(net_11517) );
SDFF_X2 inst_1159 ( .SI(net_6793), .Q(net_6793), .D(net_3892), .SE(net_3722), .CK(net_8259) );
CLKBUF_X2 inst_8740 ( .A(net_8701), .Z(net_8702) );
CLKBUF_X2 inst_9550 ( .A(net_9511), .Z(net_9512) );
CLKBUF_X2 inst_8659 ( .A(net_8620), .Z(net_8621) );
SDFF_X2 inst_402 ( .SI(net_7345), .Q(net_7345), .D(net_4776), .SE(net_3856), .CK(net_12750) );
NAND2_X2 inst_3136 ( .ZN(net_4827), .A2(net_4153), .A1(net_2182) );
DFF_X1 inst_6394 ( .QN(net_6113), .D(net_5694), .CK(net_11183) );
CLKBUF_X2 inst_10962 ( .A(net_9919), .Z(net_10924) );
CLKBUF_X2 inst_11259 ( .A(net_11220), .Z(net_11221) );
CLKBUF_X2 inst_9835 ( .A(net_9796), .Z(net_9797) );
CLKBUF_X2 inst_13025 ( .A(net_11267), .Z(net_12987) );
SDFF_X2 inst_938 ( .SI(net_7180), .Q(net_7180), .SE(net_3817), .D(net_3808), .CK(net_7846) );
INV_X2 inst_5832 ( .A(net_1302), .ZN(net_904) );
CLKBUF_X2 inst_12815 ( .A(net_11808), .Z(net_12777) );
CLKBUF_X2 inst_11189 ( .A(net_11150), .Z(net_11151) );
AOI22_X2 inst_7350 ( .B2(net_3105), .ZN(net_3100), .A2(net_2712), .A1(net_1121), .B1(net_696) );
CLKBUF_X2 inst_12552 ( .A(net_12513), .Z(net_12514) );
SDFF_X2 inst_1288 ( .D(net_7799), .SE(net_3256), .SI(net_136), .Q(net_136), .CK(net_8470) );
NAND2_X2 inst_3844 ( .A1(net_7103), .A2(net_1675), .ZN(net_1493) );
CLKBUF_X2 inst_12742 ( .A(net_12703), .Z(net_12704) );
DFF_X1 inst_6646 ( .QN(net_7620), .D(net_5207), .CK(net_13069) );
CLKBUF_X2 inst_9698 ( .A(net_8942), .Z(net_9660) );
AOI222_X1 inst_7610 ( .C1(net_5941), .B1(net_2970), .ZN(net_2873), .A1(net_2872), .B2(net_260), .C2(net_223), .A2(net_186) );
NAND2_X2 inst_3638 ( .ZN(net_1945), .A1(net_1288), .A2(net_1136) );
CLKBUF_X2 inst_8923 ( .A(net_8304), .Z(net_8885) );
NAND2_X1 inst_4365 ( .ZN(net_4362), .A2(net_3853), .A1(net_2000) );
CLKBUF_X2 inst_11329 ( .A(net_11290), .Z(net_11291) );
CLKBUF_X2 inst_9399 ( .A(net_9000), .Z(net_9361) );
CLKBUF_X2 inst_11845 ( .A(net_11806), .Z(net_11807) );
SDFF_X2 inst_1033 ( .Q(net_7549), .D(net_7549), .SE(net_3896), .SI(net_383), .CK(net_13111) );
CLKBUF_X2 inst_8957 ( .A(net_8918), .Z(net_8919) );
CLKBUF_X2 inst_11320 ( .A(net_10914), .Z(net_11282) );
INV_X4 inst_4673 ( .ZN(net_3469), .A(net_3468) );
CLKBUF_X2 inst_14253 ( .A(net_9834), .Z(net_14215) );
CLKBUF_X2 inst_14201 ( .A(net_11837), .Z(net_14163) );
INV_X4 inst_5582 ( .ZN(net_3208), .A(net_303) );
SDFFR_X2 inst_1348 ( .D(net_3808), .SE(net_3256), .SI(net_147), .Q(net_147), .CK(net_10401), .RN(x1822) );
AOI22_X2 inst_7426 ( .A1(net_2970), .B1(net_2772), .ZN(net_2766), .A2(net_242), .B2(net_168) );
OAI21_X2 inst_2102 ( .ZN(net_3980), .A(net_3979), .B2(net_3878), .B1(net_1054) );
INV_X4 inst_5427 ( .A(net_7556), .ZN(net_1979) );
CLKBUF_X2 inst_14070 ( .A(net_13292), .Z(net_14032) );
CLKBUF_X2 inst_9762 ( .A(net_9723), .Z(net_9724) );
OAI21_X2 inst_1748 ( .ZN(net_5519), .A(net_4819), .B2(net_4153), .B1(net_1065) );
INV_X4 inst_4908 ( .A(net_3897), .ZN(net_3174) );
AOI21_X4 inst_7619 ( .B2(net_5947), .B1(net_5946), .ZN(net_5609), .A(x1034) );
CLKBUF_X2 inst_11423 ( .A(net_11384), .Z(net_11385) );
AOI22_X2 inst_7356 ( .B2(net_3105), .ZN(net_3094), .B1(net_3093), .A2(net_2712), .A1(net_1123) );
CLKBUF_X2 inst_10343 ( .A(net_10304), .Z(net_10305) );
HA_X1 inst_6168 ( .B(net_6419), .S(net_898), .CO(net_897), .A(net_896) );
CLKBUF_X2 inst_8445 ( .A(net_7950), .Z(net_8407) );
INV_X4 inst_5565 ( .A(net_6156), .ZN(net_3609) );
CLKBUF_X2 inst_11684 ( .A(net_8091), .Z(net_11646) );
CLKBUF_X2 inst_11864 ( .A(net_11825), .Z(net_11826) );
CLKBUF_X2 inst_14058 ( .A(net_13632), .Z(net_14020) );
CLKBUF_X2 inst_11182 ( .A(net_11143), .Z(net_11144) );
CLKBUF_X2 inst_10145 ( .A(net_10106), .Z(net_10107) );
CLKBUF_X2 inst_9712 ( .A(net_9500), .Z(net_9674) );
CLKBUF_X2 inst_8637 ( .A(net_8598), .Z(net_8599) );
CLKBUF_X2 inst_9216 ( .A(net_9177), .Z(net_9178) );
SDFF_X2 inst_784 ( .SI(net_6894), .Q(net_6894), .SE(net_3887), .D(net_3806), .CK(net_8926) );
NAND2_X2 inst_3237 ( .ZN(net_4277), .A1(net_4276), .A2(net_1637) );
CLKBUF_X2 inst_11088 ( .A(net_11049), .Z(net_11050) );
SDFF_X2 inst_1264 ( .D(net_6389), .SE(net_6052), .SI(net_314), .Q(net_314), .CK(net_13808) );
CLKBUF_X2 inst_12046 ( .A(net_12007), .Z(net_12008) );
SDFF_X2 inst_690 ( .Q(net_6728), .D(net_6728), .SE(net_3815), .SI(net_3802), .CK(net_8965) );
DFF_X1 inst_6397 ( .QN(net_6136), .D(net_5691), .CK(net_8180) );
CLKBUF_X2 inst_11895 ( .A(net_11856), .Z(net_11857) );
OAI21_X2 inst_2025 ( .B1(net_5907), .B2(net_4497), .ZN(net_4481), .A(net_3628) );
AOI22_X2 inst_7337 ( .B2(net_3439), .ZN(net_3305), .B1(net_3080), .A2(net_2712), .A1(net_147) );
NOR2_X2 inst_2461 ( .A2(net_6184), .ZN(net_2915), .A1(net_769) );
AND2_X4 inst_7819 ( .ZN(net_3261), .A2(net_3164), .A1(net_525) );
CLKBUF_X2 inst_10607 ( .A(net_9160), .Z(net_10569) );
CLKBUF_X2 inst_8814 ( .A(net_8775), .Z(net_8776) );
SDFF_X2 inst_732 ( .Q(net_6830), .D(net_6830), .SE(net_3893), .SI(net_3806), .CK(net_8949) );
INV_X4 inst_4717 ( .ZN(net_3028), .A(net_2871) );
CLKBUF_X2 inst_12722 ( .A(net_10560), .Z(net_12684) );
CLKBUF_X2 inst_13044 ( .A(net_10670), .Z(net_13006) );
CLKBUF_X2 inst_12183 ( .A(net_12144), .Z(net_12145) );
CLKBUF_X2 inst_10969 ( .A(net_10930), .Z(net_10931) );
CLKBUF_X2 inst_9666 ( .A(net_9627), .Z(net_9628) );
CLKBUF_X2 inst_8023 ( .A(net_7831), .Z(net_7985) );
XNOR2_X2 inst_75 ( .ZN(net_1940), .B(net_674), .A(net_632) );
INV_X2 inst_5968 ( .A(net_7289), .ZN(net_1995) );
AOI21_X2 inst_7714 ( .B1(net_6730), .ZN(net_5904), .B2(net_2581), .A(net_2340) );
DFF_X1 inst_6386 ( .QN(net_6117), .D(net_5702), .CK(net_11204) );
XNOR2_X2 inst_79 ( .ZN(net_1653), .A(net_1652), .B(net_835) );
CLKBUF_X2 inst_11250 ( .A(net_11211), .Z(net_11212) );
CLKBUF_X2 inst_8930 ( .A(net_8891), .Z(net_8892) );
CLKBUF_X2 inst_7986 ( .A(net_7947), .Z(net_7948) );
NAND3_X2 inst_2654 ( .ZN(net_3946), .A3(net_3379), .A2(net_2935), .A1(net_2832) );
DFFR_X2 inst_7088 ( .QN(net_7723), .D(net_2795), .CK(net_10338), .RN(x1822) );
CLKBUF_X2 inst_9286 ( .A(net_9247), .Z(net_9248) );
AOI222_X2 inst_7600 ( .A1(net_7541), .ZN(net_5204), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_373), .C2(net_371) );
CLKBUF_X2 inst_11662 ( .A(net_11623), .Z(net_11624) );
CLKBUF_X2 inst_7891 ( .A(net_7832), .Z(net_7853) );
CLKBUF_X2 inst_12082 ( .A(net_12043), .Z(net_12044) );
CLKBUF_X2 inst_11962 ( .A(net_8011), .Z(net_11924) );
CLKBUF_X2 inst_8838 ( .A(net_8799), .Z(net_8800) );
CLKBUF_X2 inst_7895 ( .A(net_7856), .Z(net_7857) );
CLKBUF_X2 inst_13938 ( .A(net_11447), .Z(net_13900) );
CLKBUF_X2 inst_10890 ( .A(net_10851), .Z(net_10852) );
NAND2_X1 inst_4413 ( .A2(net_5974), .A1(net_5973), .ZN(net_2879) );
OAI21_X2 inst_1741 ( .ZN(net_5534), .A(net_4826), .B2(net_4153), .B1(net_1176) );
NAND2_X2 inst_2975 ( .A1(net_7160), .ZN(net_5038), .A2(net_4954) );
CLKBUF_X2 inst_10339 ( .A(net_8478), .Z(net_10301) );
SDFF_X2 inst_1024 ( .SI(net_6519), .Q(net_6519), .SE(net_3889), .D(net_3800), .CK(net_11638) );
INV_X2 inst_5827 ( .ZN(net_926), .A(net_925) );
INV_X4 inst_5594 ( .A(net_7252), .ZN(net_2021) );
CLKBUF_X2 inst_12144 ( .A(net_9272), .Z(net_12106) );
NOR2_X4 inst_2232 ( .ZN(net_5666), .A1(net_5525), .A2(net_4494) );
INV_X8 inst_4546 ( .ZN(net_1696), .A(net_919) );
CLKBUF_X2 inst_13218 ( .A(net_13179), .Z(net_13180) );
OAI221_X2 inst_1658 ( .ZN(net_4795), .A(net_4551), .C2(net_3971), .B2(net_3960), .C1(net_3761), .B1(net_1401) );
DFF_X1 inst_6515 ( .QN(net_7446), .D(net_5441), .CK(net_9292) );
CLKBUF_X2 inst_12061 ( .A(net_12022), .Z(net_12023) );
OAI21_X2 inst_1689 ( .B1(net_5778), .ZN(net_5775), .A(net_5707), .B2(net_5706) );
CLKBUF_X2 inst_9003 ( .A(net_8964), .Z(net_8965) );
NAND2_X4 inst_2846 ( .ZN(net_5477), .A1(net_4924), .A2(net_4923) );
NAND2_X2 inst_3965 ( .A1(net_6577), .A2(net_1705), .ZN(net_1317) );
NAND2_X1 inst_4267 ( .ZN(net_4652), .A2(net_3993), .A1(net_1452) );
CLKBUF_X2 inst_8279 ( .A(net_8240), .Z(net_8241) );
NAND2_X2 inst_3584 ( .ZN(net_2420), .A1(net_2419), .A2(net_2418) );
CLKBUF_X2 inst_11408 ( .A(net_11369), .Z(net_11370) );
CLKBUF_X2 inst_9472 ( .A(net_9433), .Z(net_9434) );
OAI22_X2 inst_1448 ( .B2(net_5911), .B1(net_4644), .ZN(net_4626), .A2(net_4610), .A1(net_4039) );
CLKBUF_X2 inst_12829 ( .A(net_12790), .Z(net_12791) );
CLKBUF_X2 inst_8395 ( .A(net_8136), .Z(net_8357) );
OAI21_X2 inst_1816 ( .ZN(net_5372), .B1(net_5345), .A(net_4339), .B2(net_3859) );
SDFF_X2 inst_440 ( .Q(net_7394), .D(net_7394), .SE(net_3994), .SI(net_359), .CK(net_9632) );
CLKBUF_X2 inst_11892 ( .A(net_11853), .Z(net_11854) );
CLKBUF_X2 inst_11723 ( .A(net_10325), .Z(net_11685) );
CLKBUF_X2 inst_14386 ( .A(net_11551), .Z(net_14348) );
INV_X4 inst_5012 ( .A(net_7811), .ZN(net_3831) );
INV_X4 inst_4927 ( .ZN(net_815), .A(net_814) );
NAND2_X2 inst_3381 ( .ZN(net_3484), .A1(net_3483), .A2(net_3223) );
CLKBUF_X2 inst_14123 ( .A(net_14084), .Z(net_14085) );
OAI21_X2 inst_1887 ( .B1(net_5237), .ZN(net_5194), .A(net_4570), .B2(net_3866) );
SDFF_X2 inst_1091 ( .SI(net_6933), .Q(net_6933), .D(net_3814), .SE(net_3734), .CK(net_11781) );
CLKBUF_X2 inst_11708 ( .A(net_11669), .Z(net_11670) );
CLKBUF_X2 inst_9915 ( .A(net_9876), .Z(net_9877) );
INV_X4 inst_4837 ( .ZN(net_4874), .A(net_1073) );
INV_X4 inst_5059 ( .ZN(net_739), .A(net_638) );
CLKBUF_X2 inst_8206 ( .A(net_8003), .Z(net_8168) );
CLKBUF_X2 inst_10450 ( .A(net_9052), .Z(net_10412) );
NAND2_X2 inst_3579 ( .ZN(net_2434), .A2(net_2433), .A1(net_733) );
CLKBUF_X2 inst_13800 ( .A(net_13761), .Z(net_13762) );
NAND2_X2 inst_4154 ( .A2(net_1228), .ZN(net_1067), .A1(net_376) );
CLKBUF_X2 inst_10374 ( .A(net_10335), .Z(net_10336) );
INV_X4 inst_5688 ( .A(net_7407), .ZN(net_2111) );
INV_X4 inst_5398 ( .A(net_6044), .ZN(net_578) );
OAI221_X2 inst_1672 ( .ZN(net_4171), .B2(net_4107), .C2(net_4007), .A(net_3950), .B1(net_735), .C1(net_734) );
INV_X4 inst_4816 ( .ZN(net_4783), .A(net_1141) );
CLKBUF_X2 inst_13705 ( .A(net_10589), .Z(net_13667) );
CLKBUF_X2 inst_12120 ( .A(net_12081), .Z(net_12082) );
CLKBUF_X2 inst_8625 ( .A(net_8427), .Z(net_8587) );
OAI21_X2 inst_2015 ( .B2(net_4497), .ZN(net_4493), .B1(net_4104), .A(net_3656) );
CLKBUF_X2 inst_12108 ( .A(net_12069), .Z(net_12070) );
NAND2_X2 inst_3179 ( .ZN(net_4754), .A2(net_3941), .A1(net_2158) );
NAND2_X2 inst_3059 ( .A1(net_7124), .A2(net_4950), .ZN(net_4946) );
NAND2_X2 inst_3937 ( .A1(net_6982), .A2(net_1833), .ZN(net_1356) );
NAND2_X2 inst_2970 ( .ZN(net_5457), .A1(net_4880), .A2(net_4879) );
CLKBUF_X2 inst_11357 ( .A(net_11318), .Z(net_11319) );
CLKBUF_X2 inst_11950 ( .A(net_8322), .Z(net_11912) );
CLKBUF_X2 inst_10942 ( .A(net_10903), .Z(net_10904) );
CLKBUF_X2 inst_9281 ( .A(net_9242), .Z(net_9243) );
CLKBUF_X2 inst_8278 ( .A(net_8239), .Z(net_8240) );
NAND2_X2 inst_4085 ( .A1(net_6532), .A2(net_1645), .ZN(net_967) );
CLKBUF_X2 inst_9390 ( .A(net_9061), .Z(net_9352) );
CLKBUF_X2 inst_13183 ( .A(net_13144), .Z(net_13145) );
NAND3_X2 inst_2587 ( .ZN(net_5752), .A1(net_5647), .A2(net_5265), .A3(net_4307) );
INV_X4 inst_4990 ( .A(net_7816), .ZN(net_3803) );
INV_X4 inst_5664 ( .A(net_6059), .ZN(net_1679) );
CLKBUF_X2 inst_10317 ( .A(net_9109), .Z(net_10279) );
CLKBUF_X2 inst_12285 ( .A(net_12246), .Z(net_12247) );
DFF_X1 inst_6680 ( .QN(net_7258), .D(net_5144), .CK(net_12721) );
CLKBUF_X2 inst_8868 ( .A(net_8829), .Z(net_8830) );
CLKBUF_X2 inst_9442 ( .A(net_9202), .Z(net_9404) );
CLKBUF_X2 inst_11090 ( .A(net_11051), .Z(net_11052) );
CLKBUF_X2 inst_13072 ( .A(net_13033), .Z(net_13034) );
SDFF_X2 inst_815 ( .Q(net_6990), .D(net_6990), .SE(net_3891), .SI(net_3795), .CK(net_11022) );
CLKBUF_X2 inst_8883 ( .A(net_8844), .Z(net_8845) );
NAND2_X2 inst_3031 ( .A1(net_7020), .A2(net_4979), .ZN(net_4976) );
OAI211_X2 inst_2165 ( .B(net_2724), .ZN(net_2723), .C1(net_2382), .A(net_939), .C2(net_938) );
SDFF_X2 inst_1257 ( .D(net_7799), .SI(net_6526), .Q(net_6526), .SE(net_3755), .CK(net_8607) );
SDFF_X2 inst_875 ( .SI(net_7033), .Q(net_7033), .SE(net_3818), .D(net_3798), .CK(net_9012) );
NAND2_X2 inst_3298 ( .ZN(net_3650), .A1(net_3649), .A2(net_3229) );
NAND2_X2 inst_3081 ( .ZN(net_4922), .A2(net_4328), .A1(net_2250) );
NAND2_X2 inst_3482 ( .ZN(net_2674), .A1(net_2673), .A2(net_2672) );
CLKBUF_X2 inst_12096 ( .A(net_12057), .Z(net_12058) );
INV_X4 inst_5075 ( .A(net_1140), .ZN(net_720) );
INV_X4 inst_5187 ( .ZN(net_3230), .A(net_516) );
OAI21_X2 inst_2069 ( .B2(net_4436), .ZN(net_4425), .B1(net_4424), .A(net_3622) );
CLKBUF_X2 inst_8227 ( .A(net_8188), .Z(net_8189) );
CLKBUF_X2 inst_8888 ( .A(net_8849), .Z(net_8850) );
DFFR_X2 inst_7006 ( .QN(net_7700), .D(net_3342), .CK(net_10357), .RN(x1822) );
OAI21_X2 inst_2108 ( .ZN(net_3863), .B1(net_3862), .B2(net_3861), .A(net_3732) );
NAND2_X2 inst_3572 ( .ZN(net_2495), .A2(net_1988), .A1(net_1185) );
NAND2_X2 inst_4098 ( .A1(net_7195), .A2(net_1648), .ZN(net_954) );
CLKBUF_X2 inst_12178 ( .A(net_12139), .Z(net_12140) );
CLKBUF_X2 inst_11220 ( .A(net_11181), .Z(net_11182) );
INV_X4 inst_5703 ( .A(net_5943), .ZN(net_5939) );
AOI21_X2 inst_7761 ( .B1(net_7148), .ZN(net_4066), .B2(net_2582), .A(net_2286) );
CLKBUF_X2 inst_11177 ( .A(net_11138), .Z(net_11139) );
NAND2_X2 inst_2978 ( .A1(net_6716), .ZN(net_5035), .A2(net_5031) );
SDFF_X2 inst_413 ( .D(net_6392), .SE(net_6050), .SI(net_301), .Q(net_301), .CK(net_14214) );
CLKBUF_X2 inst_14239 ( .A(net_12796), .Z(net_14201) );
CLKBUF_X2 inst_11033 ( .A(net_8065), .Z(net_10995) );
INV_X4 inst_5094 ( .A(net_7818), .ZN(net_3898) );
CLKBUF_X2 inst_11393 ( .A(net_11354), .Z(net_11355) );
SDFF_X2 inst_859 ( .SI(net_7044), .Q(net_7044), .SE(net_3818), .D(net_3785), .CK(net_11883) );
DFF_X1 inst_6623 ( .QN(net_7584), .D(net_5264), .CK(net_12269) );
CLKBUF_X2 inst_8118 ( .A(net_8072), .Z(net_8080) );
CLKBUF_X2 inst_10269 ( .A(net_10183), .Z(net_10231) );
CLKBUF_X2 inst_13446 ( .A(net_13407), .Z(net_13408) );
CLKBUF_X2 inst_14352 ( .A(net_14313), .Z(net_14314) );
CLKBUF_X2 inst_12634 ( .A(net_12595), .Z(net_12596) );
NAND2_X2 inst_3323 ( .ZN(net_3600), .A1(net_3599), .A2(net_3228) );
CLKBUF_X2 inst_13013 ( .A(net_12974), .Z(net_12975) );
OAI21_X2 inst_2019 ( .B2(net_4497), .ZN(net_4489), .B1(net_4095), .A(net_3646) );
CLKBUF_X2 inst_13679 ( .A(net_12320), .Z(net_13641) );
CLKBUF_X2 inst_8323 ( .A(net_7941), .Z(net_8285) );
INV_X4 inst_5186 ( .ZN(net_3917), .A(net_802) );
INV_X2 inst_5938 ( .A(net_7362), .ZN(net_2074) );
CLKBUF_X2 inst_13061 ( .A(net_10897), .Z(net_13023) );
XNOR2_X2 inst_69 ( .ZN(net_2478), .A(net_1060), .B(net_540) );
INV_X2 inst_5736 ( .ZN(net_5880), .A(net_4137) );
CLKBUF_X2 inst_14448 ( .A(net_14035), .Z(net_14410) );
OAI21_X2 inst_1691 ( .B2(net_5905), .ZN(net_5603), .A(net_5305), .B1(net_4132) );
NAND3_X2 inst_2669 ( .ZN(net_3959), .A2(net_3874), .A3(net_3736), .A1(net_2237) );
CLKBUF_X2 inst_9019 ( .A(net_8980), .Z(net_8981) );
CLKBUF_X2 inst_12844 ( .A(net_12650), .Z(net_12806) );
CLKBUF_X2 inst_11156 ( .A(net_11117), .Z(net_11118) );
SDFF_X2 inst_844 ( .Q(net_7025), .D(net_7025), .SE(net_3899), .SI(net_3821), .CK(net_10994) );
NOR2_X2 inst_2489 ( .ZN(net_2415), .A1(net_2414), .A2(net_2226) );
DFFR_X2 inst_6968 ( .QN(net_5993), .D(net_4006), .CK(net_10374), .RN(x1822) );
NAND2_X2 inst_3619 ( .ZN(net_1970), .A2(net_1969), .A1(net_1723) );
NAND2_X2 inst_3688 ( .A2(net_1798), .ZN(net_1758), .A1(net_1757) );
DFF_X1 inst_6709 ( .QN(net_7325), .D(net_5362), .CK(net_10157) );
INV_X2 inst_5805 ( .ZN(net_1702), .A(net_1701) );
AOI21_X2 inst_7716 ( .B1(net_6863), .ZN(net_5896), .B2(net_2579), .A(net_2344) );
DFF_X1 inst_6939 ( .D(net_2411), .Q(net_240), .CK(net_13034) );
INV_X4 inst_4641 ( .ZN(net_4181), .A(net_4021) );
DFFR_X2 inst_7056 ( .QN(net_5990), .D(net_3145), .CK(net_9609), .RN(x1822) );
CLKBUF_X2 inst_11038 ( .A(net_10999), .Z(net_11000) );
INV_X4 inst_5476 ( .ZN(net_431), .A(net_299) );
SDFF_X2 inst_460 ( .SI(net_7807), .Q(net_6470), .D(net_6470), .SE(net_3904), .CK(net_11272) );
CLKBUF_X2 inst_10877 ( .A(net_7850), .Z(net_10839) );
OAI22_X2 inst_1455 ( .B2(net_5908), .B1(net_4650), .A2(net_4614), .ZN(net_4613), .A1(net_4035) );
INV_X2 inst_5776 ( .ZN(net_2790), .A(net_2716) );
CLKBUF_X2 inst_12149 ( .A(net_9781), .Z(net_12111) );
NOR2_X2 inst_2497 ( .ZN(net_1744), .A2(net_1743), .A1(net_1093) );
CLKBUF_X2 inst_13124 ( .A(net_9018), .Z(net_13086) );
CLKBUF_X2 inst_10186 ( .A(net_8347), .Z(net_10148) );
NAND2_X2 inst_3660 ( .A1(net_7075), .ZN(net_1803), .A2(net_791) );
CLKBUF_X2 inst_11167 ( .A(net_10442), .Z(net_11129) );
SDFF_X2 inst_560 ( .SI(net_7166), .Q(net_7166), .D(net_3892), .SE(net_3817), .CK(net_13374) );
INV_X4 inst_5393 ( .A(net_7425), .ZN(net_2150) );
CLKBUF_X2 inst_9729 ( .A(net_9690), .Z(net_9691) );
NAND2_X1 inst_4230 ( .ZN(net_4697), .A2(net_3989), .A1(net_2177) );
INV_X4 inst_5199 ( .A(net_652), .ZN(net_501) );
CLKBUF_X2 inst_12953 ( .A(net_10990), .Z(net_12915) );
AOI222_X2 inst_7479 ( .C1(net_7522), .B1(net_7490), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2145), .A1(net_2144) );
INV_X4 inst_4809 ( .ZN(net_4784), .A(net_1169) );
INV_X4 inst_5571 ( .A(net_6102), .ZN(net_3499) );
CLKBUF_X2 inst_13455 ( .A(net_13416), .Z(net_13417) );
OAI21_X2 inst_1802 ( .ZN(net_5388), .A(net_4715), .B2(net_3986), .B1(net_1174) );
SDFF_X2 inst_950 ( .SI(net_7193), .Q(net_7193), .SE(net_3817), .D(net_3801), .CK(net_10627) );
CLKBUF_X2 inst_10260 ( .A(net_9861), .Z(net_10222) );
DFF_X1 inst_6851 ( .D(net_2554), .Q(net_216), .CK(net_9810) );
NAND2_X2 inst_2982 ( .A1(net_6718), .A2(net_5031), .ZN(net_5029) );
NAND2_X2 inst_3955 ( .A1(net_7107), .A2(net_1675), .ZN(net_1330) );
CLKBUF_X2 inst_11837 ( .A(net_10852), .Z(net_11799) );
CLKBUF_X2 inst_10100 ( .A(net_10061), .Z(net_10062) );
SDFF_X2 inst_1218 ( .D(net_7807), .SI(net_7209), .Q(net_7209), .SE(net_3750), .CK(net_12128) );
NAND2_X2 inst_3359 ( .ZN(net_3527), .A2(net_3225), .A1(net_3125) );
CLKBUF_X2 inst_8458 ( .A(net_8419), .Z(net_8420) );
DFF_X1 inst_6414 ( .QN(net_6161), .D(net_5756), .CK(net_11046) );
AOI222_X2 inst_7491 ( .A2(net_2135), .B2(net_2133), .C2(net_2131), .ZN(net_2102), .A1(net_2101), .B1(net_2100), .C1(net_2099) );
CLKBUF_X2 inst_14338 ( .A(net_8880), .Z(net_14300) );
NAND2_X1 inst_4418 ( .ZN(net_2739), .A2(net_229), .A1(net_228) );
CLKBUF_X2 inst_9541 ( .A(net_9502), .Z(net_9503) );
XNOR2_X2 inst_96 ( .B(net_3000), .ZN(net_1658), .A(net_1149) );
XNOR2_X2 inst_101 ( .ZN(net_2250), .A(net_1149), .B(net_1143) );
NAND2_X1 inst_4346 ( .ZN(net_4381), .A2(net_3856), .A1(net_1757) );
CLKBUF_X2 inst_8564 ( .A(net_8525), .Z(net_8526) );
CLKBUF_X2 inst_14033 ( .A(net_10812), .Z(net_13995) );
NAND2_X2 inst_3555 ( .ZN(net_2512), .A2(net_2036), .A1(net_1753) );
CLKBUF_X2 inst_11205 ( .A(net_11166), .Z(net_11167) );
CLKBUF_X2 inst_10234 ( .A(net_10195), .Z(net_10196) );
CLKBUF_X2 inst_14377 ( .A(net_14338), .Z(net_14339) );
CLKBUF_X2 inst_9330 ( .A(net_9291), .Z(net_9292) );
CLKBUF_X2 inst_11388 ( .A(net_11349), .Z(net_11350) );
INV_X4 inst_4722 ( .ZN(net_3018), .A(net_2863) );
SDFF_X2 inst_510 ( .Q(net_6712), .D(net_6712), .SI(net_3897), .SE(net_3871), .CK(net_11360) );
CLKBUF_X2 inst_10912 ( .A(net_10726), .Z(net_10874) );
CLKBUF_X2 inst_12194 ( .A(net_11455), .Z(net_12156) );
NOR2_X2 inst_2436 ( .ZN(net_3431), .A1(net_3048), .A2(net_3047) );
DFF_X1 inst_6505 ( .QN(net_7427), .D(net_5521), .CK(net_9815) );
OAI221_X2 inst_1677 ( .C1(net_5940), .ZN(net_3938), .B2(net_3937), .A(net_3730), .B1(net_3053), .C2(net_193) );
NAND2_X4 inst_2832 ( .ZN(net_5563), .A1(net_5036), .A2(net_5035) );
SDFF_X2 inst_830 ( .Q(net_7009), .D(net_7009), .SE(net_3899), .SI(net_3811), .CK(net_11009) );
SDFF_X2 inst_603 ( .Q(net_6607), .D(net_6607), .SE(net_3830), .SI(net_3809), .CK(net_7883) );
CLKBUF_X2 inst_8433 ( .A(net_8394), .Z(net_8395) );
SDFF_X2 inst_291 ( .D(net_6395), .SE(net_5801), .SI(net_340), .Q(net_340), .CK(net_14326) );
NAND2_X4 inst_2878 ( .A1(net_5884), .ZN(net_4261), .A2(net_2583) );
NOR2_X2 inst_2494 ( .ZN(net_2417), .A2(net_1921), .A1(net_1920) );
SDFF_X2 inst_776 ( .SI(net_6904), .Q(net_6904), .D(net_3813), .SE(net_3781), .CK(net_11465) );
CLKBUF_X2 inst_9488 ( .A(net_8818), .Z(net_9450) );
NOR2_X2 inst_2526 ( .ZN(net_1649), .A2(net_770), .A1(net_448) );
INV_X4 inst_5047 ( .ZN(net_766), .A(net_646) );
CLKBUF_X2 inst_12213 ( .A(net_12174), .Z(net_12175) );
CLKBUF_X2 inst_10787 ( .A(net_10748), .Z(net_10749) );
INV_X4 inst_5313 ( .A(net_7402), .ZN(net_2182) );
OAI21_X2 inst_1972 ( .B1(net_4870), .ZN(net_4864), .A(net_4386), .B2(net_3856) );
SDFF_X2 inst_558 ( .SI(net_7053), .Q(net_7053), .D(net_3898), .SE(net_3818), .CK(net_11031) );
HA_X1 inst_6167 ( .A(net_1700), .S(net_1273), .CO(net_1272), .B(net_614) );
CLKBUF_X2 inst_12704 ( .A(net_12665), .Z(net_12666) );
CLKBUF_X2 inst_10310 ( .A(net_8819), .Z(net_10272) );
DFF_X1 inst_6849 ( .D(net_2555), .QN(net_215), .CK(net_9539) );
CLKBUF_X2 inst_9110 ( .A(net_8379), .Z(net_9072) );
CLKBUF_X2 inst_10591 ( .A(net_9676), .Z(net_10553) );
SDFF_X2 inst_389 ( .SI(net_7309), .Q(net_7309), .D(net_4778), .SE(net_3859), .CK(net_9919) );
INV_X4 inst_5179 ( .ZN(net_526), .A(net_525) );
DFF_X1 inst_6512 ( .QN(net_7443), .D(net_5447), .CK(net_10094) );
CLKBUF_X2 inst_14301 ( .A(net_8420), .Z(net_14263) );
CLKBUF_X2 inst_13460 ( .A(net_13421), .Z(net_13422) );
NAND3_X2 inst_2712 ( .ZN(net_2465), .A2(net_1806), .A3(net_1572), .A1(net_1424) );
CLKBUF_X2 inst_10252 ( .A(net_10213), .Z(net_10214) );
INV_X1 inst_6152 ( .ZN(net_3025), .A(net_3024) );
DFF_X1 inst_6925 ( .D(net_2410), .Q(net_244), .CK(net_13039) );
CLKBUF_X2 inst_8650 ( .A(net_8351), .Z(net_8612) );
AOI21_X2 inst_7745 ( .B1(net_6470), .ZN(net_4049), .B2(net_2580), .A(net_2333) );
OR2_X4 inst_1382 ( .ZN(net_2903), .A2(net_2753), .A1(net_278) );
CLKBUF_X2 inst_8841 ( .A(net_8802), .Z(net_8803) );
CLKBUF_X2 inst_8600 ( .A(net_8561), .Z(net_8562) );
OAI21_X2 inst_1807 ( .ZN(net_5381), .B1(net_5363), .A(net_4351), .B2(net_3859) );
NAND3_X2 inst_2795 ( .ZN(net_2305), .A3(net_1600), .A1(net_1350), .A2(net_968) );
CLKBUF_X2 inst_9989 ( .A(net_9950), .Z(net_9951) );
CLKBUF_X2 inst_12274 ( .A(net_12235), .Z(net_12236) );
SDFF_X2 inst_913 ( .Q(net_7150), .D(net_7150), .SE(net_3903), .SI(net_3807), .CK(net_13357) );
INV_X4 inst_5266 ( .A(net_859), .ZN(net_424) );
CLKBUF_X2 inst_12712 ( .A(net_12673), .Z(net_12674) );
INV_X4 inst_4766 ( .ZN(net_2429), .A(net_1935) );
NAND2_X1 inst_4445 ( .ZN(net_1262), .A1(net_1261), .A2(net_1256) );
INV_X2 inst_5895 ( .A(net_7283), .ZN(net_2037) );
CLKBUF_X2 inst_11785 ( .A(net_11638), .Z(net_11747) );
CLKBUF_X2 inst_9977 ( .A(net_9726), .Z(net_9939) );
CLKBUF_X2 inst_12866 ( .A(net_12827), .Z(net_12828) );
CLKBUF_X2 inst_12766 ( .A(net_12727), .Z(net_12728) );
CLKBUF_X2 inst_8365 ( .A(net_8326), .Z(net_8327) );
CLKBUF_X2 inst_14195 ( .A(net_9157), .Z(net_14157) );
DFFR_X2 inst_7105 ( .D(net_1958), .QN(net_114), .CK(net_9586), .RN(x1822) );
CLKBUF_X2 inst_10843 ( .A(net_10804), .Z(net_10805) );
CLKBUF_X2 inst_11613 ( .A(net_11574), .Z(net_11575) );
AOI21_X2 inst_7687 ( .B1(net_7131), .ZN(net_4447), .B2(net_2582), .A(net_2327) );
DFF_X1 inst_6633 ( .QN(net_7589), .D(net_5249), .CK(net_13160) );
CLKBUF_X2 inst_12004 ( .A(net_11965), .Z(net_11966) );
CLKBUF_X2 inst_11133 ( .A(net_11094), .Z(net_11095) );
CLKBUF_X2 inst_10322 ( .A(net_10283), .Z(net_10284) );
CLKBUF_X2 inst_11724 ( .A(net_10088), .Z(net_11686) );
CLKBUF_X2 inst_11214 ( .A(net_10175), .Z(net_11176) );
CLKBUF_X2 inst_9298 ( .A(net_9259), .Z(net_9260) );
NOR2_X2 inst_2483 ( .A2(net_5778), .ZN(net_2654), .A1(net_2596) );
CLKBUF_X2 inst_13321 ( .A(net_13282), .Z(net_13283) );
CLKBUF_X2 inst_9446 ( .A(net_9099), .Z(net_9408) );
OR2_X2 inst_1414 ( .ZN(net_3758), .A2(net_792), .A1(net_548) );
AOI21_X4 inst_7624 ( .B1(net_6999), .ZN(net_4621), .A(net_2461), .B2(net_1100) );
CLKBUF_X2 inst_8451 ( .A(net_8267), .Z(net_8413) );
SDFF_X2 inst_449 ( .D(net_6390), .SE(net_5799), .SI(net_375), .Q(net_375), .CK(net_13892) );
NAND2_X2 inst_3994 ( .A2(net_1910), .ZN(net_1196), .A1(net_1195) );
CLKBUF_X2 inst_13467 ( .A(net_13428), .Z(net_13429) );
NAND2_X2 inst_4212 ( .ZN(net_483), .A1(x1286), .A2(x1261) );
CLKBUF_X2 inst_10797 ( .A(net_10758), .Z(net_10759) );
CLKBUF_X2 inst_10354 ( .A(net_8470), .Z(net_10316) );
NAND3_X2 inst_2790 ( .ZN(net_2310), .A3(net_1612), .A1(net_1499), .A2(net_1018) );
OAI21_X2 inst_2138 ( .ZN(net_2812), .A(net_557), .B1(net_227), .B2(net_225) );
INV_X4 inst_5599 ( .A(net_6144), .ZN(net_3615) );
CLKBUF_X2 inst_11417 ( .A(net_11378), .Z(net_11379) );
DFF_X1 inst_6593 ( .QN(net_7500), .D(net_5110), .CK(net_12476) );
INV_X2 inst_6055 ( .A(net_7655), .ZN(net_1871) );
CLKBUF_X2 inst_13362 ( .A(net_8674), .Z(net_13324) );
CLKBUF_X2 inst_11231 ( .A(net_11192), .Z(net_11193) );
NAND2_X2 inst_3249 ( .ZN(net_5087), .A2(net_3469), .A1(net_2965) );
INV_X4 inst_4935 ( .ZN(net_1179), .A(net_758) );
CLKBUF_X2 inst_12912 ( .A(net_9848), .Z(net_12874) );
CLKBUF_X2 inst_11759 ( .A(net_11720), .Z(net_11721) );
CLKBUF_X2 inst_9594 ( .A(net_8535), .Z(net_9556) );
CLKBUF_X2 inst_8961 ( .A(net_8063), .Z(net_8923) );
AOI222_X2 inst_7498 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2080), .A1(net_2079), .B1(net_2078), .C1(net_2077) );
NOR2_X2 inst_2309 ( .A2(net_6205), .A1(net_5840), .ZN(net_5832) );
CLKBUF_X2 inst_9860 ( .A(net_9821), .Z(net_9822) );
CLKBUF_X2 inst_13369 ( .A(net_8291), .Z(net_13331) );
CLKBUF_X2 inst_12420 ( .A(net_12381), .Z(net_12382) );
CLKBUF_X2 inst_11044 ( .A(net_11005), .Z(net_11006) );
CLKBUF_X2 inst_12973 ( .A(net_12934), .Z(net_12935) );
AOI21_X2 inst_7644 ( .B1(net_5914), .ZN(net_3908), .B2(net_3907), .A(net_2597) );
CLKBUF_X2 inst_8201 ( .A(net_8162), .Z(net_8163) );
CLKBUF_X2 inst_11283 ( .A(net_10771), .Z(net_11245) );
CLKBUF_X2 inst_8893 ( .A(net_8854), .Z(net_8855) );
NAND3_X2 inst_2603 ( .ZN(net_5736), .A1(net_5631), .A2(net_5176), .A3(net_4196) );
NAND2_X2 inst_3614 ( .ZN(net_2268), .A2(net_1933), .A1(net_1334) );
CLKBUF_X2 inst_11335 ( .A(net_9551), .Z(net_11297) );
INV_X4 inst_4603 ( .ZN(net_4241), .A(net_4100) );
CLKBUF_X2 inst_9339 ( .A(net_8097), .Z(net_9301) );
OAI21_X2 inst_2153 ( .B1(net_5778), .ZN(net_2791), .A(net_2665), .B2(net_2663) );
CLKBUF_X2 inst_12776 ( .A(net_12737), .Z(net_12738) );
CLKBUF_X2 inst_10752 ( .A(net_8652), .Z(net_10714) );
SDFF_X2 inst_588 ( .Q(net_6587), .D(net_6587), .SE(net_3823), .SI(net_3788), .CK(net_9119) );
CLKBUF_X2 inst_10394 ( .A(net_10355), .Z(net_10356) );
CLKBUF_X2 inst_11411 ( .A(net_11372), .Z(net_11373) );
CLKBUF_X2 inst_11271 ( .A(net_11232), .Z(net_11233) );
CLKBUF_X2 inst_11904 ( .A(net_11865), .Z(net_11866) );
CLKBUF_X2 inst_11798 ( .A(net_11759), .Z(net_11760) );
CLKBUF_X2 inst_14015 ( .A(net_13976), .Z(net_13977) );
CLKBUF_X2 inst_10329 ( .A(net_9958), .Z(net_10291) );
CLKBUF_X2 inst_9405 ( .A(net_8776), .Z(net_9367) );
INV_X4 inst_5494 ( .A(net_7569), .ZN(net_1845) );
CLKBUF_X2 inst_11060 ( .A(net_11021), .Z(net_11022) );
CLKBUF_X2 inst_10586 ( .A(net_10547), .Z(net_10548) );
INV_X4 inst_4752 ( .A(net_2718), .ZN(net_2706) );
AOI21_X2 inst_7674 ( .B1(net_7009), .ZN(net_4222), .A(net_2466), .B2(net_1100) );
CLKBUF_X2 inst_12913 ( .A(net_12874), .Z(net_12875) );
SDFFR_X2 inst_1356 ( .D(net_3807), .SE(net_3256), .SI(net_149), .Q(net_149), .CK(net_11403), .RN(x1822) );
INV_X4 inst_5441 ( .A(net_6113), .ZN(net_3669) );
CLKBUF_X2 inst_9906 ( .A(net_9867), .Z(net_9868) );
NAND3_X2 inst_2628 ( .ZN(net_5701), .A1(net_5678), .A2(net_5312), .A3(net_4252) );
DFF_X1 inst_6447 ( .QN(net_6098), .D(net_5723), .CK(net_12060) );
DFF_X1 inst_6874 ( .D(net_2550), .Q(net_194), .CK(net_9974) );
NOR3_X2 inst_2196 ( .ZN(net_3880), .A1(net_3381), .A3(net_1159), .A2(net_776) );
NAND2_X2 inst_3485 ( .ZN(net_2665), .A1(net_2664), .A2(net_2663) );
CLKBUF_X2 inst_14159 ( .A(net_14120), .Z(net_14121) );
INV_X2 inst_5854 ( .ZN(net_670), .A(net_669) );
AOI21_X2 inst_7754 ( .B1(net_6471), .ZN(net_4047), .B2(net_2580), .A(net_2281) );
CLKBUF_X2 inst_14083 ( .A(net_8225), .Z(net_14045) );
SDFF_X2 inst_1045 ( .Q(net_7245), .D(net_7245), .SE(net_3822), .SI(net_341), .CK(net_9832) );
SDFF_X2 inst_865 ( .SI(net_7051), .Q(net_7051), .SE(net_3818), .D(net_3780), .CK(net_11868) );
SDFF_X2 inst_252 ( .Q(net_6342), .SI(net_6341), .D(net_3591), .SE(net_392), .CK(net_13498) );
SDFF_X2 inst_956 ( .D(net_7802), .SI(net_7172), .Q(net_7172), .SE(net_3819), .CK(net_13326) );
CLKBUF_X2 inst_8587 ( .A(net_8548), .Z(net_8549) );
CLKBUF_X2 inst_10959 ( .A(net_10920), .Z(net_10921) );
CLKBUF_X2 inst_8680 ( .A(net_8611), .Z(net_8642) );
CLKBUF_X2 inst_10177 ( .A(net_7849), .Z(net_10139) );
INV_X4 inst_4684 ( .ZN(net_3739), .A(net_3367) );
CLKBUF_X2 inst_12757 ( .A(net_12718), .Z(net_12719) );
SDFF_X2 inst_484 ( .SI(net_6495), .Q(net_6495), .D(net_3890), .SE(net_3889), .CK(net_8801) );
CLKBUF_X2 inst_9272 ( .A(net_9233), .Z(net_9234) );
INV_X8 inst_4474 ( .ZN(net_5033), .A(net_4271) );
DFF_X1 inst_6678 ( .QN(net_7256), .D(net_5142), .CK(net_13004) );
CLKBUF_X2 inst_9129 ( .A(net_9090), .Z(net_9091) );
XNOR2_X2 inst_32 ( .ZN(net_2479), .A(net_2478), .B(net_910) );
OAI21_X2 inst_1821 ( .ZN(net_5367), .B1(net_5335), .A(net_4334), .B2(net_3859) );
CLKBUF_X2 inst_9616 ( .A(net_9577), .Z(net_9578) );
CLKBUF_X2 inst_12798 ( .A(net_12759), .Z(net_12760) );
DFFR_X2 inst_7011 ( .D(net_3269), .QN(net_281), .CK(net_12648), .RN(x1822) );
AOI22_X2 inst_7271 ( .B1(net_7085), .A1(net_7053), .A2(net_5280), .B2(net_5279), .ZN(net_5277) );
CLKBUF_X2 inst_10683 ( .A(net_7961), .Z(net_10645) );
SDFF_X2 inst_616 ( .Q(net_6621), .D(net_6621), .SE(net_3830), .SI(net_3801), .CK(net_12016) );
INV_X4 inst_5381 ( .A(net_7383), .ZN(net_568) );
CLKBUF_X2 inst_11049 ( .A(net_11010), .Z(net_11011) );
CLKBUF_X2 inst_9649 ( .A(net_8415), .Z(net_9611) );
CLKBUF_X2 inst_9320 ( .A(net_9281), .Z(net_9282) );
SDFF_X2 inst_620 ( .SI(net_7799), .Q(net_6597), .D(net_6597), .SE(net_3830), .CK(net_9339) );
OAI21_X2 inst_1784 ( .B1(net_5444), .ZN(net_5407), .A(net_4681), .B2(net_3988) );
DFF_X1 inst_6496 ( .QN(net_7408), .D(net_5543), .CK(net_10098) );
NAND2_X2 inst_3118 ( .A1(net_6589), .A2(net_4897), .ZN(net_4883) );
DFF_X1 inst_6401 ( .QN(net_6140), .D(net_5687), .CK(net_8169) );
CLKBUF_X2 inst_8040 ( .A(net_8001), .Z(net_8002) );
DFF_X1 inst_6869 ( .D(net_2549), .Q(net_222), .CK(net_12820) );
OAI21_X2 inst_2071 ( .B1(net_5901), .B2(net_4436), .ZN(net_4422), .A(net_3648) );
OR2_X2 inst_1427 ( .A2(net_6688), .A1(net_6687), .ZN(net_673) );
CLKBUF_X2 inst_10421 ( .A(net_10382), .Z(net_10383) );
OR2_X2 inst_1409 ( .A1(net_3940), .ZN(net_1688), .A2(net_1687) );
CLKBUF_X2 inst_10757 ( .A(net_10718), .Z(net_10719) );
CLKBUF_X2 inst_11570 ( .A(net_11531), .Z(net_11532) );
CLKBUF_X2 inst_9183 ( .A(net_8593), .Z(net_9145) );
CLKBUF_X2 inst_13752 ( .A(net_13713), .Z(net_13714) );
CLKBUF_X2 inst_10056 ( .A(net_9301), .Z(net_10018) );
AOI22_X2 inst_7259 ( .B1(net_6950), .A1(net_6918), .A2(net_5298), .B2(net_5297), .ZN(net_5295) );
CLKBUF_X2 inst_14296 ( .A(net_14257), .Z(net_14258) );
INV_X4 inst_4662 ( .ZN(net_5886), .A(net_3924) );
XNOR2_X2 inst_87 ( .B(net_2244), .ZN(net_1301), .A(net_1300) );
CLKBUF_X2 inst_13509 ( .A(net_12395), .Z(net_13471) );
NAND2_X2 inst_2996 ( .A1(net_6725), .A2(net_5031), .ZN(net_5015) );
INV_X4 inst_5037 ( .A(net_7819), .ZN(net_3795) );
CLKBUF_X2 inst_10601 ( .A(net_9786), .Z(net_10563) );
NAND2_X2 inst_2918 ( .A2(net_7772), .ZN(net_5774), .A1(net_5610) );
CLKBUF_X2 inst_10036 ( .A(net_9997), .Z(net_9998) );
CLKBUF_X2 inst_11946 ( .A(net_10742), .Z(net_11908) );
NAND3_X2 inst_2721 ( .ZN(net_2380), .A1(net_1676), .A3(net_1524), .A2(net_986) );
CLKBUF_X2 inst_9576 ( .A(net_8916), .Z(net_9538) );
CLKBUF_X2 inst_9517 ( .A(net_8952), .Z(net_9479) );
SDFF_X2 inst_800 ( .D(net_7802), .SI(net_6902), .Q(net_6902), .SE(net_3781), .CK(net_11787) );
NAND2_X2 inst_3074 ( .A1(net_7120), .A2(net_4950), .ZN(net_4931) );
INV_X4 inst_5281 ( .A(net_7095), .ZN(net_816) );
CLKBUF_X2 inst_9925 ( .A(net_9886), .Z(net_9887) );
XNOR2_X2 inst_10 ( .A(net_4140), .ZN(net_3826), .B(net_720) );
CLKBUF_X2 inst_14002 ( .A(net_13963), .Z(net_13964) );
CLKBUF_X2 inst_8763 ( .A(net_8724), .Z(net_8725) );
XOR2_X2 inst_4 ( .A(net_2569), .Z(net_1246), .B(net_1245) );
NAND2_X2 inst_3795 ( .A1(net_7179), .A2(net_1637), .ZN(net_1550) );
AOI21_X2 inst_7770 ( .B1(net_6869), .ZN(net_4109), .B2(net_2579), .A(net_2356) );
NAND2_X1 inst_4337 ( .ZN(net_4390), .A2(net_3856), .A1(net_1793) );
CLKBUF_X2 inst_10475 ( .A(net_8540), .Z(net_10437) );
CLKBUF_X2 inst_7981 ( .A(net_7942), .Z(net_7943) );
NAND2_X2 inst_3272 ( .ZN(net_3702), .A1(net_3701), .A2(net_3231) );
CLKBUF_X2 inst_13555 ( .A(net_13516), .Z(net_13517) );
CLKBUF_X2 inst_13186 ( .A(net_13147), .Z(net_13148) );
CLKBUF_X2 inst_9846 ( .A(net_9807), .Z(net_9808) );
CLKBUF_X2 inst_9455 ( .A(net_9416), .Z(net_9417) );
INV_X4 inst_5459 ( .A(net_6062), .ZN(net_3372) );
CLKBUF_X2 inst_10494 ( .A(net_9296), .Z(net_10456) );
CLKBUF_X2 inst_14232 ( .A(net_14193), .Z(net_14194) );
CLKBUF_X2 inst_9867 ( .A(net_9828), .Z(net_9829) );
CLKBUF_X2 inst_10090 ( .A(net_10051), .Z(net_10052) );
OAI21_X2 inst_1866 ( .ZN(net_5248), .B1(net_5202), .A(net_4533), .B2(net_3870) );
CLKBUF_X2 inst_8795 ( .A(net_8361), .Z(net_8757) );
CLKBUF_X2 inst_11961 ( .A(net_11922), .Z(net_11923) );
OAI21_X2 inst_1878 ( .ZN(net_5221), .B1(net_5220), .A(net_4584), .B2(net_3867) );
INV_X4 inst_5136 ( .A(net_1938), .ZN(net_579) );
INV_X2 inst_6016 ( .ZN(net_1117), .A(net_123) );
DFF_X1 inst_6700 ( .QN(net_7298), .D(net_5375), .CK(net_9885) );
CLKBUF_X2 inst_10290 ( .A(net_8809), .Z(net_10252) );
INV_X4 inst_4731 ( .A(net_3200), .ZN(net_3187) );
SDFF_X2 inst_1276 ( .D(net_6388), .SE(net_6051), .SI(net_306), .Q(net_306), .CK(net_14200) );
SDFF_X2 inst_765 ( .Q(net_6889), .D(net_6889), .SE(net_3901), .SI(net_3793), .CK(net_11474) );
SDFF_X2 inst_256 ( .Q(net_6378), .SI(net_6377), .D(net_3495), .SE(net_392), .CK(net_13510) );
DFF_X2 inst_6205 ( .Q(net_6394), .D(net_6393), .CK(net_14183) );
CLKBUF_X2 inst_10790 ( .A(net_9372), .Z(net_10752) );
CLKBUF_X2 inst_9870 ( .A(net_8136), .Z(net_9832) );
CLKBUF_X2 inst_10664 ( .A(net_10625), .Z(net_10626) );
CLKBUF_X2 inst_9180 ( .A(net_9141), .Z(net_9142) );
OAI21_X2 inst_1902 ( .B1(net_5365), .ZN(net_5167), .A(net_4767), .B2(net_3941) );
CLKBUF_X2 inst_8626 ( .A(net_8587), .Z(net_8588) );
CLKBUF_X2 inst_14247 ( .A(net_14208), .Z(net_14209) );
CLKBUF_X2 inst_9635 ( .A(net_9596), .Z(net_9597) );
INV_X4 inst_5052 ( .A(net_1143), .ZN(net_758) );
INV_X2 inst_6038 ( .A(net_7623), .ZN(net_1873) );
NAND2_X2 inst_3422 ( .A2(net_5914), .ZN(net_3235), .A1(net_3234) );
CLKBUF_X2 inst_13791 ( .A(net_13752), .Z(net_13753) );
CLKBUF_X2 inst_13266 ( .A(net_11061), .Z(net_13228) );
NAND2_X2 inst_3832 ( .A2(net_1696), .ZN(net_1508), .A1(net_1507) );
NAND2_X2 inst_3978 ( .ZN(net_1292), .A1(net_885), .A2(net_312) );
DFF_X1 inst_6618 ( .QN(net_7579), .D(net_5389), .CK(net_13442) );
NAND2_X2 inst_4039 ( .A1(net_6667), .A2(net_1655), .ZN(net_1013) );
INV_X2 inst_6106 ( .A(net_7629), .ZN(net_1903) );
CLKBUF_X2 inst_11264 ( .A(net_11225), .Z(net_11226) );
NAND2_X2 inst_2967 ( .ZN(net_5460), .A1(net_4886), .A2(net_4885) );
CLKBUF_X2 inst_9354 ( .A(net_9315), .Z(net_9316) );
CLKBUF_X2 inst_13279 ( .A(net_11642), .Z(net_13241) );
CLKBUF_X2 inst_10214 ( .A(net_10175), .Z(net_10176) );
CLKBUF_X2 inst_10042 ( .A(net_10003), .Z(net_10004) );
CLKBUF_X2 inst_9161 ( .A(net_9122), .Z(net_9123) );
OAI21_X2 inst_2078 ( .B2(net_4415), .ZN(net_4412), .B1(net_4033), .A(net_3508) );
DFF_X1 inst_6555 ( .QN(net_7268), .D(net_5157), .CK(net_12735) );
INV_X4 inst_5674 ( .A(net_7259), .ZN(net_2212) );
CLKBUF_X2 inst_9029 ( .A(net_7877), .Z(net_8991) );
SDFF_X2 inst_699 ( .SI(net_6769), .Q(net_6769), .SE(net_3816), .D(net_3813), .CK(net_11149) );
CLKBUF_X2 inst_8509 ( .A(net_8362), .Z(net_8471) );
OAI22_X2 inst_1462 ( .B2(net_5912), .B1(net_4637), .A2(net_4605), .ZN(net_4604), .A1(net_4014) );
CLKBUF_X2 inst_8377 ( .A(net_8338), .Z(net_8339) );
NOR2_X4 inst_2273 ( .ZN(net_5613), .A1(net_5458), .A2(net_4407) );
CLKBUF_X2 inst_9138 ( .A(net_9078), .Z(net_9100) );
CLKBUF_X2 inst_9921 ( .A(net_9882), .Z(net_9883) );
CLKBUF_X2 inst_13944 ( .A(net_12942), .Z(net_13906) );
DFF_X1 inst_6391 ( .QN(net_6122), .D(net_5697), .CK(net_11193) );
OAI21_X2 inst_2003 ( .B2(net_4518), .ZN(net_4510), .B1(net_4122), .A(net_3688) );
CLKBUF_X2 inst_9514 ( .A(net_9475), .Z(net_9476) );
INV_X4 inst_5430 ( .A(net_7557), .ZN(net_1987) );
INV_X2 inst_6084 ( .A(net_7449), .ZN(net_1476) );
INV_X2 inst_6100 ( .A(net_7602), .ZN(net_1344) );
CLKBUF_X2 inst_13823 ( .A(net_13784), .Z(net_13785) );
INV_X4 inst_5119 ( .ZN(net_3109), .A(net_598) );
INV_X4 inst_4963 ( .A(net_3778), .ZN(net_717) );
NAND3_X2 inst_2787 ( .ZN(net_2313), .A3(net_1523), .A1(net_1380), .A2(net_1021) );
INV_X4 inst_5612 ( .A(net_7706), .ZN(net_848) );
CLKBUF_X2 inst_13638 ( .A(net_13599), .Z(net_13600) );
CLKBUF_X2 inst_13144 ( .A(net_12661), .Z(net_13106) );
CLKBUF_X2 inst_12455 ( .A(net_8889), .Z(net_12417) );
CLKBUF_X2 inst_11074 ( .A(net_11035), .Z(net_11036) );
CLKBUF_X2 inst_9386 ( .A(net_9347), .Z(net_9348) );
NOR2_X2 inst_2426 ( .ZN(net_3435), .A2(net_3124), .A1(net_3050) );
NAND3_X2 inst_2599 ( .ZN(net_5740), .A1(net_5635), .A2(net_5210), .A3(net_4199) );
DFF_X2 inst_6254 ( .QN(net_7761), .D(net_2973), .CK(net_12774) );
CLKBUF_X2 inst_14211 ( .A(net_10087), .Z(net_14173) );
NAND2_X2 inst_3971 ( .A1(net_6566), .A2(net_1705), .ZN(net_1299) );
DFF_X1 inst_6377 ( .QN(net_6285), .D(net_5807), .CK(net_14255) );
OAI22_X2 inst_1485 ( .B1(net_4666), .ZN(net_4133), .A1(net_4132), .A2(net_4131), .B2(net_4130) );
CLKBUF_X2 inst_11573 ( .A(net_11534), .Z(net_11535) );
CLKBUF_X2 inst_9858 ( .A(net_8235), .Z(net_9820) );
CLKBUF_X2 inst_13596 ( .A(net_13557), .Z(net_13558) );
CLKBUF_X2 inst_12259 ( .A(net_12220), .Z(net_12221) );
SDFF_X2 inst_750 ( .Q(net_6872), .D(net_6872), .SE(net_3901), .SI(net_3813), .CK(net_11490) );
SDFF_X2 inst_317 ( .SI(net_7460), .Q(net_7460), .D(net_5101), .SE(net_3993), .CK(net_9786) );
CLKBUF_X2 inst_10561 ( .A(net_9669), .Z(net_10523) );
SDFF_X2 inst_1123 ( .SI(net_6673), .Q(net_6673), .D(net_3831), .SE(net_3471), .CK(net_12001) );
CLKBUF_X2 inst_8947 ( .A(net_7995), .Z(net_8909) );
CLKBUF_X2 inst_8747 ( .A(net_8708), .Z(net_8709) );
CLKBUF_X2 inst_13383 ( .A(net_13344), .Z(net_13345) );
SDFF_X2 inst_278 ( .D(net_6398), .SE(net_5799), .SI(net_383), .Q(net_383), .CK(net_13907) );
NAND2_X1 inst_4429 ( .A1(net_7609), .A2(net_2131), .ZN(net_1445) );
SDFF_X2 inst_467 ( .Q(net_7152), .D(net_7152), .SE(net_3903), .SI(net_3900), .CK(net_11599) );
CLKBUF_X2 inst_11763 ( .A(net_10649), .Z(net_11725) );
NAND2_X2 inst_3677 ( .A2(net_1798), .ZN(net_1779), .A1(net_1778) );
NAND2_X2 inst_3456 ( .ZN(net_2988), .A2(net_2741), .A1(net_189) );
CLKBUF_X2 inst_8061 ( .A(net_7865), .Z(net_8023) );
OAI22_X1 inst_1628 ( .B2(net_4300), .ZN(net_3981), .A2(net_3746), .A1(net_1712), .B1(net_1085) );
NAND2_X2 inst_2963 ( .ZN(net_5464), .A1(net_4894), .A2(net_4893) );
CLKBUF_X2 inst_7923 ( .A(net_7884), .Z(net_7885) );
DFF_X1 inst_6844 ( .D(net_2556), .QN(net_193), .CK(net_9978) );
CLKBUF_X2 inst_10535 ( .A(net_10496), .Z(net_10497) );
CLKBUF_X2 inst_9640 ( .A(net_9596), .Z(net_9602) );
SDFFR_X2 inst_1329 ( .SI(net_7769), .Q(net_7769), .SE(net_4804), .D(net_4803), .CK(net_12375), .RN(x1822) );
SDFF_X2 inst_1204 ( .SI(net_7088), .Q(net_7088), .D(net_3788), .SE(net_3747), .CK(net_8187) );
CLKBUF_X2 inst_8687 ( .A(net_8648), .Z(net_8649) );
NAND2_X2 inst_4066 ( .A1(net_7201), .A2(net_1648), .ZN(net_986) );
SDFF_X2 inst_225 ( .Q(net_6329), .SI(net_6328), .D(net_3627), .SE(net_392), .CK(net_14031) );
INV_X4 inst_4840 ( .A(net_3855), .ZN(net_3044) );
AOI21_X2 inst_7669 ( .B2(net_2838), .ZN(net_2810), .B1(net_2809), .A(net_2726) );
CLKBUF_X2 inst_14261 ( .A(net_11774), .Z(net_14223) );
CLKBUF_X2 inst_13568 ( .A(net_13529), .Z(net_13530) );
CLKBUF_X2 inst_12530 ( .A(net_12491), .Z(net_12492) );
CLKBUF_X2 inst_9030 ( .A(net_8991), .Z(net_8992) );
INV_X4 inst_5020 ( .A(net_7796), .ZN(net_3892) );
CLKBUF_X2 inst_13158 ( .A(net_13119), .Z(net_13120) );
CLKBUF_X2 inst_10162 ( .A(net_9522), .Z(net_10124) );
AOI22_X2 inst_7349 ( .B2(net_3105), .ZN(net_3101), .A2(net_2712), .A1(net_1129), .B1(net_739) );
SDFF_X2 inst_508 ( .SI(net_6498), .Q(net_6498), .D(net_3894), .SE(net_3889), .CK(net_8665) );
CLKBUF_X2 inst_11015 ( .A(net_10976), .Z(net_10977) );
INV_X4 inst_4888 ( .ZN(net_2252), .A(net_879) );
CLKBUF_X2 inst_8150 ( .A(net_8111), .Z(net_8112) );
CLKBUF_X2 inst_11718 ( .A(net_11679), .Z(net_11680) );
CLKBUF_X2 inst_12611 ( .A(net_12572), .Z(net_12573) );
NAND3_X2 inst_2618 ( .ZN(net_5721), .A1(net_5616), .A2(net_5133), .A3(net_4180) );
CLKBUF_X2 inst_10952 ( .A(net_10913), .Z(net_10914) );
INV_X4 inst_4950 ( .ZN(net_735), .A(net_734) );
CLKBUF_X2 inst_8853 ( .A(net_8814), .Z(net_8815) );
CLKBUF_X2 inst_11443 ( .A(net_9657), .Z(net_11405) );
CLKBUF_X2 inst_9241 ( .A(net_9202), .Z(net_9203) );
SDFF_X2 inst_590 ( .Q(net_6561), .D(net_6561), .SE(net_3823), .SI(net_3802), .CK(net_10056) );
NOR2_X2 inst_2553 ( .A2(net_5990), .A1(net_5984), .ZN(net_2893) );
CLKBUF_X2 inst_12209 ( .A(net_11147), .Z(net_12171) );
CLKBUF_X2 inst_13051 ( .A(net_13012), .Z(net_13013) );
CLKBUF_X2 inst_12671 ( .A(net_12632), .Z(net_12633) );
CLKBUF_X2 inst_14428 ( .A(net_14389), .Z(net_14390) );
CLKBUF_X2 inst_13897 ( .A(net_12051), .Z(net_13859) );
OAI21_X2 inst_1729 ( .ZN(net_5565), .B1(net_5432), .A(net_4830), .B2(net_4153) );
CLKBUF_X2 inst_8346 ( .A(net_8307), .Z(net_8308) );
SDFF_X2 inst_1105 ( .SI(net_6660), .Q(net_6660), .D(net_3798), .SE(net_3471), .CK(net_12894) );
INV_X8 inst_4531 ( .A(net_3937), .ZN(net_2838) );
CLKBUF_X2 inst_13175 ( .A(net_13136), .Z(net_13137) );
NAND3_X2 inst_2746 ( .ZN(net_2355), .A3(net_1552), .A1(net_1516), .A2(net_1007) );
INV_X16 inst_6126 ( .ZN(net_4518), .A(net_3848) );
CLKBUF_X2 inst_14387 ( .A(net_14348), .Z(net_14349) );
DFFR_X2 inst_6996 ( .QN(net_7705), .D(net_3357), .CK(net_10362), .RN(x1822) );
CLKBUF_X2 inst_13576 ( .A(net_13537), .Z(net_13538) );
INV_X4 inst_4648 ( .ZN(net_4165), .A(net_4164) );
CLKBUF_X2 inst_10469 ( .A(net_10430), .Z(net_10431) );
DFFR_X2 inst_6961 ( .QN(net_5848), .D(net_5480), .CK(net_12425), .RN(x1822) );
CLKBUF_X2 inst_8200 ( .A(net_8161), .Z(net_8162) );
SDFF_X2 inst_330 ( .SI(net_7496), .Q(net_7496), .D(net_5099), .SE(net_3989), .CK(net_9769) );
CLKBUF_X2 inst_13345 ( .A(net_13306), .Z(net_13307) );
CLKBUF_X2 inst_10297 ( .A(net_10258), .Z(net_10259) );
CLKBUF_X2 inst_13558 ( .A(net_10300), .Z(net_13520) );
CLKBUF_X2 inst_11460 ( .A(net_11421), .Z(net_11422) );
AOI222_X2 inst_7595 ( .A1(net_7395), .ZN(net_5446), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_358), .C2(net_356) );
SDFF_X2 inst_165 ( .Q(net_6249), .SI(net_6248), .D(net_3528), .SE(net_392), .CK(net_13977) );
NAND2_X2 inst_3733 ( .A1(net_6506), .A2(net_1642), .ZN(net_1612) );
NAND2_X1 inst_4305 ( .ZN(net_4561), .A2(net_3866), .A1(net_1883) );
CLKBUF_X2 inst_12101 ( .A(net_12062), .Z(net_12063) );
CLKBUF_X2 inst_13546 ( .A(net_13507), .Z(net_13508) );
INV_X4 inst_5376 ( .A(net_6147), .ZN(net_3589) );
CLKBUF_X2 inst_8786 ( .A(net_8747), .Z(net_8748) );
SDFF_X2 inst_1176 ( .SI(net_6948), .Q(net_6948), .D(net_3780), .SE(net_3734), .CK(net_11692) );
NAND2_X2 inst_3566 ( .ZN(net_2501), .A2(net_2217), .A1(net_1760) );
CLKBUF_X2 inst_13864 ( .A(net_13825), .Z(net_13826) );
CLKBUF_X2 inst_12537 ( .A(net_8459), .Z(net_12499) );
CLKBUF_X2 inst_11803 ( .A(net_11764), .Z(net_11765) );
CLKBUF_X2 inst_8159 ( .A(net_8120), .Z(net_8121) );
CLKBUF_X2 inst_12696 ( .A(net_12657), .Z(net_12658) );
SDFF_X2 inst_1232 ( .SI(net_7226), .Q(net_7226), .D(net_3800), .SE(net_3751), .CK(net_11833) );
INV_X4 inst_5450 ( .A(net_7264), .ZN(net_2059) );
CLKBUF_X2 inst_14431 ( .A(net_14392), .Z(net_14393) );
CLKBUF_X2 inst_11340 ( .A(net_8383), .Z(net_11302) );
NAND2_X2 inst_4172 ( .ZN(net_798), .A1(net_797), .A2(net_631) );
CLKBUF_X2 inst_13388 ( .A(net_13349), .Z(net_13350) );
NAND3_X2 inst_2605 ( .ZN(net_5734), .A1(net_5629), .A2(net_5172), .A3(net_4194) );
SDFF_X2 inst_758 ( .Q(net_6862), .D(net_6862), .SE(net_3901), .SI(net_3806), .CK(net_8935) );
CLKBUF_X2 inst_14423 ( .A(net_14384), .Z(net_14385) );
CLKBUF_X2 inst_14147 ( .A(net_14108), .Z(net_14109) );
OAI21_X2 inst_2146 ( .B1(net_5778), .ZN(net_2798), .A(net_2671), .B2(net_2669) );
CLKBUF_X2 inst_13759 ( .A(net_13720), .Z(net_13721) );
CLKBUF_X2 inst_13332 ( .A(net_13293), .Z(net_13294) );
AOI22_X2 inst_7252 ( .B1(net_6820), .A1(net_6788), .A2(net_5316), .B2(net_5315), .ZN(net_5308) );
CLKBUF_X2 inst_8543 ( .A(net_7932), .Z(net_8505) );
CLKBUF_X2 inst_13717 ( .A(net_13678), .Z(net_13679) );
NAND3_X2 inst_2703 ( .A3(net_5869), .ZN(net_2702), .A1(net_2644), .A2(net_689) );
NAND2_X2 inst_3437 ( .ZN(net_3211), .A2(net_3092), .A1(net_2760) );
CLKBUF_X2 inst_13425 ( .A(net_13386), .Z(net_13387) );
DFF_X1 inst_6813 ( .D(net_3253), .CK(net_13211), .Q(x195) );
CLKBUF_X2 inst_13857 ( .A(net_13818), .Z(net_13819) );
CLKBUF_X2 inst_9784 ( .A(net_9721), .Z(net_9746) );
INV_X2 inst_5764 ( .ZN(net_3027), .A(net_3026) );
SDFF_X2 inst_143 ( .Q(net_6235), .SI(net_6234), .SE(net_392), .D(net_141), .CK(net_13617) );
AOI22_X2 inst_7442 ( .ZN(net_4870), .A2(net_1222), .B1(net_1220), .B2(net_345), .A1(net_333) );
OAI21_X2 inst_1953 ( .ZN(net_5067), .B1(net_4849), .A(net_4724), .B2(net_3986) );
INV_X8 inst_4570 ( .A(net_5939), .ZN(net_5937) );
INV_X4 inst_5286 ( .A(net_6129), .ZN(net_3635) );
NAND2_X2 inst_3016 ( .A1(net_6890), .A2(net_5006), .ZN(net_4993) );
DFF_X2 inst_6260 ( .QN(net_5979), .D(net_2732), .CK(net_12203) );
OAI21_X2 inst_1958 ( .B1(net_5202), .ZN(net_5062), .A(net_4707), .B2(net_3986) );
NAND2_X1 inst_4272 ( .ZN(net_4642), .A2(net_3993), .A1(net_1448) );
CLKBUF_X2 inst_14050 ( .A(net_14011), .Z(net_14012) );
NOR2_X2 inst_2337 ( .A2(net_6281), .A1(net_5840), .ZN(net_5804) );
NAND2_X2 inst_3250 ( .ZN(net_5077), .A1(net_3855), .A2(net_3541) );
CLKBUF_X2 inst_9403 ( .A(net_9364), .Z(net_9365) );
CLKBUF_X2 inst_9357 ( .A(net_9318), .Z(net_9319) );
OAI21_X2 inst_1778 ( .B1(net_5432), .ZN(net_5416), .A(net_4695), .B2(net_3989) );
NAND2_X2 inst_3240 ( .ZN(net_4167), .A2(net_4166), .A1(net_2938) );
DFF_X1 inst_6885 ( .D(net_2500), .Q(net_161), .CK(net_10226) );
CLKBUF_X2 inst_12132 ( .A(net_12093), .Z(net_12094) );
CLKBUF_X2 inst_8091 ( .A(net_8052), .Z(net_8053) );
OAI21_X2 inst_1736 ( .ZN(net_5549), .B1(net_5548), .A(net_4811), .B2(net_4153) );
SDFF_X2 inst_1040 ( .Q(net_7543), .D(net_7543), .SE(net_3896), .SI(net_377), .CK(net_13105) );
NAND2_X2 inst_4027 ( .A1(net_6804), .A2(net_1651), .ZN(net_1025) );
CLKBUF_X2 inst_9158 ( .A(net_8940), .Z(net_9120) );
INV_X2 inst_6009 ( .A(net_6049), .ZN(net_2605) );
INV_X4 inst_5042 ( .ZN(net_754), .A(net_289) );
CLKBUF_X2 inst_13196 ( .A(net_13157), .Z(net_13158) );
XNOR2_X2 inst_111 ( .A(net_2573), .ZN(net_830), .B(net_829) );
OAI21_X2 inst_1723 ( .ZN(net_5571), .B1(net_5444), .A(net_4836), .B2(net_4153) );
NAND2_X2 inst_3146 ( .ZN(net_4817), .A2(net_4153), .A1(net_1981) );
NAND2_X2 inst_3278 ( .ZN(net_3690), .A1(net_3689), .A2(net_3231) );
CLKBUF_X2 inst_10246 ( .A(net_10207), .Z(net_10208) );
AOI22_X2 inst_7303 ( .B1(net_6541), .A1(net_6509), .A2(net_5184), .B2(net_5183), .ZN(net_5145) );
CLKBUF_X2 inst_11651 ( .A(net_11612), .Z(net_11613) );
CLKBUF_X2 inst_11425 ( .A(net_11386), .Z(net_11387) );
OAI21_X2 inst_2056 ( .B1(net_5908), .B2(net_4457), .ZN(net_4442), .A(net_3553) );
INV_X4 inst_5145 ( .ZN(net_3003), .A(net_571) );
OAI21_X2 inst_2116 ( .ZN(net_3298), .B2(net_3297), .B1(net_3170), .A(net_3081) );
CLKBUF_X2 inst_11296 ( .A(net_8338), .Z(net_11258) );
NAND3_X2 inst_2825 ( .ZN(net_1680), .A1(net_1679), .A3(net_804), .A2(net_647) );
INV_X4 inst_5071 ( .A(net_3001), .ZN(net_775) );
CLKBUF_X2 inst_13407 ( .A(net_12695), .Z(net_13369) );
NAND2_X2 inst_4031 ( .A1(net_7207), .A2(net_1648), .ZN(net_1021) );
CLKBUF_X2 inst_8135 ( .A(net_8096), .Z(net_8097) );
SDFF_X2 inst_346 ( .SI(net_7307), .Q(net_7307), .D(net_4875), .SE(net_3859), .CK(net_9478) );
CLKBUF_X2 inst_8755 ( .A(net_8716), .Z(net_8717) );
SDFF_X2 inst_978 ( .SI(net_7799), .Q(net_6430), .D(net_6430), .SE(net_3820), .CK(net_8641) );
CLKBUF_X2 inst_13506 ( .A(net_8908), .Z(net_13468) );
CLKBUF_X2 inst_10711 ( .A(net_10672), .Z(net_10673) );
NAND2_X2 inst_2955 ( .ZN(net_5485), .A1(net_5038), .A2(net_4939) );
CLKBUF_X2 inst_12058 ( .A(net_10284), .Z(net_12020) );
NAND2_X2 inst_3926 ( .A1(net_7461), .A2(net_1696), .ZN(net_1374) );
AOI22_X2 inst_7293 ( .B1(net_6543), .A1(net_6511), .ZN(net_5185), .A2(net_5184), .B2(net_5183) );
DFF_X2 inst_6195 ( .QN(net_6554), .D(net_5044), .CK(net_8819) );
CLKBUF_X2 inst_9777 ( .A(net_7944), .Z(net_9739) );
CLKBUF_X2 inst_11347 ( .A(net_11308), .Z(net_11309) );
CLKBUF_X2 inst_13160 ( .A(net_13121), .Z(net_13122) );
CLKBUF_X2 inst_12972 ( .A(net_12933), .Z(net_12934) );
NAND2_X2 inst_3929 ( .A1(net_7458), .A2(net_1696), .ZN(net_1369) );
CLKBUF_X2 inst_8856 ( .A(net_8817), .Z(net_8818) );
CLKBUF_X2 inst_12312 ( .A(net_12273), .Z(net_12274) );
CLKBUF_X2 inst_10506 ( .A(net_10467), .Z(net_10468) );
CLKBUF_X2 inst_9745 ( .A(net_9706), .Z(net_9707) );
NAND2_X2 inst_3852 ( .A1(net_6711), .A2(net_1497), .ZN(net_1483) );
CLKBUF_X2 inst_14168 ( .A(net_14129), .Z(net_14130) );
CLKBUF_X2 inst_14366 ( .A(net_14327), .Z(net_14328) );
SDFF_X2 inst_1051 ( .Q(net_7238), .D(net_7238), .SE(net_3822), .SI(net_334), .CK(net_12659) );
SDFF_X2 inst_495 ( .Q(net_6477), .D(net_6477), .SE(net_3904), .SI(net_3900), .CK(net_8098) );
NAND3_X4 inst_2566 ( .A2(net_5933), .ZN(net_3360), .A3(net_2915), .A1(net_689) );
INV_X2 inst_6102 ( .A(net_6031), .ZN(net_394) );
DFF_X1 inst_6437 ( .QN(net_6080), .D(net_5733), .CK(net_11281) );
OAI21_X2 inst_1864 ( .ZN(net_5251), .B1(net_5206), .A(net_4535), .B2(net_3870) );
CLKBUF_X2 inst_12901 ( .A(net_12862), .Z(net_12863) );
CLKBUF_X2 inst_9632 ( .A(net_9593), .Z(net_9594) );
NAND2_X2 inst_3603 ( .ZN(net_2397), .A2(net_1886), .A1(net_1414) );
CLKBUF_X2 inst_11076 ( .A(net_11037), .Z(net_11038) );
NAND2_X2 inst_3224 ( .A2(net_7778), .ZN(net_5258), .A1(net_4298) );
CLKBUF_X2 inst_10887 ( .A(net_10848), .Z(net_10849) );
NAND2_X2 inst_3043 ( .A1(net_7026), .A2(net_4979), .ZN(net_4964) );
CLKBUF_X2 inst_8063 ( .A(net_8024), .Z(net_8025) );
CLKBUF_X2 inst_13665 ( .A(net_13626), .Z(net_13627) );
CLKBUF_X2 inst_7917 ( .A(net_7878), .Z(net_7879) );
CLKBUF_X2 inst_12616 ( .A(net_12577), .Z(net_12578) );
INV_X2 inst_5752 ( .ZN(net_3909), .A(net_3737) );
CLKBUF_X2 inst_13305 ( .A(net_13266), .Z(net_13267) );
CLKBUF_X2 inst_12644 ( .A(net_12605), .Z(net_12606) );
AOI22_X2 inst_7286 ( .B1(net_7223), .A1(net_7191), .A2(net_5244), .B2(net_5243), .ZN(net_5219) );
CLKBUF_X2 inst_10548 ( .A(net_10340), .Z(net_10510) );
CLKBUF_X2 inst_8914 ( .A(net_8875), .Z(net_8876) );
CLKBUF_X2 inst_13781 ( .A(net_13742), .Z(net_13743) );
NAND2_X4 inst_2893 ( .ZN(net_3858), .A2(net_3392), .A1(net_3245) );
CLKBUF_X2 inst_11360 ( .A(net_9766), .Z(net_11322) );
CLKBUF_X2 inst_9497 ( .A(net_9458), .Z(net_9459) );
SDFF_X2 inst_573 ( .Q(net_6559), .D(net_6559), .SE(net_3823), .SI(net_3797), .CK(net_9696) );
AOI21_X2 inst_7736 ( .B1(net_7139), .ZN(net_4082), .B2(net_2582), .A(net_2298) );
CLKBUF_X2 inst_12447 ( .A(net_12408), .Z(net_12409) );
DFF_X1 inst_6727 ( .QN(net_7361), .D(net_5328), .CK(net_12248) );
CLKBUF_X2 inst_7937 ( .A(net_7898), .Z(net_7899) );
CLKBUF_X2 inst_9041 ( .A(net_9002), .Z(net_9003) );
DFF_X1 inst_6347 ( .Q(net_6211), .D(net_5837), .CK(net_13767) );
CLKBUF_X2 inst_8088 ( .A(net_8049), .Z(net_8050) );
INV_X4 inst_5364 ( .A(net_6117), .ZN(net_3695) );
OAI22_X2 inst_1453 ( .B2(net_5898), .B1(net_4650), .ZN(net_4616), .A2(net_4614), .A1(net_4068) );
NAND2_X1 inst_4245 ( .ZN(net_4682), .A2(net_3988), .A1(net_2196) );
CLKBUF_X2 inst_12466 ( .A(net_12427), .Z(net_12428) );
CLKBUF_X2 inst_12391 ( .A(net_10109), .Z(net_12353) );
CLKBUF_X2 inst_8871 ( .A(net_7996), .Z(net_8833) );
NAND2_X2 inst_3007 ( .A1(net_6853), .A2(net_5004), .ZN(net_5002) );
CLKBUF_X2 inst_8978 ( .A(net_8939), .Z(net_8940) );
NAND2_X2 inst_4185 ( .ZN(net_812), .A2(net_797), .A1(net_522) );
CLKBUF_X2 inst_11018 ( .A(net_9455), .Z(net_10980) );
NAND2_X2 inst_3512 ( .ZN(net_2555), .A2(net_2157), .A1(net_1697) );
NAND2_X2 inst_3544 ( .ZN(net_2523), .A2(net_2092), .A1(net_1196) );
DFF_X1 inst_6358 ( .QN(net_6200), .D(net_5826), .CK(net_13640) );
CLKBUF_X2 inst_11485 ( .A(net_11330), .Z(net_11447) );
CLKBUF_X2 inst_10738 ( .A(net_10699), .Z(net_10700) );
CLKBUF_X2 inst_10973 ( .A(net_9381), .Z(net_10935) );
INV_X4 inst_5632 ( .ZN(net_624), .A(x1231) );
SDFF_X2 inst_1206 ( .SI(net_7090), .Q(net_7090), .D(net_3801), .SE(net_3747), .CK(net_8181) );
CLKBUF_X2 inst_7970 ( .A(net_7872), .Z(net_7932) );
CLKBUF_X2 inst_13607 ( .A(net_7875), .Z(net_13569) );
CLKBUF_X2 inst_9362 ( .A(net_9323), .Z(net_9324) );
DFF_X1 inst_6367 ( .QN(net_6295), .D(net_5817), .CK(net_13791) );
DFF_X1 inst_6773 ( .QN(net_6145), .D(net_4599), .CK(net_9135) );
CLKBUF_X2 inst_10328 ( .A(net_10289), .Z(net_10290) );
DFFR_X2 inst_7075 ( .QN(net_6423), .D(net_2821), .CK(net_13024), .RN(x1822) );
NAND2_X2 inst_3466 ( .A2(net_3439), .ZN(net_2854), .A1(net_2853) );
CLKBUF_X2 inst_8106 ( .A(net_8067), .Z(net_8068) );
CLKBUF_X2 inst_13907 ( .A(net_13868), .Z(net_13869) );
CLKBUF_X2 inst_8358 ( .A(net_8319), .Z(net_8320) );
INV_X4 inst_4800 ( .ZN(net_4776), .A(net_1236) );
NAND2_X1 inst_4394 ( .ZN(net_4333), .A2(net_3859), .A1(net_2160) );
CLKBUF_X2 inst_11303 ( .A(net_11264), .Z(net_11265) );
INV_X4 inst_5553 ( .A(net_6691), .ZN(net_492) );
CLKBUF_X2 inst_13086 ( .A(net_13047), .Z(net_13048) );
CLKBUF_X2 inst_12631 ( .A(net_12592), .Z(net_12593) );
CLKBUF_X2 inst_11518 ( .A(net_11111), .Z(net_11480) );
OAI22_X2 inst_1487 ( .B1(net_4666), .A1(net_4132), .B2(net_4131), .ZN(net_4127), .A2(net_4126) );
INV_X2 inst_6111 ( .A(net_5920), .ZN(net_5919) );
AND2_X4 inst_7807 ( .ZN(net_3846), .A2(net_3845), .A1(net_1147) );
CLKBUF_X2 inst_13169 ( .A(net_13130), .Z(net_13131) );
OAI21_X2 inst_1933 ( .ZN(net_5112), .A(net_4772), .B2(net_3941), .B1(net_1236) );
NAND2_X2 inst_3522 ( .ZN(net_2545), .A2(net_1984), .A1(net_1704) );
AOI22_X2 inst_7246 ( .B1(net_6814), .A1(net_6782), .A2(net_5316), .B2(net_5315), .ZN(net_5314) );
DFF_X2 inst_6306 ( .Q(net_7807), .CK(net_8683), .D(x1486) );
CLKBUF_X2 inst_14119 ( .A(net_13641), .Z(net_14081) );
AOI222_X2 inst_7511 ( .B1(net_7370), .C1(net_7306), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2032), .A1(net_2031) );
OAI21_X2 inst_1758 ( .ZN(net_5441), .B1(net_5440), .A(net_4664), .B2(net_3993) );
SDFF_X2 inst_1142 ( .SI(net_6801), .Q(net_6801), .D(net_3813), .SE(net_3729), .CK(net_8262) );
DFF_X2 inst_6280 ( .D(net_7792), .QN(net_7791), .CK(net_13201) );
CLKBUF_X2 inst_12025 ( .A(net_11986), .Z(net_11987) );
NAND2_X1 inst_4320 ( .ZN(net_4544), .A2(net_3870), .A1(net_1389) );
NAND2_X2 inst_3816 ( .A1(net_6640), .A2(net_1624), .ZN(net_1529) );
CLKBUF_X2 inst_11138 ( .A(net_8080), .Z(net_11100) );
INV_X4 inst_5418 ( .A(net_6558), .ZN(net_2571) );
OR2_X4 inst_1381 ( .ZN(net_2905), .A2(net_2754), .A1(net_267) );
SDFF_X2 inst_643 ( .SI(net_6627), .Q(net_6627), .SE(net_3850), .D(net_3799), .CK(net_12901) );
AOI222_X2 inst_7572 ( .ZN(net_5222), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_384), .C2(net_382), .A1(net_370) );
DFF_X2 inst_6313 ( .QN(net_6402), .CK(net_12960) );
AOI21_X2 inst_7680 ( .B1(net_6997), .ZN(net_4598), .A(net_2463), .B2(net_1100) );
CLKBUF_X2 inst_12471 ( .A(net_12195), .Z(net_12433) );
CLKBUF_X2 inst_13726 ( .A(net_10378), .Z(net_13688) );
CLKBUF_X2 inst_14316 ( .A(net_14277), .Z(net_14278) );
CLKBUF_X2 inst_14228 ( .A(net_13268), .Z(net_14190) );
CLKBUF_X2 inst_9430 ( .A(net_9391), .Z(net_9392) );
CLKBUF_X2 inst_14182 ( .A(net_8313), .Z(net_14144) );
CLKBUF_X2 inst_10745 ( .A(net_10706), .Z(net_10707) );
AOI21_X2 inst_7763 ( .B1(net_6466), .ZN(net_4062), .B2(net_2580), .A(net_2301) );
INV_X4 inst_4771 ( .ZN(net_2486), .A(net_1832) );
CLKBUF_X2 inst_12117 ( .A(net_12078), .Z(net_12079) );
CLKBUF_X2 inst_12220 ( .A(net_12181), .Z(net_12182) );
INV_X4 inst_4961 ( .ZN(net_903), .A(net_719) );
INV_X4 inst_4669 ( .ZN(net_3714), .A(net_3713) );
AOI21_X2 inst_7695 ( .B1(net_6465), .ZN(net_4055), .B2(net_2580), .A(net_2303) );
CLKBUF_X2 inst_8588 ( .A(net_8362), .Z(net_8550) );
CLKBUF_X2 inst_8016 ( .A(net_7977), .Z(net_7978) );
CLKBUF_X2 inst_8707 ( .A(net_8668), .Z(net_8669) );
DFF_X1 inst_6466 ( .QN(net_6151), .D(net_5593), .CK(net_11975) );
CLKBUF_X2 inst_12165 ( .A(net_11512), .Z(net_12127) );
CLKBUF_X2 inst_13204 ( .A(net_8314), .Z(net_13166) );
CLKBUF_X2 inst_8581 ( .A(net_8542), .Z(net_8543) );
INV_X4 inst_5447 ( .A(net_7097), .ZN(net_539) );
DFF_X1 inst_6371 ( .QN(net_6291), .D(net_5813), .CK(net_14279) );
NAND2_X2 inst_4146 ( .ZN(net_1687), .A2(net_892), .A1(net_882) );
CLKBUF_X2 inst_12526 ( .A(net_12487), .Z(net_12488) );
CLKBUF_X2 inst_12230 ( .A(net_7905), .Z(net_12192) );
CLKBUF_X2 inst_12959 ( .A(net_12920), .Z(net_12921) );
OAI21_X2 inst_1997 ( .B2(net_4518), .ZN(net_4516), .B1(net_4130), .A(net_3696) );
DFFR_X2 inst_6971 ( .QN(net_6026), .D(net_4003), .CK(net_10763), .RN(x1822) );
SDFF_X2 inst_1017 ( .SI(net_6511), .Q(net_6511), .SE(net_3886), .D(net_3780), .CK(net_8053) );
CLKBUF_X2 inst_12669 ( .A(net_12630), .Z(net_12631) );
NOR2_X2 inst_2297 ( .A2(net_6194), .ZN(net_5846), .A1(net_5843) );
NAND2_X2 inst_3736 ( .A1(net_6488), .A2(net_1642), .ZN(net_1609) );
CLKBUF_X2 inst_13802 ( .A(net_9590), .Z(net_13764) );
SDFF_X2 inst_281 ( .D(net_6397), .SE(net_5801), .SI(net_342), .Q(net_342), .CK(net_13905) );
NAND2_X2 inst_3341 ( .ZN(net_3565), .A1(net_3564), .A2(net_3225) );
CLKBUF_X2 inst_10306 ( .A(net_10267), .Z(net_10268) );
CLKBUF_X2 inst_8500 ( .A(net_8461), .Z(net_8462) );
DFF_X2 inst_6336 ( .QN(net_7816), .CK(net_10882), .D(x1406) );
CLKBUF_X2 inst_13411 ( .A(net_13372), .Z(net_13373) );
DFFR_X2 inst_7062 ( .QN(net_6028), .D(net_3054), .CK(net_10013), .RN(x1822) );
OAI21_X2 inst_1836 ( .ZN(net_5338), .B1(net_5337), .A(net_4353), .B2(net_3856) );
DFF_X1 inst_6374 ( .QN(net_6288), .D(net_5810), .CK(net_14267) );
DFFR_X2 inst_7005 ( .QN(net_7697), .D(net_3345), .CK(net_12873), .RN(x1822) );
NOR2_X2 inst_2508 ( .A2(net_3241), .ZN(net_1182), .A1(net_1181) );
CLKBUF_X2 inst_10207 ( .A(net_8583), .Z(net_10169) );
NOR4_X2 inst_2170 ( .ZN(net_3251), .A4(net_3121), .A1(net_2636), .A3(net_2478), .A2(net_817) );
NAND2_X1 inst_4250 ( .ZN(net_4676), .A2(net_3988), .A1(net_2164) );
NAND2_X1 inst_4274 ( .ZN(net_4639), .A2(net_3993), .A1(net_1358) );
CLKBUF_X2 inst_13322 ( .A(net_10914), .Z(net_13284) );
SDFF_X2 inst_773 ( .Q(net_6869), .D(net_6869), .SE(net_3901), .SI(net_3814), .CK(net_11804) );
AOI22_X2 inst_7414 ( .B1(net_5939), .ZN(net_2780), .A1(net_2578), .B2(net_216), .A2(net_179) );
CLKBUF_X2 inst_14149 ( .A(net_13601), .Z(net_14111) );
CLKBUF_X2 inst_9940 ( .A(net_9901), .Z(net_9902) );
NAND2_X2 inst_2946 ( .ZN(net_5500), .A1(net_4960), .A2(net_4959) );
CLKBUF_X2 inst_10776 ( .A(net_10737), .Z(net_10738) );
CLKBUF_X2 inst_13091 ( .A(net_13052), .Z(net_13053) );
CLKBUF_X2 inst_10074 ( .A(net_10035), .Z(net_10036) );
NAND2_X2 inst_3620 ( .ZN(net_1968), .A2(net_1967), .A1(net_1721) );
CLKBUF_X2 inst_13827 ( .A(net_13788), .Z(net_13789) );
CLKBUF_X2 inst_10828 ( .A(net_10789), .Z(net_10790) );
CLKBUF_X2 inst_14134 ( .A(net_12909), .Z(net_14096) );
CLKBUF_X2 inst_9798 ( .A(net_9759), .Z(net_9760) );
SDFF_X2 inst_260 ( .Q(net_6374), .SI(net_6373), .D(net_3521), .SE(net_392), .CK(net_13515) );
CLKBUF_X2 inst_11277 ( .A(net_11238), .Z(net_11239) );
CLKBUF_X2 inst_9371 ( .A(net_8756), .Z(net_9333) );
CLKBUF_X2 inst_11597 ( .A(net_11558), .Z(net_11559) );
NAND2_X2 inst_3211 ( .ZN(net_4715), .A2(net_3986), .A1(net_1879) );
INV_X4 inst_4973 ( .A(net_7810), .ZN(net_3776) );
CLKBUF_X2 inst_10364 ( .A(net_10325), .Z(net_10326) );
CLKBUF_X2 inst_12702 ( .A(net_12663), .Z(net_12664) );
AOI22_X2 inst_7270 ( .B1(net_7084), .A1(net_7052), .A2(net_5280), .B2(net_5279), .ZN(net_5278) );
NAND2_X2 inst_4139 ( .ZN(net_1107), .A1(net_920), .A2(net_891) );
DFF_X1 inst_6762 ( .QN(net_7365), .D(net_4860), .CK(net_9865) );
INV_X4 inst_4611 ( .ZN(net_4233), .A(net_4085) );
CLKBUF_X2 inst_13839 ( .A(net_13800), .Z(net_13801) );
CLKBUF_X2 inst_10906 ( .A(net_9159), .Z(net_10868) );
CLKBUF_X2 inst_10725 ( .A(net_10686), .Z(net_10687) );
INV_X8 inst_4567 ( .ZN(net_5916), .A(net_2702) );
NAND2_X2 inst_3889 ( .A1(net_6696), .A2(net_1497), .ZN(net_1427) );
NOR2_X2 inst_2386 ( .ZN(net_4147), .A1(net_4146), .A2(net_4145) );
CLKBUF_X2 inst_9880 ( .A(net_9841), .Z(net_9842) );
CLKBUF_X2 inst_8739 ( .A(net_8700), .Z(net_8701) );
SDFF_X2 inst_516 ( .Q(net_6715), .D(net_6715), .SI(net_3900), .SE(net_3871), .CK(net_10934) );
CLKBUF_X2 inst_12243 ( .A(net_12204), .Z(net_12205) );
NOR2_X4 inst_2258 ( .ZN(net_5628), .A1(net_5473), .A2(net_4431) );
CLKBUF_X2 inst_13986 ( .A(net_13947), .Z(net_13948) );
CLKBUF_X2 inst_13846 ( .A(net_13807), .Z(net_13808) );
SDFF_X2 inst_190 ( .Q(net_6264), .SI(net_6263), .D(net_3485), .SE(net_392), .CK(net_13470) );
CLKBUF_X2 inst_9602 ( .A(net_9563), .Z(net_9564) );
SDFF_X2 inst_1267 ( .Q(net_5860), .SE(net_3184), .SI(net_3183), .D(net_509), .CK(net_9476) );
NAND2_X2 inst_4103 ( .A1(net_6661), .A2(net_1655), .ZN(net_949) );
OAI22_X2 inst_1507 ( .B1(net_4660), .B2(net_4498), .A1(net_4105), .A2(net_4103), .ZN(net_4085) );
INV_X4 inst_4873 ( .ZN(net_1087), .A(net_666) );
CLKBUF_X2 inst_13484 ( .A(net_13445), .Z(net_13446) );
CLKBUF_X2 inst_9932 ( .A(net_9893), .Z(net_9894) );
AOI22_X2 inst_7301 ( .B1(net_6551), .A1(net_6519), .A2(net_5184), .B2(net_5183), .ZN(net_5168) );
DFF_X1 inst_6424 ( .QN(net_6179), .D(net_5746), .CK(net_8742) );
OAI21_X2 inst_2062 ( .B2(net_4436), .ZN(net_4433), .B1(net_4062), .A(net_3576) );
NOR2_X2 inst_2350 ( .ZN(net_5654), .A1(net_5506), .A2(net_4473) );
NAND2_X2 inst_3786 ( .A1(net_6777), .A2(net_1635), .ZN(net_1559) );
AOI22_X2 inst_7260 ( .B1(net_6951), .A1(net_6919), .A2(net_5298), .B2(net_5297), .ZN(net_5294) );
NAND2_X2 inst_3404 ( .A2(net_5929), .ZN(net_3373), .A1(net_3372) );
AOI22_X2 inst_7367 ( .B1(net_7739), .A1(net_7710), .A2(net_5916), .B2(net_2957), .ZN(net_2955) );
SDFF_X2 inst_542 ( .SI(net_7173), .Q(net_7173), .D(net_3894), .SE(net_3819), .CK(net_13378) );
INV_X4 inst_5351 ( .A(net_6150), .ZN(net_3583) );
CLKBUF_X2 inst_7878 ( .A(net_7839), .Z(net_7840) );
SDFF_X2 inst_128 ( .Q(net_6193), .SI(net_6192), .D(net_3919), .SE(net_392), .CK(net_13747) );
CLKBUF_X2 inst_13589 ( .A(net_13550), .Z(net_13551) );
CLKBUF_X2 inst_14322 ( .A(net_14283), .Z(net_14284) );
CLKBUF_X2 inst_14172 ( .A(net_8234), .Z(net_14134) );
CLKBUF_X2 inst_13100 ( .A(net_8459), .Z(net_13062) );
CLKBUF_X2 inst_13222 ( .A(net_13183), .Z(net_13184) );
CLKBUF_X2 inst_11911 ( .A(net_11872), .Z(net_11873) );
NAND2_X2 inst_4000 ( .ZN(net_1156), .A1(net_918), .A2(net_812) );
CLKBUF_X2 inst_13625 ( .A(net_11367), .Z(net_13587) );
NAND2_X2 inst_3435 ( .ZN(net_3213), .A2(net_3095), .A1(net_2762) );
DFF_X1 inst_6934 ( .D(net_2386), .Q(net_250), .CK(net_10411) );
NAND2_X2 inst_3218 ( .ZN(net_4708), .A2(net_3986), .A1(net_1987) );
CLKBUF_X2 inst_9345 ( .A(net_8844), .Z(net_9307) );
SDFF_X2 inst_829 ( .Q(net_7008), .D(net_7008), .SE(net_3899), .SI(net_3812), .CK(net_8221) );
DFF_X1 inst_6904 ( .D(net_2505), .Q(net_185), .CK(net_12406) );
CLKBUF_X2 inst_8137 ( .A(net_7944), .Z(net_8099) );
SDFF_X2 inst_197 ( .Q(net_6317), .SI(net_6316), .D(net_3617), .SE(net_392), .CK(net_13591) );
AOI22_X2 inst_7277 ( .B1(net_7091), .A1(net_7059), .A2(net_5280), .B2(net_5279), .ZN(net_5271) );
NAND2_X2 inst_2958 ( .ZN(net_5482), .A1(net_4934), .A2(net_4933) );
INV_X4 inst_4702 ( .ZN(net_3339), .A(net_3070) );
INV_X2 inst_5723 ( .ZN(net_4005), .A(net_3914) );
XNOR2_X2 inst_24 ( .ZN(net_2574), .B(net_2573), .A(net_2438) );
CLKBUF_X2 inst_10129 ( .A(net_10090), .Z(net_10091) );
SDFF_X2 inst_1209 ( .SI(net_7065), .Q(net_7065), .D(net_3798), .SE(net_3747), .CK(net_11921) );
CLKBUF_X2 inst_12830 ( .A(net_12791), .Z(net_12792) );
CLKBUF_X2 inst_8190 ( .A(net_7915), .Z(net_8152) );
CLKBUF_X2 inst_11155 ( .A(net_11116), .Z(net_11117) );
CLKBUF_X2 inst_8558 ( .A(net_8519), .Z(net_8520) );
OAI22_X2 inst_1611 ( .A1(net_3273), .A2(net_3087), .B2(net_3084), .ZN(net_3067), .B1(net_480) );
SDFF_X2 inst_150 ( .Q(net_6228), .SI(net_6227), .SE(net_392), .D(net_134), .CK(net_14100) );
DFF_X1 inst_6743 ( .QN(net_7666), .D(net_4842), .CK(net_13419) );
INV_X4 inst_5358 ( .A(net_7719), .ZN(net_855) );
INV_X8 inst_4469 ( .ZN(net_5298), .A(net_4281) );
CLKBUF_X2 inst_12764 ( .A(net_12725), .Z(net_12726) );
DFF_X1 inst_6779 ( .QN(net_6105), .D(net_4325), .CK(net_8981) );
INV_X8 inst_4540 ( .ZN(net_2582), .A(net_1282) );
SDFF_X2 inst_887 ( .Q(net_7118), .D(net_7118), .SE(net_3888), .SI(net_3807), .CK(net_7864) );
CLKBUF_X2 inst_8730 ( .A(net_7983), .Z(net_8692) );
CLKBUF_X2 inst_8466 ( .A(net_8413), .Z(net_8428) );
INV_X2 inst_5849 ( .A(net_6402), .ZN(net_688) );
INV_X4 inst_5175 ( .ZN(net_3002), .A(net_532) );
CLKBUF_X2 inst_8036 ( .A(net_7855), .Z(net_7998) );
OAI221_X2 inst_1663 ( .C2(net_5897), .ZN(net_4661), .B1(net_4660), .B2(net_4485), .C1(net_4105), .A(net_3640) );
NAND3_X2 inst_2714 ( .ZN(net_2462), .A2(net_1807), .A3(net_1621), .A1(net_1405) );
CLKBUF_X2 inst_13223 ( .A(net_12742), .Z(net_13185) );
CLKBUF_X2 inst_8547 ( .A(net_8508), .Z(net_8509) );
DFFR_X2 inst_7099 ( .D(net_1957), .QN(net_117), .CK(net_9592), .RN(x1822) );
CLKBUF_X2 inst_13647 ( .A(net_13608), .Z(net_13609) );
NAND2_X1 inst_4316 ( .ZN(net_4548), .A2(net_3870), .A1(net_1465) );
NOR2_X2 inst_2357 ( .ZN(net_5647), .A1(net_5499), .A2(net_4462) );
CLKBUF_X2 inst_13036 ( .A(net_12997), .Z(net_12998) );
CLKBUF_X2 inst_13911 ( .A(net_13872), .Z(net_13873) );
DFF_X1 inst_6541 ( .QN(net_7473), .D(net_5575), .CK(net_12105) );
CLKBUF_X2 inst_7962 ( .A(net_7923), .Z(net_7924) );
CLKBUF_X2 inst_12248 ( .A(net_12209), .Z(net_12210) );
OAI21_X2 inst_1961 ( .B1(net_5196), .ZN(net_5059), .A(net_4704), .B2(net_3986) );
CLKBUF_X2 inst_14343 ( .A(net_9710), .Z(net_14305) );
INV_X2 inst_5799 ( .A(net_2486), .ZN(net_1973) );
CLKBUF_X2 inst_11285 ( .A(net_11246), .Z(net_11247) );
INV_X2 inst_5954 ( .A(net_7319), .ZN(net_1776) );
SDFF_X2 inst_1010 ( .SI(net_6503), .Q(net_6503), .SE(net_3886), .D(net_3787), .CK(net_8852) );
CLKBUF_X2 inst_10713 ( .A(net_10674), .Z(net_10675) );
CLKBUF_X2 inst_7934 ( .A(net_7839), .Z(net_7896) );
SDFF_X2 inst_867 ( .SI(net_7054), .Q(net_7054), .D(net_3790), .SE(net_3777), .CK(net_8214) );
SDFF_X2 inst_820 ( .Q(net_6994), .D(net_6994), .SE(net_3891), .SI(net_3801), .CK(net_10869) );
INV_X2 inst_6021 ( .ZN(net_1109), .A(net_119) );
CLKBUF_X2 inst_14179 ( .A(net_7969), .Z(net_14141) );
OAI22_X2 inst_1441 ( .B2(net_5895), .B1(net_4666), .ZN(net_4635), .A2(net_4634), .A1(net_4118) );
SDFF_X2 inst_157 ( .Q(net_6257), .SI(net_6256), .D(net_3544), .SE(net_392), .CK(net_13994) );
NAND2_X2 inst_2929 ( .ZN(net_5524), .A1(net_4997), .A2(net_4996) );
CLKBUF_X2 inst_12154 ( .A(net_12115), .Z(net_12116) );
NAND2_X2 inst_3443 ( .ZN(net_3163), .A2(net_3162), .A1(net_3147) );
NAND2_X2 inst_3568 ( .ZN(net_2499), .A2(net_2002), .A1(net_1773) );
DFF_X2 inst_6202 ( .QN(net_6957), .D(net_4396), .CK(net_11411) );
INV_X1 inst_6159 ( .A(net_5851), .ZN(x77) );
NAND2_X1 inst_4287 ( .ZN(net_4580), .A2(net_3867), .A1(net_1197) );
CLKBUF_X2 inst_10986 ( .A(net_10947), .Z(net_10948) );
CLKBUF_X2 inst_10760 ( .A(net_10721), .Z(net_10722) );
NOR4_X2 inst_2177 ( .A2(net_7752), .ZN(net_3317), .A3(net_3208), .A1(net_2918), .A4(net_682) );
INV_X4 inst_5491 ( .A(net_7412), .ZN(net_2205) );
CLKBUF_X2 inst_8963 ( .A(net_8924), .Z(net_8925) );
CLKBUF_X2 inst_12364 ( .A(net_10611), .Z(net_12326) );
CLKBUF_X2 inst_9342 ( .A(net_9303), .Z(net_9304) );
CLKBUF_X2 inst_9588 ( .A(net_8533), .Z(net_9550) );
NAND2_X2 inst_4158 ( .A1(net_7680), .ZN(net_918), .A2(net_457) );
CLKBUF_X2 inst_11481 ( .A(net_11442), .Z(net_11443) );
CLKBUF_X2 inst_8348 ( .A(net_7831), .Z(net_8310) );
OAI221_X2 inst_1643 ( .ZN(net_5452), .B2(net_5057), .C2(net_5055), .A(net_4956), .C1(net_1152), .B1(net_746) );
AOI22_X2 inst_7447 ( .A2(net_2952), .B2(net_2682), .ZN(net_852), .A1(net_851), .B1(net_850) );
NAND2_X2 inst_3410 ( .A2(net_5960), .ZN(net_3453), .A1(net_2881) );
INV_X4 inst_4660 ( .ZN(net_5881), .A(net_3926) );
OAI21_X2 inst_2120 ( .B2(net_3297), .ZN(net_3292), .B1(net_3291), .A(net_3074) );
NAND3_X2 inst_2678 ( .ZN(net_3458), .A3(net_3304), .A1(net_2969), .A2(net_2955) );
INV_X4 inst_5339 ( .A(net_6116), .ZN(net_3697) );
CLKBUF_X2 inst_13478 ( .A(net_13439), .Z(net_13440) );
CLKBUF_X2 inst_11506 ( .A(net_11467), .Z(net_11468) );
CLKBUF_X2 inst_9196 ( .A(net_9157), .Z(net_9158) );
CLKBUF_X2 inst_13216 ( .A(net_13177), .Z(net_13178) );
NAND3_X2 inst_2613 ( .ZN(net_5726), .A1(net_5621), .A2(net_5140), .A3(net_4185) );
XNOR2_X2 inst_17 ( .ZN(net_2635), .B(net_2634), .A(net_2481) );
CLKBUF_X2 inst_10577 ( .A(net_10041), .Z(net_10539) );
CLKBUF_X2 inst_10105 ( .A(net_10021), .Z(net_10067) );
SDFF_X2 inst_249 ( .Q(net_6345), .SI(net_6344), .D(net_3573), .SE(net_392), .CK(net_13650) );
AND2_X4 inst_7838 ( .ZN(net_1964), .A2(net_787), .A1(net_661) );
CLKBUF_X2 inst_12239 ( .A(net_11106), .Z(net_12201) );
NAND2_X2 inst_3866 ( .A2(net_1696), .ZN(net_1464), .A1(net_1463) );
CLKBUF_X2 inst_12407 ( .A(net_12368), .Z(net_12369) );
NOR2_X4 inst_2234 ( .ZN(net_5664), .A1(net_5522), .A2(net_4492) );
CLKBUF_X2 inst_10460 ( .A(net_8416), .Z(net_10422) );
DFF_X2 inst_6251 ( .QN(net_7757), .D(net_3021), .CK(net_10511) );
CLKBUF_X2 inst_8186 ( .A(net_7922), .Z(net_8148) );
CLKBUF_X2 inst_7976 ( .A(net_7937), .Z(net_7938) );
NAND2_X1 inst_4371 ( .ZN(net_4356), .A2(net_3856), .A1(net_1772) );
INV_X4 inst_5204 ( .ZN(net_646), .A(net_495) );
INV_X4 inst_5253 ( .ZN(net_681), .A(net_437) );
OAI221_X2 inst_1649 ( .ZN(net_5058), .C2(net_5057), .B2(net_5054), .A(net_4525), .B1(net_2431), .C1(net_1061) );
AOI21_X2 inst_7756 ( .B1(net_6473), .ZN(net_4043), .B2(net_2580), .A(net_2311) );
OAI22_X2 inst_1480 ( .B1(net_4855), .A1(net_4228), .B2(net_4211), .ZN(net_4174), .A2(net_4173) );
CLKBUF_X2 inst_12921 ( .A(net_10816), .Z(net_12883) );
CLKBUF_X2 inst_13594 ( .A(net_13555), .Z(net_13556) );
INV_X2 inst_5815 ( .A(net_1642), .ZN(net_1098) );
INV_X2 inst_5873 ( .ZN(net_414), .A(x977) );
CLKBUF_X2 inst_14121 ( .A(net_14082), .Z(net_14083) );
CLKBUF_X2 inst_10676 ( .A(net_9368), .Z(net_10638) );
CLKBUF_X2 inst_8697 ( .A(net_7962), .Z(net_8659) );
CLKBUF_X2 inst_12359 ( .A(net_10661), .Z(net_12321) );
CLKBUF_X2 inst_10504 ( .A(net_10200), .Z(net_10466) );
DFF_X1 inst_6472 ( .QN(net_6069), .D(net_5587), .CK(net_8104) );
AOI22_X2 inst_7409 ( .B1(net_5939), .A2(net_2838), .ZN(net_2826), .A1(net_876), .B2(net_206) );
SDFF_X2 inst_669 ( .SI(net_7799), .Q(net_6700), .D(net_6700), .SE(net_3871), .CK(net_11105) );
CLKBUF_X2 inst_9214 ( .A(net_8360), .Z(net_9176) );
CLKBUF_X2 inst_13977 ( .A(net_13938), .Z(net_13939) );
CLKBUF_X2 inst_11638 ( .A(net_11366), .Z(net_11600) );
SDFF_X2 inst_664 ( .Q(net_6696), .D(net_6696), .SE(net_3871), .SI(net_3802), .CK(net_8971) );
CLKBUF_X2 inst_10024 ( .A(net_8594), .Z(net_9986) );
CLKBUF_X2 inst_12485 ( .A(net_10978), .Z(net_12447) );
CLKBUF_X2 inst_10486 ( .A(net_10447), .Z(net_10448) );
CLKBUF_X2 inst_8988 ( .A(net_7846), .Z(net_8950) );
CLKBUF_X2 inst_14262 ( .A(net_14223), .Z(net_14224) );
CLKBUF_X2 inst_9911 ( .A(net_9872), .Z(net_9873) );
CLKBUF_X2 inst_10532 ( .A(net_10493), .Z(net_10494) );
OAI21_X2 inst_1918 ( .B1(net_5339), .ZN(net_5146), .A(net_4746), .B2(net_3941) );
CLKBUF_X2 inst_8236 ( .A(net_8197), .Z(net_8198) );
CLKBUF_X2 inst_9466 ( .A(net_9427), .Z(net_9428) );
NAND2_X2 inst_4064 ( .A1(net_6664), .A2(net_1655), .ZN(net_988) );
NAND2_X1 inst_4427 ( .A1(net_7606), .A2(net_2131), .ZN(net_1451) );
CLKBUF_X2 inst_12543 ( .A(net_12504), .Z(net_12505) );
INV_X4 inst_4897 ( .A(net_3902), .ZN(net_3188) );
AOI222_X2 inst_7603 ( .A1(net_7249), .ZN(net_5353), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_343), .C2(net_341) );
INV_X4 inst_4635 ( .ZN(net_4187), .A(net_4036) );
OAI21_X2 inst_1844 ( .B1(net_5353), .ZN(net_5328), .A(net_4368), .B2(net_3853) );
NAND2_X2 inst_3839 ( .A1(net_6831), .A2(net_1521), .ZN(net_1500) );
OAI21_X2 inst_1913 ( .ZN(net_5155), .B1(net_4868), .A(net_4757), .B2(net_3941) );
INV_X4 inst_5209 ( .A(net_598), .ZN(net_489) );
AND2_X2 inst_7862 ( .A2(net_6421), .A1(net_6420), .ZN(net_503) );
OAI21_X2 inst_1990 ( .B1(net_4847), .ZN(net_4839), .A(net_4559), .B2(net_3866) );
NOR2_X2 inst_2368 ( .ZN(net_5268), .A2(net_4620), .A1(net_4465) );
INV_X4 inst_5700 ( .A(net_5936), .ZN(net_5935) );
XNOR2_X2 inst_36 ( .ZN(net_2452), .B(net_2272), .A(net_2271) );
NAND3_X2 inst_2735 ( .ZN(net_2366), .A3(net_1586), .A1(net_1397), .A2(net_1023) );
NAND3_X2 inst_2767 ( .ZN(net_2333), .A3(net_1643), .A1(net_1391), .A2(net_1016) );
NAND2_X2 inst_2934 ( .ZN(net_5513), .A1(net_4987), .A2(net_4986) );
OR2_X4 inst_1370 ( .ZN(net_3973), .A2(net_3737), .A1(net_617) );
NOR2_X2 inst_2512 ( .A2(net_3243), .ZN(net_1162), .A1(net_1161) );
CLKBUF_X2 inst_12770 ( .A(net_9783), .Z(net_12732) );
CLKBUF_X2 inst_12093 ( .A(net_9694), .Z(net_12055) );
CLKBUF_X2 inst_13686 ( .A(net_9026), .Z(net_13648) );
CLKBUF_X2 inst_9039 ( .A(net_9000), .Z(net_9001) );
CLKBUF_X2 inst_11948 ( .A(net_11909), .Z(net_11910) );
CLKBUF_X2 inst_9652 ( .A(net_9549), .Z(net_9614) );
CLKBUF_X2 inst_11447 ( .A(net_11408), .Z(net_11409) );
CLKBUF_X2 inst_13040 ( .A(net_13001), .Z(net_13002) );
CLKBUF_X2 inst_12568 ( .A(net_9356), .Z(net_12530) );
CLKBUF_X2 inst_10721 ( .A(net_10682), .Z(net_10683) );
CLKBUF_X2 inst_7998 ( .A(net_7959), .Z(net_7960) );
NAND2_X2 inst_4124 ( .A2(net_1228), .ZN(net_1167), .A1(net_381) );
CLKBUF_X2 inst_7954 ( .A(net_7886), .Z(net_7916) );
CLKBUF_X2 inst_13078 ( .A(net_7980), .Z(net_13040) );
CLKBUF_X2 inst_13284 ( .A(net_13245), .Z(net_13246) );
NAND2_X2 inst_3067 ( .A1(net_7161), .A2(net_4954), .ZN(net_4938) );
CLKBUF_X2 inst_13023 ( .A(net_12984), .Z(net_12985) );
CLKBUF_X2 inst_9877 ( .A(net_7947), .Z(net_9839) );
CLKBUF_X2 inst_9142 ( .A(net_8675), .Z(net_9104) );
CLKBUF_X2 inst_13737 ( .A(net_13698), .Z(net_13699) );
CLKBUF_X2 inst_10058 ( .A(net_10019), .Z(net_10020) );
INV_X4 inst_5307 ( .A(net_7703), .ZN(net_850) );
INV_X4 inst_5672 ( .A(net_6182), .ZN(net_3495) );
CLKBUF_X2 inst_13188 ( .A(net_13149), .Z(net_13150) );
CLKBUF_X2 inst_10273 ( .A(net_10234), .Z(net_10235) );
SDFF_X2 inst_676 ( .SI(net_7807), .Q(net_6740), .D(net_6740), .SE(net_3815), .CK(net_11153) );
CLKBUF_X2 inst_9755 ( .A(net_9625), .Z(net_9717) );
NAND2_X2 inst_3348 ( .ZN(net_3551), .A1(net_3550), .A2(net_3226) );
AOI21_X2 inst_7700 ( .B1(net_6731), .ZN(net_5905), .B2(net_2581), .A(net_2360) );
CLKBUF_X2 inst_7888 ( .A(net_7839), .Z(net_7850) );
NAND2_X1 inst_4222 ( .ZN(net_4737), .A2(net_3988), .A1(net_2095) );
INV_X4 inst_4848 ( .ZN(net_1061), .A(net_1060) );
DFFR_X2 inst_7044 ( .QN(net_6007), .D(net_3171), .CK(net_12418), .RN(x1822) );
CLKBUF_X2 inst_11906 ( .A(net_11867), .Z(net_11868) );
DFF_X1 inst_6669 ( .QN(net_7263), .D(net_5163), .CK(net_10188) );
OAI21_X2 inst_1684 ( .B2(net_6199), .ZN(net_5847), .B1(net_2699), .A(net_2698) );
INV_X4 inst_4820 ( .A(net_2704), .ZN(net_1093) );
INV_X4 inst_4859 ( .ZN(net_3857), .A(net_682) );
CLKBUF_X2 inst_12588 ( .A(net_12288), .Z(net_12550) );
CLKBUF_X2 inst_10193 ( .A(net_10154), .Z(net_10155) );
OR2_X4 inst_1386 ( .A2(net_2730), .ZN(net_1701), .A1(net_689) );
NOR2_X4 inst_2255 ( .ZN(net_5631), .A1(net_5476), .A2(net_4434) );
INV_X8 inst_4560 ( .A(net_3255), .ZN(net_1228) );
SDFF_X2 inst_1076 ( .SI(net_7216), .Q(net_7216), .D(net_3900), .SE(net_3750), .CK(net_11544) );
SDFF_X2 inst_217 ( .Q(net_6337), .SI(net_6336), .D(net_3651), .SE(net_392), .CK(net_14059) );
DFF_X1 inst_6360 ( .QN(net_6222), .D(net_5824), .CK(net_14123) );
INV_X4 inst_4852 ( .A(net_3849), .ZN(net_1054) );
INV_X2 inst_6078 ( .A(net_6419), .ZN(net_396) );
CLKBUF_X2 inst_13292 ( .A(net_12971), .Z(net_13254) );
CLKBUF_X2 inst_9264 ( .A(net_9225), .Z(net_9226) );
OAI21_X2 inst_2000 ( .B2(net_4518), .ZN(net_4513), .B1(net_4128), .A(net_3692) );
INV_X4 inst_4616 ( .ZN(net_4206), .A(net_4073) );
NAND2_X2 inst_3748 ( .A1(net_7041), .A2(net_1975), .ZN(net_1597) );
CLKBUF_X2 inst_9816 ( .A(net_9753), .Z(net_9778) );
DFF_X1 inst_6732 ( .QN(net_7351), .D(net_5323), .CK(net_10118) );
CLKBUF_X2 inst_10223 ( .A(net_10184), .Z(net_10185) );
NOR3_X2 inst_2213 ( .ZN(net_2223), .A3(net_2222), .A1(net_1669), .A2(net_1058) );
SDFF_X2 inst_1195 ( .SI(net_7077), .Q(net_7077), .D(net_3776), .SE(net_3742), .CK(net_11851) );
DFF_X2 inst_6222 ( .QN(net_6962), .D(net_3726), .CK(net_8533) );
SDFF_X2 inst_672 ( .Q(net_6726), .D(net_6726), .SE(net_3815), .SI(net_3792), .CK(net_11099) );
OAI22_X2 inst_1471 ( .B1(net_4855), .B2(net_4231), .ZN(net_4229), .A1(net_4228), .A2(net_4227) );
CLKBUF_X2 inst_9699 ( .A(net_9660), .Z(net_9661) );
CLKBUF_X2 inst_9610 ( .A(net_8820), .Z(net_9572) );
CLKBUF_X2 inst_12252 ( .A(net_12213), .Z(net_12214) );
NAND2_X2 inst_3826 ( .A1(net_7106), .A2(net_1675), .ZN(net_1518) );
CLKBUF_X2 inst_11829 ( .A(net_8013), .Z(net_11791) );
DFF_X1 inst_6471 ( .QN(net_6068), .D(net_5588), .CK(net_8109) );
AOI222_X2 inst_7523 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_1998), .A1(net_1997), .B1(net_1996), .C1(net_1995) );
OAI22_X2 inst_1525 ( .B1(net_4644), .A1(net_4057), .B2(net_4049), .ZN(net_4046), .A2(net_4045) );
DFF_X1 inst_6839 ( .D(net_2490), .QN(net_264), .CK(net_8027) );
NAND2_X2 inst_3230 ( .ZN(net_4525), .A2(net_4291), .A1(net_2277) );
CLKBUF_X2 inst_11820 ( .A(net_8610), .Z(net_11782) );
NOR2_X4 inst_2248 ( .ZN(net_5638), .A1(net_5484), .A2(net_4450) );
NOR2_X2 inst_2453 ( .ZN(net_2817), .A2(net_2694), .A1(net_1173) );
SDFF_X2 inst_1312 ( .D(net_6383), .SE(net_5800), .SI(net_348), .Q(net_348), .CK(net_14143) );
CLKBUF_X2 inst_9538 ( .A(net_9499), .Z(net_9500) );
NAND2_X2 inst_3281 ( .ZN(net_3684), .A1(net_3683), .A2(net_3231) );
SDFF_X2 inst_703 ( .SI(net_6774), .Q(net_6774), .SE(net_3872), .D(net_3785), .CK(net_8512) );
CLKBUF_X2 inst_11125 ( .A(net_11086), .Z(net_11087) );
CLKBUF_X2 inst_9474 ( .A(net_9435), .Z(net_9436) );
NOR2_X2 inst_2546 ( .A2(net_6962), .ZN(net_1249), .A1(net_451) );
CLKBUF_X2 inst_11112 ( .A(net_11073), .Z(net_11074) );
CLKBUF_X2 inst_9882 ( .A(net_7856), .Z(net_9844) );
INV_X4 inst_4693 ( .ZN(net_4142), .A(net_3324) );
CLKBUF_X2 inst_12504 ( .A(net_8208), .Z(net_12466) );
CLKBUF_X2 inst_10449 ( .A(net_10410), .Z(net_10411) );
CLKBUF_X2 inst_14289 ( .A(net_9494), .Z(net_14251) );
INV_X2 inst_5785 ( .ZN(net_2441), .A(net_2440) );
NAND2_X2 inst_3419 ( .A2(net_5917), .ZN(net_3329), .A1(net_648) );
CLKBUF_X2 inst_12966 ( .A(net_12927), .Z(net_12928) );
SDFF_X2 inst_1067 ( .SI(net_6550), .Q(net_6550), .D(net_3801), .SE(net_3756), .CK(net_11630) );
DFF_X1 inst_6539 ( .QN(net_7471), .D(net_5577), .CK(net_9264) );
CLKBUF_X2 inst_11970 ( .A(net_11931), .Z(net_11932) );
INV_X4 inst_4787 ( .A(net_2805), .ZN(net_1719) );
AOI22_X2 inst_7411 ( .B1(net_5939), .A2(net_2838), .ZN(net_2824), .A1(net_726), .B2(net_198) );
CLKBUF_X2 inst_13749 ( .A(net_13710), .Z(net_13711) );
CLKBUF_X2 inst_9735 ( .A(net_8355), .Z(net_9697) );
CLKBUF_X2 inst_8406 ( .A(net_8367), .Z(net_8368) );
CLKBUF_X2 inst_9231 ( .A(net_9192), .Z(net_9193) );
INV_X4 inst_4951 ( .ZN(net_1302), .A(net_733) );
OAI21_X2 inst_1824 ( .ZN(net_5362), .B1(net_5361), .A(net_4382), .B2(net_3856) );
SDFF_X2 inst_1214 ( .SI(net_7211), .Q(net_7211), .D(net_3786), .SE(net_3750), .CK(net_7900) );
CLKBUF_X2 inst_8121 ( .A(net_8082), .Z(net_8083) );
SDFF_X2 inst_971 ( .Q(net_6451), .D(net_6451), .SE(net_3820), .SI(net_3789), .CK(net_8414) );
OR2_X2 inst_1417 ( .ZN(net_2861), .A2(net_781), .A1(net_524) );
SDFF_X2 inst_1219 ( .SI(net_7210), .Q(net_7210), .D(net_3810), .SE(net_3751), .CK(net_7834) );
CLKBUF_X2 inst_11103 ( .A(net_11064), .Z(net_11065) );
CLKBUF_X2 inst_8018 ( .A(net_7898), .Z(net_7980) );
NAND2_X2 inst_3459 ( .A2(net_5962), .ZN(net_2894), .A1(net_2893) );
CLKBUF_X2 inst_11887 ( .A(net_11848), .Z(net_11849) );
INV_X8 inst_4488 ( .ZN(net_4660), .A(net_3411) );
AOI21_X2 inst_7633 ( .ZN(net_4297), .B2(net_3449), .B1(net_3177), .A(x837) );
NAND2_X2 inst_3335 ( .ZN(net_3576), .A1(net_3575), .A2(net_3226) );
NAND2_X2 inst_3073 ( .A1(net_7152), .A2(net_4954), .ZN(net_4932) );
CLKBUF_X2 inst_12716 ( .A(net_12677), .Z(net_12678) );
CLKBUF_X2 inst_11732 ( .A(net_8459), .Z(net_11694) );
CLKBUF_X2 inst_11741 ( .A(net_9747), .Z(net_11703) );
OAI21_X2 inst_1980 ( .ZN(net_4852), .B1(net_4851), .A(net_4539), .B2(net_3870) );
CLKBUF_X2 inst_10488 ( .A(net_10449), .Z(net_10450) );
INV_X2 inst_5868 ( .A(net_823), .ZN(net_519) );
CLKBUF_X2 inst_9454 ( .A(net_8353), .Z(net_9416) );
CLKBUF_X2 inst_9325 ( .A(net_9286), .Z(net_9287) );
NAND2_X4 inst_2885 ( .ZN(net_3923), .A1(net_3837), .A2(net_421) );
CLKBUF_X2 inst_12628 ( .A(net_12482), .Z(net_12590) );
CLKBUF_X2 inst_10446 ( .A(net_9941), .Z(net_10408) );
NOR2_X4 inst_2221 ( .ZN(net_5677), .A1(net_5553), .A2(net_4514) );
NAND3_X2 inst_2632 ( .ZN(net_5697), .A1(net_5674), .A2(net_5308), .A3(net_4248) );
INV_X4 inst_4795 ( .ZN(net_4801), .A(net_1265) );
CLKBUF_X2 inst_12991 ( .A(net_12952), .Z(net_12953) );
OAI21_X2 inst_2082 ( .B2(net_4415), .ZN(net_4408), .B1(net_4022), .A(net_3500) );
CLKBUF_X2 inst_12469 ( .A(net_12430), .Z(net_12431) );
INV_X2 inst_5842 ( .A(net_1148), .ZN(net_762) );
CLKBUF_X2 inst_10135 ( .A(net_10096), .Z(net_10097) );
NAND2_X2 inst_3286 ( .ZN(net_3674), .A1(net_3673), .A2(net_3231) );
CLKBUF_X2 inst_12907 ( .A(net_12868), .Z(net_12869) );
NAND2_X1 inst_4225 ( .ZN(net_4702), .A2(net_3989), .A1(net_2197) );
INV_X4 inst_5625 ( .A(net_6115), .ZN(net_3699) );
CLKBUF_X2 inst_11371 ( .A(net_10131), .Z(net_11333) );
CLKBUF_X2 inst_11421 ( .A(net_9753), .Z(net_11383) );
CLKBUF_X2 inst_9533 ( .A(net_9494), .Z(net_9495) );
NAND2_X2 inst_4141 ( .A1(net_1153), .ZN(net_914), .A2(net_775) );
CLKBUF_X2 inst_13004 ( .A(net_9703), .Z(net_12966) );
CLKBUF_X2 inst_14293 ( .A(net_14254), .Z(net_14255) );
SDFF_X2 inst_692 ( .Q(net_6757), .D(net_6757), .SE(net_3815), .SI(net_3800), .CK(net_11387) );
INV_X4 inst_4591 ( .ZN(net_4307), .A(net_4212) );
DFF_X1 inst_6800 ( .D(net_3934), .CK(net_12829), .Q(x476) );
DFF_X1 inst_6897 ( .D(net_2521), .QN(net_177), .CK(net_9857) );
OAI22_X2 inst_1517 ( .B1(net_4644), .ZN(net_4063), .A2(net_4062), .B2(net_4061), .A1(net_4057) );
INV_X4 inst_5318 ( .A(net_7255), .ZN(net_2005) );
CLKBUF_X2 inst_10529 ( .A(net_10490), .Z(net_10491) );
XNOR2_X2 inst_70 ( .ZN(net_2484), .A(net_1268), .B(net_526) );
INV_X4 inst_5480 ( .A(net_7555), .ZN(net_2136) );
DFF_X1 inst_6915 ( .D(net_2392), .Q(net_243), .CK(net_13044) );
AOI222_X2 inst_7587 ( .A1(net_7540), .ZN(net_5206), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_372), .C2(net_370) );
AOI21_X2 inst_7672 ( .B1(net_7005), .ZN(net_4211), .A(net_2468), .B2(net_1100) );
CLKBUF_X2 inst_12493 ( .A(net_12454), .Z(net_12455) );
CLKBUF_X2 inst_9865 ( .A(net_7884), .Z(net_9827) );
CLKBUF_X2 inst_9162 ( .A(net_9123), .Z(net_9124) );
CLKBUF_X2 inst_14161 ( .A(net_8838), .Z(net_14123) );
CLKBUF_X2 inst_11290 ( .A(net_11251), .Z(net_11252) );
SDFF_X2 inst_188 ( .Q(net_6266), .SI(net_6265), .D(net_3481), .SE(net_392), .CK(net_13473) );
INV_X8 inst_4528 ( .ZN(net_3755), .A(net_3113) );
CLKBUF_X2 inst_13534 ( .A(net_9427), .Z(net_13496) );
NAND2_X2 inst_3768 ( .A1(net_7163), .A2(net_1637), .ZN(net_1577) );
INV_X2 inst_6028 ( .A(net_7505), .ZN(net_2095) );
INV_X2 inst_6093 ( .A(net_7785), .ZN(net_395) );
NAND2_X2 inst_4207 ( .A2(net_6031), .A1(net_6030), .ZN(net_3234) );
CLKBUF_X2 inst_9058 ( .A(net_9019), .Z(net_9020) );
CLKBUF_X2 inst_11308 ( .A(net_11269), .Z(net_11270) );
NAND2_X2 inst_3011 ( .A1(net_6855), .A2(net_5004), .ZN(net_4998) );
DFF_X2 inst_6218 ( .QN(net_7381), .D(net_3832), .CK(net_12776) );
CLKBUF_X2 inst_13306 ( .A(net_9588), .Z(net_13268) );
NAND2_X4 inst_2848 ( .ZN(net_5475), .A1(net_4919), .A2(net_4918) );
CLKBUF_X2 inst_12686 ( .A(net_12647), .Z(net_12648) );
INV_X4 inst_4826 ( .ZN(net_1085), .A(net_1084) );
DFF_X1 inst_6695 ( .QN(net_7293), .D(net_5380), .CK(net_12713) );
OAI22_X2 inst_1537 ( .B1(net_4637), .A1(net_4030), .B2(net_4024), .ZN(net_4021), .A2(net_4020) );
OAI21_X2 inst_2041 ( .B1(net_4617), .B2(net_4476), .ZN(net_4462), .A(net_3580) );
CLKBUF_X2 inst_13866 ( .A(net_11504), .Z(net_13828) );
DFF_X2 inst_6323 ( .QN(net_7824), .CK(net_8246), .D(x1345) );
INV_X4 inst_5235 ( .A(net_851), .ZN(net_456) );
NAND2_X2 inst_3593 ( .ZN(net_2407), .A2(net_1882), .A1(net_1478) );
CLKBUF_X2 inst_8529 ( .A(net_8490), .Z(net_8491) );
INV_X4 inst_4589 ( .ZN(net_4313), .A(net_4224) );
NAND2_X2 inst_3176 ( .ZN(net_4757), .A2(net_3941), .A1(net_2039) );
AOI222_X2 inst_7509 ( .B1(net_7366), .C1(net_7302), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2036), .A1(net_2035) );
DFF_X1 inst_6768 ( .QN(net_6127), .D(net_4661), .CK(net_8982) );
CLKBUF_X2 inst_11550 ( .A(net_11495), .Z(net_11512) );
NAND2_X2 inst_3325 ( .ZN(net_3596), .A1(net_3595), .A2(net_3228) );
CLKBUF_X2 inst_13393 ( .A(net_13354), .Z(net_13355) );
CLKBUF_X2 inst_11145 ( .A(net_11106), .Z(net_11107) );
CLKBUF_X2 inst_11085 ( .A(net_9197), .Z(net_11047) );
CLKBUF_X2 inst_9083 ( .A(net_9044), .Z(net_9045) );
CLKBUF_X2 inst_13991 ( .A(net_13952), .Z(net_13953) );
CLKBUF_X2 inst_13889 ( .A(net_13850), .Z(net_13851) );
CLKBUF_X2 inst_12655 ( .A(net_12616), .Z(net_12617) );
NAND2_X2 inst_4168 ( .ZN(net_925), .A2(net_593), .A1(net_495) );
SDFF_X2 inst_195 ( .QN(net_6319), .SI(net_6318), .D(net_3687), .SE(net_392), .CK(net_13596) );
CLKBUF_X2 inst_11835 ( .A(net_11796), .Z(net_11797) );
CLKBUF_X2 inst_12839 ( .A(net_12800), .Z(net_12801) );
OAI21_X2 inst_1987 ( .B1(net_4853), .ZN(net_4842), .A(net_4562), .B2(net_3866) );
CLKBUF_X2 inst_13730 ( .A(net_13691), .Z(net_13692) );
CLKBUF_X2 inst_10821 ( .A(net_9480), .Z(net_10783) );
CLKBUF_X2 inst_13418 ( .A(net_13379), .Z(net_13380) );
SDFF_X2 inst_1150 ( .SI(net_6811), .Q(net_6811), .D(net_3900), .SE(net_3722), .CK(net_8342) );
AOI21_X2 inst_7685 ( .B1(net_6591), .ZN(net_4405), .B2(net_2583), .A(net_2295) );
CLKBUF_X2 inst_14372 ( .A(net_14333), .Z(net_14334) );
INV_X4 inst_4914 ( .A(net_3802), .ZN(net_3270) );
CLKBUF_X2 inst_11355 ( .A(net_11316), .Z(net_11317) );
CLKBUF_X2 inst_11020 ( .A(net_10981), .Z(net_10982) );
INV_X4 inst_5605 ( .A(net_6077), .ZN(net_3477) );
DFFR_X2 inst_7070 ( .QN(net_6033), .D(net_3060), .CK(net_9998), .RN(x1822) );
DFFR_X2 inst_7106 ( .D(net_1949), .QN(net_127), .CK(net_12634), .RN(x1822) );
INV_X4 inst_4780 ( .ZN(net_2634), .A(net_1663) );
CLKBUF_X2 inst_12981 ( .A(net_12942), .Z(net_12943) );
CLKBUF_X2 inst_11770 ( .A(net_11731), .Z(net_11732) );
INV_X4 inst_4658 ( .ZN(net_5885), .A(net_3928) );
INV_X2 inst_5916 ( .A(net_7514), .ZN(net_2218) );
CLKBUF_X2 inst_8715 ( .A(net_8676), .Z(net_8677) );
OAI22_X2 inst_1589 ( .B2(net_3200), .A2(net_3196), .ZN(net_3175), .A1(net_3174), .B1(net_466) );
CLKBUF_X2 inst_11994 ( .A(net_8227), .Z(net_11956) );
CLKBUF_X2 inst_8926 ( .A(net_8075), .Z(net_8888) );
INV_X8 inst_4535 ( .A(net_6054), .ZN(net_5800) );
CLKBUF_X2 inst_14114 ( .A(net_14075), .Z(net_14076) );
INV_X4 inst_5607 ( .A(net_6043), .ZN(net_547) );
CLKBUF_X2 inst_14095 ( .A(net_14056), .Z(net_14057) );
INV_X8 inst_4499 ( .ZN(net_3851), .A(net_3264) );
CLKBUF_X2 inst_12852 ( .A(net_12813), .Z(net_12814) );
CLKBUF_X2 inst_10979 ( .A(net_10940), .Z(net_10941) );
DFF_X1 inst_6825 ( .D(net_2998), .CK(net_13405), .Q(x187) );
CLKBUF_X2 inst_8704 ( .A(net_7931), .Z(net_8666) );
SDFF_X2 inst_335 ( .SI(net_7494), .Q(net_7494), .D(net_5095), .SE(net_3989), .CK(net_12522) );
CLKBUF_X2 inst_12783 ( .A(net_12744), .Z(net_12745) );
CLKBUF_X2 inst_12827 ( .A(net_10765), .Z(net_12789) );
INV_X4 inst_5508 ( .A(net_6404), .ZN(net_871) );
CLKBUF_X2 inst_12661 ( .A(net_12622), .Z(net_12623) );
CLKBUF_X2 inst_14406 ( .A(net_14367), .Z(net_14368) );
CLKBUF_X2 inst_8611 ( .A(net_8572), .Z(net_8573) );
SDFF_X2 inst_658 ( .Q(net_6716), .D(net_6716), .SE(net_3871), .SI(net_3804), .CK(net_10927) );
DFF_X2 inst_6190 ( .QN(net_6959), .D(net_5078), .CK(net_11365) );
DFF_X1 inst_6862 ( .D(net_2544), .Q(net_199), .CK(net_9229) );
CLKBUF_X2 inst_8420 ( .A(net_8135), .Z(net_8382) );
AOI21_X2 inst_7779 ( .B1(net_7144), .ZN(net_4074), .B2(net_2582), .A(net_2322) );
CLKBUF_X2 inst_12192 ( .A(net_12153), .Z(net_12154) );
CLKBUF_X2 inst_9336 ( .A(net_9297), .Z(net_9298) );
INV_X8 inst_4520 ( .ZN(net_3729), .A(net_3117) );
CLKBUF_X2 inst_11562 ( .A(net_11523), .Z(net_11524) );
CLKBUF_X2 inst_14045 ( .A(net_14006), .Z(net_14007) );
CLKBUF_X2 inst_14276 ( .A(net_14237), .Z(net_14238) );
SDFF_X2 inst_438 ( .Q(net_7392), .D(net_7392), .SE(net_3994), .SI(net_357), .CK(net_12432) );
CLKBUF_X2 inst_13311 ( .A(net_13272), .Z(net_13273) );
AOI22_X2 inst_7326 ( .ZN(net_3424), .A2(net_3423), .B2(net_3422), .A1(net_1305), .B1(net_900) );
DFF_X1 inst_6351 ( .QN(net_6207), .D(net_5833), .CK(net_13712) );
CLKBUF_X2 inst_10769 ( .A(net_10730), .Z(net_10731) );
CLKBUF_X2 inst_9626 ( .A(net_9587), .Z(net_9588) );
CLKBUF_X2 inst_14336 ( .A(net_14297), .Z(net_14298) );
CLKBUF_X2 inst_9692 ( .A(net_9653), .Z(net_9654) );
CLKBUF_X2 inst_11391 ( .A(net_10898), .Z(net_11353) );
SDFF_X2 inst_324 ( .SI(net_7489), .Q(net_7489), .D(net_5103), .SE(net_3989), .CK(net_12446) );
CLKBUF_X2 inst_11640 ( .A(net_11601), .Z(net_11602) );
NAND2_X2 inst_3550 ( .ZN(net_2517), .A2(net_2060), .A1(net_1769) );
INV_X2 inst_6046 ( .A(net_7666), .ZN(net_1860) );
NAND2_X2 inst_4083 ( .A1(net_6524), .A2(net_1645), .ZN(net_969) );
CLKBUF_X2 inst_13581 ( .A(net_11134), .Z(net_13543) );
XNOR2_X2 inst_43 ( .B(net_7095), .ZN(net_2447), .A(net_1241) );
OAI21_X2 inst_2128 ( .ZN(net_2998), .B1(net_2997), .A(net_2874), .B2(net_2624) );
INV_X2 inst_5936 ( .A(net_7330), .ZN(net_1766) );
OAI21_X2 inst_1707 ( .B2(net_5911), .ZN(net_5587), .A(net_5154), .B1(net_4057) );
DFF_X1 inst_6715 ( .QN(net_7331), .D(net_5350), .CK(net_9873) );
CLKBUF_X2 inst_10452 ( .A(net_10413), .Z(net_10414) );
CLKBUF_X2 inst_8115 ( .A(net_7927), .Z(net_8077) );
SDFF_X2 inst_375 ( .SI(net_7668), .Q(net_7668), .D(net_4792), .SE(net_3866), .CK(net_13244) );
CLKBUF_X2 inst_11241 ( .A(net_9700), .Z(net_11203) );
CLKBUF_X2 inst_9959 ( .A(net_9920), .Z(net_9921) );
CLKBUF_X2 inst_8606 ( .A(net_8567), .Z(net_8568) );
NAND2_X2 inst_3490 ( .ZN(net_2651), .A1(net_2650), .A2(net_2649) );
AOI22_X2 inst_7384 ( .A2(net_5916), .B2(net_2957), .ZN(net_2936), .B1(net_2650), .A1(net_855) );
DFFR_X2 inst_7039 ( .QN(net_5999), .D(net_3141), .CK(net_10022), .RN(x1822) );
CLKBUF_X2 inst_10933 ( .A(net_10332), .Z(net_10895) );
CLKBUF_X2 inst_10086 ( .A(net_8363), .Z(net_10048) );
SDFF_X2 inst_285 ( .D(net_6396), .SE(net_5801), .SI(net_341), .Q(net_341), .CK(net_14332) );
OAI21_X2 inst_1830 ( .ZN(net_5350), .B1(net_5349), .A(net_4388), .B2(net_3856) );
CLKBUF_X2 inst_9887 ( .A(net_9025), .Z(net_9849) );
CLKBUF_X2 inst_11780 ( .A(net_8791), .Z(net_11742) );
CLKBUF_X2 inst_11385 ( .A(net_11346), .Z(net_11347) );
CLKBUF_X2 inst_9313 ( .A(net_9274), .Z(net_9275) );
INV_X4 inst_5563 ( .A(net_7430), .ZN(net_1981) );
CLKBUF_X2 inst_8289 ( .A(net_8250), .Z(net_8251) );
OAI22_X2 inst_1563 ( .B2(net_3405), .A2(net_3360), .ZN(net_3342), .A1(net_3291), .B1(net_513) );
DFF_X1 inst_6363 ( .Q(net_6299), .D(net_5821), .CK(net_13802) );
CLKBUF_X2 inst_10833 ( .A(net_10794), .Z(net_10795) );
CLKBUF_X2 inst_11402 ( .A(net_11363), .Z(net_11364) );
NAND2_X1 inst_4455 ( .A2(net_1256), .ZN(net_1120), .A1(net_1119) );
CLKBUF_X2 inst_7911 ( .A(net_7872), .Z(net_7873) );
NAND2_X2 inst_3242 ( .A1(net_7769), .ZN(net_4164), .A2(net_4001) );
AOI22_X2 inst_7398 ( .A1(net_6024), .A2(net_3105), .B1(net_2970), .ZN(net_2842), .B2(net_261) );
CLKBUF_X2 inst_10638 ( .A(net_10599), .Z(net_10600) );
CLKBUF_X2 inst_7907 ( .A(net_7868), .Z(net_7869) );
CLKBUF_X2 inst_9895 ( .A(net_9856), .Z(net_9857) );
SDFF_X2 inst_929 ( .Q(net_7139), .D(net_7139), .SE(net_3903), .SI(net_3814), .CK(net_13345) );
SDFF_X2 inst_982 ( .Q(net_6467), .D(net_6467), .SE(net_3904), .SI(net_3813), .CK(net_11257) );
NAND2_X2 inst_3138 ( .ZN(net_4825), .A2(net_4153), .A1(net_1989) );
OR2_X4 inst_1397 ( .A2(net_6554), .A1(net_6553), .ZN(net_490) );
CLKBUF_X2 inst_10864 ( .A(net_10809), .Z(net_10826) );
SDFF_X2 inst_299 ( .SI(net_7486), .Q(net_7486), .D(net_5107), .SE(net_3989), .CK(net_9805) );
CLKBUF_X2 inst_13871 ( .A(net_9188), .Z(net_13833) );
CLKBUF_X2 inst_10567 ( .A(net_10528), .Z(net_10529) );
AOI21_X2 inst_7656 ( .B2(net_3439), .ZN(net_3389), .A(net_3217), .B1(net_748) );
OAI21_X2 inst_1798 ( .ZN(net_5392), .A(net_4719), .B2(net_3986), .B1(net_1164) );
NAND2_X2 inst_2927 ( .ZN(net_5527), .A1(net_5001), .A2(net_5000) );
CLKBUF_X2 inst_13115 ( .A(net_13076), .Z(net_13077) );
NAND2_X2 inst_3303 ( .ZN(net_3640), .A1(net_3639), .A2(net_3229) );
CLKBUF_X2 inst_10336 ( .A(net_9522), .Z(net_10298) );
DFF_X2 inst_6181 ( .QN(net_7228), .D(net_5451), .CK(net_9379) );
CLKBUF_X2 inst_12938 ( .A(net_8709), .Z(net_12900) );
INV_X2 inst_5853 ( .ZN(net_672), .A(net_671) );
CLKBUF_X2 inst_10383 ( .A(net_10344), .Z(net_10345) );
CLKBUF_X2 inst_8727 ( .A(net_7875), .Z(net_8689) );
NAND3_X2 inst_2760 ( .ZN(net_2341), .A3(net_1573), .A1(net_1475), .A2(net_975) );
OAI21_X2 inst_1938 ( .B1(net_5545), .ZN(net_5106), .A(net_4739), .B2(net_3988) );
DFF_X1 inst_6478 ( .QN(net_6091), .D(net_5581), .CK(net_9385) );
DFF_X1 inst_6452 ( .QN(net_6103), .D(net_5718), .CK(net_9211) );
CLKBUF_X2 inst_11870 ( .A(net_11831), .Z(net_11832) );
CLKBUF_X2 inst_9435 ( .A(net_9396), .Z(net_9397) );
DFFR_X2 inst_7098 ( .D(net_1945), .QN(net_125), .CK(net_12847), .RN(x1822) );
DFF_X1 inst_6888 ( .D(net_2528), .Q(net_231), .CK(net_12415) );
OAI21_X2 inst_2095 ( .B2(net_4445), .ZN(net_4321), .B1(net_4080), .A(net_3527) );
DFF_X2 inst_6288 ( .D(net_2564), .CK(net_12970), .Q(x38) );
DFFR_X2 inst_7030 ( .QN(net_5995), .D(net_3130), .CK(net_10024), .RN(x1822) );
INV_X4 inst_5129 ( .ZN(net_787), .A(net_586) );
CLKBUF_X2 inst_13524 ( .A(net_13227), .Z(net_13486) );
INV_X2 inst_5794 ( .A(net_2417), .ZN(net_2234) );
CLKBUF_X2 inst_14103 ( .A(net_14064), .Z(net_14065) );
CLKBUF_X2 inst_8896 ( .A(net_8591), .Z(net_8858) );
CLKBUF_X2 inst_10656 ( .A(net_10617), .Z(net_10618) );
INV_X4 inst_4995 ( .A(net_7821), .ZN(net_3793) );
INV_X4 inst_5652 ( .A(net_6163), .ZN(net_3595) );
NAND2_X2 inst_3260 ( .A2(net_3858), .ZN(net_3856), .A1(net_3833) );
CLKBUF_X2 inst_8262 ( .A(net_8223), .Z(net_8224) );
NAND2_X2 inst_3158 ( .ZN(net_4775), .A2(net_3941), .A1(net_2031) );
NAND2_X2 inst_4190 ( .A2(net_6043), .ZN(net_1263), .A1(net_578) );
CLKBUF_X2 inst_13894 ( .A(net_13855), .Z(net_13856) );
CLKBUF_X2 inst_11248 ( .A(net_9651), .Z(net_11210) );
INV_X4 inst_5387 ( .A(net_6119), .ZN(net_3693) );
CLKBUF_X2 inst_14067 ( .A(net_11274), .Z(net_14029) );
CLKBUF_X2 inst_11813 ( .A(net_11774), .Z(net_11775) );
SDFF_X2 inst_683 ( .Q(net_6748), .D(net_6748), .SE(net_3815), .SI(net_3804), .CK(net_10918) );
INV_X4 inst_5631 ( .A(net_6095), .ZN(net_3513) );
NOR3_X2 inst_2186 ( .ZN(net_5944), .A2(net_3956), .A3(net_3885), .A1(net_3774) );
NAND2_X2 inst_3269 ( .ZN(net_3708), .A1(net_3707), .A2(net_3225) );
CLKBUF_X2 inst_9094 ( .A(net_9055), .Z(net_9056) );
OAI21_X2 inst_1944 ( .B1(net_5235), .ZN(net_5081), .A(net_4733), .B2(net_3986) );
CLKBUF_X2 inst_9079 ( .A(net_9040), .Z(net_9041) );
SDFF_X2 inst_210 ( .Q(net_6304), .SI(net_6303), .D(net_3679), .SE(net_392), .CK(net_13554) );
CLKBUF_X2 inst_13763 ( .A(net_13724), .Z(net_13725) );
CLKBUF_X2 inst_9411 ( .A(net_9372), .Z(net_9373) );
CLKBUF_X2 inst_11675 ( .A(net_11636), .Z(net_11637) );
NAND2_X2 inst_3101 ( .A1(net_6613), .ZN(net_4902), .A2(net_4899) );
CLKBUF_X2 inst_8720 ( .A(net_8681), .Z(net_8682) );
INV_X4 inst_4942 ( .ZN(net_1138), .A(net_747) );
CLKBUF_X2 inst_12103 ( .A(net_12064), .Z(net_12065) );
INV_X2 inst_5893 ( .A(net_7444), .ZN(net_1494) );
NAND2_X2 inst_3881 ( .A1(net_7459), .A2(net_1696), .ZN(net_1438) );
INV_X4 inst_5331 ( .A(net_7560), .ZN(net_1841) );
CLKBUF_X2 inst_8164 ( .A(net_8125), .Z(net_8126) );
DFFR_X1 inst_7123 ( .Q(net_6047), .D(net_4794), .CK(net_12573), .RN(x1822) );
INV_X4 inst_4778 ( .A(net_3050), .ZN(net_1723) );
SDFF_X2 inst_1294 ( .SI(net_7764), .Q(net_7764), .SE(net_5919), .D(net_2750), .CK(net_12283) );
AOI21_X2 inst_7663 ( .B2(net_5926), .ZN(net_3314), .A(net_3313), .B1(net_1831) );
OAI21_X2 inst_1712 ( .ZN(net_5582), .A(net_5127), .B2(net_4418), .B1(net_4030) );
INV_X4 inst_5325 ( .A(net_6137), .ZN(net_3659) );
INV_X4 inst_5238 ( .ZN(net_453), .A(net_452) );
SDFF_X2 inst_747 ( .Q(net_6837), .D(net_6837), .SE(net_3893), .SI(net_3814), .CK(net_11809) );
NAND2_X2 inst_3108 ( .A1(net_6584), .A2(net_4897), .ZN(net_4893) );
INV_X4 inst_4576 ( .ZN(net_5782), .A(net_5781) );
CLKBUF_X2 inst_9070 ( .A(net_8760), .Z(net_9032) );
DFF_X1 inst_6685 ( .QN(net_7273), .D(net_5119), .CK(net_9963) );
CLKBUF_X2 inst_12626 ( .A(net_12587), .Z(net_12588) );
NAND2_X4 inst_2853 ( .ZN(net_5470), .A1(net_4909), .A2(net_4908) );
NAND2_X2 inst_3806 ( .A1(net_6495), .A2(net_1642), .ZN(net_1539) );
INV_X8 inst_4486 ( .ZN(net_4228), .A(net_3715) );
CLKBUF_X2 inst_12893 ( .A(net_12854), .Z(net_12855) );
AOI22_X2 inst_7267 ( .B1(net_6946), .A1(net_6914), .A2(net_5298), .B2(net_5297), .ZN(net_5283) );
CLKBUF_X2 inst_10291 ( .A(net_10252), .Z(net_10253) );
CLKBUF_X2 inst_11362 ( .A(net_11323), .Z(net_11324) );
DFF_X1 inst_6546 ( .QN(net_7289), .D(net_5369), .CK(net_12279) );
CLKBUF_X2 inst_12166 ( .A(net_8071), .Z(net_12128) );
NAND3_X2 inst_2775 ( .ZN(net_2325), .A3(net_1575), .A1(net_1417), .A2(net_993) );
AND2_X2 inst_7855 ( .ZN(net_3037), .A1(net_2941), .A2(net_2822) );
CLKBUF_X2 inst_8553 ( .A(net_8514), .Z(net_8515) );
INV_X4 inst_5589 ( .A(net_6092), .ZN(net_3479) );
CLKBUF_X2 inst_12334 ( .A(net_8378), .Z(net_12296) );
CLKBUF_X2 inst_11658 ( .A(net_9220), .Z(net_11620) );
SDFF_X2 inst_305 ( .SI(net_7526), .Q(net_7526), .D(net_5095), .SE(net_3988), .CK(net_12451) );
DFF_X1 inst_6795 ( .D(net_3945), .CK(net_12836), .Q(x522) );
CLKBUF_X2 inst_10853 ( .A(net_10814), .Z(net_10815) );
CLKBUF_X2 inst_13516 ( .A(net_8152), .Z(net_13478) );
OAI22_X2 inst_1595 ( .B2(net_3200), .A2(net_3187), .ZN(net_3143), .A1(net_3142), .B1(net_475) );
CLKBUF_X2 inst_7881 ( .A(net_7842), .Z(net_7843) );
INV_X4 inst_5651 ( .A(net_6177), .ZN(net_3491) );
DFF_X2 inst_6291 ( .D(net_2224), .QN(net_392), .CK(net_14344) );
CLKBUF_X2 inst_7867 ( .A(net_7828), .Z(net_7829) );
CLKBUF_X2 inst_12476 ( .A(net_12437), .Z(net_12438) );
INV_X2 inst_5740 ( .ZN(net_3725), .A(net_3427) );
CLKBUF_X2 inst_13578 ( .A(net_13539), .Z(net_13540) );
CLKBUF_X2 inst_10926 ( .A(net_10887), .Z(net_10888) );
CLKBUF_X2 inst_10602 ( .A(net_10563), .Z(net_10564) );
CLKBUF_X2 inst_12319 ( .A(net_12280), .Z(net_12281) );
CLKBUF_X2 inst_10993 ( .A(net_9970), .Z(net_10955) );
DFF_X2 inst_6227 ( .QN(net_6828), .D(net_3720), .CK(net_10785) );
CLKBUF_X2 inst_13489 ( .A(net_13450), .Z(net_13451) );
CLKBUF_X2 inst_13069 ( .A(net_13030), .Z(net_13031) );
DFF_X1 inst_6585 ( .QN(net_7555), .D(net_5065), .CK(net_12271) );
CLKBUF_X2 inst_8079 ( .A(net_8040), .Z(net_8041) );
AOI21_X2 inst_7774 ( .B1(net_6601), .ZN(net_4033), .B2(net_2583), .A(net_2292) );
CLKBUF_X2 inst_11620 ( .A(net_11581), .Z(net_11582) );
CLKBUF_X2 inst_11605 ( .A(net_11566), .Z(net_11567) );
SDFF_X2 inst_963 ( .Q(net_6441), .D(net_6441), .SE(net_3820), .SI(net_3808), .CK(net_8857) );
SDFF_X2 inst_907 ( .Q(net_7143), .D(net_7143), .SE(net_3903), .SI(net_3812), .CK(net_7858) );
SDFF_X2 inst_922 ( .Q(net_7160), .D(net_7160), .SE(net_3903), .SI(net_3821), .CK(net_8078) );
OAI22_X2 inst_1614 ( .A1(net_3287), .A2(net_3087), .B2(net_3084), .ZN(net_3058), .B1(net_877) );
CLKBUF_X2 inst_11323 ( .A(net_11284), .Z(net_11285) );
CLKBUF_X2 inst_8225 ( .A(net_8186), .Z(net_8187) );
OAI22_X2 inst_1502 ( .B1(net_4660), .A1(net_4105), .B2(net_4097), .ZN(net_4094), .A2(net_4093) );
CLKBUF_X2 inst_8773 ( .A(net_8734), .Z(net_8735) );
INV_X4 inst_5436 ( .A(net_6019), .ZN(net_552) );
CLKBUF_X2 inst_12435 ( .A(net_12396), .Z(net_12397) );
CLKBUF_X2 inst_10693 ( .A(net_10654), .Z(net_10655) );
CLKBUF_X2 inst_9475 ( .A(net_9217), .Z(net_9437) );
CLKBUF_X2 inst_14418 ( .A(net_14379), .Z(net_14380) );
INV_X2 inst_6115 ( .ZN(net_5930), .A(net_5925) );
CLKBUF_X2 inst_8516 ( .A(net_8456), .Z(net_8478) );
NAND2_X2 inst_4091 ( .A1(net_7196), .A2(net_1648), .ZN(net_961) );
CLKBUF_X2 inst_12621 ( .A(net_12582), .Z(net_12583) );
AOI222_X2 inst_7602 ( .A1(net_7399), .ZN(net_5438), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_362), .C2(net_360) );
DFFR_X2 inst_6989 ( .QN(net_7699), .D(net_3343), .CK(net_12881), .RN(x1822) );
CLKBUF_X2 inst_13231 ( .A(net_13192), .Z(net_13193) );
NAND2_X2 inst_3907 ( .A1(net_6845), .A2(net_1521), .ZN(net_1403) );
DFF_X1 inst_6807 ( .D(net_3460), .CK(net_8576), .Q(x420) );
CLKBUF_X2 inst_9619 ( .A(net_8932), .Z(net_9581) );
OAI22_X2 inst_1568 ( .A2(net_3297), .B2(net_3286), .ZN(net_3283), .A1(net_3282), .B1(net_729) );
CLKBUF_X2 inst_11439 ( .A(net_11400), .Z(net_11401) );
DFF_X2 inst_6177 ( .Q(net_6397), .D(net_6396), .CK(net_13851) );
CLKBUF_X2 inst_12383 ( .A(net_12344), .Z(net_12345) );
CLKBUF_X2 inst_8487 ( .A(net_8448), .Z(net_8449) );
CLKBUF_X2 inst_12223 ( .A(net_11228), .Z(net_12185) );
CLKBUF_X2 inst_9258 ( .A(net_9219), .Z(net_9220) );
SDFF_X2 inst_873 ( .SI(net_7059), .Q(net_7059), .D(net_3800), .SE(net_3777), .CK(net_10982) );
NAND2_X2 inst_3366 ( .ZN(net_3514), .A1(net_3513), .A2(net_3223) );
NAND2_X2 inst_3692 ( .A2(net_1798), .ZN(net_1752), .A1(net_1751) );
SDFF_X2 inst_653 ( .Q(net_6710), .D(net_6710), .SE(net_3871), .SI(net_3786), .CK(net_8523) );
DFF_X1 inst_6454 ( .QN(net_6093), .D(net_5716), .CK(net_9204) );
CLKBUF_X2 inst_13439 ( .A(net_13400), .Z(net_13401) );
CLKBUF_X2 inst_10164 ( .A(net_10125), .Z(net_10126) );
CLKBUF_X2 inst_10022 ( .A(net_9983), .Z(net_9984) );
CLKBUF_X2 inst_8563 ( .A(net_8524), .Z(net_8525) );
CLKBUF_X2 inst_8304 ( .A(net_8265), .Z(net_8266) );
CLKBUF_X2 inst_10282 ( .A(net_10243), .Z(net_10244) );
NAND2_X2 inst_3767 ( .A1(net_7043), .A2(net_1975), .ZN(net_1578) );
OAI21_X2 inst_1746 ( .ZN(net_5523), .A(net_4821), .B2(net_4153), .B1(net_1178) );
CLKBUF_X2 inst_11099 ( .A(net_11060), .Z(net_11061) );
CLKBUF_X2 inst_8839 ( .A(net_8800), .Z(net_8801) );
CLKBUF_X2 inst_8679 ( .A(net_8640), .Z(net_8641) );
NAND2_X1 inst_4431 ( .A2(net_2131), .ZN(net_1429), .A1(net_1428) );
NAND2_X2 inst_3371 ( .ZN(net_3504), .A1(net_3503), .A2(net_3223) );
NAND2_X2 inst_3052 ( .A1(net_7153), .ZN(net_4955), .A2(net_4954) );
CLKBUF_X2 inst_13406 ( .A(net_13367), .Z(net_13368) );
CLKBUF_X2 inst_8233 ( .A(net_8194), .Z(net_8195) );
DFFR_X2 inst_6982 ( .QN(net_6049), .D(net_3443), .CK(net_10529), .RN(x1822) );
NAND2_X2 inst_3649 ( .A1(net_7070), .ZN(net_1814), .A2(net_791) );
CLKBUF_X2 inst_13548 ( .A(net_11631), .Z(net_13510) );
NAND2_X2 inst_2907 ( .ZN(net_5791), .A2(net_5774), .A1(net_404) );
INV_X4 inst_4609 ( .ZN(net_4235), .A(net_4088) );
NAND2_X2 inst_4072 ( .A1(net_6805), .A2(net_1651), .ZN(net_980) );
DFF_X1 inst_6526 ( .QN(net_7442), .D(net_5425), .CK(net_10086) );
CLKBUF_X2 inst_11843 ( .A(net_11213), .Z(net_11805) );
NAND3_X2 inst_2656 ( .ZN(net_3944), .A3(net_3390), .A2(net_2951), .A1(net_2826) );
INV_X2 inst_5901 ( .A(net_7599), .ZN(net_1455) );
NAND2_X2 inst_3000 ( .A1(net_6715), .A2(net_5031), .ZN(net_5011) );
CLKBUF_X2 inst_9668 ( .A(net_9629), .Z(net_9630) );
SDFF_X2 inst_1163 ( .SI(net_6797), .Q(net_6797), .D(net_3883), .SE(net_3729), .CK(net_11288) );
CLKBUF_X2 inst_10641 ( .A(net_10602), .Z(net_10603) );
CLKBUF_X2 inst_8282 ( .A(net_8243), .Z(net_8244) );
OAI22_X2 inst_1604 ( .A1(net_3275), .B2(net_3200), .A2(net_3193), .ZN(net_3130), .B1(net_1724) );
CLKBUF_X2 inst_8301 ( .A(net_8243), .Z(net_8263) );
NAND2_X2 inst_3239 ( .ZN(net_4273), .A1(net_4272), .A2(net_1624) );
NOR2_X2 inst_2314 ( .A2(net_6200), .A1(net_5843), .ZN(net_5827) );
CLKBUF_X2 inst_9426 ( .A(net_9387), .Z(net_9388) );
CLKBUF_X2 inst_12885 ( .A(net_12846), .Z(net_12847) );
CLKBUF_X2 inst_13854 ( .A(net_11922), .Z(net_13816) );
NAND3_X2 inst_2812 ( .ZN(net_2286), .A3(net_1571), .A1(net_1354), .A2(net_964) );
CLKBUF_X2 inst_14441 ( .A(net_14402), .Z(net_14403) );
INV_X4 inst_4743 ( .A(net_2753), .ZN(net_2750) );
CLKBUF_X2 inst_8592 ( .A(net_8553), .Z(net_8554) );
NAND2_X2 inst_3197 ( .ZN(net_4729), .A2(net_3986), .A1(net_1898) );
INV_X4 inst_4651 ( .ZN(net_4629), .A(net_4280) );
CLKBUF_X2 inst_10126 ( .A(net_10087), .Z(net_10088) );
XNOR2_X2 inst_7 ( .A(net_4151), .ZN(net_3829), .B(net_759) );
CLKBUF_X2 inst_13640 ( .A(net_13601), .Z(net_13602) );
CLKBUF_X2 inst_9672 ( .A(net_9633), .Z(net_9634) );
NAND2_X2 inst_3450 ( .A2(net_5925), .ZN(net_2922), .A1(net_1215) );
CLKBUF_X2 inst_8006 ( .A(net_7870), .Z(net_7968) );
CLKBUF_X2 inst_9707 ( .A(net_8234), .Z(net_9669) );
CLKBUF_X2 inst_13742 ( .A(net_13703), .Z(net_13704) );
SDFF_X2 inst_1083 ( .SI(net_6947), .Q(net_6947), .D(net_3775), .SE(net_3741), .CK(net_11451) );
INV_X4 inst_5408 ( .A(net_6153), .ZN(net_3579) );
NAND2_X2 inst_4073 ( .A1(net_6530), .A2(net_1645), .ZN(net_979) );
INV_X16 inst_6123 ( .ZN(net_4950), .A(net_4264) );
CLKBUF_X2 inst_12036 ( .A(net_10609), .Z(net_11998) );
SDFF_X2 inst_1136 ( .SI(net_6659), .Q(net_6659), .D(net_3799), .SE(net_3471), .CK(net_10039) );
NOR2_X2 inst_2466 ( .ZN(net_2731), .A1(net_2730), .A2(net_2729) );
CLKBUF_X2 inst_11979 ( .A(net_11940), .Z(net_11941) );
CLKBUF_X2 inst_11877 ( .A(net_8573), .Z(net_11839) );
CLKBUF_X2 inst_12070 ( .A(net_9329), .Z(net_12032) );
CLKBUF_X2 inst_10402 ( .A(net_10363), .Z(net_10364) );
CLKBUF_X2 inst_13615 ( .A(net_13576), .Z(net_13577) );
CLKBUF_X2 inst_13360 ( .A(net_13321), .Z(net_13322) );
CLKBUF_X2 inst_11262 ( .A(net_11223), .Z(net_11224) );
SDFF_X2 inst_696 ( .Q(net_6734), .D(net_6734), .SE(net_3815), .SI(net_3814), .CK(net_8962) );
CLKBUF_X2 inst_9719 ( .A(net_8370), .Z(net_9681) );
CLKBUF_X2 inst_9621 ( .A(net_9582), .Z(net_9583) );
NAND2_X2 inst_3311 ( .ZN(net_3624), .A1(net_3623), .A2(net_3226) );
CLKBUF_X2 inst_13598 ( .A(net_11332), .Z(net_13560) );
CLKBUF_X2 inst_11890 ( .A(net_11018), .Z(net_11852) );
CLKBUF_X2 inst_13339 ( .A(net_9253), .Z(net_13301) );
CLKBUF_X2 inst_12059 ( .A(net_12020), .Z(net_12021) );
CLKBUF_X2 inst_10755 ( .A(net_9885), .Z(net_10717) );
INV_X4 inst_5055 ( .ZN(net_872), .A(net_278) );
INV_X4 inst_5081 ( .ZN(net_719), .A(net_267) );
INV_X4 inst_5117 ( .A(net_769), .ZN(net_637) );
INV_X4 inst_4929 ( .ZN(net_1304), .A(net_799) );
INV_X4 inst_5114 ( .ZN(net_604), .A(net_603) );
CLKBUF_X2 inst_13942 ( .A(net_13780), .Z(net_13904) );
INV_X16 inst_6128 ( .ZN(net_4476), .A(net_3844) );
CLKBUF_X2 inst_10778 ( .A(net_10739), .Z(net_10740) );
CLKBUF_X2 inst_11712 ( .A(net_10437), .Z(net_11674) );
NAND2_X2 inst_3969 ( .A1(net_2382), .A2(net_1820), .ZN(net_1311) );
CLKBUF_X2 inst_9909 ( .A(net_8413), .Z(net_9871) );
NOR2_X2 inst_2363 ( .ZN(net_5287), .A2(net_4630), .A1(net_4486) );
INV_X2 inst_6014 ( .A(net_7364), .ZN(net_2046) );
CLKBUF_X2 inst_10423 ( .A(net_10384), .Z(net_10385) );
DFF_X2 inst_6257 ( .Q(net_6387), .D(net_6386), .CK(net_13687) );
NAND2_X2 inst_4029 ( .A1(net_6808), .A2(net_1651), .ZN(net_1023) );
OAI22_X1 inst_1629 ( .B2(net_4107), .ZN(net_3860), .A2(net_3442), .A1(net_1708), .B1(net_1091) );
AOI22_X2 inst_7341 ( .ZN(net_3182), .A2(net_2988), .B2(net_2906), .A1(net_1748), .B1(net_922) );
NAND2_X2 inst_3424 ( .A2(net_5891), .ZN(net_3324), .A1(net_627) );
DFF_X2 inst_6268 ( .QN(net_5974), .D(net_2639), .CK(net_8556) );
CLKBUF_X2 inst_12138 ( .A(net_12099), .Z(net_12100) );
CLKBUF_X2 inst_13923 ( .A(net_13884), .Z(net_13885) );
NAND2_X2 inst_3713 ( .A1(net_6766), .A2(net_1635), .ZN(net_1633) );
NAND3_X2 inst_2580 ( .ZN(net_5759), .A1(net_5654), .A2(net_5276), .A3(net_4314) );
INV_X4 inst_5681 ( .A(net_6148), .ZN(net_3587) );
NOR2_X2 inst_2394 ( .A2(net_3996), .ZN(net_3991), .A1(net_888) );
CLKBUF_X2 inst_11342 ( .A(net_11303), .Z(net_11304) );
INV_X4 inst_4574 ( .ZN(net_5786), .A(net_5785) );
CLKBUF_X2 inst_14213 ( .A(net_14174), .Z(net_14175) );
CLKBUF_X2 inst_8562 ( .A(net_8299), .Z(net_8524) );
CLKBUF_X2 inst_12268 ( .A(net_12229), .Z(net_12230) );
CLKBUF_X2 inst_9404 ( .A(net_8647), .Z(net_9366) );
CLKBUF_X2 inst_10681 ( .A(net_10319), .Z(net_10643) );
CLKBUF_X2 inst_10612 ( .A(net_10355), .Z(net_10574) );
INV_X2 inst_5840 ( .ZN(net_777), .A(net_776) );
OAI21_X2 inst_2054 ( .B1(net_5898), .B2(net_4457), .ZN(net_4444), .A(net_3557) );
CLKBUF_X2 inst_12216 ( .A(net_12177), .Z(net_12178) );
CLKBUF_X2 inst_13448 ( .A(net_11229), .Z(net_13410) );
INV_X4 inst_5294 ( .A(net_6142), .ZN(net_3649) );
INV_X4 inst_5251 ( .A(net_472), .ZN(net_439) );
SDFF_X2 inst_1259 ( .SI(net_6528), .Q(net_6528), .D(net_3814), .SE(net_3755), .CK(net_11214) );
NAND2_X1 inst_4422 ( .A1(net_7610), .A2(net_2131), .ZN(net_1510) );
CLKBUF_X2 inst_12578 ( .A(net_12539), .Z(net_12540) );
CLKBUF_X2 inst_12219 ( .A(net_12180), .Z(net_12181) );
CLKBUF_X2 inst_14056 ( .A(net_14017), .Z(net_14018) );
CLKBUF_X2 inst_11905 ( .A(net_11866), .Z(net_11867) );
CLKBUF_X2 inst_8623 ( .A(net_8317), .Z(net_8585) );
AND2_X4 inst_7821 ( .ZN(net_3257), .A2(net_3158), .A1(net_597) );
INV_X4 inst_5092 ( .A(net_7803), .ZN(net_3894) );
CLKBUF_X2 inst_10702 ( .A(net_10663), .Z(net_10664) );
OAI21_X2 inst_1796 ( .ZN(net_5394), .A(net_4720), .B2(net_3986), .B1(net_1067) );
CLKBUF_X2 inst_12318 ( .A(net_8122), .Z(net_12280) );
AOI21_X2 inst_7649 ( .B2(net_3439), .ZN(net_3398), .A(net_3221), .B1(net_1224) );
CLKBUF_X2 inst_11341 ( .A(net_11302), .Z(net_11303) );
SDFF_X2 inst_535 ( .Q(net_6566), .D(net_6566), .SI(net_3883), .SE(net_3823), .CK(net_7889) );
INV_X4 inst_5342 ( .A(net_7227), .ZN(net_433) );
CLKBUF_X2 inst_12970 ( .A(net_12931), .Z(net_12932) );
OAI221_X2 inst_1670 ( .ZN(net_4529), .C2(net_4301), .B2(net_4300), .A(net_4159), .B1(net_870), .C1(net_869) );
CLKBUF_X2 inst_12932 ( .A(net_12893), .Z(net_12894) );
CLKBUF_X2 inst_11491 ( .A(net_11452), .Z(net_11453) );
CLKBUF_X2 inst_10059 ( .A(net_10020), .Z(net_10021) );
AND2_X2 inst_7853 ( .ZN(net_3745), .A1(net_3452), .A2(net_113) );
CLKBUF_X2 inst_11670 ( .A(net_11631), .Z(net_11632) );
CLKBUF_X2 inst_10352 ( .A(net_7943), .Z(net_10314) );
CLKBUF_X2 inst_8646 ( .A(net_7953), .Z(net_8608) );
NOR2_X2 inst_2427 ( .ZN(net_3429), .A2(net_3123), .A1(net_3044) );
CLKBUF_X2 inst_9028 ( .A(net_8989), .Z(net_8990) );
CLKBUF_X2 inst_10496 ( .A(net_10457), .Z(net_10458) );
CLKBUF_X2 inst_8603 ( .A(net_8447), .Z(net_8565) );
CLKBUF_X2 inst_10677 ( .A(net_10638), .Z(net_10639) );
NAND2_X2 inst_3317 ( .ZN(net_3612), .A1(net_3611), .A2(net_3228) );
CLKBUF_X2 inst_10327 ( .A(net_9266), .Z(net_10289) );
INV_X4 inst_5027 ( .ZN(net_885), .A(net_663) );
INV_X2 inst_5883 ( .A(net_7442), .ZN(net_1358) );
NAND2_X2 inst_3113 ( .A1(net_6619), .A2(net_4899), .ZN(net_4888) );
CLKBUF_X2 inst_13500 ( .A(net_10359), .Z(net_13462) );
INV_X2 inst_6079 ( .A(net_7293), .ZN(net_2013) );
CLKBUF_X2 inst_13245 ( .A(net_13206), .Z(net_13207) );
CLKBUF_X2 inst_11348 ( .A(net_8650), .Z(net_11310) );
NAND2_X2 inst_3695 ( .ZN(net_1735), .A1(net_1279), .A2(net_1096) );
CLKBUF_X2 inst_12309 ( .A(net_12270), .Z(net_12271) );
NAND2_X2 inst_3168 ( .ZN(net_4765), .A2(net_3941), .A1(net_2015) );
DFF_X1 inst_6687 ( .QN(net_7276), .D(net_5116), .CK(net_9961) );
NOR2_X2 inst_2385 ( .ZN(net_4294), .A1(net_4149), .A2(net_4148) );
NOR2_X2 inst_2336 ( .A2(net_6282), .A1(net_5843), .ZN(net_5805) );
NAND2_X2 inst_3855 ( .A1(net_6703), .A2(net_1497), .ZN(net_1480) );
INV_X2 inst_5927 ( .A(net_7515), .ZN(net_2168) );
CLKBUF_X2 inst_8589 ( .A(net_8447), .Z(net_8551) );
CLKBUF_X2 inst_8574 ( .A(net_8289), .Z(net_8536) );
CLKBUF_X2 inst_13549 ( .A(net_11009), .Z(net_13511) );
CLKBUF_X2 inst_10594 ( .A(net_8208), .Z(net_10556) );
CLKBUF_X2 inst_9482 ( .A(net_8126), .Z(net_9444) );
NAND2_X2 inst_3318 ( .ZN(net_3610), .A1(net_3609), .A2(net_3228) );
CLKBUF_X2 inst_12771 ( .A(net_12732), .Z(net_12733) );
SDFF_X2 inst_223 ( .Q(net_6331), .SI(net_6330), .D(net_3663), .SE(net_392), .CK(net_14041) );
CLKBUF_X2 inst_10299 ( .A(net_10260), .Z(net_10261) );
DFF_X1 inst_6814 ( .D(net_3254), .CK(net_13209), .Q(x264) );
INV_X4 inst_5278 ( .ZN(net_611), .A(net_415) );
INV_X2 inst_6042 ( .A(net_7601), .ZN(net_1398) );
CLKBUF_X2 inst_13811 ( .A(net_13772), .Z(net_13773) );
NOR2_X2 inst_2420 ( .A2(net_5917), .ZN(net_3231), .A1(net_3230) );
NAND2_X2 inst_3564 ( .ZN(net_2503), .A2(net_2018), .A1(net_1756) );
INV_X4 inst_5176 ( .ZN(net_661), .A(net_530) );
CLKBUF_X2 inst_12672 ( .A(net_12633), .Z(net_12634) );
NAND2_X2 inst_4205 ( .A2(net_6042), .A1(net_6041), .ZN(net_3236) );
SDFF_X2 inst_1322 ( .D(net_6382), .SE(net_5801), .SI(net_327), .Q(net_327), .CK(net_14290) );
CLKBUF_X2 inst_11862 ( .A(net_11823), .Z(net_11824) );
CLKBUF_X2 inst_11452 ( .A(net_11413), .Z(net_11414) );
CLKBUF_X2 inst_9633 ( .A(net_9085), .Z(net_9595) );
CLKBUF_X2 inst_10954 ( .A(net_10915), .Z(net_10916) );
CLKBUF_X2 inst_14004 ( .A(net_13965), .Z(net_13966) );
CLKBUF_X2 inst_10712 ( .A(net_10267), .Z(net_10674) );
CLKBUF_X2 inst_14237 ( .A(net_14198), .Z(net_14199) );
CLKBUF_X2 inst_10248 ( .A(net_10209), .Z(net_10210) );
CLKBUF_X2 inst_12027 ( .A(net_11988), .Z(net_11989) );
AOI21_X2 inst_7668 ( .ZN(net_3009), .B1(net_2860), .B2(net_2744), .A(net_921) );
CLKBUF_X2 inst_11063 ( .A(net_11024), .Z(net_11025) );
CLKBUF_X2 inst_9408 ( .A(net_8513), .Z(net_9370) );
CLKBUF_X2 inst_10156 ( .A(net_10117), .Z(net_10118) );
CLKBUF_X2 inst_8379 ( .A(net_8140), .Z(net_8341) );
NAND2_X2 inst_3493 ( .ZN(net_2729), .A2(net_2628), .A1(net_2591) );
INV_X1 inst_6156 ( .A(net_5850), .ZN(x63) );
CLKBUF_X2 inst_13151 ( .A(net_13112), .Z(net_13113) );
CLKBUF_X2 inst_10413 ( .A(net_7881), .Z(net_10375) );
CLKBUF_X2 inst_9776 ( .A(net_9737), .Z(net_9738) );
NAND2_X2 inst_3019 ( .A1(net_6859), .A2(net_5004), .ZN(net_4990) );
INV_X4 inst_4622 ( .ZN(net_4200), .A(net_4060) );
NOR2_X2 inst_2327 ( .A2(net_6291), .A1(net_5843), .ZN(net_5814) );
CLKBUF_X2 inst_13430 ( .A(net_12036), .Z(net_13392) );
NAND2_X2 inst_3487 ( .ZN(net_2659), .A1(net_2658), .A2(net_2657) );
INV_X4 inst_5078 ( .A(net_7810), .ZN(net_3808) );
DFF_X1 inst_6866 ( .D(net_2540), .Q(net_200), .CK(net_10066) );
CLKBUF_X2 inst_14421 ( .A(net_14382), .Z(net_14383) );
CLKBUF_X2 inst_11783 ( .A(net_11744), .Z(net_11745) );
NAND2_X2 inst_3597 ( .ZN(net_2403), .A2(net_1859), .A1(net_1517) );
CLKBUF_X2 inst_8210 ( .A(net_8171), .Z(net_8172) );
CLKBUF_X2 inst_10661 ( .A(net_7952), .Z(net_10623) );
CLKBUF_X2 inst_11757 ( .A(net_11521), .Z(net_11719) );
CLKBUF_X2 inst_13422 ( .A(net_8902), .Z(net_13384) );
NAND3_X2 inst_2607 ( .ZN(net_5732), .A1(net_5627), .A2(net_5170), .A3(net_4192) );
CLKBUF_X2 inst_11579 ( .A(net_11540), .Z(net_11541) );
XNOR2_X2 inst_113 ( .A(net_2565), .ZN(net_824), .B(net_823) );
CLKBUF_X2 inst_13893 ( .A(net_8134), .Z(net_13855) );
CLKBUF_X2 inst_8133 ( .A(net_8094), .Z(net_8095) );
CLKBUF_X2 inst_11395 ( .A(net_11356), .Z(net_11357) );
CLKBUF_X2 inst_10433 ( .A(net_10394), .Z(net_10395) );
AND4_X4 inst_7791 ( .A3(net_7688), .ZN(net_1664), .A2(net_1219), .A4(net_1218), .A1(net_411) );
CLKBUF_X2 inst_14023 ( .A(net_13984), .Z(net_13985) );
NAND3_X2 inst_2690 ( .ZN(net_3151), .A2(net_3150), .A3(net_3043), .A1(net_3004) );
CLKBUF_X2 inst_9680 ( .A(net_9028), .Z(net_9642) );
CLKBUF_X2 inst_9106 ( .A(net_9067), .Z(net_9068) );
CLKBUF_X2 inst_8479 ( .A(net_8207), .Z(net_8441) );
CLKBUF_X2 inst_8689 ( .A(net_8597), .Z(net_8651) );
CLKBUF_X2 inst_10849 ( .A(net_8719), .Z(net_10811) );
CLKBUF_X2 inst_10467 ( .A(net_10428), .Z(net_10429) );
AOI22_X2 inst_7298 ( .B1(net_6548), .A1(net_6516), .A2(net_5184), .B2(net_5183), .ZN(net_5171) );
OAI22_X2 inst_1544 ( .B2(net_3405), .ZN(net_3362), .A2(net_3360), .A1(net_3273), .B1(net_454) );
NAND2_X2 inst_4063 ( .A1(net_6807), .A2(net_1651), .ZN(net_989) );
CLKBUF_X2 inst_10069 ( .A(net_10030), .Z(net_10031) );
CLKBUF_X2 inst_8340 ( .A(net_8231), .Z(net_8302) );
DFF_X2 inst_6261 ( .QN(net_5971), .D(net_2734), .CK(net_11410) );
CLKBUF_X2 inst_9016 ( .A(net_8977), .Z(net_8978) );
NAND3_X2 inst_2625 ( .ZN(net_5704), .A1(net_5681), .A2(net_5317), .A3(net_4255) );
CLKBUF_X2 inst_9771 ( .A(net_9732), .Z(net_9733) );
NAND2_X2 inst_3148 ( .ZN(net_4815), .A2(net_4153), .A1(net_2093) );
CLKBUF_X2 inst_14088 ( .A(net_14049), .Z(net_14050) );
INV_X2 inst_6064 ( .A(net_7591), .ZN(net_1320) );
CLKBUF_X2 inst_12652 ( .A(net_10015), .Z(net_12614) );
CLKBUF_X2 inst_9244 ( .A(net_9205), .Z(net_9206) );
NAND2_X2 inst_3329 ( .ZN(net_3588), .A1(net_3587), .A2(net_3228) );
INV_X4 inst_4761 ( .ZN(net_2564), .A(net_2263) );
INV_X4 inst_5180 ( .ZN(net_524), .A(net_523) );
NAND2_X2 inst_3026 ( .ZN(net_4983), .A2(net_4330), .A1(net_2260) );
INV_X2 inst_5769 ( .ZN(net_2996), .A(net_2900) );
CLKBUF_X2 inst_13844 ( .A(net_8020), .Z(net_13806) );
NAND2_X4 inst_2847 ( .ZN(net_5476), .A1(net_4921), .A2(net_4920) );
OAI22_X2 inst_1442 ( .B2(net_5904), .B1(net_4666), .A2(net_4634), .ZN(net_4633), .A1(net_4116) );
CLKBUF_X2 inst_8573 ( .A(net_8534), .Z(net_8535) );
DFFS_X2 inst_6952 ( .QN(net_6409), .D(net_2720), .CK(net_14400), .SN(x1822) );
NAND2_X2 inst_3639 ( .ZN(net_1944), .A1(net_1297), .A2(net_1110) );
SDFF_X2 inst_332 ( .D(net_6393), .SE(net_5800), .SI(net_358), .Q(net_358), .CK(net_13670) );
CLKBUF_X2 inst_14192 ( .A(net_8120), .Z(net_14154) );
NAND2_X2 inst_4013 ( .ZN(net_1236), .A2(net_1222), .A1(net_345) );
OAI21_X2 inst_2132 ( .ZN(net_2902), .A(net_2901), .B2(net_2896), .B1(net_902) );
SDFF_X2 inst_1289 ( .D(net_3883), .SE(net_3256), .SI(net_137), .Q(net_137), .CK(net_8467) );
CLKBUF_X2 inst_13646 ( .A(net_13607), .Z(net_13608) );
INV_X4 inst_4979 ( .A(net_7816), .ZN(net_3782) );
CLKBUF_X2 inst_10411 ( .A(net_10372), .Z(net_10373) );
CLKBUF_X2 inst_9194 ( .A(net_9155), .Z(net_9156) );
INV_X4 inst_4686 ( .ZN(net_3737), .A(net_3365) );
CLKBUF_X2 inst_14241 ( .A(net_14202), .Z(net_14203) );
CLKBUF_X2 inst_13130 ( .A(net_11726), .Z(net_13092) );
INV_X4 inst_4869 ( .A(net_3042), .ZN(net_1092) );
CLKBUF_X2 inst_12769 ( .A(net_12730), .Z(net_12731) );
NAND2_X2 inst_3245 ( .A2(net_3992), .ZN(net_3989), .A1(net_3982) );
SDFF_X2 inst_752 ( .Q(net_6874), .D(net_6874), .SE(net_3901), .SI(net_3811), .CK(net_8878) );
NAND2_X2 inst_3202 ( .ZN(net_4724), .A2(net_3986), .A1(net_2101) );
NAND2_X1 inst_4279 ( .ZN(net_4588), .A2(net_3867), .A1(net_1903) );
OAI21_X2 inst_1951 ( .ZN(net_5069), .B1(net_4853), .A(net_4726), .B2(net_3986) );
SDFF_X2 inst_378 ( .SI(net_7673), .Q(net_7673), .D(net_4797), .SE(net_3866), .CK(net_13238) );
AOI22_X2 inst_7444 ( .A2(net_2938), .B2(net_2670), .ZN(net_860), .A1(net_859), .B1(net_858) );
OR2_X4 inst_1384 ( .A2(net_6184), .A1(net_2997), .ZN(net_2743) );
CLKBUF_X2 inst_8151 ( .A(net_8112), .Z(net_8113) );
OAI21_X2 inst_2118 ( .B2(net_3297), .ZN(net_3295), .B1(net_3142), .A(net_3078) );
CLKBUF_X2 inst_11302 ( .A(net_11113), .Z(net_11264) );
CLKBUF_X2 inst_8750 ( .A(net_8711), .Z(net_8712) );
NOR3_X2 inst_2200 ( .ZN(net_3449), .A3(net_3173), .A2(net_3010), .A1(net_2859) );
AOI21_X2 inst_7749 ( .B1(net_6861), .ZN(net_4487), .B2(net_2579), .A(net_2328) );
CLKBUF_X2 inst_8817 ( .A(net_8150), .Z(net_8779) );
INV_X4 inst_4937 ( .ZN(net_756), .A(net_755) );
INV_X4 inst_5048 ( .A(net_2999), .ZN(net_883) );
CLKBUF_X2 inst_10320 ( .A(net_9500), .Z(net_10282) );
CLKBUF_X2 inst_8284 ( .A(net_8245), .Z(net_8246) );
CLKBUF_X2 inst_8080 ( .A(net_7901), .Z(net_8042) );
CLKBUF_X2 inst_11470 ( .A(net_10217), .Z(net_11432) );
CLKBUF_X2 inst_9948 ( .A(net_9909), .Z(net_9910) );
CLKBUF_X2 inst_12693 ( .A(net_12171), .Z(net_12655) );
SDFF_X2 inst_250 ( .Q(net_6344), .SI(net_6343), .D(net_3587), .SE(net_392), .CK(net_13648) );
NAND2_X1 inst_4356 ( .ZN(net_4371), .A2(net_3853), .A1(net_2078) );
CLKBUF_X2 inst_9275 ( .A(net_9236), .Z(net_9237) );
CLKBUF_X2 inst_11707 ( .A(net_10743), .Z(net_11669) );
AOI21_X2 inst_7708 ( .B1(net_6871), .ZN(net_4110), .B2(net_2579), .A(net_2355) );
INV_X2 inst_5762 ( .ZN(net_3033), .A(net_2975) );
CLKBUF_X2 inst_12250 ( .A(net_12080), .Z(net_12212) );
CLKBUF_X2 inst_9975 ( .A(net_9936), .Z(net_9937) );
DFF_X1 inst_6595 ( .QN(net_7484), .D(net_5415), .CK(net_9811) );
CLKBUF_X2 inst_9384 ( .A(net_9345), .Z(net_9346) );
INV_X4 inst_5329 ( .A(net_6110), .ZN(net_3675) );
NOR2_X2 inst_2539 ( .A2(net_7758), .A1(net_3208), .ZN(net_655) );
OAI22_X2 inst_1523 ( .B1(net_4644), .A1(net_4057), .B2(net_4053), .ZN(net_4050), .A2(net_4049) );
CLKBUF_X2 inst_10141 ( .A(net_10102), .Z(net_10103) );
CLKBUF_X2 inst_9941 ( .A(net_8129), .Z(net_9903) );
SDFF_X2 inst_1048 ( .Q(net_7249), .D(net_7249), .SE(net_3822), .SI(net_345), .CK(net_9826) );
DFFR_X1 inst_7120 ( .QN(net_5850), .D(net_5684), .CK(net_10255), .RN(x1822) );
CLKBUF_X2 inst_13496 ( .A(net_13457), .Z(net_13458) );
NAND3_X2 inst_2797 ( .ZN(net_2303), .A3(net_1595), .A1(net_1318), .A2(net_958) );
NAND2_X2 inst_3431 ( .ZN(net_3217), .A2(net_3101), .A1(net_2766) );
CLKBUF_X2 inst_13537 ( .A(net_8089), .Z(net_13499) );
CLKBUF_X2 inst_13193 ( .A(net_13154), .Z(net_13155) );
NOR2_X4 inst_2270 ( .ZN(net_5616), .A1(net_5461), .A2(net_4410) );
OAI21_X2 inst_2085 ( .B2(net_4415), .ZN(net_4404), .B1(net_4403), .A(net_3484) );
CLKBUF_X2 inst_11624 ( .A(net_11585), .Z(net_11586) );
NOR2_X2 inst_2401 ( .ZN(net_3771), .A1(net_3770), .A2(net_3769) );
CLKBUF_X2 inst_11097 ( .A(net_9887), .Z(net_11059) );
CLKBUF_X2 inst_12979 ( .A(net_12940), .Z(net_12941) );
INV_X4 inst_5264 ( .A(net_835), .ZN(net_426) );
CLKBUF_X2 inst_10092 ( .A(net_10053), .Z(net_10054) );
CLKBUF_X2 inst_12649 ( .A(net_12610), .Z(net_12611) );
CLKBUF_X2 inst_9356 ( .A(net_9317), .Z(net_9318) );
CLKBUF_X2 inst_8367 ( .A(net_8328), .Z(net_8329) );
CLKBUF_X2 inst_8015 ( .A(net_7976), .Z(net_7977) );
CLKBUF_X2 inst_12910 ( .A(net_7875), .Z(net_12872) );
INV_X1 inst_6150 ( .A(net_3403), .ZN(net_3327) );
DFFR_X2 inst_7069 ( .QN(net_6031), .D(net_3063), .CK(net_9999), .RN(x1822) );
CLKBUF_X2 inst_14230 ( .A(net_14191), .Z(net_14192) );
CLKBUF_X2 inst_8196 ( .A(net_7899), .Z(net_8158) );
CLKBUF_X2 inst_11779 ( .A(net_11740), .Z(net_11741) );
SDFF_X2 inst_556 ( .SI(net_7192), .Q(net_7192), .D(net_3821), .SE(net_3819), .CK(net_10671) );
INV_X2 inst_6050 ( .ZN(net_397), .A(x1006) );
CLKBUF_X2 inst_14287 ( .A(net_14248), .Z(net_14249) );
NAND2_X2 inst_3632 ( .A2(net_5931), .ZN(net_2727), .A1(net_1951) );
DFF_X2 inst_6204 ( .QN(net_6552), .D(net_4393), .CK(net_7935) );
CLKBUF_X2 inst_8618 ( .A(net_7902), .Z(net_8580) );
CLKBUF_X2 inst_9710 ( .A(net_9671), .Z(net_9672) );
SDFF_X2 inst_420 ( .Q(net_6363), .SI(net_6362), .D(net_3562), .SE(net_392), .CK(net_13739) );
INV_X4 inst_5147 ( .ZN(net_683), .A(net_569) );
CLKBUF_X2 inst_13758 ( .A(net_13719), .Z(net_13720) );
NAND2_X2 inst_3992 ( .ZN(net_1230), .A2(net_860), .A1(net_857) );
CLKBUF_X2 inst_12522 ( .A(net_9625), .Z(net_12484) );
NAND2_X2 inst_3265 ( .ZN(net_4141), .A1(net_3852), .A2(net_3463) );
CLKBUF_X2 inst_12573 ( .A(net_12534), .Z(net_12535) );
CLKBUF_X2 inst_9650 ( .A(net_9611), .Z(net_9612) );
NAND2_X2 inst_3300 ( .ZN(net_3646), .A1(net_3645), .A2(net_3229) );
AOI222_X2 inst_7558 ( .A1(net_7397), .ZN(net_5442), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_360), .C2(net_358) );
SDFF_X2 inst_1305 ( .D(net_6386), .SE(net_6052), .SI(net_311), .Q(net_311), .CK(net_13722) );
CLKBUF_X2 inst_7997 ( .A(net_7958), .Z(net_7959) );
SDFF_X2 inst_314 ( .SI(net_7456), .Q(net_7456), .D(net_5104), .SE(net_3993), .CK(net_12072) );
CLKBUF_X2 inst_8713 ( .A(net_7971), .Z(net_8675) );
NAND2_X2 inst_3225 ( .A2(net_7779), .ZN(net_5255), .A1(net_4296) );
CLKBUF_X2 inst_13367 ( .A(net_13328), .Z(net_13329) );
AOI222_X2 inst_7597 ( .A1(net_7235), .ZN(net_4868), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_329), .C2(net_327) );
CLKBUF_X2 inst_12728 ( .A(net_12689), .Z(net_12690) );
CLKBUF_X2 inst_8757 ( .A(net_8018), .Z(net_8719) );
NAND2_X2 inst_3822 ( .A1(net_7175), .A2(net_1637), .ZN(net_1523) );
CLKBUF_X2 inst_9603 ( .A(net_8591), .Z(net_9565) );
SDFF_X2 inst_597 ( .SI(net_7802), .Q(net_6568), .D(net_6568), .SE(net_3823), .CK(net_9178) );
INV_X1 inst_6161 ( .A(net_5855), .ZN(x106) );
AOI222_X2 inst_7522 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2002), .A1(net_2001), .B1(net_2000), .C1(net_1999) );
INV_X4 inst_4593 ( .ZN(net_4305), .A(net_4172) );
INV_X4 inst_5524 ( .A(net_6006), .ZN(net_516) );
AOI22_X2 inst_7257 ( .B1(net_6948), .A1(net_6916), .ZN(net_5299), .A2(net_5298), .B2(net_5297) );
INV_X2 inst_6070 ( .A(net_7589), .ZN(net_1985) );
NAND2_X2 inst_3307 ( .ZN(net_3632), .A1(net_3631), .A2(net_3229) );
CLKBUF_X2 inst_11859 ( .A(net_9647), .Z(net_11821) );
DFF_X1 inst_6927 ( .D(net_2401), .Q(net_237), .CK(net_13132) );
CLKBUF_X2 inst_12272 ( .A(net_12142), .Z(net_12234) );
OAI22_X2 inst_1587 ( .B2(net_3200), .A2(net_3187), .ZN(net_3186), .A1(net_822), .B1(net_501) );
SDFF_X2 inst_1185 ( .SI(net_6930), .Q(net_6930), .D(net_3798), .SE(net_3741), .CK(net_8905) );
INV_X4 inst_5452 ( .A(net_7276), .ZN(net_2117) );
CLKBUF_X2 inst_8742 ( .A(net_8703), .Z(net_8704) );
SDFF_X2 inst_472 ( .Q(net_7540), .D(net_7540), .SE(net_3896), .SI(net_374), .CK(net_13124) );
SDFF_X2 inst_447 ( .D(net_6390), .SE(net_5801), .SI(net_335), .Q(net_335), .CK(net_14307) );
INV_X8 inst_4533 ( .A(net_6055), .ZN(net_5799) );
CLKBUF_X2 inst_13715 ( .A(net_13676), .Z(net_13677) );
SDFF_X2 inst_457 ( .Q(net_6056), .SI(net_3917), .SE(net_3310), .D(net_3309), .CK(net_10509) );
INV_X2 inst_5987 ( .A(net_7484), .ZN(net_2141) );
OAI21_X2 inst_1738 ( .ZN(net_5543), .B1(net_5542), .A(net_4809), .B2(net_4153) );
CLKBUF_X2 inst_12872 ( .A(net_12833), .Z(net_12834) );
NAND3_X2 inst_2802 ( .ZN(net_2296), .A3(net_1574), .A1(net_1518), .A2(net_959) );
NAND3_X2 inst_2623 ( .ZN(net_5716), .A1(net_5611), .A2(net_5124), .A3(net_4175) );
OR2_X4 inst_1391 ( .A2(net_7766), .ZN(net_2807), .A1(net_289) );
NAND2_X2 inst_4171 ( .A1(net_891), .ZN(net_808), .A2(net_612) );
SDFF_X2 inst_665 ( .Q(net_6724), .D(net_6724), .SE(net_3871), .SI(net_3801), .CK(net_11393) );
INV_X4 inst_4843 ( .ZN(net_4791), .A(net_1067) );
CLKBUF_X2 inst_12929 ( .A(net_12890), .Z(net_12891) );
CLKBUF_X2 inst_12014 ( .A(net_9429), .Z(net_11976) );
CLKBUF_X2 inst_11276 ( .A(net_11237), .Z(net_11238) );
CLKBUF_X2 inst_10219 ( .A(net_10180), .Z(net_10181) );
NAND2_X2 inst_3538 ( .ZN(net_2529), .A2(net_2130), .A1(net_1194) );
INV_X4 inst_5529 ( .A(net_6406), .ZN(net_437) );
CLKBUF_X2 inst_10250 ( .A(net_10211), .Z(net_10212) );
CLKBUF_X2 inst_8953 ( .A(net_8299), .Z(net_8915) );
INV_X2 inst_6103 ( .A(net_7509), .ZN(net_2192) );
NAND2_X2 inst_3755 ( .A1(net_7168), .A2(net_1637), .ZN(net_1590) );
SDFF_X2 inst_146 ( .Q(net_6232), .SI(net_6231), .SE(net_392), .D(net_138), .CK(net_14112) );
CLKBUF_X2 inst_8718 ( .A(net_7905), .Z(net_8680) );
CLKBUF_X2 inst_9810 ( .A(net_9771), .Z(net_9772) );
NAND2_X2 inst_3999 ( .A2(net_1910), .ZN(net_1185), .A1(net_1184) );
SDFF_X2 inst_1196 ( .SI(net_7078), .Q(net_7078), .D(net_3831), .SE(net_3747), .CK(net_11923) );
CLKBUF_X2 inst_12501 ( .A(net_12462), .Z(net_12463) );
CLKBUF_X2 inst_13815 ( .A(net_10493), .Z(net_13777) );
CLKBUF_X2 inst_10589 ( .A(net_10502), .Z(net_10551) );
SDFF_X2 inst_817 ( .Q(net_6992), .D(net_6992), .SE(net_3891), .SI(net_3793), .CK(net_11018) );
SDFF_X2 inst_326 ( .SI(net_7491), .Q(net_7491), .D(net_5102), .SE(net_3989), .CK(net_9774) );
CLKBUF_X2 inst_12550 ( .A(net_12511), .Z(net_12512) );
NAND2_X2 inst_3428 ( .ZN(net_3220), .A2(net_3108), .A1(net_2774) );
NOR3_X2 inst_2194 ( .ZN(net_3882), .A1(net_3385), .A3(net_1157), .A2(net_805) );
CLKBUF_X2 inst_10789 ( .A(net_10750), .Z(net_10751) );
CLKBUF_X2 inst_10510 ( .A(net_10471), .Z(net_10472) );
NAND2_X2 inst_3336 ( .ZN(net_3574), .A1(net_3573), .A2(net_3228) );
CLKBUF_X2 inst_7963 ( .A(net_7924), .Z(net_7925) );
CLKBUF_X2 inst_9034 ( .A(net_8995), .Z(net_8996) );
NAND2_X2 inst_3293 ( .ZN(net_3660), .A1(net_3659), .A2(net_3229) );
NAND2_X2 inst_3793 ( .A1(net_6903), .A2(net_1639), .ZN(net_1552) );
NAND2_X4 inst_2837 ( .ZN(net_5553), .A1(net_5024), .A2(net_5023) );
DFFR_X1 inst_7115 ( .QN(net_5855), .D(net_5795), .CK(net_10465), .RN(x1822) );
CLKBUF_X2 inst_11143 ( .A(net_11104), .Z(net_11105) );
OAI21_X2 inst_1845 ( .B1(net_5351), .ZN(net_5327), .A(net_4377), .B2(net_3853) );
XNOR2_X2 inst_108 ( .ZN(net_2414), .B(net_1204), .A(net_835) );
NAND2_X2 inst_3778 ( .A1(net_7037), .A2(net_1975), .ZN(net_1567) );
INV_X4 inst_4799 ( .ZN(net_5105), .A(net_1255) );
CLKBUF_X2 inst_9296 ( .A(net_8070), .Z(net_9258) );
DFF_X1 inst_6905 ( .D(net_2504), .Q(net_158), .CK(net_12223) );
NAND2_X2 inst_3940 ( .A1(net_6972), .A2(net_1833), .ZN(net_1351) );
DFF_X1 inst_6503 ( .QN(net_7425), .D(net_5526), .CK(net_12502) );
OR2_X2 inst_1429 ( .A2(net_6823), .A1(net_6822), .ZN(net_671) );
CLKBUF_X2 inst_8439 ( .A(net_8350), .Z(net_8401) );
CLKBUF_X2 inst_11937 ( .A(net_11376), .Z(net_11899) );
SDFF_X2 inst_638 ( .SI(net_6651), .Q(net_6651), .SE(net_3850), .D(net_3793), .CK(net_9108) );
AOI21_X2 inst_7786 ( .ZN(net_2423), .A(net_2232), .B1(net_1941), .B2(net_1684) );
CLKBUF_X2 inst_10311 ( .A(net_10272), .Z(net_10273) );
CLKBUF_X2 inst_12919 ( .A(net_12880), .Z(net_12881) );
SDFF_X2 inst_586 ( .Q(net_6585), .D(net_6585), .SE(net_3823), .SI(net_3790), .CK(net_12035) );
INV_X4 inst_5220 ( .ZN(net_796), .A(net_472) );
CLKBUF_X2 inst_9828 ( .A(net_9789), .Z(net_9790) );
CLKBUF_X2 inst_10563 ( .A(net_10524), .Z(net_10525) );
NAND3_X2 inst_2591 ( .ZN(net_5748), .A1(net_5643), .A2(net_5234), .A3(net_4207) );
CLKBUF_X2 inst_9237 ( .A(net_9198), .Z(net_9199) );
NAND2_X2 inst_3275 ( .ZN(net_3696), .A1(net_3695), .A2(net_3231) );
INV_X4 inst_5008 ( .A(net_7820), .ZN(net_3789) );
OAI22_X2 inst_1466 ( .B2(net_5077), .ZN(net_4396), .A1(net_4143), .A2(net_3827), .B1(net_1138) );
NAND2_X4 inst_2841 ( .ZN(net_5541), .A1(net_5016), .A2(net_5015) );
OAI21_X2 inst_1726 ( .ZN(net_5568), .B1(net_5438), .A(net_4833), .B2(net_4153) );
NAND3_X2 inst_2652 ( .A3(net_5959), .A2(net_5958), .ZN(net_3948), .A1(net_2831) );
INV_X4 inst_5221 ( .ZN(net_632), .A(net_471) );
SDFF_X2 inst_1203 ( .SI(net_7087), .Q(net_7087), .D(net_3789), .SE(net_3747), .CK(net_10977) );
CLKBUF_X2 inst_14251 ( .A(net_8479), .Z(net_14213) );
SDFF_X2 inst_802 ( .Q(net_6975), .D(net_6975), .SE(net_3891), .SI(net_3813), .CK(net_8421) );
SDFF_X2 inst_296 ( .D(net_6394), .SE(net_5799), .SI(net_379), .Q(net_379), .CK(net_14322) );
DFFR_X1 inst_7118 ( .QN(net_5852), .D(net_5686), .CK(net_12808), .RN(x1822) );
CLKBUF_X2 inst_10892 ( .A(net_8219), .Z(net_10854) );
SDFF_X2 inst_905 ( .Q(net_7131), .D(net_7131), .SE(net_3903), .SI(net_3797), .CK(net_13358) );
CLKBUF_X2 inst_11571 ( .A(net_11532), .Z(net_11533) );
NAND2_X1 inst_4370 ( .ZN(net_4357), .A2(net_3856), .A1(net_1776) );
CLKBUF_X2 inst_11218 ( .A(net_11179), .Z(net_11180) );
CLKBUF_X2 inst_9185 ( .A(net_9146), .Z(net_9147) );
NAND2_X2 inst_4214 ( .ZN(net_3255), .A2(net_292), .A1(net_291) );
CLKBUF_X2 inst_12753 ( .A(net_12714), .Z(net_12715) );
CLKBUF_X2 inst_11047 ( .A(net_11008), .Z(net_11009) );
NAND2_X2 inst_3834 ( .A1(net_7100), .A2(net_1675), .ZN(net_1505) );
NAND2_X2 inst_3943 ( .A1(net_6574), .A2(net_1705), .ZN(net_1348) );
NAND2_X2 inst_3651 ( .A1(net_7063), .ZN(net_1812), .A2(net_791) );
CLKBUF_X2 inst_14280 ( .A(net_14241), .Z(net_14242) );
OAI21_X2 inst_1759 ( .ZN(net_5439), .B1(net_5438), .A(net_4662), .B2(net_3993) );
CLKBUF_X2 inst_11792 ( .A(net_11753), .Z(net_11754) );
NAND3_X2 inst_2615 ( .ZN(net_5724), .A1(net_5619), .A2(net_5136), .A3(net_4183) );
NOR2_X2 inst_2532 ( .ZN(net_3983), .A1(net_1730), .A2(net_527) );
INV_X4 inst_5485 ( .A(net_6085), .ZN(net_3493) );
CLKBUF_X2 inst_13859 ( .A(net_11811), .Z(net_13821) );
CLKBUF_X2 inst_13263 ( .A(net_7862), .Z(net_13225) );
NAND2_X2 inst_3463 ( .A2(net_5978), .ZN(net_2886), .A1(net_2885) );
NOR2_X2 inst_2463 ( .ZN(net_2736), .A1(net_2735), .A2(net_2733) );
DFFR_X2 inst_7017 ( .D(net_3272), .QN(net_291), .CK(net_11440), .RN(x1822) );
CLKBUF_X2 inst_11206 ( .A(net_10537), .Z(net_11168) );
CLKBUF_X2 inst_10907 ( .A(net_9773), .Z(net_10869) );
AOI221_X2 inst_7617 ( .C2(net_3105), .B1(net_2970), .ZN(net_2962), .A(net_2781), .C1(net_474), .B2(net_252) );
CLKBUF_X2 inst_12492 ( .A(net_12453), .Z(net_12454) );
CLKBUF_X2 inst_11115 ( .A(net_8993), .Z(net_11077) );
INV_X4 inst_5610 ( .A(net_6041), .ZN(net_479) );
DFF_X1 inst_6375 ( .QN(net_6287), .D(net_5809), .CK(net_14262) );
NAND2_X2 inst_4055 ( .A1(net_6799), .A2(net_1651), .ZN(net_997) );
OAI22_X2 inst_1464 ( .B2(net_5383), .ZN(net_4398), .A1(net_4150), .A2(net_3829), .B1(net_1161) );
SDFF_X2 inst_1247 ( .SI(net_6542), .Q(net_6542), .D(net_3775), .SE(net_3756), .CK(net_8397) );
CLKBUF_X2 inst_12778 ( .A(net_11323), .Z(net_12740) );
INV_X4 inst_5284 ( .A(net_6687), .ZN(net_421) );
CLKBUF_X2 inst_8490 ( .A(net_8451), .Z(net_8452) );
INV_X4 inst_5031 ( .ZN(net_763), .A(net_661) );
CLKBUF_X2 inst_13275 ( .A(net_13236), .Z(net_13237) );
CLKBUF_X2 inst_13498 ( .A(net_13459), .Z(net_13460) );
CLKBUF_X2 inst_13215 ( .A(net_13176), .Z(net_13177) );
OAI22_X2 inst_1493 ( .B1(net_4666), .A1(net_4132), .B2(net_4118), .ZN(net_4115), .A2(net_4114) );
DFF_X1 inst_6441 ( .QN(net_6072), .D(net_5729), .CK(net_10891) );
SDFF_X2 inst_1308 ( .SE(net_7680), .Q(net_7680), .D(net_2925), .SI(net_2924), .CK(net_10768) );
NAND2_X2 inst_3070 ( .A1(net_7130), .A2(net_4950), .ZN(net_4935) );
XNOR2_X2 inst_85 ( .B(net_2249), .ZN(net_1305), .A(net_1304) );
INV_X4 inst_4733 ( .A(net_5966), .ZN(net_3877) );
NAND2_X2 inst_2998 ( .A1(net_6714), .A2(net_5031), .ZN(net_5013) );
CLKBUF_X2 inst_11734 ( .A(net_11695), .Z(net_11696) );
CLKBUF_X2 inst_14116 ( .A(net_14077), .Z(net_14078) );
CLKBUF_X2 inst_13348 ( .A(net_9730), .Z(net_13310) );
NAND3_X2 inst_2612 ( .ZN(net_5727), .A1(net_5622), .A2(net_5141), .A3(net_4186) );
INV_X2 inst_5963 ( .A(net_7592), .ZN(net_1363) );
CLKBUF_X2 inst_9681 ( .A(net_8674), .Z(net_9643) );
CLKBUF_X2 inst_11850 ( .A(net_11811), .Z(net_11812) );
CLKBUF_X2 inst_12598 ( .A(net_12559), .Z(net_12560) );
CLKBUF_X2 inst_11314 ( .A(net_11275), .Z(net_11276) );
NAND2_X2 inst_4022 ( .A1(net_6790), .A2(net_1651), .ZN(net_1030) );
SDFFR_X2 inst_1362 ( .SI(net_7744), .Q(net_7744), .D(net_4596), .SE(net_2602), .CK(net_13175), .RN(x1822) );
CLKBUF_X2 inst_13798 ( .A(net_13759), .Z(net_13760) );
CLKBUF_X2 inst_12888 ( .A(net_12849), .Z(net_12850) );
CLKBUF_X2 inst_8881 ( .A(net_8054), .Z(net_8843) );
OAI21_X2 inst_1978 ( .B1(net_4866), .ZN(net_4858), .A(net_4391), .B2(net_3853) );
SDFF_X2 inst_290 ( .Q(net_6365), .SI(net_6364), .D(net_3571), .SE(net_392), .CK(net_13606) );
CLKBUF_X2 inst_14311 ( .A(net_8069), .Z(net_14273) );
SDFF_X2 inst_272 ( .D(net_6399), .SE(net_5801), .SI(net_344), .Q(net_344), .CK(net_13909) );
INV_X4 inst_4718 ( .ZN(net_3026), .A(net_2870) );
CLKBUF_X2 inst_14122 ( .A(net_13973), .Z(net_14084) );
OAI21_X2 inst_2112 ( .ZN(net_3438), .B1(net_3337), .B2(net_2747), .A(net_432) );
AOI21_X2 inst_7743 ( .B1(net_7146), .ZN(net_4070), .B2(net_2582), .A(net_2334) );
NAND2_X2 inst_3036 ( .A1(net_6990), .A2(net_4977), .ZN(net_4971) );
SDFF_X2 inst_814 ( .Q(net_6988), .D(net_6988), .SE(net_3891), .SI(net_3796), .CK(net_11904) );
CLKBUF_X2 inst_13441 ( .A(net_13402), .Z(net_13403) );
CLKBUF_X2 inst_9465 ( .A(net_9426), .Z(net_9427) );
CLKBUF_X2 inst_9213 ( .A(net_9174), .Z(net_9175) );
INV_X4 inst_5203 ( .ZN(net_497), .A(net_496) );
CLKBUF_X2 inst_8973 ( .A(net_8934), .Z(net_8935) );
NAND2_X2 inst_3471 ( .ZN(net_2744), .A1(net_2705), .A2(net_192) );
OAI22_X2 inst_1458 ( .B2(net_5901), .B1(net_4644), .A2(net_4610), .ZN(net_4609), .A1(net_4043) );
NAND2_X2 inst_4133 ( .ZN(net_1259), .A2(net_1225), .A1(net_357) );
CLKBUF_X2 inst_11332 ( .A(net_11293), .Z(net_11294) );
NOR2_X4 inst_2275 ( .ZN(net_5611), .A1(net_5456), .A2(net_4399) );
OAI21_X2 inst_1860 ( .ZN(net_5257), .B1(net_5225), .A(net_4543), .B2(net_3870) );
OAI21_X2 inst_1810 ( .ZN(net_5378), .B1(net_5357), .A(net_4348), .B2(net_3859) );
OAI21_X2 inst_1806 ( .ZN(net_5382), .B1(net_5365), .A(net_4333), .B2(net_3859) );
SDFF_X2 inst_789 ( .SI(net_6919), .Q(net_6919), .D(net_3790), .SE(net_3781), .CK(net_8136) );
OAI21_X2 inst_1885 ( .ZN(net_5197), .B1(net_5196), .A(net_4572), .B2(net_3867) );
CLKBUF_X2 inst_13232 ( .A(net_13193), .Z(net_13194) );
CLKBUF_X2 inst_10212 ( .A(net_10173), .Z(net_10174) );
CLKBUF_X2 inst_11184 ( .A(net_11145), .Z(net_11146) );
CLKBUF_X2 inst_7926 ( .A(net_7887), .Z(net_7888) );
SDFF_X2 inst_822 ( .Q(net_6968), .D(net_6968), .SE(net_3891), .SI(net_3799), .CK(net_11962) );
CLKBUF_X2 inst_14136 ( .A(net_14097), .Z(net_14098) );
CLKBUF_X2 inst_12053 ( .A(net_12014), .Z(net_12015) );
SDFF_X2 inst_1125 ( .SI(net_6675), .Q(net_6675), .D(net_3783), .SE(net_3471), .CK(net_9082) );
NAND2_X1 inst_4341 ( .ZN(net_4386), .A2(net_3856), .A1(net_1749) );
INV_X2 inst_5996 ( .A(net_6005), .ZN(net_2595) );
CLKBUF_X2 inst_13189 ( .A(net_13150), .Z(net_13151) );
INV_X4 inst_4885 ( .ZN(net_2241), .A(net_883) );
CLKBUF_X2 inst_10984 ( .A(net_8701), .Z(net_10946) );
SDFF_X2 inst_609 ( .Q(net_6614), .D(net_6614), .SE(net_3830), .SI(net_3803), .CK(net_10665) );
CLKBUF_X2 inst_11521 ( .A(net_11208), .Z(net_11483) );
NOR2_X2 inst_2496 ( .ZN(net_1746), .A2(net_1745), .A1(net_1266) );
SDFF_X2 inst_795 ( .SI(net_6924), .Q(net_6924), .D(net_3800), .SE(net_3781), .CK(net_8356) );
CLKBUF_X2 inst_8261 ( .A(net_8222), .Z(net_8223) );
CLKBUF_X2 inst_8393 ( .A(net_8354), .Z(net_8355) );
NOR2_X2 inst_2491 ( .ZN(net_2390), .A1(net_2389), .A2(net_2228) );
CLKBUF_X2 inst_13466 ( .A(net_8038), .Z(net_13428) );
NAND2_X1 inst_4381 ( .ZN(net_4346), .A2(net_3859), .A1(net_2053) );
DFF_X1 inst_6668 ( .QN(net_7262), .D(net_5164), .CK(net_13005) );
CLKBUF_X2 inst_14127 ( .A(net_10684), .Z(net_14089) );
CLKBUF_X2 inst_11406 ( .A(net_11367), .Z(net_11368) );
CLKBUF_X2 inst_11179 ( .A(net_11140), .Z(net_11141) );
CLKBUF_X2 inst_12848 ( .A(net_12809), .Z(net_12810) );
CLKBUF_X2 inst_11280 ( .A(net_11241), .Z(net_11242) );
CLKBUF_X2 inst_8215 ( .A(net_8176), .Z(net_8177) );
CLKBUF_X2 inst_8229 ( .A(net_8190), .Z(net_8191) );
SDFF_X2 inst_619 ( .Q(net_6596), .D(net_6596), .SE(net_3830), .SI(net_3798), .CK(net_12904) );
NAND3_X2 inst_2671 ( .ZN(net_3864), .A3(net_3334), .A1(net_2848), .A2(net_2810) );
CLKBUF_X2 inst_9638 ( .A(net_9132), .Z(net_9600) );
CLKBUF_X2 inst_12139 ( .A(net_12100), .Z(net_12101) );
OAI221_X2 inst_1654 ( .ZN(net_4800), .A(net_4595), .C2(net_3979), .B2(net_3968), .C1(net_3773), .B1(net_1968) );
CLKBUF_X2 inst_13068 ( .A(net_13029), .Z(net_13030) );
INV_X8 inst_4547 ( .ZN(net_2131), .A(net_918) );
AND2_X4 inst_7831 ( .ZN(net_3013), .A2(net_2816), .A1(net_2246) );
SDFFR_X2 inst_1355 ( .D(net_3810), .SE(net_3297), .SI(net_285), .Q(net_285), .CK(net_9552), .RN(x1822) );
CLKBUF_X2 inst_10545 ( .A(net_10506), .Z(net_10507) );
SDFF_X2 inst_877 ( .SI(net_7036), .Q(net_7036), .D(net_3814), .SE(net_3777), .CK(net_8203) );
DFF_X1 inst_6612 ( .QN(net_7573), .D(net_5395), .CK(net_8041) );
CLKBUF_X2 inst_10553 ( .A(net_10514), .Z(net_10515) );
CLKBUF_X2 inst_10267 ( .A(net_10228), .Z(net_10229) );
CLKBUF_X2 inst_10704 ( .A(net_9631), .Z(net_10666) );
DFF_X1 inst_6563 ( .QN(net_7499), .D(net_5111), .CK(net_12096) );
CLKBUF_X2 inst_12698 ( .A(net_11915), .Z(net_12660) );
AOI22_X2 inst_7372 ( .A2(net_5916), .B2(net_2957), .ZN(net_2950), .B1(net_2949), .A1(net_842) );
CLKBUF_X2 inst_10265 ( .A(net_9407), .Z(net_10227) );
DFF_X1 inst_6486 ( .QN(net_7417), .D(net_5566), .CK(net_9688) );
OAI21_X2 inst_2076 ( .B2(net_4415), .ZN(net_4414), .B1(net_4032), .A(net_3512) );
INV_X2 inst_5879 ( .A(net_7436), .ZN(net_1471) );
DFF_X1 inst_6384 ( .QN(net_6115), .D(net_5704), .CK(net_8387) );
NOR2_X2 inst_2481 ( .A2(net_5778), .ZN(net_2646), .A1(net_2600) );
AND2_X4 inst_7824 ( .ZN(net_3116), .A2(net_3043), .A1(net_1249) );
CLKBUF_X2 inst_11474 ( .A(net_8879), .Z(net_11436) );
INV_X2 inst_5829 ( .ZN(net_922), .A(net_921) );
CLKBUF_X2 inst_13385 ( .A(net_13346), .Z(net_13347) );
NAND2_X1 inst_4285 ( .ZN(net_4582), .A2(net_3867), .A1(net_1885) );
SDFF_X2 inst_1162 ( .SI(net_6798), .Q(net_6798), .D(net_3814), .SE(net_3722), .CK(net_11058) );
CLKBUF_X2 inst_10274 ( .A(net_10235), .Z(net_10236) );
INV_X2 inst_5904 ( .A(net_7658), .ZN(net_1905) );
AOI222_X2 inst_7485 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2122), .A1(net_2121), .B1(net_2120), .C1(net_2119) );
CLKBUF_X2 inst_14384 ( .A(net_14345), .Z(net_14346) );
INV_X2 inst_6108 ( .A(net_7507), .ZN(net_2196) );
DFF_X1 inst_6572 ( .QN(net_7562), .D(net_5082), .CK(net_10596) );
CLKBUF_X2 inst_13123 ( .A(net_13084), .Z(net_13085) );
AOI22_X2 inst_7449 ( .A2(net_2685), .B2(net_2655), .ZN(net_846), .A1(net_845), .B1(net_844) );
CLKBUF_X2 inst_10734 ( .A(net_10337), .Z(net_10696) );
NAND2_X2 inst_2973 ( .ZN(net_5495), .A2(net_5255), .A1(net_410) );
CLKBUF_X2 inst_11013 ( .A(net_9984), .Z(net_10975) );
CLKBUF_X2 inst_11454 ( .A(net_8852), .Z(net_11416) );
OAI22_X2 inst_1433 ( .B1(net_5856), .ZN(net_5796), .A2(net_5788), .B2(net_5787), .A1(net_5772) );
SDFF_X2 inst_793 ( .SI(net_6895), .Q(net_6895), .D(net_3802), .SE(net_3781), .CK(net_11798) );
CLKBUF_X2 inst_9206 ( .A(net_9167), .Z(net_9168) );
OAI21_X2 inst_1894 ( .B1(net_5220), .ZN(net_5187), .A(net_4563), .B2(net_3866) );
CLKBUF_X2 inst_13960 ( .A(net_13921), .Z(net_13922) );
INV_X4 inst_4815 ( .ZN(net_4797), .A(net_1163) );
DFF_X1 inst_6707 ( .QN(net_7291), .D(net_5367), .CK(net_12986) );
OAI21_X2 inst_1999 ( .B2(net_4518), .ZN(net_4514), .B1(net_4131), .A(net_3694) );
INV_X4 inst_4643 ( .ZN(net_4179), .A(net_4017) );
CLKBUF_X2 inst_14379 ( .A(net_14340), .Z(net_14341) );
NAND3_X2 inst_2733 ( .ZN(net_2368), .A3(net_1627), .A1(net_1487), .A2(net_1024) );
CLKBUF_X2 inst_12405 ( .A(net_12366), .Z(net_12367) );
CLKBUF_X2 inst_11750 ( .A(net_11711), .Z(net_11712) );
DFF_X1 inst_6636 ( .QN(net_7592), .D(net_5246), .CK(net_13158) );
CLKBUF_X2 inst_13677 ( .A(net_11544), .Z(net_13639) );
CLKBUF_X2 inst_8808 ( .A(net_8769), .Z(net_8770) );
SDFF_X2 inst_475 ( .Q(net_7141), .D(net_7141), .SE(net_3903), .SI(net_3894), .CK(net_7895) );
CLKBUF_X2 inst_13253 ( .A(net_13214), .Z(net_13215) );
CLKBUF_X2 inst_9436 ( .A(net_8213), .Z(net_9398) );
INV_X4 inst_4738 ( .A(net_5970), .ZN(net_3876) );
CLKBUF_X2 inst_9412 ( .A(net_9373), .Z(net_9374) );
NAND3_X2 inst_2701 ( .ZN(net_2691), .A3(net_2566), .A2(net_2426), .A1(net_2265) );
NAND2_X1 inst_4412 ( .A2(net_5978), .A1(net_5977), .ZN(net_2880) );
CLKBUF_X2 inst_9171 ( .A(net_8882), .Z(net_9133) );
CLKBUF_X2 inst_8321 ( .A(net_8276), .Z(net_8283) );
CLKBUF_X2 inst_12595 ( .A(net_12033), .Z(net_12557) );
CLKBUF_X2 inst_10385 ( .A(net_10346), .Z(net_10347) );
NAND2_X2 inst_3165 ( .ZN(net_4768), .A2(net_3941), .A1(net_1993) );
CLKBUF_X2 inst_9564 ( .A(net_9525), .Z(net_9526) );
CLKBUF_X2 inst_12804 ( .A(net_12765), .Z(net_12766) );
CLKBUF_X2 inst_11222 ( .A(net_11017), .Z(net_11184) );
SDFF_X2 inst_575 ( .Q(net_6571), .D(net_6571), .SE(net_3823), .SI(net_3812), .CK(net_12928) );
CLKBUF_X2 inst_11738 ( .A(net_11699), .Z(net_11700) );
INV_X2 inst_5724 ( .ZN(net_4004), .A(net_3912) );
CLKBUF_X2 inst_10151 ( .A(net_9252), .Z(net_10113) );
CLKBUF_X2 inst_8276 ( .A(net_8237), .Z(net_8238) );
NAND2_X1 inst_4331 ( .ZN(net_4533), .A2(net_3870), .A1(net_2089) );
CLKBUF_X2 inst_11054 ( .A(net_11015), .Z(net_11016) );
CLKBUF_X2 inst_8049 ( .A(net_8010), .Z(net_8011) );
INV_X4 inst_4705 ( .ZN(net_3258), .A(net_3007) );
CLKBUF_X2 inst_10940 ( .A(net_7896), .Z(net_10902) );
SDFF_X2 inst_627 ( .SI(net_6638), .Q(net_6638), .SE(net_3850), .D(net_3787), .CK(net_7874) );
INV_X4 inst_4725 ( .A(net_5979), .ZN(net_3045) );
DFF_X1 inst_6831 ( .D(net_2588), .QN(net_262), .CK(net_10815) );
NAND2_X2 inst_3352 ( .ZN(net_3543), .A1(net_3542), .A2(net_3226) );
SDFF_X2 inst_344 ( .SI(net_7339), .Q(net_7339), .D(net_4875), .SE(net_3856), .CK(net_9482) );
CLKBUF_X2 inst_11543 ( .A(net_11504), .Z(net_11505) );
DFF_X1 inst_6928 ( .D(net_2416), .Q(net_242), .CK(net_13036) );
NAND2_X2 inst_3580 ( .ZN(net_2432), .A2(net_2431), .A1(net_699) );
NAND2_X2 inst_3818 ( .A1(net_6642), .A2(net_1624), .ZN(net_1527) );
CLKBUF_X2 inst_12321 ( .A(net_12282), .Z(net_12283) );
INV_X2 inst_5975 ( .A(net_7476), .ZN(net_2203) );
SDFFR_X2 inst_1338 ( .Q(net_7715), .D(net_7715), .SI(net_3796), .SE(net_3405), .CK(net_10719), .RN(x1822) );
CLKBUF_X2 inst_11531 ( .A(net_11492), .Z(net_11493) );
CLKBUF_X2 inst_10004 ( .A(net_8938), .Z(net_9966) );
NOR2_X2 inst_2430 ( .ZN(net_3420), .A2(net_3120), .A1(net_3052) );
NAND2_X2 inst_3080 ( .A1(net_6448), .A2(net_4925), .ZN(net_4923) );
DFF_X1 inst_6857 ( .D(net_2537), .QN(net_221), .CK(net_9738) );
CLKBUF_X2 inst_13093 ( .A(net_8571), .Z(net_13055) );
NOR2_X2 inst_2434 ( .ZN(net_3419), .A1(net_3052), .A2(net_3051) );
INV_X4 inst_4952 ( .ZN(net_3985), .A(net_732) );
AOI22_X2 inst_7432 ( .A1(net_2970), .B1(net_2772), .ZN(net_2760), .A2(net_234), .B2(net_160) );
NAND2_X2 inst_3731 ( .A1(net_7177), .A2(net_1637), .ZN(net_1614) );
SDFF_X2 inst_1107 ( .SI(net_6682), .Q(net_6682), .D(net_3789), .SE(net_3471), .CK(net_12005) );
CLKBUF_X2 inst_13932 ( .A(net_13893), .Z(net_13894) );
CLKBUF_X2 inst_10039 ( .A(net_8038), .Z(net_10001) );
DFF_X1 inst_6899 ( .D(net_2508), .QN(net_180), .CK(net_9423) );
OAI21_X2 inst_2028 ( .B2(net_4476), .ZN(net_4475), .B1(net_4230), .A(net_3610) );
INV_X4 inst_4839 ( .ZN(net_5095), .A(net_1070) );
CLKBUF_X2 inst_12909 ( .A(net_12870), .Z(net_12871) );
INV_X2 inst_5930 ( .A(net_7751), .ZN(net_5875) );
CLKBUF_X2 inst_9916 ( .A(net_9877), .Z(net_9878) );
CLKBUF_X2 inst_8381 ( .A(net_8052), .Z(net_8343) );
NAND2_X1 inst_4253 ( .ZN(net_4673), .A2(net_3988), .A1(net_2140) );
NAND3_X2 inst_2776 ( .ZN(net_2324), .A3(net_1548), .A1(net_1349), .A2(net_978) );
SDFF_X2 inst_722 ( .D(net_7802), .SI(net_6767), .Q(net_6767), .SE(net_3816), .CK(net_8273) );
CLKBUF_X2 inst_9646 ( .A(net_9607), .Z(net_9608) );
CLKBUF_X2 inst_8612 ( .A(net_8573), .Z(net_8574) );
SDFF_X2 inst_746 ( .SI(net_7799), .Q(net_6835), .D(net_6835), .SE(net_3893), .CK(net_11812) );
INV_X2 inst_6019 ( .A(net_7586), .ZN(net_2146) );
CLKBUF_X2 inst_8093 ( .A(net_8054), .Z(net_8055) );
CLKBUF_X2 inst_13016 ( .A(net_12977), .Z(net_12978) );
DFF_X1 inst_6553 ( .QN(net_7275), .D(net_5117), .CK(net_9549) );
CLKBUF_X2 inst_9502 ( .A(net_9463), .Z(net_9464) );
NAND2_X1 inst_4232 ( .ZN(net_4695), .A2(net_3989), .A1(net_2219) );
CLKBUF_X2 inst_8660 ( .A(net_7922), .Z(net_8622) );
NOR2_X4 inst_2267 ( .ZN(net_5619), .A1(net_5464), .A2(net_4413) );
NAND2_X1 inst_4270 ( .ZN(net_4646), .A2(net_3993), .A1(net_1411) );
NAND2_X2 inst_3010 ( .A1(net_6887), .A2(net_5006), .ZN(net_4999) );
CLKBUF_X2 inst_8010 ( .A(net_7971), .Z(net_7972) );
DFFR_X1 inst_7127 ( .D(net_3371), .Q(net_275), .CK(net_12805), .RN(x1822) );
CLKBUF_X2 inst_12282 ( .A(net_12243), .Z(net_12244) );
NAND2_X2 inst_3133 ( .ZN(net_4830), .A2(net_4153), .A1(net_2220) );
INV_X4 inst_5662 ( .A(net_7510), .ZN(net_2083) );
CLKBUF_X2 inst_8207 ( .A(net_8168), .Z(net_8169) );
DFF_X1 inst_6412 ( .QN(net_6159), .D(net_5758), .CK(net_11050) );
CLKBUF_X2 inst_7893 ( .A(net_7829), .Z(net_7855) );
CLKBUF_X2 inst_10050 ( .A(net_10011), .Z(net_10012) );
INV_X2 inst_5820 ( .ZN(net_1049), .A(net_1048) );
CLKBUF_X2 inst_8721 ( .A(net_8682), .Z(net_8683) );
OAI22_X2 inst_1577 ( .A2(net_3297), .B2(net_3286), .ZN(net_3267), .A1(net_3194), .B1(net_422) );
AOI21_X2 inst_7722 ( .B1(net_6738), .ZN(net_4128), .B2(net_2581), .A(net_2370) );
NAND3_X2 inst_2588 ( .ZN(net_5751), .A1(net_5646), .A2(net_5250), .A3(net_4210) );
SDFF_X2 inst_1110 ( .SI(net_6678), .Q(net_6678), .D(net_3780), .SE(net_3465), .CK(net_10618) );
INV_X2 inst_5778 ( .ZN(net_2895), .A(net_192) );
DFF_X1 inst_6547 ( .Q(net_7772), .D(net_5610), .CK(net_10429) );
NAND2_X4 inst_2873 ( .A1(net_5886), .ZN(net_4266), .A2(net_1100) );
AOI21_X2 inst_7724 ( .B1(net_6464), .ZN(net_4061), .B2(net_2580), .A(net_2326) );
DFFR_X2 inst_6994 ( .QN(net_7702), .D(net_3361), .CK(net_10366), .RN(x1822) );
INV_X4 inst_4665 ( .ZN(net_4301), .A(net_3865) );
CLKBUF_X2 inst_8468 ( .A(net_8359), .Z(net_8430) );
NOR2_X2 inst_2442 ( .A2(net_5979), .ZN(net_3162), .A1(net_3002) );
CLKBUF_X2 inst_9676 ( .A(net_9637), .Z(net_9638) );
OAI21_X2 inst_2066 ( .B2(net_4436), .ZN(net_4429), .B1(net_4049), .A(net_3543) );
CLKBUF_X2 inst_12126 ( .A(net_12087), .Z(net_12088) );
INV_X2 inst_5712 ( .ZN(net_4254), .A(net_4129) );
OAI21_X2 inst_1742 ( .ZN(net_5532), .A(net_4825), .B2(net_4153), .B1(net_1166) );
INV_X8 inst_4466 ( .ZN(net_5183), .A(net_4285) );
INV_X4 inst_5374 ( .A(net_7405), .ZN(net_2121) );
INV_X4 inst_5562 ( .A(net_7717), .ZN(net_859) );
CLKBUF_X2 inst_12085 ( .A(net_12046), .Z(net_12047) );
CLKBUF_X2 inst_11058 ( .A(net_11019), .Z(net_11020) );
CLKBUF_X2 inst_13603 ( .A(net_13206), .Z(net_13565) );
CLKBUF_X2 inst_12091 ( .A(net_12052), .Z(net_12053) );
CLKBUF_X2 inst_11035 ( .A(net_10996), .Z(net_10997) );
DFF_X2 inst_6236 ( .Q(net_6390), .D(net_6389), .CK(net_14342) );
CLKBUF_X2 inst_8447 ( .A(net_8408), .Z(net_8409) );
NAND2_X4 inst_2875 ( .A1(net_4276), .ZN(net_4264), .A2(net_1675) );
INV_X4 inst_4779 ( .ZN(net_1832), .A(net_1664) );
CLKBUF_X2 inst_9522 ( .A(net_9483), .Z(net_9484) );
CLKBUF_X2 inst_9067 ( .A(net_9028), .Z(net_9029) );
CLKBUF_X2 inst_11084 ( .A(net_11045), .Z(net_11046) );
CLKBUF_X2 inst_10341 ( .A(net_9530), .Z(net_10303) );
CLKBUF_X2 inst_9396 ( .A(net_9357), .Z(net_9358) );
NAND2_X2 inst_3175 ( .ZN(net_4758), .A2(net_3941), .A1(net_2043) );
NOR2_X2 inst_2302 ( .A2(net_6185), .A1(net_5843), .ZN(net_5839) );
CLKBUF_X2 inst_11021 ( .A(net_8221), .Z(net_10983) );
NAND2_X2 inst_3389 ( .ZN(net_3772), .A2(net_3368), .A1(net_2893) );
DFF_X2 inst_6248 ( .QN(net_7755), .D(net_3023), .CK(net_8564) );
CLKBUF_X2 inst_9967 ( .A(net_9928), .Z(net_9929) );
NOR2_X2 inst_2447 ( .ZN(net_2869), .A1(net_2868), .A2(net_2867) );
SDFF_X2 inst_782 ( .SI(net_6910), .Q(net_6910), .SE(net_3887), .D(net_3808), .CK(net_8865) );
INV_X2 inst_5744 ( .ZN(net_3720), .A(net_3417) );
CLKBUF_X2 inst_12043 ( .A(net_12004), .Z(net_12005) );
NAND2_X4 inst_2869 ( .A1(net_4282), .ZN(net_4270), .A2(net_1497) );
CLKBUF_X2 inst_10546 ( .A(net_9808), .Z(net_10508) );
CLKBUF_X2 inst_10603 ( .A(net_8933), .Z(net_10565) );
XOR2_X2 inst_6 ( .Z(net_1203), .B(net_899), .A(net_642) );
NOR2_X2 inst_2486 ( .A2(net_5778), .ZN(net_2660), .A1(net_2594) );
CLKBUF_X2 inst_11648 ( .A(net_11609), .Z(net_11610) );
INV_X4 inst_5461 ( .ZN(net_3341), .A(net_153) );
NOR2_X2 inst_2410 ( .ZN(net_3732), .A2(net_3437), .A1(net_2703) );
CLKBUF_X2 inst_11151 ( .A(net_11112), .Z(net_11113) );
CLKBUF_X2 inst_11832 ( .A(net_11793), .Z(net_11794) );
CLKBUF_X2 inst_10914 ( .A(net_10875), .Z(net_10876) );
CLKBUF_X2 inst_9695 ( .A(net_8171), .Z(net_9657) );
CLKBUF_X2 inst_8927 ( .A(net_8888), .Z(net_8889) );
AOI21_X4 inst_7622 ( .B2(net_5955), .B1(net_5954), .ZN(net_5605), .A(x906) );
CLKBUF_X2 inst_8728 ( .A(net_8689), .Z(net_8690) );
INV_X16 inst_6141 ( .ZN(net_1624), .A(net_813) );
CLKBUF_X2 inst_7921 ( .A(net_7882), .Z(net_7883) );
CLKBUF_X2 inst_13303 ( .A(net_13264), .Z(net_13265) );
CLKBUF_X2 inst_12760 ( .A(net_8573), .Z(net_12722) );
INV_X4 inst_4803 ( .ZN(net_4793), .A(net_1183) );
SDFF_X2 inst_935 ( .D(net_7807), .SI(net_7177), .Q(net_7177), .SE(net_3819), .CK(net_12149) );
DFF_X1 inst_6619 ( .QN(net_7580), .D(net_5388), .CK(net_13162) );
CLKBUF_X2 inst_11726 ( .A(net_11687), .Z(net_11688) );
INV_X4 inst_5699 ( .A(net_5934), .ZN(net_5933) );
CLKBUF_X2 inst_13030 ( .A(net_12991), .Z(net_12992) );
INV_X4 inst_4772 ( .ZN(net_1724), .A(net_1723) );
CLKBUF_X2 inst_12781 ( .A(net_12742), .Z(net_12743) );
INV_X4 inst_4634 ( .ZN(net_4188), .A(net_4037) );
CLKBUF_X2 inst_8108 ( .A(net_7977), .Z(net_8070) );
CLKBUF_X2 inst_8211 ( .A(net_7930), .Z(net_8173) );
INV_X2 inst_6031 ( .ZN(net_3077), .A(net_295) );
CLKBUF_X2 inst_11255 ( .A(net_11216), .Z(net_11217) );
AOI21_X2 inst_7729 ( .B1(net_6468), .ZN(net_4053), .B2(net_2580), .A(net_2378) );
CLKBUF_X2 inst_9284 ( .A(net_7960), .Z(net_9246) );
CLKBUF_X2 inst_11587 ( .A(net_8396), .Z(net_11549) );
NAND2_X2 inst_2944 ( .ZN(net_5502), .A1(net_4964), .A2(net_4963) );
SDFF_X2 inst_1320 ( .D(net_6385), .SE(net_5799), .SI(net_370), .Q(net_370), .CK(net_13857) );
SDFF_X2 inst_1026 ( .D(net_7799), .SI(net_6494), .Q(net_6494), .SE(net_3886), .CK(net_8632) );
INV_X4 inst_5011 ( .ZN(net_730), .A(net_677) );
CLKBUF_X2 inst_11289 ( .A(net_11250), .Z(net_11251) );
DFF_X2 inst_6250 ( .Q(net_6389), .D(net_6388), .CK(net_14250) );
CLKBUF_X2 inst_12826 ( .A(net_12787), .Z(net_12788) );
INV_X4 inst_5576 ( .A(net_6124), .ZN(net_3667) );
NAND2_X2 inst_3376 ( .ZN(net_3494), .A1(net_3493), .A2(net_3223) );
XNOR2_X2 inst_95 ( .B(net_3003), .ZN(net_1663), .A(net_1150) );
INV_X4 inst_5246 ( .ZN(net_3000), .A(net_445) );
NAND2_X2 inst_2921 ( .A2(net_7775), .ZN(net_5771), .A1(net_5607) );
CLKBUF_X2 inst_13690 ( .A(net_13651), .Z(net_13652) );
CLKBUF_X2 inst_13058 ( .A(net_13019), .Z(net_13020) );
CLKBUF_X2 inst_10622 ( .A(net_10583), .Z(net_10584) );
CLKBUF_X2 inst_10499 ( .A(net_8839), .Z(net_10461) );
CLKBUF_X2 inst_8314 ( .A(net_8275), .Z(net_8276) );
NAND2_X4 inst_2862 ( .ZN(net_4289), .A1(net_4282), .A2(net_1651) );
CLKBUF_X2 inst_7949 ( .A(net_7910), .Z(net_7911) );
CLKBUF_X2 inst_8391 ( .A(net_8352), .Z(net_8353) );
NAND2_X2 inst_4009 ( .ZN(net_1255), .A2(net_1225), .A1(net_356) );
CLKBUF_X2 inst_13397 ( .A(net_12321), .Z(net_13359) );
CLKBUF_X2 inst_10870 ( .A(net_10831), .Z(net_10832) );
CLKBUF_X2 inst_9766 ( .A(net_9727), .Z(net_9728) );
CLKBUF_X2 inst_8071 ( .A(net_8032), .Z(net_8033) );
CLKBUF_X2 inst_8297 ( .A(net_8258), .Z(net_8259) );
INV_X4 inst_4900 ( .A(net_3900), .ZN(net_3139) );
DFF_X1 inst_6510 ( .QN(net_7432), .D(net_5511), .CK(net_12621) );
CLKBUF_X2 inst_13325 ( .A(net_12647), .Z(net_13287) );
INV_X2 inst_5808 ( .A(net_1693), .ZN(net_1209) );
INV_X4 inst_5394 ( .A(net_6000), .ZN(net_541) );
INV_X2 inst_5837 ( .ZN(net_806), .A(net_805) );
CLKBUF_X2 inst_13883 ( .A(net_9152), .Z(net_13845) );
CLKBUF_X2 inst_12181 ( .A(net_12142), .Z(net_12143) );
CLKBUF_X2 inst_13390 ( .A(net_13257), .Z(net_13352) );
CLKBUF_X2 inst_11268 ( .A(net_8746), .Z(net_11230) );
DFF_X1 inst_6859 ( .D(net_2542), .Q(net_196), .CK(net_9735) );
AOI22_X2 inst_7439 ( .ZN(net_4872), .A2(net_1222), .B1(net_1220), .B2(net_344), .A1(net_332) );
AOI222_X2 inst_7537 ( .C1(net_7672), .A1(net_7640), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1890), .B1(net_1889) );
CLKBUF_X2 inst_10407 ( .A(net_10368), .Z(net_10369) );
NAND2_X1 inst_4454 ( .A2(net_1256), .ZN(net_1122), .A1(net_1121) );
CLKBUF_X2 inst_12369 ( .A(net_11487), .Z(net_12331) );
CLKBUF_X2 inst_8955 ( .A(net_8916), .Z(net_8917) );
INV_X4 inst_4901 ( .ZN(net_1308), .A(net_868) );
CLKBUF_X2 inst_12813 ( .A(net_10679), .Z(net_12775) );
NAND2_X2 inst_3590 ( .ZN(net_2410), .A2(net_1853), .A1(net_1390) );
CLKBUF_X2 inst_8709 ( .A(net_8670), .Z(net_8671) );
NAND2_X1 inst_4315 ( .ZN(net_4549), .A2(net_3870), .A1(net_2127) );
SDFF_X2 inst_365 ( .SI(net_7615), .Q(net_7615), .D(net_4793), .SE(net_3870), .CK(net_7994) );
XNOR2_X2 inst_67 ( .ZN(net_2474), .A(net_1087), .B(net_595) );
SDFF_X2 inst_954 ( .D(net_7799), .SI(net_7169), .Q(net_7169), .SE(net_3817), .CK(net_13330) );
CLKBUF_X2 inst_13162 ( .A(net_13123), .Z(net_13124) );
CLKBUF_X2 inst_9252 ( .A(net_9213), .Z(net_9214) );
CLKBUF_X2 inst_8145 ( .A(net_8106), .Z(net_8107) );
INV_X4 inst_4974 ( .ZN(net_882), .A(net_691) );
CLKBUF_X2 inst_10836 ( .A(net_9902), .Z(net_10798) );
CLKBUF_X2 inst_8582 ( .A(net_8543), .Z(net_8544) );
CLKBUF_X2 inst_14186 ( .A(net_14147), .Z(net_14148) );
CLKBUF_X2 inst_11216 ( .A(net_11177), .Z(net_11178) );
CLKBUF_X2 inst_8569 ( .A(net_8530), .Z(net_8531) );
NOR2_X2 inst_2476 ( .A2(net_5778), .ZN(net_2604), .A1(net_517) );
CLKBUF_X2 inst_11685 ( .A(net_11646), .Z(net_11647) );
CLKBUF_X2 inst_12078 ( .A(net_12039), .Z(net_12040) );
OAI21_X2 inst_1823 ( .ZN(net_5364), .B1(net_5363), .A(net_4383), .B2(net_3856) );
INV_X4 inst_5084 ( .A(net_3236), .ZN(net_627) );
SDFF_X2 inst_202 ( .Q(net_6312), .SI(net_6311), .D(net_3697), .SE(net_392), .CK(net_13575) );
CLKBUF_X2 inst_8116 ( .A(net_8077), .Z(net_8078) );
AOI22_X2 inst_7359 ( .B2(net_3105), .ZN(net_3032), .A2(net_2712), .A1(net_1113), .B1(net_606) );
CLKBUF_X2 inst_9154 ( .A(net_8428), .Z(net_9116) );
NOR3_X2 inst_2212 ( .ZN(net_2264), .A3(net_1207), .A1(net_408), .A2(x1155) );
CLKBUF_X2 inst_13786 ( .A(net_12170), .Z(net_13748) );
OR2_X4 inst_1401 ( .A1(net_7530), .A2(net_7529), .ZN(net_690) );
INV_X8 inst_4502 ( .ZN(net_3872), .A(net_3262) );
INV_X4 inst_4830 ( .ZN(net_1080), .A(net_1079) );
CLKBUF_X2 inst_14258 ( .A(net_11507), .Z(net_14220) );
CLKBUF_X2 inst_13444 ( .A(net_11398), .Z(net_13406) );
OAI21_X2 inst_2030 ( .B2(net_4476), .ZN(net_4473), .B1(net_4231), .A(net_3604) );
INV_X4 inst_5624 ( .A(net_6109), .ZN(net_3677) );
CLKBUF_X2 inst_8254 ( .A(net_8083), .Z(net_8216) );
AOI22_X2 inst_7451 ( .B2(net_2847), .A2(net_2661), .ZN(net_840), .A1(net_839), .B1(net_838) );
CLKBUF_X2 inst_11172 ( .A(net_11133), .Z(net_11134) );
AOI222_X2 inst_7458 ( .A1(net_7714), .A2(net_5916), .C2(net_3439), .ZN(net_2977), .B1(net_2970), .C1(net_296), .B2(net_253) );
CLKBUF_X2 inst_14072 ( .A(net_14033), .Z(net_14034) );
XNOR2_X2 inst_30 ( .ZN(net_2483), .A(net_2482), .B(net_913) );
SDFF_X2 inst_610 ( .Q(net_6615), .D(net_6615), .SE(net_3830), .SI(net_3796), .CK(net_7879) );
SDFF_X2 inst_1036 ( .Q(net_7538), .D(net_7538), .SE(net_3896), .SI(net_372), .CK(net_10265) );
DFF_X2 inst_6271 ( .QN(net_6413), .D(net_2690), .CK(net_10205) );
SDFF_X2 inst_233 ( .Q(net_6321), .SI(net_6320), .D(net_3643), .SE(net_392), .CK(net_14008) );
CLKBUF_X2 inst_9704 ( .A(net_9665), .Z(net_9666) );
CLKBUF_X2 inst_8639 ( .A(net_7831), .Z(net_8601) );
CLKBUF_X2 inst_10094 ( .A(net_8512), .Z(net_10056) );
CLKBUF_X2 inst_8595 ( .A(net_8273), .Z(net_8557) );
CLKBUF_X2 inst_10334 ( .A(net_10295), .Z(net_10296) );
CLKBUF_X2 inst_12296 ( .A(net_12257), .Z(net_12258) );
CLKBUF_X2 inst_9527 ( .A(net_9488), .Z(net_9489) );
CLKBUF_X2 inst_9127 ( .A(net_9088), .Z(net_9089) );
CLKBUF_X2 inst_8653 ( .A(net_7949), .Z(net_8615) );
XNOR2_X2 inst_60 ( .B(net_3940), .ZN(net_1925), .A(net_1687) );
INV_X4 inst_5694 ( .A(net_7578), .ZN(net_1848) );
CLKBUF_X2 inst_8939 ( .A(net_8560), .Z(net_8901) );
DFF_X1 inst_6651 ( .QN(net_7648), .D(net_5195), .CK(net_12264) );
CLKBUF_X2 inst_13540 ( .A(net_13501), .Z(net_13502) );
CLKBUF_X2 inst_12141 ( .A(net_8968), .Z(net_12103) );
INV_X4 inst_4613 ( .ZN(net_4209), .A(net_4081) );
INV_X2 inst_5852 ( .ZN(net_674), .A(net_673) );
AOI21_X2 inst_7752 ( .B1(net_6874), .ZN(net_4099), .B2(net_2579), .A(net_2351) );
NOR2_X2 inst_2376 ( .ZN(net_5153), .A2(net_4608), .A1(net_4423) );
CLKBUF_X2 inst_13285 ( .A(net_13246), .Z(net_13247) );
AOI222_X2 inst_7496 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2086), .A1(net_2085), .B1(net_2084), .C1(net_2083) );
CLKBUF_X2 inst_7925 ( .A(net_7868), .Z(net_7887) );
CLKBUF_X2 inst_12862 ( .A(net_12823), .Z(net_12824) );
NAND2_X1 inst_4360 ( .ZN(net_4367), .A2(net_3853), .A1(net_2050) );
DFFR_X2 inst_7050 ( .QN(net_6020), .D(net_3202), .CK(net_8591), .RN(x1822) );
AOI22_X2 inst_7339 ( .B2(net_3439), .ZN(net_3303), .A2(net_2712), .B1(net_737), .A1(net_151) );
CLKBUF_X2 inst_12189 ( .A(net_12150), .Z(net_12151) );
SDFF_X2 inst_860 ( .SI(net_7045), .Q(net_7045), .SE(net_3818), .D(net_3776), .CK(net_11879) );
SDFF_X2 inst_563 ( .SI(net_7181), .Q(net_7181), .D(net_3831), .SE(net_3817), .CK(net_7920) );
CLKBUF_X2 inst_14074 ( .A(net_14035), .Z(net_14036) );
NAND2_X2 inst_3962 ( .A1(net_6836), .A2(net_1521), .ZN(net_1322) );
CLKBUF_X2 inst_10392 ( .A(net_7887), .Z(net_10354) );
CLKBUF_X2 inst_8389 ( .A(net_8350), .Z(net_8351) );
SDFF_X2 inst_943 ( .SI(net_7186), .Q(net_7186), .SE(net_3817), .D(net_3803), .CK(net_8699) );
CLKBUF_X2 inst_14397 ( .A(net_9928), .Z(net_14359) );
NAND2_X2 inst_3478 ( .ZN(net_2686), .A1(net_2685), .A2(net_2684) );
CLKBUF_X2 inst_11252 ( .A(net_11213), .Z(net_11214) );
CLKBUF_X2 inst_10181 ( .A(net_7861), .Z(net_10143) );
INV_X4 inst_5314 ( .ZN(net_1657), .A(x1322) );
NAND3_X2 inst_2782 ( .ZN(net_2318), .A3(net_1611), .A1(net_1336), .A2(net_965) );
INV_X4 inst_4711 ( .ZN(net_3124), .A(net_3049) );
AOI22_X2 inst_7248 ( .B1(net_6816), .A1(net_6784), .A2(net_5316), .B2(net_5315), .ZN(net_5312) );
CLKBUF_X2 inst_12151 ( .A(net_12112), .Z(net_12113) );
OAI21_X2 inst_1964 ( .B1(net_5412), .ZN(net_5046), .A(net_4653), .B2(net_3993) );
OAI21_X2 inst_1765 ( .B1(net_5548), .ZN(net_5429), .A(net_4646), .B2(net_3993) );
AOI222_X2 inst_7464 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2195), .A1(net_2194), .B1(net_2193), .C1(net_2192) );
INV_X4 inst_5475 ( .A(net_7535), .ZN(net_835) );
CLKBUF_X2 inst_13887 ( .A(net_10975), .Z(net_13849) );
CLKBUF_X2 inst_11191 ( .A(net_11152), .Z(net_11153) );
NAND2_X2 inst_3720 ( .A1(net_6773), .A2(net_1635), .ZN(net_1626) );
CLKBUF_X2 inst_11964 ( .A(net_11925), .Z(net_11926) );
CLKBUF_X2 inst_12444 ( .A(net_12405), .Z(net_12406) );
OAI21_X2 inst_2005 ( .B2(net_4518), .ZN(net_4507), .B1(net_4506), .A(net_3678) );
CLKBUF_X2 inst_11988 ( .A(net_10790), .Z(net_11950) );
CLKBUF_X2 inst_13377 ( .A(net_13338), .Z(net_13339) );
SDFF_X2 inst_736 ( .Q(net_6853), .D(net_6853), .SE(net_3893), .SI(net_3791), .CK(net_8151) );
SDFF_X2 inst_544 ( .Q(net_7138), .D(net_7138), .SE(net_3903), .SI(net_3890), .CK(net_11592) );
CLKBUF_X2 inst_13525 ( .A(net_13486), .Z(net_13487) );
INV_X2 inst_5865 ( .A(net_833), .ZN(net_561) );
CLKBUF_X2 inst_8021 ( .A(net_7982), .Z(net_7983) );
INV_X4 inst_5465 ( .A(net_7094), .ZN(net_569) );
CLKBUF_X2 inst_11944 ( .A(net_8570), .Z(net_11906) );
DFF_X1 inst_6357 ( .QN(net_6201), .D(net_5827), .CK(net_13933) );
CLKBUF_X2 inst_8232 ( .A(net_8128), .Z(net_8194) );
SDFF_X2 inst_178 ( .Q(net_6276), .SI(net_6275), .D(net_3503), .SE(net_392), .CK(net_13482) );
CLKBUF_X2 inst_9179 ( .A(net_8188), .Z(net_9141) );
NAND2_X1 inst_4402 ( .A2(net_3297), .ZN(net_3076), .A1(net_3075) );
SDFF_X2 inst_734 ( .Q(net_6851), .D(net_6851), .SE(net_3893), .SI(net_3804), .CK(net_10901) );
AOI22_X2 inst_7352 ( .B2(net_3105), .ZN(net_3098), .A2(net_2712), .A1(net_1257), .B1(net_442) );
SDFF_X2 inst_1282 ( .D(net_3811), .SE(net_3256), .SI(net_143), .Q(net_143), .CK(net_10695) );
CLKBUF_X2 inst_8528 ( .A(net_8489), .Z(net_8490) );
CLKBUF_X2 inst_8257 ( .A(net_8218), .Z(net_8219) );
INV_X2 inst_5941 ( .A(net_7649), .ZN(net_2100) );
CLKBUF_X2 inst_13562 ( .A(net_12172), .Z(net_13524) );
NAND2_X2 inst_3919 ( .A1(net_7463), .A2(net_1696), .ZN(net_1384) );
SDFF_X2 inst_1148 ( .SI(net_6809), .Q(net_6809), .D(net_3807), .SE(net_3722), .CK(net_11296) );
AOI21_X2 inst_7661 ( .B2(net_5926), .ZN(net_3318), .A(net_3317), .B1(net_1827) );
CLKBUF_X2 inst_10425 ( .A(net_8281), .Z(net_10387) );
CLKBUF_X2 inst_8898 ( .A(net_8859), .Z(net_8860) );
CLKBUF_X2 inst_10292 ( .A(net_10253), .Z(net_10254) );
NAND2_X1 inst_4350 ( .ZN(net_4377), .A2(net_3853), .A1(net_2074) );
CLKBUF_X2 inst_8270 ( .A(net_8231), .Z(net_8232) );
INV_X4 inst_5634 ( .A(net_6415), .ZN(net_2421) );
CLKBUF_X2 inst_9597 ( .A(net_9558), .Z(net_9559) );
NAND2_X2 inst_3587 ( .ZN(net_2413), .A2(net_1915), .A1(net_1514) );
CLKBUF_X2 inst_8777 ( .A(net_8738), .Z(net_8739) );
CLKBUF_X2 inst_10139 ( .A(net_10100), .Z(net_10101) );
CLKBUF_X2 inst_13003 ( .A(net_12964), .Z(net_12965) );
CLKBUF_X2 inst_10147 ( .A(net_10108), .Z(net_10109) );
CLKBUF_X2 inst_9659 ( .A(net_8458), .Z(net_9621) );
INV_X4 inst_5543 ( .ZN(net_1220), .A(net_270) );
INV_X2 inst_6004 ( .A(net_7475), .ZN(net_2197) );
DFF_X1 inst_6392 ( .QN(net_6123), .D(net_5696), .CK(net_8383) );
SDFF_X2 inst_842 ( .Q(net_7023), .D(net_7023), .SE(net_3899), .SI(net_3789), .CK(net_10998) );
INV_X4 inst_5588 ( .A(net_6828), .ZN(net_2575) );
CLKBUF_X2 inst_11427 ( .A(net_11388), .Z(net_11389) );
OAI21_X2 inst_2068 ( .B2(net_4436), .ZN(net_4427), .B1(net_4426), .A(net_3710) );
CLKBUF_X2 inst_9897 ( .A(net_9505), .Z(net_9859) );
DFF_X2 inst_6183 ( .QN(net_6823), .D(net_5454), .CK(net_10802) );
CLKBUF_X2 inst_9697 ( .A(net_9658), .Z(net_9659) );
SDFF_X2 inst_551 ( .Q(net_6427), .D(net_6427), .SI(net_3892), .SE(net_3820), .CK(net_8788) );
OAI21_X2 inst_2101 ( .ZN(net_3984), .B1(net_3983), .B2(net_3982), .A(net_3865) );
CLKBUF_X2 inst_11529 ( .A(net_9829), .Z(net_11491) );
CLKBUF_X2 inst_8542 ( .A(net_8503), .Z(net_8504) );
SDFF_X2 inst_353 ( .SI(net_7605), .Q(net_7605), .D(net_4801), .SE(net_3870), .CK(net_8005) );
NAND2_X2 inst_3808 ( .A1(net_6634), .A2(net_1624), .ZN(net_1537) );
OAI21_X2 inst_1940 ( .B1(net_5539), .ZN(net_5093), .A(net_4737), .B2(net_3988) );
DFF_X2 inst_6286 ( .D(net_2390), .QN(net_189), .CK(net_12287) );
CLKBUF_X2 inst_8492 ( .A(net_8453), .Z(net_8454) );
INV_X4 inst_4632 ( .ZN(net_4190), .A(net_4040) );
CLKBUF_X2 inst_10400 ( .A(net_10361), .Z(net_10362) );
CLKBUF_X2 inst_13456 ( .A(net_13417), .Z(net_13418) );
CLKBUF_X2 inst_13917 ( .A(net_9911), .Z(net_13879) );
DFF_X2 inst_6212 ( .QN(net_7685), .D(net_4108), .CK(net_10793) );
NAND2_X2 inst_4041 ( .A1(net_7197), .A2(net_1648), .ZN(net_1011) );
CLKBUF_X2 inst_13761 ( .A(net_12355), .Z(net_13723) );
NAND2_X2 inst_3701 ( .A1(net_7455), .ZN(net_1697), .A2(net_1696) );
NAND2_X2 inst_3357 ( .ZN(net_3531), .A1(net_3530), .A2(net_3225) );
CLKBUF_X2 inst_9559 ( .A(net_9520), .Z(net_9521) );
CLKBUF_X2 inst_14184 ( .A(net_11758), .Z(net_14146) );
DFFR_X2 inst_7082 ( .QN(net_7735), .D(net_2800), .CK(net_10342), .RN(x1822) );
CLKBUF_X2 inst_11822 ( .A(net_11783), .Z(net_11784) );
XNOR2_X2 inst_8 ( .A(net_4149), .ZN(net_3828), .B(net_875) );
CLKBUF_X2 inst_13869 ( .A(net_13830), .Z(net_13831) );
CLKBUF_X2 inst_11321 ( .A(net_11282), .Z(net_11283) );
DFF_X1 inst_6745 ( .QN(net_7602), .D(net_4854), .CK(net_8030) );
CLKBUF_X2 inst_8925 ( .A(net_8886), .Z(net_8887) );
CLKBUF_X2 inst_14064 ( .A(net_10172), .Z(net_14026) );
DFFR_X2 inst_6984 ( .QN(net_6027), .D(net_3445), .CK(net_10755), .RN(x1822) );
OAI21_X2 inst_2090 ( .B2(net_4508), .ZN(net_4326), .B1(net_4132), .A(net_3704) );
SDFF_X2 inst_965 ( .Q(net_6425), .D(net_6425), .SE(net_3820), .SI(net_3778), .CK(net_11553) );
CLKBUF_X2 inst_13980 ( .A(net_10775), .Z(net_13942) );
CLKBUF_X2 inst_12624 ( .A(net_10344), .Z(net_12586) );
NAND2_X2 inst_3370 ( .ZN(net_3506), .A1(net_3505), .A2(net_3223) );
CLKBUF_X2 inst_8228 ( .A(net_8167), .Z(net_8190) );
CLKBUF_X2 inst_10168 ( .A(net_10129), .Z(net_10130) );
CLKBUF_X2 inst_12267 ( .A(net_12228), .Z(net_12229) );
CLKBUF_X2 inst_8677 ( .A(net_8638), .Z(net_8639) );
CLKBUF_X2 inst_11991 ( .A(net_11952), .Z(net_11953) );
CLKBUF_X2 inst_8993 ( .A(net_8954), .Z(net_8955) );
CLKBUF_X2 inst_12284 ( .A(net_12245), .Z(net_12246) );
CLKBUF_X2 inst_11976 ( .A(net_8814), .Z(net_11938) );
DFF_X1 inst_6579 ( .QN(net_7568), .D(net_5071), .CK(net_13458) );
INV_X4 inst_5392 ( .A(net_6029), .ZN(net_2809) );
SDFF_X2 inst_901 ( .Q(net_7104), .D(net_7104), .SE(net_3888), .SI(net_3798), .CK(net_13368) );
DFF_X2 inst_6179 ( .QN(net_6958), .D(net_5453), .CK(net_11415) );
CLKBUF_X2 inst_10992 ( .A(net_10953), .Z(net_10954) );
INV_X2 inst_6094 ( .A(net_7326), .ZN(net_1751) );
AOI22_X2 inst_7261 ( .B1(net_6952), .A1(net_6920), .A2(net_5298), .B2(net_5297), .ZN(net_5293) );
CLKBUF_X2 inst_13821 ( .A(net_13782), .Z(net_13783) );
CLKBUF_X2 inst_7913 ( .A(net_7849), .Z(net_7875) );
CLKBUF_X2 inst_9957 ( .A(net_9918), .Z(net_9919) );
CLKBUF_X2 inst_13288 ( .A(net_8042), .Z(net_13250) );
CLKBUF_X2 inst_10863 ( .A(net_10824), .Z(net_10825) );
CLKBUF_X2 inst_14013 ( .A(net_13974), .Z(net_13975) );
NOR2_X2 inst_2403 ( .ZN(net_3765), .A1(net_3764), .A2(net_3763) );
INV_X4 inst_4948 ( .A(net_2384), .ZN(net_1941) );
CLKBUF_X2 inst_9104 ( .A(net_9065), .Z(net_9066) );
OAI21_X2 inst_1934 ( .B1(net_5410), .ZN(net_5111), .A(net_4743), .B2(net_3988) );
DFF_X1 inst_6759 ( .QN(net_7333), .D(net_4864), .CK(net_9868) );
CLKBUF_X2 inst_9429 ( .A(net_9390), .Z(net_9391) );
NAND2_X2 inst_3098 ( .A1(net_6477), .A2(net_4927), .ZN(net_4905) );
NAND2_X2 inst_3916 ( .A1(net_6964), .A2(net_1833), .ZN(net_1388) );
INV_X2 inst_5739 ( .ZN(net_3726), .A(net_3430) );
INV_X4 inst_5401 ( .ZN(net_769), .A(x1261) );
CLKBUF_X2 inst_13834 ( .A(net_8439), .Z(net_13796) );
CLKBUF_X2 inst_10679 ( .A(net_8648), .Z(net_10641) );
CLKBUF_X2 inst_9970 ( .A(net_9931), .Z(net_9932) );
CLKBUF_X2 inst_8319 ( .A(net_8265), .Z(net_8281) );
INV_X16 inst_6144 ( .ZN(net_1639), .A(net_773) );
CLKBUF_X2 inst_8539 ( .A(net_8086), .Z(net_8501) );
INV_X4 inst_5013 ( .A(net_7809), .ZN(net_718) );
CLKBUF_X2 inst_13359 ( .A(net_13320), .Z(net_13321) );
CLKBUF_X2 inst_12034 ( .A(net_11995), .Z(net_11996) );
CLKBUF_X2 inst_8464 ( .A(net_8425), .Z(net_8426) );
CLKBUF_X2 inst_10968 ( .A(net_10929), .Z(net_10930) );
OAI21_X2 inst_2097 ( .B2(net_4424), .ZN(net_4319), .B1(net_4057), .A(net_3537) );
CLKBUF_X2 inst_12943 ( .A(net_12265), .Z(net_12905) );
SDFF_X2 inst_928 ( .SI(net_7799), .Q(net_7137), .D(net_7137), .SE(net_3903), .CK(net_11567) );
INV_X8 inst_4484 ( .ZN(net_4278), .A(net_3924) );
INV_X2 inst_5910 ( .ZN(net_410), .A(x868) );
CLKBUF_X2 inst_10695 ( .A(net_10656), .Z(net_10657) );
NAND3_X2 inst_2662 ( .ZN(net_3934), .A3(net_3395), .A2(net_2950), .A1(net_2835) );
OAI22_X2 inst_1539 ( .B1(net_4637), .A1(net_4030), .B2(net_4020), .ZN(net_4017), .A2(net_4016) );
CLKBUF_X2 inst_8053 ( .A(net_8014), .Z(net_8015) );
DFF_X2 inst_6215 ( .Q(net_6393), .D(net_6392), .CK(net_13692) );
OAI21_X2 inst_1718 ( .ZN(net_5576), .B1(net_5542), .A(net_4686), .B2(net_3989) );
CLKBUF_X2 inst_12225 ( .A(net_12186), .Z(net_12187) );
SDFF_X2 inst_1050 ( .Q(net_7237), .D(net_7237), .SE(net_3822), .SI(net_333), .CK(net_9386) );
DFF_X1 inst_6476 ( .QN(net_6089), .D(net_5583), .CK(net_12954) );
CLKBUF_X2 inst_9424 ( .A(net_9041), .Z(net_9386) );
CLKBUF_X2 inst_8549 ( .A(net_8510), .Z(net_8511) );
CLKBUF_X2 inst_11126 ( .A(net_11087), .Z(net_11088) );
AOI21_X2 inst_7654 ( .B2(net_3439), .ZN(net_3391), .A(net_3220), .B1(net_274) );
SDFF_X2 inst_1296 ( .D(net_6387), .SE(net_5801), .SI(net_332), .Q(net_332), .CK(net_13878) );
INV_X4 inst_4661 ( .ZN(net_5883), .A(net_3925) );
CLKBUF_X2 inst_14443 ( .A(net_14404), .Z(net_14405) );
OAI21_X2 inst_1852 ( .B1(net_5337), .ZN(net_5320), .A(net_4354), .B2(net_3853) );
DFF_X1 inst_6809 ( .D(net_3752), .CK(net_10823), .Q(x342) );
DFF_X2 inst_6273 ( .QN(net_5924), .D(net_391), .CK(net_8011) );
NAND2_X2 inst_3671 ( .A1(net_7335), .A2(net_1798), .ZN(net_1787) );
CLKBUF_X2 inst_7978 ( .A(net_7939), .Z(net_7940) );
NAND2_X2 inst_3282 ( .ZN(net_3682), .A1(net_3681), .A2(net_3226) );
CLKBUF_X2 inst_12667 ( .A(net_12628), .Z(net_12629) );
CLKBUF_X2 inst_13121 ( .A(net_10921), .Z(net_13083) );
NAND2_X2 inst_4074 ( .A1(net_6531), .A2(net_1645), .ZN(net_978) );
NAND2_X2 inst_3783 ( .A1(net_7029), .A2(net_1975), .ZN(net_1562) );
INV_X8 inst_4513 ( .ZN(net_3820), .A(net_3160) );
CLKBUF_X2 inst_13613 ( .A(net_13574), .Z(net_13575) );
OAI22_X2 inst_1557 ( .B2(net_3405), .A2(net_3360), .ZN(net_3348), .A1(net_3265), .B1(net_455) );
NOR2_X2 inst_2399 ( .A1(net_5778), .ZN(net_4166), .A2(net_297) );
CLKBUF_X2 inst_12207 ( .A(net_12168), .Z(net_12169) );
NAND2_X2 inst_3412 ( .A2(net_5964), .ZN(net_3386), .A1(net_2878) );
INV_X4 inst_4698 ( .A(net_5972), .ZN(net_3365) );
CLKBUF_X2 inst_10855 ( .A(net_10816), .Z(net_10817) );
CLKBUF_X2 inst_9620 ( .A(net_9581), .Z(net_9582) );
CLKBUF_X2 inst_8485 ( .A(net_8283), .Z(net_8447) );
DFF_X2 inst_6290 ( .QN(net_7687), .D(net_2264), .CK(net_9493) );
NAND2_X1 inst_4452 ( .A2(net_1256), .ZN(net_1126), .A1(net_1125) );
CLKBUF_X2 inst_11326 ( .A(net_11287), .Z(net_11288) );
CLKBUF_X2 inst_10633 ( .A(net_9515), .Z(net_10595) );
OAI22_X2 inst_1616 ( .A1(net_3128), .A2(net_3087), .B2(net_3084), .ZN(net_3054), .B1(net_3053) );
CLKBUF_X2 inst_14090 ( .A(net_13563), .Z(net_14052) );
CLKBUF_X2 inst_8813 ( .A(net_8774), .Z(net_8775) );
INV_X4 inst_5646 ( .A(net_6557), .ZN(net_597) );
CLKBUF_X2 inst_13167 ( .A(net_13128), .Z(net_13129) );
CLKBUF_X2 inst_11295 ( .A(net_10507), .Z(net_11257) );
CLKBUF_X2 inst_11403 ( .A(net_11364), .Z(net_11365) );
CLKBUF_X2 inst_9954 ( .A(net_9915), .Z(net_9916) );
OAI21_X2 inst_1825 ( .ZN(net_5360), .B1(net_5359), .A(net_4380), .B2(net_3856) );
NAND2_X2 inst_4151 ( .A2(net_1225), .ZN(net_1176), .A1(net_354) );
NAND2_X4 inst_2851 ( .ZN(net_5472), .A1(net_4913), .A2(net_4912) );
OAI22_X2 inst_1606 ( .A1(net_3277), .B2(net_3200), .A2(net_3193), .ZN(net_3127), .B1(net_1080) );
INV_X4 inst_5356 ( .A(net_7270), .ZN(net_2035) );
CLKBUF_X2 inst_13110 ( .A(net_13071), .Z(net_13072) );
INV_X4 inst_5619 ( .A(net_7786), .ZN(net_546) );
INV_X4 inst_5126 ( .A(net_850), .ZN(net_590) );
SDFF_X2 inst_410 ( .SI(net_7375), .Q(net_7375), .D(net_4876), .SE(net_3853), .CK(net_9397) );
SDFF_X2 inst_316 ( .SI(net_7459), .Q(net_7459), .D(net_5102), .SE(net_3993), .CK(net_9788) );
CLKBUF_X2 inst_8690 ( .A(net_8013), .Z(net_8652) );
CLKBUF_X2 inst_12860 ( .A(net_12821), .Z(net_12822) );
CLKBUF_X2 inst_11786 ( .A(net_11747), .Z(net_11748) );
CLKBUF_X2 inst_11621 ( .A(net_11582), .Z(net_11583) );
SDFF_X2 inst_1174 ( .SI(net_6945), .Q(net_6945), .D(net_3783), .SE(net_3741), .CK(net_8126) );
SDFF_X2 inst_1023 ( .SI(net_6518), .Q(net_6518), .SE(net_3886), .D(net_3801), .CK(net_11639) );
NAND2_X2 inst_3186 ( .ZN(net_4747), .A2(net_3941), .A1(net_2005) );
CLKBUF_X2 inst_8515 ( .A(net_8476), .Z(net_8477) );
SDFF_X2 inst_678 ( .Q(net_6742), .D(net_6742), .SE(net_3815), .SI(net_3786), .CK(net_11343) );
NAND2_X2 inst_3762 ( .A1(net_7032), .A2(net_1975), .ZN(net_1583) );
INV_X4 inst_5653 ( .A(net_6135), .ZN(net_3663) );
CLKBUF_X2 inst_10925 ( .A(net_9029), .Z(net_10887) );
NAND2_X2 inst_3259 ( .ZN(net_4150), .A1(net_3857), .A2(net_3466) );
SDFF_X2 inst_854 ( .SI(net_7039), .Q(net_7039), .D(net_3813), .SE(net_3777), .CK(net_10859) );
CLKBUF_X2 inst_12464 ( .A(net_10306), .Z(net_12426) );
CLKBUF_X2 inst_13293 ( .A(net_13254), .Z(net_13255) );
CLKBUF_X2 inst_13796 ( .A(net_13757), .Z(net_13758) );
NAND2_X1 inst_4359 ( .ZN(net_4368), .A2(net_3853), .A1(net_2054) );
AOI22_X2 inst_7310 ( .B1(net_6683), .A1(net_6651), .A2(net_5139), .B2(net_5138), .ZN(net_5133) );
CLKBUF_X2 inst_13177 ( .A(net_12640), .Z(net_13139) );
NAND2_X2 inst_3678 ( .A2(net_1798), .ZN(net_1777), .A1(net_1776) );
NAND2_X2 inst_3979 ( .ZN(net_1291), .A1(net_885), .A2(net_310) );
DFF_X2 inst_6297 ( .QN(net_5961), .D(net_1662), .CK(net_10724) );
CLKBUF_X2 inst_8033 ( .A(net_7913), .Z(net_7995) );
CLKBUF_X2 inst_12191 ( .A(net_11156), .Z(net_12153) );
OAI21_X2 inst_1946 ( .B1(net_5230), .ZN(net_5079), .A(net_4731), .B2(net_3986) );
CLKBUF_X2 inst_7865 ( .A(net_7826), .Z(net_7827) );
CLKBUF_X2 inst_10478 ( .A(net_10439), .Z(net_10440) );
CLKBUF_X2 inst_10472 ( .A(net_10433), .Z(net_10434) );
CLKBUF_X2 inst_12006 ( .A(net_11967), .Z(net_11968) );
CLKBUF_X2 inst_8686 ( .A(net_8647), .Z(net_8648) );
CLKBUF_X2 inst_9226 ( .A(net_9187), .Z(net_9188) );
INV_X4 inst_5322 ( .A(net_6057), .ZN(net_803) );
CLKBUF_X2 inst_8008 ( .A(net_7969), .Z(net_7970) );
CLKBUF_X2 inst_13401 ( .A(net_13362), .Z(net_13363) );
CLKBUF_X2 inst_9786 ( .A(net_9747), .Z(net_9748) );
CLKBUF_X2 inst_9073 ( .A(net_9034), .Z(net_9035) );
CLKBUF_X2 inst_10861 ( .A(net_10822), .Z(net_10823) );
NAND2_X2 inst_3457 ( .ZN(net_2986), .A2(net_2739), .A1(net_226) );
CLKBUF_X2 inst_12996 ( .A(net_12957), .Z(net_12958) );
CLKBUF_X2 inst_9464 ( .A(net_9425), .Z(net_9426) );
SDFF_X2 inst_688 ( .Q(net_6754), .D(net_6754), .SE(net_3815), .SI(net_3788), .CK(net_8368) );
NOR2_X2 inst_2549 ( .A2(net_7756), .A1(net_3208), .ZN(net_616) );
OAI21_X2 inst_1749 ( .ZN(net_5517), .A(net_4818), .B2(net_4153), .B1(net_1063) );
CLKBUF_X2 inst_9717 ( .A(net_9678), .Z(net_9679) );
NAND2_X2 inst_3641 ( .ZN(net_1922), .A2(net_1921), .A1(net_1683) );
DFF_X1 inst_6519 ( .QN(net_7450), .D(net_5433), .CK(net_9673) );
CLKBUF_X2 inst_14105 ( .A(net_14066), .Z(net_14067) );
INV_X4 inst_4894 ( .A(net_3796), .ZN(net_873) );
INV_X4 inst_5514 ( .A(net_6959), .ZN(net_566) );
CLKBUF_X2 inst_12518 ( .A(net_12479), .Z(net_12480) );
CLKBUF_X2 inst_9071 ( .A(net_9032), .Z(net_9033) );
NOR2_X2 inst_2387 ( .ZN(net_4293), .A1(net_4144), .A2(net_4143) );
CLKBUF_X2 inst_14416 ( .A(net_14377), .Z(net_14378) );
CLKBUF_X2 inst_13351 ( .A(net_13312), .Z(net_13313) );
CLKBUF_X2 inst_12980 ( .A(net_12853), .Z(net_12942) );
CLKBUF_X2 inst_12474 ( .A(net_12435), .Z(net_12436) );
CLKBUF_X2 inst_11872 ( .A(net_11362), .Z(net_11834) );
CLKBUF_X2 inst_9017 ( .A(net_8978), .Z(net_8979) );
NAND2_X1 inst_4391 ( .ZN(net_4336), .A2(net_3859), .A1(net_1995) );
CLKBUF_X2 inst_10137 ( .A(net_9211), .Z(net_10099) );
CLKBUF_X2 inst_10017 ( .A(net_8675), .Z(net_9979) );
CLKBUF_X2 inst_10163 ( .A(net_10124), .Z(net_10125) );
NAND2_X2 inst_3156 ( .ZN(net_4807), .A2(net_4153), .A1(net_2190) );
DFF_X1 inst_6423 ( .QN(net_6178), .D(net_5747), .CK(net_8743) );
NAND3_X2 inst_2747 ( .ZN(net_2354), .A3(net_1605), .A1(net_1322), .A2(net_963) );
CLKBUF_X2 inst_13744 ( .A(net_8797), .Z(net_13706) );
SDFF_X2 inst_840 ( .Q(net_7020), .D(net_7020), .SE(net_3899), .SI(net_3791), .CK(net_11892) );
SDFF_X2 inst_1220 ( .SI(net_7212), .Q(net_7212), .D(net_3776), .SE(net_3751), .CK(net_7833) );
CLKBUF_X2 inst_8554 ( .A(net_8515), .Z(net_8516) );
NOR4_X2 inst_2181 ( .A2(net_7760), .ZN(net_3309), .A4(net_3224), .A3(net_3208), .A1(net_2919) );
OAI22_X2 inst_1456 ( .B2(net_5909), .B1(net_4650), .A2(net_4614), .ZN(net_4612), .A1(net_4064) );
CLKBUF_X2 inst_11900 ( .A(net_10646), .Z(net_11862) );
CLKBUF_X2 inst_13523 ( .A(net_13484), .Z(net_13485) );
CLKBUF_X2 inst_12498 ( .A(net_12459), .Z(net_12460) );
CLKBUF_X2 inst_8909 ( .A(net_8870), .Z(net_8871) );
INV_X2 inst_6117 ( .A(net_5933), .ZN(net_5932) );
CLKBUF_X2 inst_10736 ( .A(net_10697), .Z(net_10698) );
CLKBUF_X2 inst_8965 ( .A(net_7840), .Z(net_8927) );
INV_X4 inst_5154 ( .A(net_563), .ZN(net_562) );
INV_X2 inst_5876 ( .A(net_7439), .ZN(net_1409) );
AOI222_X2 inst_7497 ( .C1(net_7517), .B1(net_7485), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2082), .A1(net_2081) );
CLKBUF_X2 inst_10593 ( .A(net_8458), .Z(net_10555) );
NAND2_X2 inst_4195 ( .A1(net_2809), .ZN(net_1213), .A2(net_305) );
NAND2_X1 inst_4294 ( .ZN(net_4572), .A2(net_3867), .A1(net_1869) );
CLKBUF_X2 inst_8473 ( .A(net_8434), .Z(net_8435) );
CLKBUF_X2 inst_9305 ( .A(net_9266), .Z(net_9267) );
CLKBUF_X2 inst_13605 ( .A(net_13566), .Z(net_13567) );
AOI222_X2 inst_7589 ( .ZN(net_5220), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_385), .C2(net_383), .A1(net_371) );
NAND2_X1 inst_4440 ( .A1(net_7607), .A2(net_2131), .ZN(net_1346) );
CLKBUF_X2 inst_14302 ( .A(net_14263), .Z(net_14264) );
CLKBUF_X2 inst_10799 ( .A(net_10119), .Z(net_10761) );
INV_X2 inst_5710 ( .ZN(net_4256), .A(net_4136) );
CLKBUF_X2 inst_11607 ( .A(net_11568), .Z(net_11569) );
INV_X2 inst_5959 ( .A(net_7323), .ZN(net_1761) );
DFFR_X2 inst_7072 ( .QN(net_6039), .D(net_3056), .CK(net_9993), .RN(x1822) );
CLKBUF_X2 inst_9536 ( .A(net_9031), .Z(net_9498) );
INV_X2 inst_5939 ( .A(net_7689), .ZN(net_836) );
CLKBUF_X2 inst_9149 ( .A(net_8399), .Z(net_9111) );
CLKBUF_X2 inst_11846 ( .A(net_11556), .Z(net_11808) );
NAND2_X2 inst_4199 ( .ZN(net_1830), .A1(net_645), .A2(net_306) );
CLKBUF_X2 inst_13588 ( .A(net_13549), .Z(net_13550) );
INV_X4 inst_5679 ( .A(net_7722), .ZN(net_2934) );
AOI22_X2 inst_7272 ( .B1(net_7086), .A1(net_7054), .A2(net_5280), .B2(net_5279), .ZN(net_5276) );
CLKBUF_X2 inst_14370 ( .A(net_14331), .Z(net_14332) );
CLKBUF_X2 inst_11141 ( .A(net_11102), .Z(net_11103) );
CLKBUF_X2 inst_9200 ( .A(net_9161), .Z(net_9162) );
CLKBUF_X2 inst_12718 ( .A(net_11974), .Z(net_12680) );
SDFF_X2 inst_617 ( .Q(net_6622), .D(net_6622), .SE(net_3830), .SI(net_3800), .CK(net_9165) );
CLKBUF_X2 inst_9167 ( .A(net_9128), .Z(net_9129) );
CLKBUF_X2 inst_8902 ( .A(net_8863), .Z(net_8864) );
INV_X2 inst_5734 ( .ZN(net_5888), .A(net_4148) );
INV_X2 inst_5749 ( .ZN(net_3915), .A(net_3740) );
DFF_X2 inst_6225 ( .QN(net_6557), .D(net_3723), .CK(net_8811) );
CLKBUF_X2 inst_12754 ( .A(net_12715), .Z(net_12716) );
CLKBUF_X2 inst_10823 ( .A(net_10784), .Z(net_10785) );
CLKBUF_X2 inst_14209 ( .A(net_14170), .Z(net_14171) );
NAND2_X1 inst_4420 ( .A1(net_7615), .A2(net_2131), .ZN(net_1517) );
CLKBUF_X2 inst_13795 ( .A(net_13756), .Z(net_13757) );
SDFF_X2 inst_1057 ( .Q(net_6744), .D(net_6744), .SI(net_3897), .SE(net_3815), .CK(net_11315) );
CLKBUF_X2 inst_8123 ( .A(net_8084), .Z(net_8085) );
CLKBUF_X2 inst_14097 ( .A(net_14058), .Z(net_14059) );
DFF_X1 inst_6614 ( .QN(net_7575), .D(net_5393), .CK(net_8033) );
CLKBUF_X2 inst_10359 ( .A(net_10320), .Z(net_10321) );
CLKBUF_X2 inst_8843 ( .A(net_8804), .Z(net_8805) );
INV_X4 inst_5191 ( .A(net_853), .ZN(net_512) );
INV_X2 inst_6029 ( .A(net_6031), .ZN(net_2830) );
INV_X4 inst_5602 ( .A(net_6079), .ZN(net_3548) );
CLKBUF_X2 inst_10743 ( .A(net_10704), .Z(net_10705) );
CLKBUF_X2 inst_11956 ( .A(net_11132), .Z(net_11918) );
CLKBUF_X2 inst_10610 ( .A(net_10571), .Z(net_10572) );
SDFF_X2 inst_748 ( .SI(net_7802), .Q(net_6838), .D(net_6838), .SE(net_3893), .CK(net_11808) );
CLKBUF_X2 inst_8609 ( .A(net_8570), .Z(net_8571) );
NAND2_X4 inst_2839 ( .ZN(net_5547), .A1(net_5020), .A2(net_5019) );
DFF_X1 inst_6730 ( .QN(net_7349), .D(net_5325), .CK(net_9438) );
CLKBUF_X2 inst_11373 ( .A(net_11334), .Z(net_11335) );
CLKBUF_X2 inst_9266 ( .A(net_9227), .Z(net_9228) );
INV_X4 inst_4582 ( .A(net_5074), .ZN(net_4330) );
INV_X4 inst_5482 ( .A(net_7250), .ZN(net_2162) );
DFF_X1 inst_6739 ( .QN(net_7284), .D(net_4867), .CK(net_10112) );
INV_X8 inst_4526 ( .ZN(net_3750), .A(net_3114) );
INV_X4 inst_5532 ( .A(net_7429), .ZN(net_2103) );
CLKBUF_X2 inst_8916 ( .A(net_8877), .Z(net_8878) );
CLKBUF_X2 inst_11070 ( .A(net_10600), .Z(net_11032) );
CLKBUF_X2 inst_9818 ( .A(net_9779), .Z(net_9780) );
CLKBUF_X2 inst_8798 ( .A(net_8759), .Z(net_8760) );
NAND2_X2 inst_2909 ( .ZN(net_5787), .A2(net_5772), .A1(net_397) );
OAI21_X2 inst_1986 ( .B1(net_4847), .ZN(net_4843), .A(net_4580), .B2(net_3867) );
INV_X4 inst_4587 ( .ZN(net_4315), .A(net_4229) );
OAI21_X2 inst_1949 ( .B1(net_5222), .ZN(net_5071), .A(net_4728), .B2(net_3986) );
CLKBUF_X2 inst_12636 ( .A(net_11358), .Z(net_12598) );
INV_X2 inst_5726 ( .ZN(net_4000), .A(net_3908) );
HA_X1 inst_6170 ( .S(net_1692), .CO(net_893), .A(net_892), .B(net_891) );
CLKBUF_X2 inst_12163 ( .A(net_12124), .Z(net_12125) );
CLKBUF_X2 inst_10644 ( .A(net_10173), .Z(net_10606) );
NAND2_X2 inst_3135 ( .ZN(net_4828), .A2(net_4153), .A1(net_2142) );
INV_X2 inst_5867 ( .A(net_1657), .ZN(net_531) );
SDFF_X2 inst_701 ( .SI(net_6771), .Q(net_6771), .SE(net_3872), .D(net_3811), .CK(net_11144) );
CLKBUF_X2 inst_8243 ( .A(net_8204), .Z(net_8205) );
NAND2_X2 inst_2911 ( .ZN(net_5783), .A2(net_5770), .A1(net_400) );
CLKBUF_X2 inst_13770 ( .A(net_13731), .Z(net_13732) );
NOR2_X2 inst_2380 ( .ZN(net_5127), .A2(net_4604), .A1(net_4402) );
CLKBUF_X2 inst_12337 ( .A(net_12298), .Z(net_12299) );
AOI222_X2 inst_7583 ( .A1(net_7240), .ZN(net_5341), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_334), .C2(net_332) );
INV_X4 inst_5261 ( .ZN(net_1068), .A(net_429) );
AOI21_X2 inst_7739 ( .B1(net_7140), .ZN(net_4078), .B2(net_2582), .A(net_2297) );
OAI21_X2 inst_1859 ( .ZN(net_5259), .B1(net_5227), .A(net_4544), .B2(net_3870) );
AOI21_X2 inst_7734 ( .B1(net_6743), .ZN(net_4118), .B2(net_2581), .A(net_2330) );
DFF_X1 inst_6933 ( .D(net_2399), .Q(net_239), .CK(net_10538) );
CLKBUF_X2 inst_8238 ( .A(net_8199), .Z(net_8200) );
NAND3_X2 inst_2815 ( .ZN(net_2283), .A3(net_1527), .A1(net_1503), .A2(net_995) );
SDFF_X2 inst_1007 ( .SI(net_6499), .Q(net_6499), .SE(net_3889), .D(net_3813), .CK(net_8637) );
CLKBUF_X2 inst_11011 ( .A(net_10972), .Z(net_10973) );
CLKBUF_X2 inst_8267 ( .A(net_8117), .Z(net_8229) );
INV_X2 inst_5754 ( .ZN(net_3905), .A(net_3735) );
CLKBUF_X2 inst_11674 ( .A(net_11635), .Z(net_11636) );
CLKBUF_X2 inst_8426 ( .A(net_8158), .Z(net_8388) );
NAND2_X2 inst_4208 ( .ZN(net_3222), .A2(net_270), .A1(net_269) );
NAND2_X2 inst_3605 ( .ZN(net_2395), .A2(net_1866), .A1(net_1450) );
CLKBUF_X2 inst_11932 ( .A(net_11893), .Z(net_11894) );
CLKBUF_X2 inst_9617 ( .A(net_8986), .Z(net_9579) );
SDFF_X2 inst_651 ( .Q(net_6707), .D(net_6707), .SE(net_3871), .SI(net_3811), .CK(net_11163) );
INV_X4 inst_5066 ( .A(net_1728), .ZN(net_734) );
CLKBUF_X2 inst_11998 ( .A(net_11959), .Z(net_11960) );
CLKBUF_X2 inst_11392 ( .A(net_11353), .Z(net_11354) );
NAND2_X4 inst_2883 ( .ZN(net_3925), .A1(net_3839), .A2(net_447) );
CLKBUF_X2 inst_11560 ( .A(net_11521), .Z(net_11522) );
CLKBUF_X2 inst_11313 ( .A(net_9340), .Z(net_11275) );
SDFF_X2 inst_1157 ( .SI(net_6792), .Q(net_6792), .D(net_3802), .SE(net_3722), .CK(net_11069) );
CLKBUF_X2 inst_8065 ( .A(net_8026), .Z(net_8027) );
CLKBUF_X2 inst_9993 ( .A(net_9954), .Z(net_9955) );
CLKBUF_X2 inst_11108 ( .A(net_9693), .Z(net_11070) );
CLKBUF_X2 inst_13395 ( .A(net_13356), .Z(net_13357) );
CLKBUF_X2 inst_8408 ( .A(net_8369), .Z(net_8370) );
NAND2_X2 inst_3528 ( .ZN(net_2539), .A2(net_2086), .A1(net_1362) );
CLKBUF_X2 inst_10083 ( .A(net_10044), .Z(net_10045) );
OAI21_X2 inst_2061 ( .B2(net_4436), .ZN(net_4434), .B1(net_4055), .A(net_3478) );
NAND2_X2 inst_3685 ( .A1(net_7341), .A2(net_1798), .ZN(net_1763) );
CLKBUF_X2 inst_10527 ( .A(net_10070), .Z(net_10489) );
CLKBUF_X2 inst_13486 ( .A(net_13447), .Z(net_13448) );
NAND2_X1 inst_4255 ( .ZN(net_4671), .A2(net_3993), .A1(net_1459) );
DFF_X1 inst_6891 ( .D(net_2520), .Q(net_166), .CK(net_10223) );
CLKBUF_X2 inst_11301 ( .A(net_11262), .Z(net_11263) );
OAI22_X2 inst_1472 ( .B1(net_4855), .A1(net_4228), .B2(net_4227), .ZN(net_4226), .A2(net_4225) );
NAND2_X1 inst_4261 ( .ZN(net_4659), .A2(net_3993), .A1(net_1463) );
AOI221_X2 inst_7616 ( .C2(net_3105), .B1(net_2970), .ZN(net_2963), .A(net_2782), .C1(net_863), .B2(net_251) );
CLKBUF_X2 inst_12511 ( .A(net_12472), .Z(net_12473) );
INV_X16 inst_6138 ( .ZN(net_1521), .A(net_789) );
NAND2_X2 inst_3784 ( .A1(net_6490), .A2(net_1642), .ZN(net_1561) );
SDFF_X2 inst_1183 ( .SI(net_6956), .Q(net_6956), .D(net_3800), .SE(net_3734), .CK(net_8330) );
CLKBUF_X2 inst_9577 ( .A(net_9538), .Z(net_9539) );
OAI22_X2 inst_1489 ( .B1(net_4666), .A1(net_4132), .B2(net_4126), .ZN(net_4123), .A2(net_4122) );
NOR2_X2 inst_2415 ( .A1(net_6041), .ZN(net_3408), .A2(net_3400) );
INV_X4 inst_5272 ( .ZN(net_3921), .A(net_800) );
CLKBUF_X2 inst_12353 ( .A(net_12314), .Z(net_12315) );
NAND2_X2 inst_3288 ( .ZN(net_3670), .A1(net_3669), .A2(net_3231) );
NOR2_X4 inst_2262 ( .ZN(net_5624), .A1(net_5469), .A2(net_4421) );
INV_X4 inst_4981 ( .ZN(net_862), .A(net_685) );
CLKBUF_X2 inst_8352 ( .A(net_8313), .Z(net_8314) );
INV_X4 inst_5506 ( .A(net_7263), .ZN(net_2063) );
CLKBUF_X2 inst_9131 ( .A(net_8060), .Z(net_9093) );
OR2_X4 inst_1394 ( .A2(net_7681), .A1(net_797), .ZN(net_779) );
SDFF_X2 inst_1160 ( .SI(net_6794), .Q(net_6794), .D(net_3799), .SE(net_3722), .CK(net_11067) );
CLKBUF_X2 inst_13724 ( .A(net_13685), .Z(net_13686) );
DFFR_X2 inst_7102 ( .D(net_1954), .QN(net_122), .CK(net_12325), .RN(x1822) );
CLKBUF_X2 inst_10767 ( .A(net_10370), .Z(net_10729) );
OAI21_X2 inst_1808 ( .ZN(net_5380), .B1(net_5361), .A(net_4350), .B2(net_3859) );
CLKBUF_X2 inst_8440 ( .A(net_8112), .Z(net_8402) );
OAI21_X2 inst_1876 ( .ZN(net_5226), .B1(net_5225), .A(net_4586), .B2(net_3867) );
SDFF_X2 inst_988 ( .Q(net_6475), .D(net_6475), .SE(net_3904), .SI(net_3807), .CK(net_8773) );
CLKBUF_X2 inst_10288 ( .A(net_10249), .Z(net_10250) );
CLKBUF_X2 inst_9333 ( .A(net_9294), .Z(net_9295) );
CLKBUF_X2 inst_12869 ( .A(net_11194), .Z(net_12831) );
SDFF_X2 inst_1315 ( .D(net_6385), .SE(net_5800), .SI(net_350), .Q(net_350), .CK(net_14137) );
INV_X4 inst_4954 ( .ZN(net_729), .A(net_728) );
INV_X4 inst_5035 ( .A(net_7809), .ZN(net_3809) );
NOR2_X2 inst_2392 ( .ZN(net_3997), .A2(net_3996), .A1(net_1931) );
INV_X4 inst_4759 ( .ZN(net_3252), .A(net_2872) );
NAND2_X1 inst_4308 ( .ZN(net_4558), .A2(net_3866), .A1(net_2134) );
INV_X4 inst_4678 ( .ZN(net_3387), .A(net_3386) );
CLKBUF_X2 inst_11026 ( .A(net_10987), .Z(net_10988) );
CLKBUF_X2 inst_9531 ( .A(net_9492), .Z(net_9493) );
CLKBUF_X2 inst_13513 ( .A(net_13474), .Z(net_13475) );
NAND2_X2 inst_3667 ( .A1(net_7339), .A2(net_1798), .ZN(net_1792) );
AOI222_X2 inst_7569 ( .A1(net_7547), .ZN(net_5235), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_379), .C2(net_377) );
CLKBUF_X2 inst_7972 ( .A(net_7933), .Z(net_7934) );
NAND2_X1 inst_4434 ( .A2(net_2131), .ZN(net_1399), .A1(net_1398) );
DFF_X1 inst_6380 ( .QN(net_6282), .D(net_5804), .CK(net_14252) );
CLKBUF_X2 inst_10049 ( .A(net_10010), .Z(net_10011) );
INV_X4 inst_4967 ( .A(net_3892), .ZN(net_3265) );
CLKBUF_X2 inst_9808 ( .A(net_8502), .Z(net_9770) );
DFF_X1 inst_6785 ( .Q(net_7778), .D(net_4298), .CK(net_12788) );
CLKBUF_X2 inst_10792 ( .A(net_10753), .Z(net_10754) );
INV_X4 inst_5527 ( .A(net_7414), .ZN(net_2085) );
DFFR_X2 inst_7007 ( .QN(net_7695), .D(net_3347), .CK(net_10353), .RN(x1822) );
CLKBUF_X2 inst_13993 ( .A(net_13954), .Z(net_13955) );
CLKBUF_X2 inst_10866 ( .A(net_10827), .Z(net_10828) );
SDFF_X2 inst_656 ( .Q(net_6695), .D(net_6695), .SE(net_3871), .SI(net_3778), .CK(net_8293) );
CLKBUF_X2 inst_9690 ( .A(net_9117), .Z(net_9652) );
DFF_X1 inst_6718 ( .QN(net_7319), .D(net_5344), .CK(net_10232) );
DFF_X1 inst_6900 ( .D(net_2507), .Q(net_181), .CK(net_9943) );
CLKBUF_X2 inst_12562 ( .A(net_12523), .Z(net_12524) );
INV_X2 inst_5919 ( .A(net_7516), .ZN(net_2140) );
XNOR2_X2 inst_45 ( .B(net_6555), .ZN(net_2442), .A(net_1237) );
CLKBUF_X2 inst_13471 ( .A(net_7903), .Z(net_13433) );
CLKBUF_X2 inst_9551 ( .A(net_9512), .Z(net_9513) );
CLKBUF_X2 inst_12500 ( .A(net_12461), .Z(net_12462) );
NAND2_X2 inst_3093 ( .A1(net_6454), .A2(net_4925), .ZN(net_4910) );
SDFF_X2 inst_458 ( .Q(net_6463), .D(net_6463), .SE(net_3904), .SI(net_3883), .CK(net_8809) );
CLKBUF_X2 inst_9934 ( .A(net_8310), .Z(net_9896) );
OAI22_X2 inst_1562 ( .B2(net_3405), .A2(net_3360), .ZN(net_3343), .A1(net_3275), .B1(net_2959) );
NAND2_X2 inst_4148 ( .A2(net_1222), .ZN(net_1086), .A1(net_344) );
CLKBUF_X2 inst_11814 ( .A(net_11775), .Z(net_11776) );
CLKBUF_X2 inst_8644 ( .A(net_8605), .Z(net_8606) );
INV_X4 inst_4618 ( .ZN(net_4204), .A(net_4069) );
INV_X4 inst_5539 ( .ZN(net_1226), .A(net_292) );
DFF_X1 inst_6827 ( .Q(net_6360), .D(net_2701), .CK(net_13763) );
OAI21_X2 inst_1922 ( .ZN(net_5123), .A(net_4752), .B2(net_3941), .B1(net_1064) );
NAND2_X2 inst_3361 ( .ZN(net_3524), .A1(net_3523), .A2(net_3228) );
NAND2_X2 inst_3170 ( .ZN(net_4763), .A2(net_3941), .A1(net_2063) );
SDFF_X2 inst_741 ( .Q(net_6831), .D(net_6831), .SE(net_3893), .SI(net_3802), .CK(net_8945) );
NAND2_X2 inst_3232 ( .ZN(net_4523), .A2(net_4290), .A1(net_1736) );
CLKBUF_X2 inst_8335 ( .A(net_8296), .Z(net_8297) );
CLKBUF_X2 inst_13062 ( .A(net_13023), .Z(net_13024) );
CLKBUF_X2 inst_9377 ( .A(net_8198), .Z(net_9339) );
CLKBUF_X2 inst_10524 ( .A(net_10485), .Z(net_10486) );
CLKBUF_X2 inst_10444 ( .A(net_10405), .Z(net_10406) );
INV_X2 inst_5973 ( .A(net_7635), .ZN(net_1885) );
CLKBUF_X2 inst_8700 ( .A(net_8245), .Z(net_8662) );
DFF_X1 inst_6942 ( .D(net_1942), .Q(net_388), .CK(net_14363) );
CLKBUF_X2 inst_9338 ( .A(net_9299), .Z(net_9300) );
SDFFR_X2 inst_1350 ( .D(net_3900), .SE(net_3256), .SI(net_151), .Q(net_151), .CK(net_8547), .RN(x1822) );
CLKBUF_X2 inst_12156 ( .A(net_12117), .Z(net_12118) );
CLKBUF_X2 inst_10178 ( .A(net_10139), .Z(net_10140) );
CLKBUF_X2 inst_12964 ( .A(net_12925), .Z(net_12926) );
NAND2_X2 inst_3012 ( .A1(net_6888), .A2(net_5006), .ZN(net_4997) );
CLKBUF_X2 inst_11369 ( .A(net_11330), .Z(net_11331) );
NAND3_X2 inst_2635 ( .ZN(net_5694), .A1(net_5671), .A2(net_5301), .A3(net_4245) );
CLKBUF_X2 inst_8124 ( .A(net_8085), .Z(net_8086) );
NAND3_X2 inst_2828 ( .A2(net_3854), .ZN(net_1214), .A3(net_1213), .A1(net_655) );
CLKBUF_X2 inst_14014 ( .A(net_13975), .Z(net_13976) );
CLKBUF_X2 inst_8673 ( .A(net_8634), .Z(net_8635) );
CLKBUF_X2 inst_13560 ( .A(net_13521), .Z(net_13522) );
AOI21_X2 inst_7769 ( .B1(net_7150), .ZN(net_4064), .B2(net_2582), .A(net_2318) );
NAND2_X2 inst_3877 ( .A1(net_6848), .A2(net_1521), .ZN(net_1443) );
NAND2_X2 inst_3363 ( .ZN(net_3520), .A1(net_3519), .A2(net_3223) );
INV_X4 inst_4745 ( .A(net_2752), .ZN(net_2746) );
CLKBUF_X2 inst_9859 ( .A(net_9820), .Z(net_9821) );
NAND3_X2 inst_2666 ( .ZN(net_3965), .A2(net_3877), .A3(net_3739), .A1(net_2240) );
AOI22_X2 inst_7320 ( .ZN(net_4551), .B2(net_3972), .A2(net_3380), .A1(net_1160), .B1(net_930) );
SDFF_X2 inst_1131 ( .SI(net_6683), .Q(net_6683), .D(net_3788), .SE(net_3471), .CK(net_9071) );
SDFFR_X2 inst_1357 ( .Q(net_6013), .D(net_6013), .SI(net_3782), .SE(net_3200), .CK(net_13182), .RN(x1822) );
SDFF_X2 inst_691 ( .Q(net_6756), .D(net_6756), .SE(net_3815), .SI(net_3801), .CK(net_8366) );
CLKBUF_X2 inst_11769 ( .A(net_11730), .Z(net_11731) );
CLKBUF_X2 inst_10938 ( .A(net_10899), .Z(net_10900) );
CLKBUF_X2 inst_9547 ( .A(net_9508), .Z(net_9509) );
DFF_X1 inst_6402 ( .QN(net_6141), .D(net_5768), .CK(net_11762) );
CLKBUF_X2 inst_12845 ( .A(net_12806), .Z(net_12807) );
SDFF_X2 inst_770 ( .Q(net_6865), .D(net_6865), .SE(net_3901), .SI(net_3799), .CK(net_11807) );
SDFF_X2 inst_565 ( .Q(net_6577), .D(net_6577), .SI(net_3897), .SE(net_3823), .CK(net_9188) );
OAI21_X2 inst_1971 ( .B1(net_4872), .ZN(net_4865), .A(net_4387), .B2(net_3856) );
SDFF_X2 inst_622 ( .SI(net_7802), .Q(net_6600), .D(net_6600), .SE(net_3830), .CK(net_9162) );
INV_X4 inst_5302 ( .A(net_7092), .ZN(net_502) );
AOI22_X2 inst_7418 ( .B1(net_5939), .A1(net_2872), .ZN(net_2775), .B2(net_224), .A2(net_187) );
CLKBUF_X2 inst_14345 ( .A(net_14306), .Z(net_14307) );
CLKBUF_X2 inst_12342 ( .A(net_12151), .Z(net_12304) );
INV_X8 inst_4476 ( .ZN(net_5006), .A(net_4268) );
CLKBUF_X2 inst_11307 ( .A(net_11268), .Z(net_11269) );
DFF_X1 inst_6861 ( .D(net_2546), .Q(net_198), .CK(net_12076) );
CLKBUF_X2 inst_11679 ( .A(net_10176), .Z(net_11641) );
SDFF_X2 inst_409 ( .SI(net_7373), .Q(net_7373), .D(net_4778), .SE(net_3853), .CK(net_9894) );
CLKBUF_X2 inst_12323 ( .A(net_12284), .Z(net_12285) );
NOR2_X4 inst_2288 ( .A2(net_7791), .ZN(net_2871), .A1(net_801) );
CLKBUF_X2 inst_13644 ( .A(net_8698), .Z(net_13606) );
CLKBUF_X2 inst_11505 ( .A(net_11466), .Z(net_11467) );
DFF_X1 inst_6672 ( .QN(net_7267), .D(net_5158), .CK(net_9965) );
INV_X2 inst_5813 ( .ZN(net_1102), .A(net_1101) );
INV_X4 inst_4841 ( .A(net_3857), .ZN(net_3050) );
CLKBUF_X2 inst_9368 ( .A(net_8245), .Z(net_9330) );
OAI21_X2 inst_1834 ( .ZN(net_5342), .B1(net_5341), .A(net_4356), .B2(net_3856) );
CLKBUF_X2 inst_12933 ( .A(net_12757), .Z(net_12895) );
CLKBUF_X2 inst_8013 ( .A(net_7974), .Z(net_7975) );
NAND2_X2 inst_3506 ( .ZN(net_2561), .A2(net_1990), .A1(net_1343) );
NAND2_X2 inst_3574 ( .ZN(net_2493), .A2(net_2028), .A1(net_1763) );
NOR2_X4 inst_2228 ( .ZN(net_5670), .A1(net_5533), .A2(net_4501) );
CLKBUF_X2 inst_9220 ( .A(net_9181), .Z(net_9182) );
CLKBUF_X2 inst_11947 ( .A(net_11908), .Z(net_11909) );
DFFR_X2 inst_7092 ( .QN(net_6418), .D(net_2719), .CK(net_13022), .RN(x1822) );
AOI22_X2 inst_7396 ( .A2(net_3105), .B1(net_2970), .ZN(net_2845), .A1(net_552), .B2(net_256) );
CLKBUF_X2 inst_11389 ( .A(net_11350), .Z(net_11351) );
SDFF_X2 inst_768 ( .Q(net_6891), .D(net_6891), .SE(net_3901), .SI(net_3801), .CK(net_11726) );
AND4_X2 inst_7795 ( .ZN(net_804), .A1(net_803), .A2(net_802), .A3(net_801), .A4(net_800) );
SDFF_X2 inst_663 ( .Q(net_6722), .D(net_6722), .SE(net_3871), .SI(net_3788), .CK(net_8377) );
OAI21_X2 inst_2121 ( .B1(net_3291), .ZN(net_3090), .B2(net_3087), .A(net_2913) );
INV_X4 inst_4850 ( .ZN(net_1058), .A(net_1057) );
NAND2_X2 inst_3227 ( .ZN(net_4528), .A2(net_4295), .A1(net_1732) );
CLKBUF_X2 inst_12067 ( .A(net_12028), .Z(net_12029) );
CLKBUF_X2 inst_8949 ( .A(net_8910), .Z(net_8911) );
DFF_X1 inst_6639 ( .QN(net_7627), .D(net_5236), .CK(net_10564) );
CLKBUF_X2 inst_11001 ( .A(net_10962), .Z(net_10963) );
CLKBUF_X2 inst_13225 ( .A(net_8690), .Z(net_13187) );
DFF_X1 inst_6774 ( .QN(net_6144), .D(net_4601), .CK(net_9132) );
NAND2_X2 inst_3494 ( .A2(net_2644), .ZN(net_2625), .A1(net_2590) );
NAND2_X1 inst_4224 ( .ZN(net_4703), .A2(net_3989), .A1(net_2173) );
OAI21_X2 inst_1867 ( .ZN(net_5247), .B1(net_5200), .A(net_4532), .B2(net_3870) );
CLKBUF_X2 inst_13627 ( .A(net_13588), .Z(net_13589) );
DFF_X2 inst_6314 ( .QN(net_7811), .CK(net_8435), .D(x1451) );
AOI222_X2 inst_7580 ( .A1(net_7389), .ZN(net_5551), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_352), .C2(net_350) );
DFFR_X2 inst_7046 ( .QN(net_6010), .D(net_3134), .CK(net_10443), .RN(x1822) );
AOI22_X2 inst_7279 ( .B1(net_7081), .A1(net_7049), .A2(net_5280), .B2(net_5279), .ZN(net_5265) );
NOR2_X4 inst_2290 ( .A2(net_7791), .ZN(net_2866), .A1(net_1679) );
CLKBUF_X2 inst_13782 ( .A(net_9746), .Z(net_13744) );
CLKBUF_X2 inst_7909 ( .A(net_7853), .Z(net_7871) );
CLKBUF_X2 inst_11913 ( .A(net_11874), .Z(net_11875) );
INV_X4 inst_5670 ( .ZN(net_1227), .A(net_291) );
DFF_X1 inst_6791 ( .D(net_3949), .CK(net_12840), .Q(x538) );
INV_X4 inst_5070 ( .ZN(net_1142), .A(net_631) );
CLKBUF_X2 inst_13695 ( .A(net_9871), .Z(net_13657) );
CLKBUF_X2 inst_12575 ( .A(net_12536), .Z(net_12537) );
INV_X2 inst_5797 ( .ZN(net_2227), .A(net_2226) );
CLKBUF_X2 inst_14143 ( .A(net_14104), .Z(net_14105) );
INV_X4 inst_4912 ( .ZN(net_1043), .A(net_862) );
NAND2_X2 inst_3342 ( .ZN(net_3563), .A1(net_3562), .A2(net_3225) );
INV_X4 inst_4825 ( .ZN(net_4777), .A(net_1086) );
CLKBUF_X2 inst_9832 ( .A(net_9793), .Z(net_9794) );
NAND3_X2 inst_2621 ( .ZN(net_5718), .A1(net_5613), .A2(net_5130), .A3(net_4177) );
CLKBUF_X2 inst_8175 ( .A(net_8097), .Z(net_8137) );
CLKBUF_X2 inst_9159 ( .A(net_9120), .Z(net_9121) );
CLKBUF_X2 inst_10815 ( .A(net_10776), .Z(net_10777) );
CLKBUF_X2 inst_14454 ( .A(net_14415), .Z(net_14416) );
NAND2_X2 inst_3895 ( .A1(net_6434), .A2(net_1677), .ZN(net_1419) );
CLKBUF_X2 inst_11928 ( .A(net_11889), .Z(net_11890) );
CLKBUF_X2 inst_9358 ( .A(net_9319), .Z(net_9320) );
SDFF_X2 inst_303 ( .SI(net_7521), .Q(net_7521), .D(net_5103), .SE(net_3988), .CK(net_12458) );
CLKBUF_X2 inst_13518 ( .A(net_13479), .Z(net_13480) );
CLKBUF_X2 inst_14324 ( .A(net_14285), .Z(net_14286) );
AOI21_X2 inst_7699 ( .B1(net_6728), .ZN(net_5894), .B2(net_2581), .A(net_2364) );
NAND2_X2 inst_3263 ( .ZN(net_4139), .A1(net_3854), .A2(net_3713) );
OAI221_X2 inst_1647 ( .ZN(net_5088), .C2(net_5087), .B2(net_5084), .A(net_4527), .B1(net_2435), .C1(net_1078) );
CLKBUF_X2 inst_12114 ( .A(net_9628), .Z(net_12076) );
SDFF_X2 inst_1275 ( .D(net_6388), .SE(net_5801), .SI(net_333), .Q(net_333), .CK(net_13883) );
XNOR2_X2 inst_26 ( .ZN(net_2570), .B(net_2569), .A(net_2447) );
CLKBUF_X2 inst_13052 ( .A(net_11586), .Z(net_13014) );
CLKBUF_X2 inst_10480 ( .A(net_10441), .Z(net_10442) );
CLKBUF_X2 inst_8104 ( .A(net_7912), .Z(net_8066) );
CLKBUF_X2 inst_10198 ( .A(net_10159), .Z(net_10160) );
NAND2_X4 inst_2882 ( .ZN(net_3926), .A1(net_3845), .A2(net_567) );
OR2_X4 inst_1376 ( .ZN(net_3445), .A2(net_3247), .A1(net_2610) );
CLKBUF_X2 inst_12731 ( .A(net_12692), .Z(net_12693) );
CLKBUF_X2 inst_14038 ( .A(net_13999), .Z(net_14000) );
CLKBUF_X2 inst_12605 ( .A(net_8366), .Z(net_12567) );
CLKBUF_X2 inst_10507 ( .A(net_8649), .Z(net_10469) );
CLKBUF_X2 inst_10001 ( .A(net_9962), .Z(net_9963) );
DFF_X1 inst_6530 ( .QN(net_7477), .D(net_5421), .CK(net_9275) );
AOI222_X2 inst_7490 ( .C1(net_7525), .B1(net_7493), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2104), .A1(net_2103) );
CLKBUF_X2 inst_12895 ( .A(net_11460), .Z(net_12857) );
CLKBUF_X2 inst_11483 ( .A(net_8843), .Z(net_11445) );
CLKBUF_X2 inst_8182 ( .A(net_8143), .Z(net_8144) );
INV_X4 inst_4864 ( .A(net_2222), .ZN(net_1820) );
CLKBUF_X2 inst_10654 ( .A(net_10615), .Z(net_10616) );
DFF_X2 inst_6188 ( .QN(net_6824), .D(net_5088), .CK(net_10798) );
NAND2_X2 inst_3765 ( .A1(net_6767), .A2(net_1635), .ZN(net_1580) );
CLKBUF_X2 inst_10742 ( .A(net_10703), .Z(net_10704) );
OAI221_X2 inst_1659 ( .ZN(net_4794), .A(net_4550), .C2(net_3969), .B2(net_3958), .C1(net_3758), .B1(net_1485) );
NAND2_X1 inst_4218 ( .ZN(net_4742), .A2(net_3988), .A1(net_2123) );
AOI21_X2 inst_7718 ( .B1(net_6865), .ZN(net_5906), .B2(net_2579), .A(net_2342) );
CLKBUF_X2 inst_10062 ( .A(net_10023), .Z(net_10024) );
DFF_X1 inst_6456 ( .QN(net_6109), .D(net_5603), .CK(net_11180) );
SDFF_X2 inst_398 ( .SI(net_7340), .Q(net_7340), .D(net_4779), .SE(net_3856), .CK(net_9913) );
INV_X4 inst_5702 ( .ZN(net_5940), .A(net_5939) );
CLKBUF_X2 inst_8184 ( .A(net_8145), .Z(net_8146) );
SDFF_X2 inst_436 ( .Q(net_7389), .D(net_7389), .SE(net_3994), .SI(net_354), .CK(net_9639) );
DFFR_X2 inst_7064 ( .QN(net_6043), .D(net_3085), .CK(net_10012), .RN(x1822) );
CLKBUF_X2 inst_13265 ( .A(net_11868), .Z(net_13227) );
CLKBUF_X2 inst_11766 ( .A(net_8623), .Z(net_11728) );
CLKBUF_X2 inst_9852 ( .A(net_8116), .Z(net_9814) );
DFF_X1 inst_6529 ( .QN(net_7476), .D(net_5422), .CK(net_10080) );
CLKBUF_X2 inst_11636 ( .A(net_11597), .Z(net_11598) );
CLKBUF_X2 inst_13702 ( .A(net_9784), .Z(net_13664) );
NAND2_X2 inst_3705 ( .A1(net_2299), .ZN(net_1671), .A2(net_1670) );
AOI21_X4 inst_7623 ( .ZN(net_4162), .A(net_3745), .B1(net_937), .B2(net_113) );
CLKBUF_X2 inst_11469 ( .A(net_11430), .Z(net_11431) );
INV_X4 inst_5053 ( .A(net_3232), .ZN(net_644) );
DFF_X1 inst_6746 ( .QN(net_7585), .D(net_4850), .CK(net_10297) );
NOR2_X4 inst_2231 ( .ZN(net_5667), .A1(net_5527), .A2(net_4495) );
SDFF_X2 inst_144 ( .Q(net_6234), .SI(net_6233), .SE(net_392), .D(net_140), .CK(net_13616) );
OAI22_X2 inst_1438 ( .B1(net_5851), .ZN(net_5685), .A2(net_5496), .B2(net_5495), .A1(net_5255) );
CLKBUF_X2 inst_9750 ( .A(net_9711), .Z(net_9712) );
CLKBUF_X2 inst_10454 ( .A(net_10415), .Z(net_10416) );
CLKBUF_X2 inst_10565 ( .A(net_7882), .Z(net_10527) );
DFF_X1 inst_6373 ( .QN(net_6289), .D(net_5811), .CK(net_14272) );
CLKBUF_X2 inst_13660 ( .A(net_13621), .Z(net_13622) );
CLKBUF_X2 inst_12681 ( .A(net_11810), .Z(net_12643) );
SDFF_X2 inst_880 ( .Q(net_7110), .D(net_7110), .SE(net_3888), .SI(net_3813), .CK(net_13373) );
DFF_X1 inst_6912 ( .D(net_2423), .Q(net_387), .CK(net_14376) );
INV_X4 inst_4857 ( .ZN(net_1090), .A(net_1043) );
CLKBUF_X2 inst_9763 ( .A(net_9607), .Z(net_9725) );
CLKBUF_X2 inst_12241 ( .A(net_11570), .Z(net_12203) );
CLKBUF_X2 inst_11437 ( .A(net_10396), .Z(net_11399) );
NAND3_X2 inst_2681 ( .ZN(net_3205), .A2(net_2940), .A3(net_2846), .A1(net_2779) );
NAND2_X2 inst_3445 ( .ZN(net_3155), .A2(net_3154), .A1(net_3152) );
CLKBUF_X2 inst_10026 ( .A(net_9451), .Z(net_9988) );
INV_X4 inst_5555 ( .A(net_6963), .ZN(net_2573) );
NAND2_X1 inst_4447 ( .A2(net_1256), .ZN(net_1136), .A1(net_1135) );
CLKBUF_X2 inst_9118 ( .A(net_9079), .Z(net_9080) );
CLKBUF_X2 inst_12370 ( .A(net_10957), .Z(net_12332) );
DFF_X2 inst_6194 ( .QN(net_7230), .D(net_5051), .CK(net_9370) );
CLKBUF_X2 inst_8493 ( .A(net_8454), .Z(net_8455) );
CLKBUF_X2 inst_9044 ( .A(net_9005), .Z(net_9006) );
NAND2_X2 inst_3972 ( .ZN(net_1298), .A1(net_885), .A2(net_317) );
DFF_X1 inst_6670 ( .QN(net_7265), .D(net_5160), .CK(net_12259) );
CLKBUF_X2 inst_11633 ( .A(net_11035), .Z(net_11595) );
OR2_X4 inst_1388 ( .A2(net_7762), .ZN(net_2851), .A1(net_267) );
NAND3_X2 inst_2699 ( .ZN(net_2693), .A3(net_2568), .A2(net_2428), .A1(net_2266) );
CLKBUF_X2 inst_12470 ( .A(net_12431), .Z(net_12432) );
DFF_X2 inst_6329 ( .QN(net_7818), .CK(net_11032), .D(x1390) );
NAND2_X2 inst_3517 ( .ZN(net_2550), .A2(net_2183), .A1(net_1422) );
CLKBUF_X2 inst_9291 ( .A(net_9252), .Z(net_9253) );
CLKBUF_X2 inst_8506 ( .A(net_8105), .Z(net_8468) );
NAND2_X2 inst_3396 ( .ZN(net_3463), .A2(net_3324), .A1(net_3237) );
OR2_X4 inst_1372 ( .ZN(net_3969), .A2(net_3735), .A1(net_3224) );
SDFFR_X2 inst_1360 ( .SI(net_6046), .Q(net_6046), .D(net_3810), .SE(net_3087), .CK(net_12815), .RN(x1822) );
AOI22_X2 inst_7332 ( .A2(net_3423), .B2(net_3422), .ZN(net_3414), .B1(net_2567), .A1(net_1248) );
CLKBUF_X2 inst_12109 ( .A(net_8024), .Z(net_12071) );
CLKBUF_X2 inst_10631 ( .A(net_10592), .Z(net_10593) );
CLKBUF_X2 inst_9759 ( .A(net_9720), .Z(net_9721) );
SDFF_X2 inst_466 ( .Q(net_6882), .D(net_6882), .SE(net_3901), .SI(net_3900), .CK(net_10938) );
INV_X2 inst_6081 ( .A(net_6034), .ZN(net_2828) );
NAND2_X2 inst_3981 ( .ZN(net_1289), .A1(net_885), .A2(net_320) );
NAND3_X2 inst_2761 ( .ZN(net_2340), .A3(net_1620), .A1(net_1482), .A2(net_1017) );
SDFF_X2 inst_989 ( .Q(net_6457), .D(net_6457), .SE(net_3904), .SI(net_3806), .CK(net_11548) );
INV_X4 inst_5205 ( .ZN(net_494), .A(net_493) );
NOR2_X4 inst_2283 ( .ZN(net_5893), .A2(net_5875), .A1(net_3026) );
CLKBUF_X2 inst_10073 ( .A(net_10034), .Z(net_10035) );
NAND2_X2 inst_3038 ( .A1(net_6991), .A2(net_4977), .ZN(net_4969) );
CLKBUF_X2 inst_14154 ( .A(net_14115), .Z(net_14116) );
SDFF_X2 inst_858 ( .SI(net_7043), .Q(net_7043), .SE(net_3818), .D(net_3787), .CK(net_11887) );
AOI222_X2 inst_7605 ( .A1(net_7400), .ZN(net_5436), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_363), .C2(net_361) );
AOI222_X2 inst_7542 ( .C1(net_7677), .A1(net_7645), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1878), .B1(net_1877) );
NAND2_X2 inst_3864 ( .A1(net_6830), .A2(net_1521), .ZN(net_1468) );
CLKBUF_X2 inst_9111 ( .A(net_9072), .Z(net_9073) );
CLKBUF_X2 inst_13779 ( .A(net_13740), .Z(net_13741) );
CLKBUF_X2 inst_12060 ( .A(net_12021), .Z(net_12022) );
CLKBUF_X2 inst_12735 ( .A(net_12696), .Z(net_12697) );
NAND2_X2 inst_2936 ( .ZN(net_5510), .A1(net_4982), .A2(net_4981) );
NOR2_X2 inst_2468 ( .ZN(net_2925), .A1(net_2703), .A2(net_264) );
XNOR2_X2 inst_54 ( .ZN(net_2247), .A(net_1918), .B(net_893) );
CLKBUF_X2 inst_12610 ( .A(net_12571), .Z(net_12572) );
CLKBUF_X2 inst_10556 ( .A(net_10517), .Z(net_10518) );
OAI22_X2 inst_1482 ( .A1(net_7782), .ZN(net_4163), .A2(net_4162), .B2(net_4161), .B1(net_1041) );
OR2_X2 inst_1420 ( .ZN(net_3773), .A2(net_784), .A1(net_428) );
CLKBUF_X2 inst_9757 ( .A(net_9718), .Z(net_9719) );
AOI22_X2 inst_7406 ( .B1(net_5939), .A2(net_2838), .ZN(net_2831), .A1(net_2830), .B2(net_196) );
CLKBUF_X2 inst_12177 ( .A(net_12138), .Z(net_12139) );
CLKBUF_X2 inst_12988 ( .A(net_9603), .Z(net_12950) );
INV_X4 inst_5214 ( .A(net_573), .ZN(net_481) );
AOI22_X2 inst_7283 ( .B1(net_7220), .A1(net_7188), .A2(net_5244), .B2(net_5243), .ZN(net_5234) );
INV_X4 inst_5337 ( .A(net_6105), .ZN(net_3685) );
NAND2_X2 inst_4062 ( .A1(net_6929), .A2(net_1654), .ZN(net_990) );
CLKBUF_X2 inst_13331 ( .A(net_13292), .Z(net_13293) );
INV_X2 inst_5730 ( .ZN(net_3964), .A(net_3963) );
NAND2_X2 inst_4108 ( .A1(net_6672), .A2(net_1655), .ZN(net_944) );
INV_X4 inst_4626 ( .ZN(net_4196), .A(net_4052) );
CLKBUF_X2 inst_8780 ( .A(net_8741), .Z(net_8742) );
CLKBUF_X2 inst_13838 ( .A(net_13799), .Z(net_13800) );
INV_X4 inst_4794 ( .A(net_2855), .ZN(net_1266) );
CLKBUF_X2 inst_13688 ( .A(net_13649), .Z(net_13650) );
CLKBUF_X2 inst_10804 ( .A(net_8064), .Z(net_10766) );
CLKBUF_X2 inst_9491 ( .A(net_7884), .Z(net_9453) );
CLKBUF_X2 inst_11595 ( .A(net_11482), .Z(net_11557) );
NAND2_X2 inst_3829 ( .A1(net_6573), .A2(net_1705), .ZN(net_1512) );
CLKBUF_X2 inst_7883 ( .A(net_7844), .Z(net_7845) );
CLKBUF_X2 inst_13414 ( .A(net_13375), .Z(net_13376) );
CLKBUF_X2 inst_9012 ( .A(net_8821), .Z(net_8974) );
SDFF_X2 inst_497 ( .Q(net_6982), .D(net_6982), .SI(net_3897), .SE(net_3891), .CK(net_11968) );
CLKBUF_X2 inst_10971 ( .A(net_10148), .Z(net_10933) );
CLKBUF_X2 inst_10325 ( .A(net_10286), .Z(net_10287) );
CLKBUF_X2 inst_13918 ( .A(net_13879), .Z(net_13880) );
CLKBUF_X2 inst_13826 ( .A(net_13787), .Z(net_13788) );
AOI222_X2 inst_7517 ( .B1(net_7376), .C1(net_7312), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2018), .A1(net_2017) );
NOR3_X2 inst_2195 ( .ZN(net_3881), .A1(net_3383), .A3(net_1739), .A2(net_700) );
CLKBUF_X2 inst_8161 ( .A(net_8122), .Z(net_8123) );
CLKBUF_X2 inst_8787 ( .A(net_8589), .Z(net_8749) );
OAI211_X2 inst_2168 ( .B(net_2724), .ZN(net_2720), .A(net_2420), .C1(net_2419), .C2(net_2418) );
SDFFR_X2 inst_1335 ( .SI(net_6417), .Q(net_6417), .SE(net_3753), .D(net_1929), .CK(net_10203), .RN(x1822) );
CLKBUF_X2 inst_9924 ( .A(net_8841), .Z(net_9886) );
NAND2_X2 inst_3845 ( .A1(net_6705), .A2(net_1497), .ZN(net_1492) );
CLKBUF_X2 inst_10124 ( .A(net_9024), .Z(net_10086) );
INV_X4 inst_5168 ( .ZN(net_788), .A(net_541) );
NAND2_X2 inst_3128 ( .ZN(net_4835), .A2(net_4153), .A1(net_2194) );
CLKBUF_X2 inst_10715 ( .A(net_8938), .Z(net_10677) );
SDFF_X2 inst_1078 ( .SI(net_7064), .Q(net_7064), .D(net_3799), .SE(net_3747), .CK(net_11928) );
NAND2_X1 inst_4322 ( .ZN(net_4542), .A2(net_3870), .A1(net_1352) );
NOR2_X2 inst_2517 ( .A1(net_6421), .ZN(net_1937), .A2(net_1071) );
DFF_X1 inst_6497 ( .QN(net_7409), .D(net_5540), .CK(net_12119) );
NAND2_X2 inst_4183 ( .A1(net_6688), .ZN(net_698), .A2(net_632) );
CLKBUF_X2 inst_10806 ( .A(net_10767), .Z(net_10768) );
NAND2_X2 inst_3557 ( .ZN(net_2510), .A2(net_2034), .A1(net_1783) );
OAI21_X2 inst_1992 ( .ZN(net_4601), .B2(net_4600), .B1(net_4228), .A(net_3616) );
SDFF_X2 inst_1039 ( .Q(net_7542), .D(net_7542), .SE(net_3896), .SI(net_376), .CK(net_10257) );
SDFF_X2 inst_714 ( .SI(net_6787), .Q(net_6787), .D(net_3821), .SE(net_3816), .CK(net_11321) );
NAND2_X2 inst_3005 ( .A1(net_6852), .ZN(net_5005), .A2(net_5004) );
NAND2_X4 inst_2895 ( .ZN(net_3437), .A1(net_3258), .A2(net_3255) );
INV_X4 inst_5449 ( .A(net_7563), .ZN(net_1913) );
CLKBUF_X2 inst_9005 ( .A(net_8966), .Z(net_8967) );
NAND2_X2 inst_4048 ( .A1(net_6520), .A2(net_1645), .ZN(net_1004) );
AOI222_X2 inst_7549 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1857), .A1(net_1856), .B1(net_1855), .C1(net_1854) );
NAND2_X2 inst_4003 ( .ZN(net_1281), .A1(net_678), .A2(net_639) );
DFF_X1 inst_6868 ( .D(net_2536), .Q(net_195), .CK(net_12075) );
SDFF_X2 inst_1061 ( .SI(net_7046), .Q(net_7046), .D(net_3831), .SE(net_3818), .CK(net_11930) );
INV_X4 inst_5033 ( .A(net_7821), .ZN(net_3788) );
CLKBUF_X2 inst_8306 ( .A(net_8267), .Z(net_8268) );
CLKBUF_X2 inst_13966 ( .A(net_10420), .Z(net_13928) );
CLKBUF_X2 inst_11201 ( .A(net_11162), .Z(net_11163) );
NOR2_X2 inst_2326 ( .A2(net_6292), .A1(net_5840), .ZN(net_5815) );
CLKBUF_X2 inst_8846 ( .A(net_8807), .Z(net_8808) );
INV_X4 inst_5363 ( .A(net_6026), .ZN(net_2611) );
DFF_X1 inst_6657 ( .QN(net_7664), .D(net_5188), .CK(net_13424) );
XNOR2_X2 inst_72 ( .ZN(net_1932), .B(net_672), .A(net_630) );
DFFR_X2 inst_6967 ( .QN(net_6048), .D(net_3999), .CK(net_10533), .RN(x1822) );
CLKBUF_X2 inst_11703 ( .A(net_10165), .Z(net_11665) );
NAND2_X2 inst_3542 ( .ZN(net_2525), .A2(net_2137), .A1(net_1189) );
OAI222_X2 inst_1634 ( .A1(net_5863), .C2(net_5057), .ZN(net_5056), .A2(net_5055), .B2(net_5054), .B1(net_2448), .C1(net_507) );
CLKBUF_X2 inst_8998 ( .A(net_7991), .Z(net_8960) );
DFF_X2 inst_6300 ( .D(net_1693), .QN(net_228), .CK(net_9489) );
XNOR2_X2 inst_115 ( .A(net_2575), .ZN(net_819), .B(net_818) );
CLKBUF_X2 inst_7980 ( .A(net_7881), .Z(net_7942) );
CLKBUF_X2 inst_10619 ( .A(net_8999), .Z(net_10581) );
DFF_X1 inst_6729 ( .QN(net_7363), .D(net_5326), .CK(net_9957) );
DFF_X1 inst_6650 ( .QN(net_7625), .D(net_5197), .CK(net_10557) );
CLKBUF_X2 inst_9485 ( .A(net_8354), .Z(net_9447) );
INV_X4 inst_4691 ( .ZN(net_4149), .A(net_3329) );
NAND2_X2 inst_3726 ( .A1(net_6763), .A2(net_1635), .ZN(net_1619) );
CLKBUF_X2 inst_12415 ( .A(net_12376), .Z(net_12377) );
CLKBUF_X2 inst_12357 ( .A(net_12318), .Z(net_12319) );
INV_X4 inst_4638 ( .ZN(net_4184), .A(net_4027) );
NAND2_X2 inst_3045 ( .A1(net_7027), .A2(net_4979), .ZN(net_4962) );
CLKBUF_X2 inst_11487 ( .A(net_9452), .Z(net_11449) );
CLKBUF_X2 inst_9801 ( .A(net_9762), .Z(net_9763) );
CLKBUF_X2 inst_13426 ( .A(net_7907), .Z(net_13388) );
OAI22_X2 inst_1582 ( .B1(net_6023), .B2(net_3200), .ZN(net_3197), .A2(net_3196), .A1(net_828) );
CLKBUF_X2 inst_13202 ( .A(net_13163), .Z(net_13164) );
CLKBUF_X2 inst_12741 ( .A(net_10787), .Z(net_12703) );
DFF_X2 inst_6334 ( .QN(net_7806), .CK(net_8674), .D(x1494) );
CLKBUF_X2 inst_13905 ( .A(net_13866), .Z(net_13867) );
INV_X2 inst_5846 ( .A(net_1153), .ZN(net_723) );
OAI21_X2 inst_1840 ( .B1(net_5361), .ZN(net_5332), .A(net_4372), .B2(net_3853) );
DFF_X1 inst_6345 ( .QN(net_6186), .D(net_5839), .CK(net_13642) );
SDFF_X2 inst_133 ( .Q(net_6217), .SI(net_6216), .SE(net_392), .D(net_151), .CK(net_14238) );
SDFF_X2 inst_1263 ( .D(net_6389), .SE(net_6051), .SI(net_307), .Q(net_307), .CK(net_14207) );
INV_X2 inst_6113 ( .A(net_5924), .ZN(net_5923) );
CLKBUF_X2 inst_13847 ( .A(net_9196), .Z(net_13809) );
NAND2_X2 inst_3330 ( .ZN(net_3586), .A1(net_3585), .A2(net_3226) );
CLKBUF_X2 inst_8047 ( .A(net_8008), .Z(net_8009) );
CLKBUF_X2 inst_9988 ( .A(net_9949), .Z(net_9950) );
CLKBUF_X2 inst_10225 ( .A(net_10186), .Z(net_10187) );
OAI21_X2 inst_1721 ( .ZN(net_5573), .B1(net_5448), .A(net_4838), .B2(net_4153) );
AOI22_X2 inst_7374 ( .A2(net_5916), .B2(net_2957), .ZN(net_2947), .B1(net_2682), .A1(net_850) );
OAI22_X2 inst_1445 ( .B2(net_5897), .B1(net_4660), .ZN(net_4630), .A2(net_4629), .A1(net_4091) );
CLKBUF_X2 inst_11907 ( .A(net_8563), .Z(net_11869) );
CLKBUF_X2 inst_9744 ( .A(net_9705), .Z(net_9706) );
CLKBUF_X2 inst_10884 ( .A(net_10845), .Z(net_10846) );
NAND2_X2 inst_3990 ( .A1(net_6635), .A2(net_1624), .ZN(net_1274) );
CLKBUF_X2 inst_8976 ( .A(net_8788), .Z(net_8938) );
CLKBUF_X2 inst_13156 ( .A(net_11543), .Z(net_13118) );
CLKBUF_X2 inst_12854 ( .A(net_9621), .Z(net_12816) );
CLKBUF_X2 inst_12115 ( .A(net_8152), .Z(net_12077) );
SDFF_X2 inst_126 ( .Q(net_6196), .SI(net_6195), .D(net_3921), .SE(net_392), .CK(net_13754) );
INV_X2 inst_5982 ( .A(net_7593), .ZN(net_1315) );
CLKBUF_X2 inst_7931 ( .A(net_7892), .Z(net_7893) );
OAI22_X2 inst_1512 ( .B1(net_4650), .A1(net_4080), .B2(net_4076), .ZN(net_4073), .A2(net_4072) );
CLKBUF_X2 inst_7932 ( .A(net_7893), .Z(net_7894) );
NAND2_X2 inst_3887 ( .A2(net_1696), .ZN(net_1432), .A1(net_1431) );
CLKBUF_X2 inst_10366 ( .A(net_10327), .Z(net_10328) );
CLKBUF_X2 inst_14163 ( .A(net_14124), .Z(net_14125) );
INV_X4 inst_5160 ( .ZN(net_553), .A(net_552) );
CLKBUF_X2 inst_8733 ( .A(net_8694), .Z(net_8695) );
OAI222_X2 inst_1631 ( .A1(net_5864), .C2(net_5383), .ZN(net_5091), .A2(net_5090), .B2(net_5089), .B1(net_2446), .C1(net_519) );
CLKBUF_X2 inst_13209 ( .A(net_13170), .Z(net_13171) );
CLKBUF_X2 inst_12651 ( .A(net_12612), .Z(net_12613) );
AOI222_X2 inst_7510 ( .B1(net_7368), .C1(net_7304), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2034), .A1(net_2033) );
CLKBUF_X2 inst_14395 ( .A(net_14356), .Z(net_14357) );
CLKBUF_X2 inst_13106 ( .A(net_8165), .Z(net_13068) );
SDFF_X2 inst_1086 ( .SI(net_7086), .Q(net_7086), .D(net_3790), .SE(net_3747), .CK(net_10980) );
CLKBUF_X2 inst_14360 ( .A(net_14321), .Z(net_14322) );
CLKBUF_X2 inst_10727 ( .A(net_10246), .Z(net_10689) );
NAND3_X2 inst_2643 ( .ZN(net_5945), .A3(net_3967), .A2(net_1967), .A1(net_794) );
CLKBUF_X2 inst_12088 ( .A(net_11740), .Z(net_12050) );
CLKBUF_X2 inst_13950 ( .A(net_13911), .Z(net_13912) );
CLKBUF_X2 inst_12615 ( .A(net_12576), .Z(net_12577) );
AOI21_X2 inst_7692 ( .B1(net_6733), .ZN(net_4519), .B2(net_2581), .A(net_2372) );
CLKBUF_X2 inst_12713 ( .A(net_9979), .Z(net_12675) );
OAI21_X2 inst_1688 ( .B1(net_5778), .ZN(net_5776), .A(net_5709), .B2(net_5708) );
CLKBUF_X2 inst_11691 ( .A(net_11652), .Z(net_11653) );
NOR2_X2 inst_2299 ( .A2(net_6188), .ZN(net_5844), .A1(net_5843) );
CLKBUF_X2 inst_13651 ( .A(net_13612), .Z(net_13613) );
CLKBUF_X2 inst_12441 ( .A(net_8455), .Z(net_12403) );
CLKBUF_X2 inst_13732 ( .A(net_13693), .Z(net_13694) );
CLKBUF_X2 inst_12146 ( .A(net_12107), .Z(net_12108) );
AOI222_X2 inst_7504 ( .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2056), .A1(net_2055), .B1(net_2054), .C1(net_2053) );
INV_X4 inst_5292 ( .A(net_7580), .ZN(net_1879) );
CLKBUF_X2 inst_13084 ( .A(net_13045), .Z(net_13046) );
SDFF_X2 inst_914 ( .Q(net_7132), .D(net_7132), .SE(net_3903), .SI(net_3806), .CK(net_7912) );
DFF_X1 inst_6364 ( .QN(net_6298), .D(net_5820), .CK(net_13797) );
INV_X4 inst_5170 ( .ZN(net_3224), .A(net_538) );
AOI222_X2 inst_7578 ( .A1(net_7545), .ZN(net_5196), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_377), .C2(net_375) );
INV_X4 inst_5182 ( .A(net_712), .ZN(net_521) );
CLKBUF_X2 inst_12366 ( .A(net_12327), .Z(net_12328) );
CLKBUF_X2 inst_12198 ( .A(net_12159), .Z(net_12160) );
CLKBUF_X2 inst_8166 ( .A(net_8127), .Z(net_8128) );
CLKBUF_X2 inst_11588 ( .A(net_11549), .Z(net_11550) );
OAI221_X2 inst_1642 ( .ZN(net_5453), .B2(net_5077), .C2(net_5075), .A(net_4983), .C1(net_1148), .B1(net_762) );
SDFF_X2 inst_384 ( .SI(net_7302), .Q(net_7302), .D(net_4783), .SE(net_3859), .CK(net_9930) );
SDFF_X2 inst_1252 ( .SI(net_6549), .Q(net_6549), .D(net_3821), .SE(net_3756), .CK(net_11217) );
CLKBUF_X2 inst_12773 ( .A(net_12734), .Z(net_12735) );
NAND2_X2 inst_3800 ( .A1(net_7034), .A2(net_1975), .ZN(net_1545) );
CLKBUF_X2 inst_12703 ( .A(net_8404), .Z(net_12665) );
CLKBUF_X2 inst_13434 ( .A(net_13395), .Z(net_13396) );
SDFF_X2 inst_199 ( .Q(net_6315), .SI(net_6314), .D(net_3693), .SE(net_392), .CK(net_13586) );
INV_X2 inst_6086 ( .A(net_7595), .ZN(net_1513) );
CLKBUF_X2 inst_12540 ( .A(net_12501), .Z(net_12502) );
CLKBUF_X2 inst_13259 ( .A(net_10794), .Z(net_13221) );
CLKBUF_X2 inst_12989 ( .A(net_12950), .Z(net_12951) );
CLKBUF_X2 inst_10271 ( .A(net_8971), .Z(net_10233) );
NOR3_X2 inst_2209 ( .A3(net_2384), .ZN(net_2383), .A2(net_2382), .A1(net_1822) );
NAND3_X2 inst_2722 ( .ZN(net_2379), .A3(net_1531), .A1(net_1474), .A2(net_972) );
CLKBUF_X2 inst_13034 ( .A(net_9660), .Z(net_12996) );
SDFF_X2 inst_1238 ( .SI(net_6531), .Q(net_6531), .D(net_3813), .SE(net_3755), .CK(net_8614) );
DFF_X1 inst_6764 ( .QN(net_6166), .D(net_4654), .CK(net_7952) );
AOI22_X2 inst_7361 ( .ZN(net_2992), .A2(net_2991), .B2(net_2990), .A1(net_1310), .B1(net_920) );
NOR4_X2 inst_2171 ( .ZN(net_3250), .A4(net_3122), .A1(net_2634), .A3(net_2480), .A2(net_819) );
CLKBUF_X2 inst_13313 ( .A(net_13274), .Z(net_13275) );
DFFR_X2 inst_6976 ( .QN(net_7787), .D(net_3997), .CK(net_13027), .RN(x1822) );
CLKBUF_X2 inst_9031 ( .A(net_8992), .Z(net_8993) );
CLKBUF_X2 inst_7941 ( .A(net_7875), .Z(net_7903) );
CLKBUF_X2 inst_14274 ( .A(net_13389), .Z(net_14236) );
CLKBUF_X2 inst_8527 ( .A(net_8142), .Z(net_8489) );
INV_X4 inst_4875 ( .ZN(net_1055), .A(net_611) );
NAND2_X2 inst_3402 ( .A2(net_5980), .ZN(net_3377), .A1(net_2882) );
CLKBUF_X2 inst_14252 ( .A(net_14213), .Z(net_14214) );
CLKBUF_X2 inst_14318 ( .A(net_8878), .Z(net_14280) );
SDFF_X2 inst_1011 ( .SI(net_6504), .Q(net_6504), .SE(net_3886), .D(net_3785), .CK(net_8768) );
SDFF_X2 inst_540 ( .Q(net_7243), .D(net_7243), .SE(net_3822), .SI(net_339), .CK(net_9838) );
NAND2_X2 inst_4114 ( .A2(net_1222), .ZN(net_1066), .A1(net_340) );
NOR2_X2 inst_2356 ( .ZN(net_5648), .A1(net_5500), .A2(net_4463) );
SDFF_X2 inst_404 ( .SI(net_7368), .Q(net_7368), .D(net_4782), .SE(net_3853), .CK(net_9904) );
SDFF_X2 inst_998 ( .Q(net_6458), .D(net_6458), .SE(net_3904), .SI(net_3802), .CK(net_11659) );
INV_X2 inst_6044 ( .A(net_7585), .ZN(net_2099) );
CLKBUF_X2 inst_7989 ( .A(net_7950), .Z(net_7951) );
NAND2_X2 inst_3209 ( .ZN(net_4717), .A2(net_3986), .A1(net_1848) );
INV_X2 inst_5952 ( .ZN(net_1125), .A(net_116) );
INV_X2 inst_5838 ( .ZN(net_794), .A(net_793) );
NAND2_X2 inst_3615 ( .ZN(net_2267), .A2(net_1935), .A1(net_1300) );
CLKBUF_X2 inst_9628 ( .A(net_9589), .Z(net_9590) );
CLKBUF_X2 inst_13989 ( .A(net_13950), .Z(net_13951) );
CLKBUF_X2 inst_14042 ( .A(net_12648), .Z(net_14004) );
CLKBUF_X2 inst_12298 ( .A(net_9273), .Z(net_12260) );
CLKBUF_X2 inst_9730 ( .A(net_9691), .Z(net_9692) );
NAND2_X2 inst_3216 ( .ZN(net_4710), .A2(net_3986), .A1(net_2136) );
CLKBUF_X2 inst_8748 ( .A(net_8709), .Z(net_8710) );
CLKBUF_X2 inst_9792 ( .A(net_9753), .Z(net_9754) );
CLKBUF_X2 inst_11442 ( .A(net_9488), .Z(net_11404) );
CLKBUF_X2 inst_10205 ( .A(net_10166), .Z(net_10167) );
CLKBUF_X2 inst_9242 ( .A(net_9203), .Z(net_9204) );
INV_X4 inst_5090 ( .A(net_2883), .ZN(net_805) );
CLKBUF_X2 inst_14400 ( .A(net_14361), .Z(net_14362) );
SDFF_X2 inst_192 ( .Q(net_6262), .SI(net_6261), .D(net_3489), .SE(net_392), .CK(net_13776) );
DFF_X1 inst_6720 ( .QN(net_7322), .D(net_5338), .CK(net_12706) );
NAND3_X2 inst_2715 ( .ZN(net_2461), .A2(net_1812), .A3(net_1569), .A1(net_1435) );
CLKBUF_X2 inst_13059 ( .A(net_13020), .Z(net_13021) );
NAND2_X1 inst_4242 ( .ZN(net_4685), .A2(net_3989), .A1(net_2096) );
NAND2_X2 inst_3540 ( .ZN(net_2527), .A2(net_2118), .A1(net_1780) );
AOI21_X2 inst_7701 ( .B1(net_7137), .ZN(net_4460), .B2(net_2582), .A(net_2380) );
NAND2_X2 inst_4126 ( .A2(net_1228), .ZN(net_1164), .A1(net_378) );
AOI22_X2 inst_7434 ( .ZN(net_2716), .A2(net_2715), .B2(net_2714), .B1(net_1700), .A1(net_1273) );
CLKBUF_X2 inst_14005 ( .A(net_13966), .Z(net_13967) );
CLKBUF_X2 inst_10904 ( .A(net_10203), .Z(net_10866) );
CLKBUF_X2 inst_8741 ( .A(net_8328), .Z(net_8703) );
NAND2_X2 inst_3547 ( .ZN(net_2520), .A2(net_2068), .A1(net_1775) );
NAND2_X2 inst_4178 ( .A2(net_6958), .ZN(net_773), .A1(net_566) );
CLKBUF_X2 inst_12720 ( .A(net_12681), .Z(net_12682) );
NOR2_X2 inst_2413 ( .A1(net_6030), .ZN(net_3410), .A2(net_3403) );
OAI22_X2 inst_1574 ( .A2(net_3297), .B2(net_3286), .ZN(net_3272), .A1(net_3174), .B1(net_555) );
DFF_X1 inst_6558 ( .QN(net_7451), .D(net_5048), .CK(net_12102) );
AOI222_X2 inst_7528 ( .C1(net_7526), .B1(net_7494), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_1982), .A1(net_1981) );
CLKBUF_X2 inst_9739 ( .A(net_9700), .Z(net_9701) );
SDFF_X2 inst_228 ( .Q(net_6326), .SI(net_6325), .D(net_3633), .SE(net_392), .CK(net_14025) );
SDFF_X2 inst_486 ( .Q(net_7544), .D(net_7544), .SE(net_3896), .SI(net_378), .CK(net_13120) );
CLKBUF_X2 inst_12977 ( .A(net_12721), .Z(net_12939) );
CLKBUF_X2 inst_14034 ( .A(net_13995), .Z(net_13996) );
DFF_X1 inst_6872 ( .D(net_2531), .QN(net_209), .CK(net_12608) );
CLKBUF_X2 inst_13365 ( .A(net_11655), .Z(net_13327) );
CLKBUF_X2 inst_12008 ( .A(net_11969), .Z(net_11970) );
SDFF_X2 inst_1240 ( .D(net_7807), .SI(net_6534), .Q(net_6534), .SE(net_3755), .CK(net_8611) );
INV_X4 inst_5445 ( .A(net_6096), .ZN(net_3511) );
DFF_X1 inst_6597 ( .QN(net_7466), .D(net_5413), .CK(net_9982) );
CLKBUF_X2 inst_12279 ( .A(net_12240), .Z(net_12241) );
CLKBUF_X2 inst_8759 ( .A(net_8720), .Z(net_8721) );
SDFF_X2 inst_244 ( .Q(net_6350), .SI(net_6349), .D(net_3613), .SE(net_392), .CK(net_13940) );
CLKBUF_X2 inst_13514 ( .A(net_13475), .Z(net_13476) );
INV_X4 inst_5262 ( .ZN(net_428), .A(net_427) );
CLKBUF_X2 inst_11472 ( .A(net_8036), .Z(net_11434) );
CLKBUF_X2 inst_13464 ( .A(net_13425), .Z(net_13426) );
CLKBUF_X2 inst_12136 ( .A(net_11670), .Z(net_12098) );
CLKBUF_X2 inst_11794 ( .A(net_11755), .Z(net_11756) );
INV_X4 inst_5537 ( .A(net_6100), .ZN(net_3503) );
CLKBUF_X2 inst_9186 ( .A(net_9147), .Z(net_9148) );
OAI22_X2 inst_1521 ( .B1(net_4644), .B2(net_4062), .A1(net_4057), .ZN(net_4054), .A2(net_4053) );
CLKBUF_X2 inst_11339 ( .A(net_11300), .Z(net_11301) );
DFF_X1 inst_6620 ( .QN(net_7581), .D(net_5387), .CK(net_10307) );
CLKBUF_X2 inst_13692 ( .A(net_9476), .Z(net_13654) );
CLKBUF_X2 inst_9679 ( .A(net_9640), .Z(net_9641) );
NAND2_X2 inst_3079 ( .A1(net_6480), .A2(net_4927), .ZN(net_4924) );
CLKBUF_X2 inst_12976 ( .A(net_12937), .Z(net_12938) );
CLKBUF_X2 inst_11208 ( .A(net_11169), .Z(net_11170) );
CLKBUF_X2 inst_10766 ( .A(net_10554), .Z(net_10728) );
NAND4_X2 inst_2563 ( .ZN(net_1674), .A3(net_852), .A1(net_849), .A4(net_846), .A2(net_843) );
SDFF_X2 inst_1306 ( .D(net_6386), .SE(net_6051), .SI(net_304), .Q(net_304), .CK(net_13718) );
INV_X4 inst_4845 ( .ZN(net_5101), .A(net_1065) );
CLKBUF_X2 inst_10143 ( .A(net_9906), .Z(net_10105) );
CLKBUF_X2 inst_12529 ( .A(net_12490), .Z(net_12491) );
CLKBUF_X2 inst_9931 ( .A(net_9892), .Z(net_9893) );
CLKBUF_X2 inst_12916 ( .A(net_12877), .Z(net_12878) );
OR2_X2 inst_1407 ( .A1(net_6408), .ZN(net_2418), .A2(net_1921) );
INV_X4 inst_5487 ( .A(net_7274), .ZN(net_2031) );
CLKBUF_X2 inst_8096 ( .A(net_7832), .Z(net_8058) );
CLKBUF_X2 inst_13803 ( .A(net_13764), .Z(net_13765) );
CLKBUF_X2 inst_13128 ( .A(net_10373), .Z(net_13090) );
AOI222_X2 inst_7599 ( .A1(net_7239), .ZN(net_5343), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_333), .C2(net_331) );
DFFR_X2 inst_7018 ( .D(net_3285), .QN(net_293), .CK(net_13295), .RN(x1822) );
CLKBUF_X2 inst_11789 ( .A(net_11750), .Z(net_11751) );
CLKBUF_X2 inst_9132 ( .A(net_9093), .Z(net_9094) );
INV_X2 inst_6052 ( .ZN(net_1257), .A(net_129) );
CLKBUF_X2 inst_10303 ( .A(net_9408), .Z(net_10265) );
CLKBUF_X2 inst_11526 ( .A(net_11487), .Z(net_11488) );
NAND2_X2 inst_3606 ( .ZN(net_2392), .A2(net_1904), .A1(net_1373) );
XNOR2_X2 inst_93 ( .B(net_3002), .ZN(net_1661), .A(net_1152) );
INV_X4 inst_4832 ( .ZN(net_1078), .A(net_1077) );
DFFR_X2 inst_7026 ( .D(net_3296), .QN(net_268), .CK(net_12422), .RN(x1822) );
DFFR_X2 inst_6965 ( .QN(net_7783), .D(net_4160), .CK(net_10251), .RN(x1822) );
CLKBUF_X2 inst_11051 ( .A(net_11012), .Z(net_11013) );
CLKBUF_X2 inst_12105 ( .A(net_10556), .Z(net_12067) );
CLKBUF_X2 inst_10217 ( .A(net_9648), .Z(net_10179) );
CLKBUF_X2 inst_9687 ( .A(net_9648), .Z(net_9649) );
AOI21_X2 inst_7784 ( .B1(net_6596), .ZN(net_5913), .B2(net_2583), .A(net_2278) );
INV_X4 inst_4595 ( .ZN(net_5085), .A(net_4294) );
INV_X4 inst_5099 ( .A(net_3238), .ZN(net_619) );
CLKBUF_X2 inst_11116 ( .A(net_11077), .Z(net_11078) );
INV_X16 inst_6134 ( .ZN(net_3105), .A(net_2627) );
OAI221_X2 inst_1675 ( .ZN(net_4108), .C2(net_4107), .B2(net_4008), .C1(net_3985), .A(net_3863), .B1(net_1926) );
CLKBUF_X2 inst_9561 ( .A(net_9411), .Z(net_9523) );
SDFF_X2 inst_584 ( .Q(net_6582), .D(net_6582), .SE(net_3823), .SI(net_3803), .CK(net_10669) );
CLKBUF_X2 inst_11086 ( .A(net_11047), .Z(net_11048) );
NAND2_X2 inst_3433 ( .ZN(net_3215), .A2(net_3099), .A1(net_2764) );
CLKBUF_X2 inst_8668 ( .A(net_8105), .Z(net_8630) );
SDFF_X2 inst_470 ( .Q(net_7017), .D(net_7017), .SI(net_3900), .SE(net_3899), .CK(net_11912) );
CLKBUF_X2 inst_11274 ( .A(net_11235), .Z(net_11236) );
INV_X4 inst_5149 ( .ZN(net_1147), .A(net_567) );
CLKBUF_X2 inst_8958 ( .A(net_8222), .Z(net_8920) );
CLKBUF_X2 inst_12917 ( .A(net_11775), .Z(net_12879) );
CLKBUF_X2 inst_13713 ( .A(net_13674), .Z(net_13675) );
NAND2_X1 inst_4237 ( .ZN(net_4690), .A2(net_3989), .A1(net_2124) );
CLKBUF_X2 inst_10709 ( .A(net_10670), .Z(net_10671) );
CLKBUF_X2 inst_8138 ( .A(net_8099), .Z(net_8100) );
SDFF_X2 inst_148 ( .Q(net_6230), .SI(net_6229), .SE(net_392), .D(net_136), .CK(net_14105) );
INV_X8 inst_4490 ( .ZN(net_4644), .A(net_3409) );
SDFF_X2 inst_554 ( .Q(net_6445), .D(net_6445), .SI(net_3900), .SE(net_3820), .CK(net_10873) );
OAI21_X2 inst_1752 ( .ZN(net_5511), .A(net_4814), .B2(net_4153), .B1(net_1235) );
CLKBUF_X2 inst_13675 ( .A(net_13636), .Z(net_13637) );
CLKBUF_X2 inst_13621 ( .A(net_13582), .Z(net_13583) );
SDFF_X2 inst_1187 ( .SI(net_6932), .Q(net_6932), .D(net_3890), .SE(net_3741), .CK(net_11684) );
INV_X2 inst_6000 ( .A(net_7477), .ZN(net_2193) );
NAND2_X1 inst_4333 ( .ZN(net_4531), .A2(net_3870), .A1(net_1363) );
DFF_X1 inst_6816 ( .D(net_3205), .CK(net_13409), .Q(x249) );
SDFF_X2 inst_1063 ( .Q(net_6864), .D(net_6864), .SE(net_3901), .SI(net_3892), .CK(net_8922) );
INV_X4 inst_5499 ( .A(net_7694), .ZN(net_839) );
NAND3_X2 inst_2700 ( .ZN(net_2692), .A3(net_2572), .A2(net_2430), .A1(net_2267) );
CLKBUF_X2 inst_10740 ( .A(net_10701), .Z(net_10702) );
CLKBUF_X2 inst_8951 ( .A(net_8379), .Z(net_8913) );
OAI21_X2 inst_1917 ( .B1(net_5343), .ZN(net_5147), .A(net_4747), .B2(net_3941) );
NAND2_X2 inst_3252 ( .ZN(net_5052), .A1(net_3852), .A2(net_3464) );
CLKBUF_X2 inst_13542 ( .A(net_8086), .Z(net_13504) );
INV_X8 inst_4565 ( .ZN(net_1655), .A(net_528) );
CLKBUF_X2 inst_12695 ( .A(net_12656), .Z(net_12657) );
INV_X4 inst_4755 ( .ZN(net_2715), .A(net_2687) );
INV_X4 inst_4955 ( .ZN(net_727), .A(net_726) );
CLKBUF_X2 inst_11553 ( .A(net_11514), .Z(net_11515) );
CLKBUF_X2 inst_12386 ( .A(net_12347), .Z(net_12348) );
INV_X4 inst_5276 ( .ZN(net_795), .A(net_592) );
CLKBUF_X2 inst_9452 ( .A(net_9413), .Z(net_9414) );
SDFF_X2 inst_1167 ( .SI(net_6937), .Q(net_6937), .D(net_3812), .SE(net_3734), .CK(net_11448) );
OAI21_X2 inst_2087 ( .B1(net_5903), .B2(net_4415), .ZN(net_4401), .A(net_3520) );
DFF_X1 inst_6879 ( .D(net_2529), .Q(net_230), .CK(net_9431) );
CLKBUF_X2 inst_8767 ( .A(net_8728), .Z(net_8729) );
CLKBUF_X2 inst_13891 ( .A(net_13852), .Z(net_13853) );
CLKBUF_X2 inst_9881 ( .A(net_9842), .Z(net_9843) );
SDFF_X2 inst_1303 ( .SI(net_7762), .Q(net_7762), .SE(net_5921), .D(net_2748), .CK(net_12739) );
OAI22_X2 inst_1623 ( .B1(net_5937), .A1(net_2784), .ZN(net_2781), .B2(net_215), .A2(net_178) );
CLKBUF_X2 inst_8571 ( .A(net_8532), .Z(net_8533) );
CLKBUF_X2 inst_12788 ( .A(net_12749), .Z(net_12750) );
NAND2_X2 inst_4088 ( .A1(net_7212), .A2(net_1648), .ZN(net_964) );
INV_X1 inst_6163 ( .A(net_5929), .ZN(net_5928) );
INV_X4 inst_4922 ( .A(net_3778), .ZN(net_822) );
DFF_X1 inst_6501 ( .QN(net_7423), .D(net_5530), .CK(net_12624) );
SDFF_X2 inst_819 ( .Q(net_6966), .D(net_6966), .SE(net_3891), .SI(net_3802), .CK(net_9099) );
INV_X8 inst_4464 ( .ZN(net_5279), .A(net_4287) );
NAND2_X2 inst_3320 ( .ZN(net_3606), .A1(net_3605), .A2(net_3228) );
CLKBUF_X2 inst_8369 ( .A(net_8128), .Z(net_8331) );
OAI22_X2 inst_1468 ( .B2(net_5052), .ZN(net_4394), .A1(net_4141), .A2(net_3825), .B1(net_1179) );
CLKBUF_X2 inst_10183 ( .A(net_10144), .Z(net_10145) );
CLKBUF_X2 inst_9663 ( .A(net_9624), .Z(net_9625) );
NAND2_X2 inst_3452 ( .A2(net_5925), .ZN(net_2920), .A1(net_1213) );
NAND2_X2 inst_3776 ( .A1(net_7031), .A2(net_1975), .ZN(net_1569) );
OAI22_X2 inst_1516 ( .B1(net_4650), .A1(net_4080), .B2(net_4066), .ZN(net_4065), .A2(net_4064) );
CLKBUF_X2 inst_14046 ( .A(net_14007), .Z(net_14008) );
SDFF_X2 inst_386 ( .SI(net_7305), .Q(net_7305), .D(net_4781), .SE(net_3859), .CK(net_12766) );
CLKBUF_X2 inst_12372 ( .A(net_12333), .Z(net_12334) );
CLKBUF_X2 inst_8497 ( .A(net_8458), .Z(net_8459) );
CLKBUF_X2 inst_8857 ( .A(net_8818), .Z(net_8819) );
INV_X2 inst_5859 ( .ZN(net_622), .A(net_621) );
AOI22_X2 inst_7255 ( .B1(net_6811), .A1(net_6779), .A2(net_5316), .B2(net_5315), .ZN(net_5301) );
NAND3_X2 inst_2617 ( .ZN(net_5722), .A1(net_5617), .A2(net_5134), .A3(net_4181) );
CLKBUF_X2 inst_10543 ( .A(net_10504), .Z(net_10505) );
CLKBUF_X2 inst_9863 ( .A(net_9824), .Z(net_9825) );
CLKBUF_X2 inst_8089 ( .A(net_8050), .Z(net_8051) );
NAND2_X2 inst_3942 ( .A1(net_6435), .A2(net_1677), .ZN(net_1349) );
AND2_X4 inst_7826 ( .ZN(net_3114), .A2(net_3041), .A1(net_1247) );
CLKBUF_X2 inst_11040 ( .A(net_11001), .Z(net_11002) );
CLKBUF_X2 inst_9459 ( .A(net_8511), .Z(net_9421) );
NAND2_X2 inst_3068 ( .A1(net_7129), .A2(net_4950), .ZN(net_4937) );
INV_X4 inst_5225 ( .A(net_1220), .ZN(net_464) );
INV_X2 inst_5850 ( .A(net_681), .ZN(net_679) );
CLKBUF_X2 inst_10173 ( .A(net_10134), .Z(net_10135) );
CLKBUF_X2 inst_9826 ( .A(net_9787), .Z(net_9788) );
NAND3_X2 inst_2778 ( .ZN(net_2322), .A3(net_1534), .A1(net_1402), .A2(net_946) );
NOR2_X4 inst_2277 ( .ZN(net_3845), .A1(net_3404), .A2(net_3238) );
INV_X4 inst_5320 ( .A(net_7280), .ZN(net_2017) );
CLKBUF_X2 inst_9518 ( .A(net_9479), .Z(net_9480) );
CLKBUF_X2 inst_11883 ( .A(net_11844), .Z(net_11845) );
CLKBUF_X2 inst_8245 ( .A(net_8114), .Z(net_8207) );
INV_X4 inst_5223 ( .ZN(net_468), .A(net_467) );
INV_X4 inst_5468 ( .ZN(net_542), .A(net_277) );
CLKBUF_X2 inst_9599 ( .A(net_9172), .Z(net_9561) );
NAND2_X2 inst_2962 ( .ZN(net_5465), .A1(net_4896), .A2(net_4895) );
CLKBUF_X2 inst_10060 ( .A(net_10021), .Z(net_10022) );
CLKBUF_X2 inst_8716 ( .A(net_8677), .Z(net_8678) );
CLKBUF_X2 inst_11064 ( .A(net_11025), .Z(net_11026) );
CLKBUF_X2 inst_12375 ( .A(net_12336), .Z(net_12337) );
SDFF_X2 inst_811 ( .Q(net_6984), .D(net_6984), .SE(net_3891), .SI(net_3805), .CK(net_9033) );
CLKBUF_X2 inst_13973 ( .A(net_13934), .Z(net_13935) );
CLKBUF_X2 inst_10605 ( .A(net_10566), .Z(net_10567) );
CLKBUF_X2 inst_9973 ( .A(net_8802), .Z(net_9935) );
SDFF_X2 inst_208 ( .Q(net_6306), .SI(net_6305), .D(net_3675), .SE(net_392), .CK(net_13559) );
CLKBUF_X2 inst_13756 ( .A(net_13717), .Z(net_13718) );
CLKBUF_X2 inst_14272 ( .A(net_11705), .Z(net_14234) );
NAND2_X2 inst_4202 ( .ZN(net_1745), .A1(net_608), .A2(net_282) );
CLKBUF_X2 inst_9591 ( .A(net_7991), .Z(net_9553) );
NAND2_X2 inst_3774 ( .A1(net_7180), .A2(net_1637), .ZN(net_1571) );
DFFR_X2 inst_7101 ( .D(net_1952), .QN(net_115), .CK(net_9590), .RN(x1822) );
NAND2_X2 inst_3909 ( .ZN(net_1401), .A2(net_1400), .A1(net_1076) );
INV_X4 inst_5282 ( .ZN(net_1221), .A(net_269) );
OAI21_X2 inst_1869 ( .ZN(net_5242), .B1(net_5196), .A(net_4530), .B2(net_3870) );
SDFF_X2 inst_897 ( .Q(net_7101), .D(net_7101), .SE(net_3888), .SI(net_3802), .CK(net_10499) );
CLKBUF_X2 inst_12751 ( .A(net_12712), .Z(net_12713) );
CLKBUF_X2 inst_11935 ( .A(net_11896), .Z(net_11897) );
CLKBUF_X2 inst_10294 ( .A(net_10066), .Z(net_10256) );
NAND2_X2 inst_3945 ( .A1(net_7454), .A2(net_1696), .ZN(net_1343) );
CLKBUF_X2 inst_11656 ( .A(net_11617), .Z(net_11618) );
SDFF_X2 inst_1201 ( .SI(net_7084), .Q(net_7084), .D(net_3779), .SE(net_3742), .CK(net_8986) );
CLKBUF_X2 inst_8760 ( .A(net_8721), .Z(net_8722) );
INV_X2 inst_5899 ( .A(net_7659), .ZN(net_1912) );
CLKBUF_X2 inst_9294 ( .A(net_9216), .Z(net_9256) );
SDFF_X2 inst_636 ( .SI(net_6649), .Q(net_6649), .SE(net_3851), .D(net_3795), .CK(net_9110) );
OAI21_X2 inst_1927 ( .ZN(net_5118), .A(net_4775), .B2(net_3941), .B1(net_1175) );
SDFF_X2 inst_184 ( .Q(net_6270), .SI(net_6269), .D(net_3515), .SE(net_392), .CK(net_13916) );
OAI21_X2 inst_1847 ( .B1(net_5347), .ZN(net_5325), .A(net_4364), .B2(net_3853) );
CLKBUF_X2 inst_12499 ( .A(net_12460), .Z(net_12461) );
CLKBUF_X2 inst_8878 ( .A(net_8839), .Z(net_8840) );
CLKBUF_X2 inst_12270 ( .A(net_8156), .Z(net_12232) );
CLKBUF_X2 inst_11777 ( .A(net_11738), .Z(net_11739) );
OAI21_X2 inst_1907 ( .B1(net_5355), .ZN(net_5162), .A(net_4762), .B2(net_3941) );
DFF_X1 inst_6921 ( .D(net_2391), .Q(net_256), .CK(net_10810) );
DFFR_X2 inst_7015 ( .D(net_3278), .QN(net_289), .CK(net_11444), .RN(x1822) );
CLKBUF_X2 inst_8775 ( .A(net_8713), .Z(net_8737) );
CLKBUF_X2 inst_8384 ( .A(net_8345), .Z(net_8346) );
CLKBUF_X2 inst_10313 ( .A(net_9486), .Z(net_10275) );
NAND2_X2 inst_3836 ( .A1(net_6578), .A2(net_1705), .ZN(net_1503) );
DFFR_X2 inst_6999 ( .QN(net_7716), .D(net_3353), .CK(net_13226), .RN(x1822) );
CLKBUF_X2 inst_13461 ( .A(net_13422), .Z(net_13423) );
CLKBUF_X2 inst_9409 ( .A(net_8752), .Z(net_9371) );
CLKBUF_X2 inst_8472 ( .A(net_8433), .Z(net_8434) );
AOI21_X2 inst_7742 ( .B1(net_6598), .ZN(net_4416), .B2(net_2583), .A(net_2291) );
CLKBUF_X2 inst_9125 ( .A(net_9086), .Z(net_9087) );
CLKBUF_X2 inst_10919 ( .A(net_10880), .Z(net_10881) );
NOR3_X2 inst_2192 ( .ZN(net_3885), .A1(net_3454), .A3(net_1737), .A2(net_793) );
INV_X2 inst_5980 ( .A(net_6413), .ZN(net_405) );
AND2_X4 inst_7806 ( .ZN(net_3848), .A2(net_3847), .A1(net_1144) );
OAI21_X2 inst_2114 ( .B1(net_7767), .A(net_5925), .ZN(net_3455), .B2(net_155) );
NAND3_X2 inst_2784 ( .ZN(net_2316), .A3(net_1587), .A1(net_1441), .A2(net_987) );
CLKBUF_X2 inst_13817 ( .A(net_13778), .Z(net_13779) );
NAND2_X2 inst_4216 ( .ZN(net_1040), .A2(x1126), .A1(x1101) );
DFF_X2 inst_6330 ( .QN(net_7804), .CK(net_11524), .D(x1511) );
XNOR2_X2 inst_106 ( .B(net_7782), .A(net_7781), .ZN(net_1041) );
CLKBUF_X2 inst_13001 ( .A(net_12962), .Z(net_12963) );
NAND3_X2 inst_2583 ( .ZN(net_5756), .A1(net_5651), .A2(net_5273), .A3(net_4311) );
CLKBUF_X2 inst_10753 ( .A(net_10714), .Z(net_10715) );
CLKBUF_X2 inst_9036 ( .A(net_8997), .Z(net_8998) );
CLKBUF_X2 inst_10538 ( .A(net_10284), .Z(net_10500) );
NAND2_X2 inst_3997 ( .A2(net_1910), .ZN(net_1189), .A1(net_1188) );
CLKBUF_X2 inst_13458 ( .A(net_12346), .Z(net_13420) );
CLKBUF_X2 inst_13697 ( .A(net_10099), .Z(net_13659) );
CLKBUF_X2 inst_11344 ( .A(net_8556), .Z(net_11306) );
NAND2_X1 inst_4377 ( .ZN(net_4350), .A2(net_3859), .A1(net_2013) );
INV_X4 inst_5241 ( .ZN(net_770), .A(net_449) );
CLKBUF_X2 inst_9903 ( .A(net_9864), .Z(net_9865) );
NAND2_X1 inst_4383 ( .ZN(net_4344), .A2(net_3859), .A1(net_2049) );
NAND2_X1 inst_4301 ( .ZN(net_4565), .A2(net_3866), .A1(net_1897) );
CLKBUF_X2 inst_13432 ( .A(net_13393), .Z(net_13394) );
CLKBUF_X2 inst_8537 ( .A(net_8498), .Z(net_8499) );
CLKBUF_X2 inst_9208 ( .A(net_9169), .Z(net_9170) );
OR2_X2 inst_1410 ( .A1(net_3985), .ZN(net_1686), .A2(net_1685) );
INV_X4 inst_5106 ( .A(net_6553), .ZN(net_613) );
CLKBUF_X2 inst_10675 ( .A(net_10636), .Z(net_10637) );
INV_X4 inst_5434 ( .A(net_7704), .ZN(net_841) );
CLKBUF_X2 inst_10418 ( .A(net_10379), .Z(net_10380) );
NAND2_X2 inst_3756 ( .A1(net_6628), .A2(net_1624), .ZN(net_1589) );
INV_X4 inst_4991 ( .A(net_7228), .ZN(net_1149) );
NAND2_X1 inst_4424 ( .A2(net_2131), .ZN(net_1466), .A1(net_1465) );
CLKBUF_X2 inst_10811 ( .A(net_8104), .Z(net_10773) );
OAI21_X2 inst_1733 ( .ZN(net_5558), .B1(net_5410), .A(net_4816), .B2(net_4153) );
CLKBUF_X2 inst_9489 ( .A(net_9450), .Z(net_9451) );
CLKBUF_X2 inst_8832 ( .A(net_8709), .Z(net_8794) );
CLKBUF_X2 inst_11714 ( .A(net_8439), .Z(net_11676) );
DFFR_X2 inst_7028 ( .D(net_3267), .QN(net_292), .CK(net_11433), .RN(x1822) );
CLKBUF_X2 inst_8911 ( .A(net_8777), .Z(net_8873) );
NAND2_X2 inst_3900 ( .A2(net_1696), .ZN(net_1412), .A1(net_1411) );
NOR3_X2 inst_2199 ( .ZN(net_3450), .A3(net_3149), .A2(net_3011), .A1(net_2869) );
SDFF_X2 inst_918 ( .Q(net_7155), .D(net_7155), .SE(net_3903), .SI(net_3791), .CK(net_8707) );
INV_X4 inst_4751 ( .ZN(net_2629), .A(net_263) );
INV_X2 inst_5994 ( .A(net_7480), .ZN(net_2177) );
DFF_X1 inst_6588 ( .QN(net_7558), .D(net_5062), .CK(net_10588) );
AOI21_X2 inst_7678 ( .B1(net_7015), .ZN(net_4214), .A(net_2464), .B2(net_1100) );
CLKBUF_X2 inst_10210 ( .A(net_10171), .Z(net_10172) );
CLKBUF_X2 inst_13921 ( .A(net_13882), .Z(net_13883) );
DFF_X1 inst_6653 ( .QN(net_7660), .D(net_5192), .CK(net_13067) );
CLKBUF_X2 inst_9177 ( .A(net_9138), .Z(net_9139) );
OAI21_X2 inst_2074 ( .ZN(net_4419), .B1(net_4418), .B2(net_4415), .A(net_3516) );
NAND2_X2 inst_4035 ( .A1(net_6794), .A2(net_1651), .ZN(net_1017) );
CLKBUF_X2 inst_11330 ( .A(net_9128), .Z(net_11292) );
OAI21_X2 inst_1862 ( .ZN(net_5254), .B1(net_5220), .A(net_4541), .B2(net_3870) );
INV_X4 inst_4823 ( .A(net_3857), .ZN(net_1089) );
AOI22_X2 inst_7296 ( .B1(net_6546), .A1(net_6514), .A2(net_5184), .B2(net_5183), .ZN(net_5173) );
SDFF_X2 inst_221 ( .Q(net_6333), .SI(net_6332), .D(net_3659), .SE(net_392), .CK(net_14046) );
SDFF_X2 inst_1236 ( .SI(net_6520), .Q(net_6520), .D(net_3797), .SE(net_3755), .CK(net_8757) );
CLKBUF_X2 inst_14108 ( .A(net_10107), .Z(net_14070) );
CLKBUF_X2 inst_12928 ( .A(net_12280), .Z(net_12890) );
INV_X4 inst_5112 ( .ZN(net_607), .A(net_606) );
CLKBUF_X2 inst_12640 ( .A(net_12601), .Z(net_12602) );
NAND2_X2 inst_3313 ( .ZN(net_3620), .A1(net_3619), .A2(net_3228) );
INV_X2 inst_5929 ( .A(net_7533), .ZN(net_409) );
CLKBUF_X2 inst_9545 ( .A(net_9506), .Z(net_9507) );
NAND2_X2 inst_3562 ( .ZN(net_2505), .A2(net_2024), .A1(net_1791) );
CLKBUF_X2 inst_13502 ( .A(net_13463), .Z(net_13464) );
AOI222_X2 inst_7466 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2187), .A1(net_2186), .B1(net_2185), .C1(net_2184) );
CLKBUF_X2 inst_11967 ( .A(net_8872), .Z(net_11929) );
NOR2_X2 inst_2334 ( .A2(net_6284), .A1(net_5840), .ZN(net_5807) );
NOR2_X2 inst_2429 ( .ZN(net_3426), .A2(net_3121), .A1(net_3046) );
NOR3_X2 inst_2210 ( .A3(net_2384), .ZN(net_2381), .A1(net_1825), .A2(net_878) );
CLKBUF_X2 inst_10596 ( .A(net_8981), .Z(net_10558) );
CLKBUF_X2 inst_10463 ( .A(net_10411), .Z(net_10425) );
SDFF_X2 inst_754 ( .Q(net_6876), .D(net_6876), .SE(net_3901), .SI(net_3787), .CK(net_11741) );
INV_X2 inst_6040 ( .A(net_7625), .ZN(net_1869) );
CLKBUF_X2 inst_10531 ( .A(net_10492), .Z(net_10493) );
CLKBUF_X2 inst_10030 ( .A(net_9991), .Z(net_9992) );
INV_X4 inst_5028 ( .A(net_7817), .ZN(net_3796) );
NAND3_X2 inst_2590 ( .ZN(net_5749), .A1(net_5644), .A2(net_5239), .A3(net_4208) );
CLKBUF_X2 inst_10332 ( .A(net_10293), .Z(net_10294) );
NAND2_X2 inst_2913 ( .ZN(net_5715), .A2(net_5714), .A1(net_2952) );
AOI21_X2 inst_7647 ( .ZN(net_5956), .B2(net_3439), .A(net_3218), .B1(net_1223) );
CLKBUF_X2 inst_11577 ( .A(net_11538), .Z(net_11539) );
CLKBUF_X2 inst_10949 ( .A(net_10887), .Z(net_10911) );
CLKBUF_X2 inst_10435 ( .A(net_8159), .Z(net_10397) );
CLKBUF_X2 inst_8783 ( .A(net_8576), .Z(net_8745) );
INV_X4 inst_5025 ( .A(net_3152), .ZN(net_868) );
NAND2_X2 inst_3295 ( .ZN(net_3656), .A1(net_3655), .A2(net_3229) );
CLKBUF_X2 inst_8792 ( .A(net_8003), .Z(net_8754) );
CLKBUF_X2 inst_13341 ( .A(net_13302), .Z(net_13303) );
INV_X4 inst_5057 ( .ZN(net_742), .A(net_640) );
CLKBUF_X2 inst_8828 ( .A(net_8549), .Z(net_8790) );
AOI22_X2 inst_7394 ( .A2(net_2957), .B1(net_2872), .ZN(net_2848), .A1(net_2847), .B2(net_157) );
CLKBUF_X2 inst_13997 ( .A(net_13958), .Z(net_13959) );
CLKBUF_X2 inst_13140 ( .A(net_12715), .Z(net_13102) );
CLKBUF_X2 inst_12451 ( .A(net_12412), .Z(net_12413) );
CLKBUF_X2 inst_12998 ( .A(net_12959), .Z(net_12960) );
NAND2_X1 inst_4459 ( .A2(net_1256), .ZN(net_1112), .A1(net_1111) );
NAND2_X2 inst_2923 ( .A2(net_7777), .ZN(net_5769), .A1(net_5605) );
CLKBUF_X2 inst_14028 ( .A(net_13989), .Z(net_13990) );
CLKBUF_X2 inst_7957 ( .A(net_7853), .Z(net_7919) );
NAND3_X2 inst_2707 ( .ZN(net_2470), .A2(net_1802), .A3(net_1551), .A1(net_1351) );
SDFF_X2 inst_1117 ( .SI(net_6665), .Q(net_6665), .D(net_3894), .SE(net_3465), .CK(net_9142) );
NAND2_X2 inst_4015 ( .A1(net_6936), .A2(net_1654), .ZN(net_1037) );
AOI22_X2 inst_7343 ( .ZN(net_3180), .A2(net_2978), .B2(net_2902), .A1(net_1744), .B1(net_934) );
CLKBUF_X2 inst_13909 ( .A(net_13870), .Z(net_13871) );
CLKBUF_X2 inst_11374 ( .A(net_11335), .Z(net_11336) );
NAND2_X2 inst_3958 ( .A1(net_6567), .A2(net_1705), .ZN(net_1326) );
DFF_X1 inst_6887 ( .D(net_2499), .Q(net_162), .CK(net_13054) );
NAND3_X2 inst_2725 ( .ZN(net_2376), .A3(net_1590), .A1(net_1496), .A2(net_983) );
INV_X4 inst_5141 ( .A(net_3106), .ZN(net_575) );
DFF_X1 inst_6681 ( .QN(net_7259), .D(net_5143), .CK(net_13000) );
CLKBUF_X2 inst_8204 ( .A(net_8165), .Z(net_8166) );
SDFF_X2 inst_334 ( .D(net_6393), .SE(net_6052), .SI(net_318), .Q(net_318), .CK(net_13820) );
OAI22_X2 inst_1610 ( .A1(net_3289), .A2(net_3087), .ZN(net_3085), .B2(net_3084), .B1(net_751) );
CLKBUF_X2 inst_10465 ( .A(net_10426), .Z(net_10427) );
CLKBUF_X2 inst_10166 ( .A(net_10127), .Z(net_10128) );
INV_X4 inst_4620 ( .ZN(net_4202), .A(net_4065) );
CLKBUF_X2 inst_12674 ( .A(net_12635), .Z(net_12636) );
CLKBUF_X2 inst_9277 ( .A(net_9238), .Z(net_9239) );
NAND2_X2 inst_3707 ( .A1(net_6502), .ZN(net_1643), .A2(net_1642) );
CLKBUF_X2 inst_13337 ( .A(net_13298), .Z(net_13299) );
CLKBUF_X2 inst_11869 ( .A(net_11830), .Z(net_11831) );
CLKBUF_X2 inst_14243 ( .A(net_14204), .Z(net_14205) );
SDFF_X2 inst_1042 ( .SI(net_6911), .Q(net_6911), .D(net_3897), .SE(net_3887), .CK(net_8843) );
CLKBUF_X2 inst_14190 ( .A(net_14151), .Z(net_14152) );
CLKBUF_X2 inst_12431 ( .A(net_12392), .Z(net_12393) );
CLKBUF_X2 inst_10158 ( .A(net_10119), .Z(net_10120) );
INV_X2 inst_5961 ( .A(net_7438), .ZN(net_1411) );
CLKBUF_X2 inst_8131 ( .A(net_8092), .Z(net_8093) );
INV_X4 inst_5388 ( .A(net_6007), .ZN(net_650) );
INV_X4 inst_5595 ( .A(net_6407), .ZN(net_484) );
INV_X8 inst_4492 ( .ZN(net_4637), .A(net_3407) );
CLKBUF_X2 inst_13551 ( .A(net_13512), .Z(net_13513) );
CLKBUF_X2 inst_8153 ( .A(net_7968), .Z(net_8115) );
CLKBUF_X2 inst_9773 ( .A(net_9734), .Z(net_9735) );
NAND2_X2 inst_3056 ( .A1(net_7155), .A2(net_4954), .ZN(net_4949) );
CLKBUF_X2 inst_12214 ( .A(net_9108), .Z(net_12176) );
CLKBUF_X2 inst_8058 ( .A(net_8004), .Z(net_8020) );
CLKBUF_X2 inst_13255 ( .A(net_13194), .Z(net_13217) );
SDFF_X2 inst_595 ( .SI(net_7799), .Q(net_6565), .D(net_6565), .SE(net_3823), .CK(net_12919) );
NAND3_X2 inst_2609 ( .ZN(net_5730), .A1(net_5625), .A2(net_5168), .A3(net_4190) );
NOR2_X2 inst_2556 ( .A2(net_6023), .A1(net_6017), .ZN(net_2889) );
INV_X4 inst_5002 ( .A(net_6958), .ZN(net_678) );
INV_X4 inst_5371 ( .A(net_6183), .ZN(net_3532) );
CLKBUF_X2 inst_8222 ( .A(net_8183), .Z(net_8184) );
OAI21_X2 inst_1704 ( .ZN(net_5590), .A(net_5213), .B2(net_4460), .B1(net_4080) );
DFF_X1 inst_6343 ( .QN(net_6188), .D(net_5842), .CK(net_13646) );
CLKBUF_X2 inst_13554 ( .A(net_12493), .Z(net_13516) );
CLKBUF_X2 inst_9014 ( .A(net_8975), .Z(net_8976) );
INV_X4 inst_4604 ( .ZN(net_4240), .A(net_4098) );
SDFF_X2 inst_161 ( .Q(net_6253), .SI(net_6252), .D(net_3477), .SE(net_392), .CK(net_13535) );
INV_X4 inst_4688 ( .ZN(net_3735), .A(net_3363) );
CLKBUF_X2 inst_12658 ( .A(net_12241), .Z(net_12620) );
CLKBUF_X2 inst_10956 ( .A(net_10917), .Z(net_10918) );
INV_X4 inst_4798 ( .ZN(net_5104), .A(net_1259) );
NAND2_X2 inst_3849 ( .A1(net_6707), .A2(net_1497), .ZN(net_1487) );
INV_X2 inst_6118 ( .A(net_5936), .ZN(net_5934) );
CLKBUF_X2 inst_12205 ( .A(net_12166), .Z(net_12167) );
CLKBUF_X2 inst_11287 ( .A(net_11248), .Z(net_11249) );
SDFF_X2 inst_1029 ( .SI(net_6492), .Q(net_6492), .SE(net_3886), .D(net_3799), .CK(net_8847) );
CLKBUF_X2 inst_9624 ( .A(net_9585), .Z(net_9586) );
INV_X4 inst_5413 ( .A(net_7697), .ZN(net_713) );
CLKBUF_X2 inst_11764 ( .A(net_11725), .Z(net_11726) );
CLKBUF_X2 inst_9246 ( .A(net_8214), .Z(net_9208) );
DFF_X1 inst_6666 ( .QN(net_7260), .D(net_5166), .CK(net_13008) );
DFF_X1 inst_6841 ( .D(net_2516), .QN(net_172), .CK(net_9863) );
NOR2_X2 inst_2408 ( .ZN(net_3731), .A2(net_3336), .A1(net_2960) );
CLKBUF_X2 inst_10519 ( .A(net_10480), .Z(net_10481) );
CLKBUF_X2 inst_9778 ( .A(net_9739), .Z(net_9740) );
SDFF_X2 inst_1324 ( .D(net_6383), .SE(net_5801), .SI(net_328), .Q(net_328), .CK(net_13854) );
DFF_X2 inst_6245 ( .QN(net_7682), .D(net_3030), .CK(net_8315) );
DFFR_X2 inst_7032 ( .QN(net_5986), .D(net_3192), .CK(net_9613), .RN(x1822) );
DFF_X1 inst_6551 ( .Q(net_7776), .D(net_5606), .CK(net_9987) );
CLKBUF_X2 inst_11848 ( .A(net_8598), .Z(net_11810) );
CLKBUF_X2 inst_10646 ( .A(net_10607), .Z(net_10608) );
SDFF_X2 inst_342 ( .SI(net_7367), .Q(net_7367), .D(net_4874), .SE(net_3853), .CK(net_9849) );
CLKBUF_X2 inst_13048 ( .A(net_8025), .Z(net_13010) );
INV_X2 inst_5767 ( .ZN(net_3019), .A(net_3018) );
CLKBUF_X2 inst_10067 ( .A(net_10028), .Z(net_10029) );
DFF_X1 inst_6443 ( .QN(net_6094), .D(net_5727), .CK(net_9226) );
CLKBUF_X2 inst_14404 ( .A(net_14365), .Z(net_14366) );
SDFF_X2 inst_463 ( .Q(net_7156), .D(net_7156), .SE(net_3903), .SI(net_3902), .CK(net_8735) );
OAI22_X2 inst_1534 ( .B1(net_4637), .B2(net_4033), .A1(net_4030), .ZN(net_4027), .A2(net_4026) );
CLKBUF_X2 inst_10667 ( .A(net_10628), .Z(net_10629) );
CLKBUF_X2 inst_9985 ( .A(net_9946), .Z(net_9947) );
CLKBUF_X2 inst_13571 ( .A(net_13532), .Z(net_13533) );
NAND2_X2 inst_3820 ( .A1(net_6627), .A2(net_1624), .ZN(net_1525) );
INV_X4 inst_4667 ( .A(net_4008), .ZN(net_3733) );
CLKBUF_X2 inst_9108 ( .A(net_9069), .Z(net_9070) );
SDFF_X2 inst_319 ( .SI(net_7463), .Q(net_7463), .D(net_5097), .SE(net_3993), .CK(net_9702) );
NOR2_X2 inst_2422 ( .A2(net_5914), .ZN(net_3228), .A1(net_3227) );
CLKBUF_X2 inst_12762 ( .A(net_12723), .Z(net_12724) );
DFFR_X2 inst_6992 ( .QN(net_7701), .D(net_3362), .CK(net_10369), .RN(x1822) );
CLKBUF_X2 inst_12745 ( .A(net_8883), .Z(net_12707) );
CLKBUF_X2 inst_10688 ( .A(net_10649), .Z(net_10650) );
INV_X2 inst_5923 ( .A(net_7652), .ZN(net_1978) );
SDFF_X2 inst_649 ( .Q(net_6705), .D(net_6705), .SE(net_3871), .SI(net_3813), .CK(net_8301) );
OAI21_X2 inst_2158 ( .A(net_2419), .ZN(net_1684), .B1(net_1683), .B2(net_1682) );
INV_X2 inst_5790 ( .A(net_5981), .ZN(net_2238) );
INV_X4 inst_5560 ( .A(net_7426), .ZN(net_2144) );
OAI21_X2 inst_1711 ( .B2(net_5913), .ZN(net_5583), .A(net_5128), .B1(net_4030) );
CLKBUF_X2 inst_10660 ( .A(net_8945), .Z(net_10622) );
CLKBUF_X2 inst_8504 ( .A(net_8465), .Z(net_8466) );
NAND2_X2 inst_3426 ( .A2(net_5892), .ZN(net_3233), .A1(net_3232) );
NAND3_X2 inst_2597 ( .ZN(net_5742), .A1(net_5637), .A2(net_5216), .A3(net_4202) );
CLKBUF_X2 inst_14269 ( .A(net_14230), .Z(net_14231) );
CLKBUF_X2 inst_12227 ( .A(net_11897), .Z(net_12189) );
INV_X4 inst_5185 ( .ZN(net_518), .A(net_517) );
INV_X4 inst_5569 ( .A(net_7269), .ZN(net_2043) );
OAI21_X2 inst_2052 ( .B2(net_4457), .ZN(net_4448), .B1(net_4447), .A(net_3561) );
SDFF_X2 inst_995 ( .Q(net_6483), .D(net_6483), .SE(net_3904), .SI(net_3789), .CK(net_8409) );
OAI22_X2 inst_1575 ( .A2(net_3297), .B2(net_3286), .ZN(net_3271), .A1(net_3270), .B1(net_584) );
INV_X2 inst_6059 ( .A(net_7621), .ZN(net_1184) );
CLKBUF_X2 inst_9644 ( .A(net_7844), .Z(net_9606) );
CLKBUF_X2 inst_8850 ( .A(net_8175), .Z(net_8812) );
AOI21_X2 inst_7726 ( .B1(net_6727), .ZN(net_4506), .B2(net_2581), .A(net_2338) );
CLKBUF_X2 inst_13948 ( .A(net_11901), .Z(net_13910) );
CLKBUF_X2 inst_10697 ( .A(net_10658), .Z(net_10659) );
NOR2_X2 inst_2470 ( .A2(net_5778), .ZN(net_2684), .A1(net_2612) );
INV_X2 inst_6049 ( .A(net_7620), .ZN(net_1191) );
INV_X4 inst_5522 ( .A(net_7562), .ZN(net_1906) );
SDFF_X2 inst_1258 ( .SI(net_6527), .Q(net_6527), .D(net_3890), .SE(net_3756), .CK(net_8751) );
CLKBUF_X2 inst_10148 ( .A(net_10109), .Z(net_10110) );
NAND2_X2 inst_3141 ( .ZN(net_4822), .A2(net_4153), .A1(net_2150) );
NAND2_X2 inst_3921 ( .A2(net_1696), .ZN(net_1382), .A1(net_1381) );
OAI21_X2 inst_1957 ( .B1(net_5204), .ZN(net_5063), .A(net_4708), .B2(net_3986) );
NAND2_X2 inst_3857 ( .A2(net_1696), .ZN(net_1477), .A1(net_1476) );
INV_X4 inst_5151 ( .ZN(net_781), .A(net_565) );
CLKBUF_X2 inst_13860 ( .A(net_13821), .Z(net_13822) );
CLKBUF_X2 inst_9524 ( .A(net_9485), .Z(net_9486) );
SDFF_X2 inst_1060 ( .Q(net_6701), .D(net_6701), .SI(net_3883), .SE(net_3871), .CK(net_11708) );
INV_X2 inst_5920 ( .A(net_7356), .ZN(net_2066) );
AOI22_X2 inst_7446 ( .B2(net_2757), .A2(net_2658), .ZN(net_854), .A1(net_853), .B1(net_438) );
CLKBUF_X2 inst_10456 ( .A(net_10417), .Z(net_10418) );
SDFF_X2 inst_900 ( .Q(net_7103), .D(net_7103), .SE(net_3888), .SI(net_3799), .CK(net_10494) );
DFFS_X2 inst_6950 ( .QN(net_6405), .D(net_2713), .CK(net_14409), .SN(x1822) );
CLKBUF_X2 inst_10568 ( .A(net_9217), .Z(net_10530) );
INV_X4 inst_4949 ( .ZN(net_5869), .A(net_736) );
CLKBUF_X2 inst_13813 ( .A(net_13774), .Z(net_13775) );
CLKBUF_X2 inst_12677 ( .A(net_12638), .Z(net_12639) );
INV_X4 inst_4624 ( .ZN(net_4198), .A(net_4058) );
NAND3_X2 inst_2807 ( .ZN(net_2291), .A3(net_1592), .A1(net_1299), .A2(net_1026) );
CLKBUF_X2 inst_12458 ( .A(net_12419), .Z(net_12420) );
AND2_X4 inst_7811 ( .ZN(net_3838), .A2(net_3837), .A1(net_1145) );
CLKBUF_X2 inst_11257 ( .A(net_11218), .Z(net_11219) );
CLKBUF_X2 inst_13608 ( .A(net_13569), .Z(net_13570) );
CLKBUF_X2 inst_9254 ( .A(net_8108), .Z(net_9216) );
INV_X2 inst_6062 ( .ZN(net_1127), .A(net_115) );
AOI22_X2 inst_7428 ( .A1(net_2970), .B1(net_2772), .ZN(net_2764), .A2(net_244), .B2(net_170) );
NAND2_X2 inst_2983 ( .A1(net_6751), .A2(net_5033), .ZN(net_5028) );
INV_X4 inst_5327 ( .A(net_7380), .ZN(net_1201) );
DFF_X1 inst_6608 ( .QN(net_7515), .D(net_5400), .CK(net_12082) );
AOI21_X2 inst_7778 ( .B1(net_6604), .ZN(net_4024), .B2(net_2583), .A(net_2359) );
INV_X4 inst_5423 ( .A(net_5991), .ZN(net_493) );
CLKBUF_X2 inst_9995 ( .A(net_9956), .Z(net_9957) );
CLKBUF_X2 inst_8803 ( .A(net_8764), .Z(net_8765) );
CLKBUF_X2 inst_8651 ( .A(net_8612), .Z(net_8613) );
AOI22_X2 inst_7421 ( .A1(net_2970), .B1(net_2772), .ZN(net_2771), .A2(net_239), .B2(net_165) );
CLKBUF_X2 inst_13584 ( .A(net_8221), .Z(net_13546) );
CLKBUF_X2 inst_13233 ( .A(net_13194), .Z(net_13195) );
CLKBUF_X2 inst_9969 ( .A(net_9183), .Z(net_9931) );
CLKBUF_X2 inst_8862 ( .A(net_8823), .Z(net_8824) );
CLKBUF_X2 inst_12881 ( .A(net_12842), .Z(net_12843) );
CLKBUF_X2 inst_10470 ( .A(net_10310), .Z(net_10432) );
SDFF_X2 inst_1120 ( .D(net_7807), .SI(net_6669), .Q(net_6669), .SE(net_3465), .CK(net_9316) );
CLKBUF_X2 inst_12986 ( .A(net_11883), .Z(net_12948) );
DFF_X2 inst_6238 ( .QN(net_7530), .D(net_3036), .CK(net_12597) );
CLKBUF_X2 inst_8545 ( .A(net_8506), .Z(net_8507) );
CLKBUF_X2 inst_7882 ( .A(net_7843), .Z(net_7844) );
CLKBUF_X2 inst_11617 ( .A(net_11578), .Z(net_11579) );
CLKBUF_X2 inst_12161 ( .A(net_12122), .Z(net_12123) );
NAND2_X2 inst_3184 ( .ZN(net_4749), .A2(net_3941), .A1(net_2009) );
DFF_X1 inst_6767 ( .QN(net_6106), .D(net_4669), .CK(net_11125) );
CLKBUF_X2 inst_9715 ( .A(net_9676), .Z(net_9677) );
DFF_X1 inst_6398 ( .QN(net_6137), .D(net_5690), .CK(net_8177) );
CLKBUF_X2 inst_8084 ( .A(net_8045), .Z(net_8046) );
SDFF_X2 inst_731 ( .Q(net_6848), .D(net_6848), .SE(net_3893), .SI(net_3807), .CK(net_11751) );
SDFF_X2 inst_947 ( .SI(net_7190), .Q(net_7190), .SE(net_3817), .D(net_3794), .CK(net_10634) );
SDFF_X2 inst_1225 ( .SI(net_7218), .Q(net_7218), .D(net_3803), .SE(net_3751), .CK(net_8688) );
CLKBUF_X2 inst_10909 ( .A(net_8987), .Z(net_10871) );
CLKBUF_X2 inst_13788 ( .A(net_8886), .Z(net_13750) );
AOI222_X2 inst_7535 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1896), .A1(net_1895), .B1(net_1894), .C1(net_1893) );
CLKBUF_X2 inst_12411 ( .A(net_10095), .Z(net_12373) );
NOR2_X2 inst_2459 ( .ZN(net_2991), .A1(net_2804), .A2(net_190) );
CLKBUF_X2 inst_14256 ( .A(net_14217), .Z(net_14218) );
SDFF_X2 inst_363 ( .SI(net_7612), .Q(net_7612), .D(net_4786), .SE(net_3870), .CK(net_7997) );
SDFF_X2 inst_301 ( .SI(net_7519), .Q(net_7519), .D(net_5105), .SE(net_3988), .CK(net_9798) );
INV_X4 inst_5316 ( .A(net_7582), .ZN(net_1875) );
OAI21_X2 inst_2141 ( .B1(net_5778), .ZN(net_2803), .A(net_2686), .B2(net_2684) );
INV_X4 inst_5530 ( .ZN(net_556), .A(net_287) );
CLKBUF_X2 inst_14427 ( .A(net_12801), .Z(net_14389) );
CLKBUF_X2 inst_14215 ( .A(net_14176), .Z(net_14177) );
CLKBUF_X2 inst_12041 ( .A(net_12002), .Z(net_12003) );
INV_X8 inst_4551 ( .ZN(net_2211), .A(net_808) );
CLKBUF_X2 inst_11397 ( .A(net_11358), .Z(net_11359) );
NAND2_X1 inst_4313 ( .ZN(net_4553), .A2(net_3866), .A1(net_1840) );
DFF_X1 inst_6609 ( .QN(net_7516), .D(net_5398), .CK(net_9650) );
CLKBUF_X2 inst_13213 ( .A(net_13174), .Z(net_13175) );
DFFR_X2 inst_7079 ( .QN(net_7726), .D(net_2794), .CK(net_12556), .RN(x1822) );
CLKBUF_X2 inst_13153 ( .A(net_13114), .Z(net_13115) );
INV_X4 inst_4714 ( .ZN(net_3122), .A(net_3047) );
CLKBUF_X2 inst_7870 ( .A(net_7830), .Z(net_7832) );
CLKBUF_X2 inst_14021 ( .A(net_13457), .Z(net_13983) );
CLKBUF_X2 inst_12898 ( .A(net_12859), .Z(net_12860) );
NAND2_X1 inst_4348 ( .ZN(net_4379), .A2(net_3856), .A1(net_1768) );
INV_X4 inst_4706 ( .ZN(net_3240), .A(net_2974) );
NAND2_X2 inst_2956 ( .ZN(net_5484), .A1(net_4938), .A2(net_4937) );
INV_X4 inst_4713 ( .ZN(net_3121), .A(net_3045) );
CLKBUF_X2 inst_14312 ( .A(net_14273), .Z(net_14274) );
NAND2_X2 inst_3729 ( .A1(net_6894), .A2(net_1639), .ZN(net_1616) );
CLKBUF_X2 inst_8521 ( .A(net_8482), .Z(net_8483) );
SDFF_X2 inst_412 ( .SI(net_7377), .Q(net_7377), .D(net_4776), .SE(net_3853), .CK(net_12746) );
CLKBUF_X2 inst_10430 ( .A(net_8011), .Z(net_10392) );
AOI222_X2 inst_7548 ( .C1(net_7679), .A1(net_7647), .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1859), .B1(net_1858) );
CLKBUF_X2 inst_9282 ( .A(net_9243), .Z(net_9244) );
CLKBUF_X2 inst_8345 ( .A(net_8306), .Z(net_8307) );
CLKBUF_X2 inst_11687 ( .A(net_11648), .Z(net_11649) );
NAND3_X2 inst_2650 ( .ZN(net_3986), .A1(net_3985), .A3(net_3869), .A2(net_1728) );
INV_X4 inst_5463 ( .ZN(net_586), .A(net_294) );
INV_X8 inst_4508 ( .ZN(net_3886), .A(net_3257) );
CLKBUF_X2 inst_7943 ( .A(net_7864), .Z(net_7905) );
CLKBUF_X2 inst_13022 ( .A(net_12983), .Z(net_12984) );
CLKBUF_X2 inst_11626 ( .A(net_9728), .Z(net_11588) );
CLKBUF_X2 inst_9490 ( .A(net_9451), .Z(net_9452) );
CLKBUF_X2 inst_11666 ( .A(net_11627), .Z(net_11628) );
CLKBUF_X2 inst_8295 ( .A(net_8216), .Z(net_8257) );
CLKBUF_X2 inst_13969 ( .A(net_10412), .Z(net_13931) );
NAND2_X2 inst_3189 ( .ZN(net_4744), .A2(net_3941), .A1(net_2001) );
NAND2_X2 inst_3163 ( .ZN(net_4770), .A2(net_3941), .A1(net_2025) );
NOR2_X2 inst_2504 ( .ZN(net_1241), .A1(net_1240), .A2(net_621) );
CLKBUF_X2 inst_8918 ( .A(net_8879), .Z(net_8880) );
CLKBUF_X2 inst_13511 ( .A(net_13472), .Z(net_13473) );
CLKBUF_X2 inst_12818 ( .A(net_11435), .Z(net_12780) );
INV_X4 inst_5548 ( .A(net_7421), .ZN(net_2081) );
INV_X2 inst_5985 ( .ZN(net_404), .A(x1062) );
DFF_X1 inst_6855 ( .D(net_2534), .Q(net_219), .CK(net_9534) );
CLKBUF_X2 inst_14076 ( .A(net_14037), .Z(net_14038) );
CLKBUF_X2 inst_14188 ( .A(net_8658), .Z(net_14150) );
CLKBUF_X2 inst_10902 ( .A(net_10863), .Z(net_10864) );
SDFF_X2 inst_684 ( .Q(net_6749), .D(net_6749), .SE(net_3815), .SI(net_3803), .CK(net_8376) );
DFF_X2 inst_6263 ( .QN(net_5983), .D(net_2728), .CK(net_10510) );
NAND2_X2 inst_3374 ( .ZN(net_3498), .A1(net_3497), .A2(net_3223) );
NAND2_X1 inst_4354 ( .ZN(net_4373), .A2(net_3853), .A1(net_2066) );
NAND2_X1 inst_4400 ( .A2(net_3297), .ZN(net_3079), .A1(net_2927) );
NAND2_X2 inst_3438 ( .ZN(net_3210), .A2(net_3091), .A1(net_2759) );
NAND2_X2 inst_3177 ( .ZN(net_4756), .A2(net_3941), .A1(net_2035) );
CLKBUF_X2 inst_12187 ( .A(net_12148), .Z(net_12149) );
CLKBUF_X2 inst_12541 ( .A(net_10685), .Z(net_12503) );
CLKBUF_X2 inst_10437 ( .A(net_8135), .Z(net_10399) );
INV_X4 inst_4930 ( .ZN(net_2244), .A(net_775) );
CLKBUF_X2 inst_7965 ( .A(net_7919), .Z(net_7927) );
NAND2_X2 inst_3811 ( .A1(net_7176), .A2(net_1637), .ZN(net_1534) );
CLKBUF_X2 inst_11857 ( .A(net_11818), .Z(net_11819) );
NAND2_X2 inst_3653 ( .A1(net_7061), .ZN(net_1810), .A2(net_791) );
DFFR_X2 inst_6959 ( .QN(net_7725), .D(net_5776), .CK(net_12882), .RN(x1822) );
CLKBUF_X2 inst_8213 ( .A(net_8174), .Z(net_8175) );
CLKBUF_X2 inst_10700 ( .A(net_10661), .Z(net_10662) );
SDFF_X2 inst_1138 ( .SI(net_6662), .Q(net_6662), .D(net_3890), .SE(net_3471), .CK(net_7836) );
SDFF_X2 inst_1241 ( .SI(net_6535), .Q(net_6535), .D(net_3787), .SE(net_3755), .CK(net_8832) );
SDFF_X2 inst_1038 ( .Q(net_7541), .D(net_7541), .SE(net_3896), .SI(net_375), .CK(net_10262) );
DFF_X1 inst_6568 ( .QN(net_7504), .D(net_5096), .CK(net_10075) );
SDFF_X2 inst_940 ( .SI(net_7164), .Q(net_7164), .SE(net_3817), .D(net_3806), .CK(net_7904) );
SDFF_X2 inst_1004 ( .Q(net_6464), .D(net_6464), .SE(net_3904), .SI(net_3814), .CK(net_11651) );
CLKBUF_X2 inst_9417 ( .A(net_9378), .Z(net_9379) );
CLKBUF_X2 inst_11705 ( .A(net_11666), .Z(net_11667) );
CLKBUF_X2 inst_11641 ( .A(net_11602), .Z(net_11603) );
NAND2_X2 inst_3595 ( .ZN(net_2405), .A2(net_1878), .A1(net_1420) );
CLKBUF_X2 inst_11830 ( .A(net_11791), .Z(net_11792) );
CLKBUF_X2 inst_9316 ( .A(net_9277), .Z(net_9278) );
SDFF_X2 inst_189 ( .Q(net_6265), .SI(net_6264), .D(net_3483), .SE(net_392), .CK(net_13471) );
INV_X4 inst_4876 ( .ZN(net_3855), .A(net_617) );
CLKBUF_X2 inst_8103 ( .A(net_8064), .Z(net_8065) );
AOI21_X2 inst_7732 ( .B1(net_6879), .ZN(net_4089), .B2(net_2579), .A(net_2285) );
CLKBUF_X2 inst_9008 ( .A(net_8969), .Z(net_8970) );
NOR2_X2 inst_2450 ( .ZN(net_2859), .A1(net_2858), .A2(net_2857) );
CLKBUF_X2 inst_13248 ( .A(net_12340), .Z(net_13210) );
CLKBUF_X2 inst_8597 ( .A(net_8558), .Z(net_8559) );
NAND2_X1 inst_4362 ( .ZN(net_4365), .A2(net_3853), .A1(net_2042) );
AOI22_X2 inst_7437 ( .B1(net_7007), .A1(net_6975), .ZN(net_1834), .A2(net_1833), .B2(net_1100) );
CLKBUF_X2 inst_9581 ( .A(net_9542), .Z(net_9543) );
AOI22_X2 inst_7430 ( .A1(net_2970), .B1(net_2772), .ZN(net_2762), .A2(net_232), .B2(net_158) );
CLKBUF_X2 inst_11006 ( .A(net_10967), .Z(net_10968) );
CLKBUF_X2 inst_9529 ( .A(net_9490), .Z(net_9491) );
XNOR2_X2 inst_62 ( .ZN(net_1731), .B(net_1730), .A(net_1084) );
CLKBUF_X2 inst_12608 ( .A(net_12569), .Z(net_12570) );
NAND2_X1 inst_4369 ( .ZN(net_4358), .A2(net_3856), .A1(net_1770) );
INV_X4 inst_4696 ( .A(net_5964), .ZN(net_3367) );
NAND2_X2 inst_3743 ( .A1(net_6895), .A2(net_1639), .ZN(net_1602) );
NAND2_X4 inst_2860 ( .A1(net_5879), .ZN(net_5049), .A2(net_4142) );
CLKBUF_X2 inst_11899 ( .A(net_9839), .Z(net_11861) );
INV_X4 inst_5194 ( .ZN(net_509), .A(net_508) );
CLKBUF_X2 inst_11236 ( .A(net_11197), .Z(net_11198) );
CLKBUF_X2 inst_13076 ( .A(net_13037), .Z(net_13038) );
CLKBUF_X2 inst_8387 ( .A(net_8348), .Z(net_8349) );
NAND2_X2 inst_4007 ( .A2(net_2232), .ZN(net_1916), .A1(net_1823) );
SDFF_X2 inst_879 ( .Q(net_7099), .D(net_7099), .SE(net_3888), .SI(net_3792), .CK(net_10501) );
CLKBUF_X2 inst_11266 ( .A(net_8248), .Z(net_11228) );
INV_X2 inst_5888 ( .A(net_7448), .ZN(net_1463) );
CLKBUF_X2 inst_13956 ( .A(net_13917), .Z(net_13918) );
CLKBUF_X2 inst_11162 ( .A(net_11123), .Z(net_11124) );
CLKBUF_X2 inst_12416 ( .A(net_12377), .Z(net_12378) );
AOI22_X2 inst_7344 ( .ZN(net_3108), .B2(net_3105), .A2(net_2712), .A1(net_1261), .B1(net_493) );
CLKBUF_X2 inst_8252 ( .A(net_8213), .Z(net_8214) );
INV_X8 inst_4482 ( .ZN(net_4280), .A(net_3926) );
NAND2_X1 inst_4291 ( .ZN(net_4576), .A2(net_3867), .A1(net_1195) );
INV_X4 inst_5692 ( .A(net_6066), .ZN(net_3534) );
SDFF_X2 inst_629 ( .SI(net_6640), .Q(net_6640), .SE(net_3850), .D(net_3776), .CK(net_12163) );
INV_X4 inst_4903 ( .ZN(net_2256), .A(net_866) );
SDFF_X2 inst_1100 ( .SI(net_6817), .Q(net_6817), .D(net_3789), .SE(net_3722), .CK(net_11309) );
CLKBUF_X2 inst_7903 ( .A(net_7852), .Z(net_7865) );
CLKBUF_X2 inst_10872 ( .A(net_10833), .Z(net_10834) );
SDFF_X2 inst_791 ( .SI(net_6921), .Q(net_6921), .SE(net_3887), .D(net_3788), .CK(net_11456) );
CLKBUF_X2 inst_13371 ( .A(net_9087), .Z(net_13333) );
CLKBUF_X2 inst_10427 ( .A(net_10388), .Z(net_10389) );
OAI21_X2 inst_2021 ( .B2(net_4497), .ZN(net_4486), .B1(net_4485), .A(net_3636) );
CLKBUF_X2 inst_9631 ( .A(net_8753), .Z(net_9593) );
NAND2_X2 inst_3383 ( .ZN(net_3480), .A1(net_3479), .A2(net_3223) );
NAND2_X1 inst_4379 ( .ZN(net_4348), .A2(net_3859), .A1(net_2061) );
SDFF_X2 inst_1191 ( .SI(net_7072), .Q(net_7072), .D(net_3812), .SE(net_3742), .CK(net_8994) );
INV_X4 inst_5668 ( .A(net_7418), .ZN(net_2220) );
CLKBUF_X2 inst_13326 ( .A(net_9456), .Z(net_13288) );
SDFF_X2 inst_533 ( .Q(net_6601), .D(net_6601), .SI(net_3894), .SE(net_3830), .CK(net_9195) );
INV_X4 inst_5086 ( .A(net_7812), .ZN(net_3784) );
CLKBUF_X2 inst_12811 ( .A(net_12765), .Z(net_12773) );
NOR2_X2 inst_2478 ( .A2(net_5778), .ZN(net_2602), .A1(net_556) );
INV_X4 inst_4972 ( .A(net_3808), .ZN(net_3170) );
NAND3_X2 inst_2751 ( .ZN(net_2350), .A3(net_1532), .A1(net_1325), .A2(net_1005) );
CLKBUF_X2 inst_14399 ( .A(net_14360), .Z(net_14361) );
CLKBUF_X2 inst_8576 ( .A(net_8537), .Z(net_8538) );
CLKBUF_X2 inst_13020 ( .A(net_12981), .Z(net_12982) );
CLKBUF_X2 inst_11924 ( .A(net_11885), .Z(net_11886) );
OAI21_X2 inst_1760 ( .ZN(net_5437), .B1(net_5436), .A(net_4659), .B2(net_3993) );
OAI21_X2 inst_1874 ( .ZN(net_5231), .B1(net_5230), .A(net_4588), .B2(net_3867) );
CLKBUF_X2 inst_11888 ( .A(net_11849), .Z(net_11850) );
OAI21_X2 inst_2022 ( .B1(net_5896), .B2(net_4497), .ZN(net_4484), .A(net_3634) );
NAND2_X2 inst_3960 ( .A1(net_6568), .A2(net_1705), .ZN(net_1324) );
NAND3_X2 inst_2821 ( .A2(net_3855), .ZN(net_1831), .A3(net_1830), .A1(net_616) );
SDFF_X2 inst_1095 ( .SI(net_6936), .Q(net_6936), .D(net_3813), .SE(net_3734), .CK(net_8627) );
CLKBUF_X2 inst_8042 ( .A(net_8003), .Z(net_8004) );
CLKBUF_X2 inst_10516 ( .A(net_10266), .Z(net_10478) );
CLKBUF_X2 inst_10096 ( .A(net_10057), .Z(net_10058) );
CLKBUF_X2 inst_9052 ( .A(net_9013), .Z(net_9014) );
NOR2_X2 inst_2439 ( .ZN(net_3422), .A1(net_3042), .A2(net_3041) );
SDFF_X2 inst_176 ( .Q(net_6278), .SI(net_6277), .D(net_3499), .SE(net_392), .CK(net_13490) );
NAND3_X2 inst_2826 ( .ZN(net_1669), .A3(net_1668), .A1(net_1665), .A2(net_1068) );
AND2_X4 inst_7848 ( .ZN(net_1971), .A2(net_781), .A1(net_634) );
INV_X16 inst_6143 ( .ZN(net_1642), .A(net_774) );
CLKBUF_X2 inst_8142 ( .A(net_7924), .Z(net_8104) );
AOI22_X2 inst_7304 ( .B1(net_6677), .A1(net_6645), .ZN(net_5141), .A2(net_5139), .B2(net_5138) );
CLKBUF_X2 inst_9069 ( .A(net_9030), .Z(net_9031) );
CLKBUF_X2 inst_10894 ( .A(net_10855), .Z(net_10856) );
CLKBUF_X2 inst_12864 ( .A(net_12825), .Z(net_12826) );
SDFFR_X2 inst_1336 ( .SE(net_3895), .SI(net_113), .CK(net_10201), .RN(x1822), .Q(x0), .D(x0) );
INV_X4 inst_5472 ( .A(net_7403), .ZN(net_2071) );
CLKBUF_X2 inst_10387 ( .A(net_8986), .Z(net_10349) );
NAND2_X1 inst_4404 ( .A2(net_3087), .ZN(net_2914), .A1(net_2830) );
CLKBUF_X2 inst_8937 ( .A(net_8898), .Z(net_8899) );
OAI221_X2 inst_1665 ( .C2(net_5899), .ZN(net_4651), .B1(net_4650), .B2(net_4445), .C1(net_4080), .A(net_3563) );
INV_X8 inst_4500 ( .ZN(net_3818), .A(net_3263) );
CLKBUF_X2 inst_13962 ( .A(net_13669), .Z(net_13924) );
INV_X4 inst_4763 ( .ZN(net_2786), .A(net_2772) );
SDFF_X2 inst_780 ( .SI(net_6908), .Q(net_6908), .SE(net_3887), .D(net_3810), .CK(net_8868) );
INV_X4 inst_5626 ( .A(net_6174), .ZN(net_3568) );
CLKBUF_X2 inst_9054 ( .A(net_9015), .Z(net_9016) );
DFF_X1 inst_6581 ( .QN(net_7569), .D(net_5070), .CK(net_13287) );
CLKBUF_X2 inst_8154 ( .A(net_8115), .Z(net_8116) );
DFF_X1 inst_6783 ( .QN(net_6085), .D(net_4317), .CK(net_12941) );
CLKBUF_X2 inst_8255 ( .A(net_8216), .Z(net_8217) );
CLKBUF_X2 inst_11261 ( .A(net_10358), .Z(net_11223) );
CLKBUF_X2 inst_12016 ( .A(net_11977), .Z(net_11978) );
DFF_X1 inst_6716 ( .QN(net_7317), .D(net_5348), .CK(net_9443) );
NAND2_X2 inst_3967 ( .A1(net_6563), .A2(net_1705), .ZN(net_1313) );
INV_X4 inst_5541 ( .A(net_7716), .ZN(net_858) );
CLKBUF_X2 inst_8722 ( .A(net_8186), .Z(net_8684) );
NAND2_X2 inst_4018 ( .A1(net_6926), .A2(net_1654), .ZN(net_1034) );
NAND2_X2 inst_3669 ( .A1(net_7342), .A2(net_1798), .ZN(net_1790) );
OAI21_X2 inst_1767 ( .B1(net_5542), .ZN(net_5427), .A(net_4642), .B2(net_3993) );
INV_X4 inst_5636 ( .A(net_7747), .ZN(net_2667) );
NOR2_X4 inst_2219 ( .ZN(net_5679), .A1(net_5557), .A2(net_4516) );
CLKBUF_X2 inst_8884 ( .A(net_8845), .Z(net_8846) );
CLKBUF_X2 inst_8331 ( .A(net_8292), .Z(net_8293) );
SDFF_X2 inst_546 ( .Q(net_6459), .D(net_6459), .SE(net_3904), .SI(net_3892), .CK(net_8789) );
SDFF_X2 inst_1284 ( .D(net_3810), .SE(net_3256), .SI(net_145), .Q(net_145), .CK(net_10688) );
CLKBUF_X2 inst_13564 ( .A(net_13525), .Z(net_13526) );
NOR2_X2 inst_2465 ( .A2(net_2733), .ZN(net_2732), .A1(net_2727) );
NOR2_X2 inst_2361 ( .ZN(net_5303), .A2(net_4632), .A1(net_4504) );
SDFF_X2 inst_704 ( .SI(net_6775), .Q(net_6775), .SE(net_3872), .D(net_3808), .CK(net_8507) );
CLKBUF_X2 inst_11497 ( .A(net_11458), .Z(net_11459) );
CLKBUF_X2 inst_10237 ( .A(net_10198), .Z(net_10199) );
CLKBUF_X2 inst_9301 ( .A(net_9262), .Z(net_9263) );
INV_X2 inst_6006 ( .A(net_7465), .ZN(net_2173) );
INV_X8 inst_4542 ( .ZN(net_2583), .A(net_1280) );
INV_X4 inst_5558 ( .A(net_6554), .ZN(net_581) );
DFFR_X2 inst_7084 ( .QN(net_7745), .D(net_2798), .CK(net_9601), .RN(x1822) );
DFF_X1 inst_6802 ( .D(net_3936), .CK(net_12544), .Q(x638) );
CLKBUF_X2 inst_8285 ( .A(net_8140), .Z(net_8247) );
NOR2_X4 inst_2226 ( .ZN(net_5672), .A1(net_5536), .A2(net_4503) );
INV_X4 inst_5467 ( .A(net_6693), .ZN(net_2565) );
SDFF_X2 inst_694 ( .Q(net_6731), .D(net_6731), .SE(net_3815), .SI(net_3798), .CK(net_8282) );
INV_X4 inst_5574 ( .A(net_7686), .ZN(net_820) );
DFF_X1 inst_6382 ( .QN(net_6280), .D(net_5802), .CK(net_13635) );
NOR2_X2 inst_2498 ( .A1(net_3050), .ZN(net_1742), .A2(net_1741) );
CLKBUF_X2 inst_12402 ( .A(net_9879), .Z(net_12364) );
NAND2_X2 inst_3154 ( .ZN(net_4809), .A2(net_4153), .A1(net_2107) );
DFFR_X2 inst_6986 ( .QN(net_6005), .D(net_3447), .CK(net_10029), .RN(x1822) );
CLKBUF_X2 inst_11476 ( .A(net_11437), .Z(net_11438) );
CLKBUF_X2 inst_11523 ( .A(net_11484), .Z(net_11485) );
CLKBUF_X2 inst_8983 ( .A(net_8944), .Z(net_8945) );
INV_X4 inst_5396 ( .A(net_7576), .ZN(net_1889) );
CLKBUF_X2 inst_13885 ( .A(net_8577), .Z(net_13847) );
CLKBUF_X2 inst_11467 ( .A(net_11428), .Z(net_11429) );
INV_X4 inst_5211 ( .ZN(net_615), .A(net_486) );
CLKBUF_X2 inst_9394 ( .A(net_9124), .Z(net_9356) );
NAND2_X2 inst_2971 ( .ZN(net_5456), .A1(net_4878), .A2(net_4877) );
SDFFR_X2 inst_1342 ( .Q(net_7709), .D(net_7709), .SI(net_3897), .SE(net_3405), .CK(net_10713), .RN(x1822) );
AND2_X4 inst_7814 ( .ZN(net_3896), .A2(net_3258), .A1(net_685) );
CLKBUF_X2 inst_12071 ( .A(net_12032), .Z(net_12033) );
SDFF_X2 inst_787 ( .SI(net_6916), .Q(net_6916), .SE(net_3887), .D(net_3780), .CK(net_11718) );
NAND2_X1 inst_4396 ( .A2(net_5890), .ZN(net_3239), .A1(net_3238) );
CLKBUF_X2 inst_11211 ( .A(net_11172), .Z(net_11173) );
INV_X8 inst_4549 ( .ZN(net_2135), .A(net_798) );
CLKBUF_X2 inst_12958 ( .A(net_9370), .Z(net_12920) );
AOI222_X2 inst_7483 ( .A2(net_2135), .B2(net_2133), .C2(net_2131), .ZN(net_2130), .A1(net_2129), .B1(net_2128), .C1(net_2127) );
CLKBUF_X2 inst_14439 ( .A(net_10655), .Z(net_14401) );
CLKBUF_X2 inst_10551 ( .A(net_10512), .Z(net_10513) );
INV_X2 inst_6012 ( .ZN(net_402), .A(net_155) );
NAND2_X2 inst_3933 ( .A2(net_1696), .ZN(net_1362), .A1(net_1361) );
SDFF_X2 inst_825 ( .Q(net_6972), .D(net_6972), .SE(net_3891), .SI(net_3814), .CK(net_11955) );
NAND3_X2 inst_2586 ( .ZN(net_5753), .A1(net_5648), .A2(net_5266), .A3(net_4308) );
OAI221_X2 inst_1656 ( .ZN(net_4798), .A(net_4590), .C2(net_3975), .B2(net_3964), .C1(net_3767), .B1(net_1387) );
INV_X2 inst_5881 ( .A(net_7618), .ZN(net_1197) );
CLKBUF_X2 inst_7928 ( .A(net_7867), .Z(net_7890) );
OAI21_X2 inst_1881 ( .ZN(net_5205), .B1(net_5204), .A(net_4577), .B2(net_3867) );
CLKBUF_X2 inst_12886 ( .A(net_11850), .Z(net_12848) );
NAND2_X2 inst_3034 ( .A1(net_6989), .A2(net_4977), .ZN(net_4973) );
OAI21_X2 inst_1892 ( .B1(net_5225), .ZN(net_5189), .A(net_4565), .B2(net_3866) );
INV_X4 inst_5590 ( .A(net_7683), .ZN(net_499) );
AND2_X2 inst_7860 ( .ZN(net_2271), .A1(net_1699), .A2(net_1698) );
CLKBUF_X2 inst_11404 ( .A(net_9764), .Z(net_11366) );
SDFF_X2 inst_295 ( .D(net_6394), .SE(net_5800), .SI(net_359), .Q(net_359), .CK(net_14153) );
SDFF_X2 inst_726 ( .Q(net_6842), .D(net_6842), .SE(net_3893), .SI(net_3811), .CK(net_8887) );
CLKBUF_X2 inst_10583 ( .A(net_10544), .Z(net_10545) );
CLKBUF_X2 inst_13018 ( .A(net_8976), .Z(net_12980) );
CLKBUF_X2 inst_8971 ( .A(net_8141), .Z(net_8933) );
INV_X4 inst_4726 ( .A(net_5971), .ZN(net_3047) );
CLKBUF_X2 inst_8073 ( .A(net_8034), .Z(net_8035) );
SDFF_X2 inst_320 ( .SI(net_7464), .Q(net_7464), .D(net_5099), .SE(net_3993), .CK(net_9967) );
SDFF_X2 inst_607 ( .Q(net_6611), .D(net_6611), .SE(net_3830), .SI(net_3805), .CK(net_12167) );
DFF_X1 inst_6484 ( .QN(net_7415), .D(net_5568), .CK(net_9310) );
NOR2_X2 inst_2432 ( .ZN(net_3072), .A1(net_3071), .A2(net_3068) );
NAND2_X1 inst_4263 ( .ZN(net_4657), .A2(net_3993), .A1(net_1365) );
XOR2_X2 inst_1 ( .A(net_2575), .Z(net_1252), .B(net_1251) );
INV_X4 inst_5061 ( .A(net_7818), .ZN(net_3902) );
DFF_X1 inst_6693 ( .QN(net_7282), .D(net_5382), .CK(net_12717) );
CLKBUF_X2 inst_8273 ( .A(net_8234), .Z(net_8235) );
OAI21_X2 inst_1891 ( .B1(net_5227), .ZN(net_5190), .A(net_4566), .B2(net_3866) );
AOI221_X2 inst_7614 ( .C2(net_3105), .B1(net_2970), .ZN(net_2966), .C1(net_2965), .A(net_2788), .B2(net_246) );
CLKBUF_X2 inst_10130 ( .A(net_10091), .Z(net_10092) );
CLKBUF_X2 inst_8560 ( .A(net_8521), .Z(net_8522) );
NAND2_X1 inst_4343 ( .ZN(net_4384), .A2(net_3853), .A1(net_2215) );
CLKBUF_X2 inst_12794 ( .A(net_12224), .Z(net_12756) );
INV_X4 inst_5684 ( .A(net_6056), .ZN(net_802) );
CLKBUF_X2 inst_11537 ( .A(net_11498), .Z(net_11499) );
INV_X8 inst_4558 ( .ZN(net_2202), .A(net_690) );
DFF_X1 inst_6627 ( .QN(net_7597), .D(net_5260), .CK(net_13078) );
CLKBUF_X2 inst_11841 ( .A(net_11802), .Z(net_11803) );
CLKBUF_X2 inst_11493 ( .A(net_11454), .Z(net_11455) );
SDFF_X2 inst_235 ( .Q(net_6359), .SI(net_6358), .D(net_3595), .SE(net_392), .CK(net_13964) );
NAND2_X2 inst_3063 ( .A1(net_7126), .A2(net_4950), .ZN(net_4942) );
CLKBUF_X2 inst_13881 ( .A(net_13842), .Z(net_13843) );
CLKBUF_X2 inst_8610 ( .A(net_8085), .Z(net_8572) );
OAI21_X2 inst_1812 ( .ZN(net_5376), .B1(net_5353), .A(net_4346), .B2(net_3859) );
AOI222_X2 inst_7608 ( .ZN(net_5349), .A2(net_1222), .B1(net_1221), .C1(net_1220), .B2(net_345), .C2(net_343), .A1(net_331) );
CLKBUF_X2 inst_12257 ( .A(net_12115), .Z(net_12219) );
INV_X4 inst_5643 ( .A(net_7411), .ZN(net_2198) );
DFF_X1 inst_6750 ( .QN(net_7617), .D(net_4844), .CK(net_10290) );
CLKBUF_X2 inst_12555 ( .A(net_12516), .Z(net_12517) );
CLKBUF_X2 inst_8217 ( .A(net_8178), .Z(net_8179) );
CLKBUF_X2 inst_8370 ( .A(net_8092), .Z(net_8332) );
CLKBUF_X2 inst_12051 ( .A(net_12012), .Z(net_12013) );
NAND2_X1 inst_4338 ( .ZN(net_4389), .A2(net_3856), .A1(net_1766) );
CLKBUF_X2 inst_8806 ( .A(net_8671), .Z(net_8768) );
CLKBUF_X2 inst_12726 ( .A(net_12687), .Z(net_12688) );
CLKBUF_X2 inst_13066 ( .A(net_8596), .Z(net_13028) );
INV_X4 inst_4721 ( .ZN(net_3020), .A(net_2864) );
CLKBUF_X2 inst_13601 ( .A(net_8219), .Z(net_13563) );
CLKBUF_X2 inst_8194 ( .A(net_8155), .Z(net_8156) );
CLKBUF_X2 inst_12846 ( .A(net_12807), .Z(net_12808) );
NAND2_X4 inst_2835 ( .ZN(net_5557), .A1(net_5028), .A2(net_5027) );
DFF_X1 inst_6638 ( .QN(net_7616), .D(net_5241), .CK(net_9461) );
CLKBUF_X2 inst_11136 ( .A(net_9496), .Z(net_11098) );
CLKBUF_X2 inst_10399 ( .A(net_10360), .Z(net_10361) );
NAND3_X2 inst_2731 ( .ZN(net_2370), .A3(net_1628), .A1(net_1407), .A2(net_977) );
CLKBUF_X2 inst_13019 ( .A(net_12980), .Z(net_12981) );
CLKBUF_X2 inst_8663 ( .A(net_8624), .Z(net_8625) );
NOR3_X2 inst_2207 ( .ZN(net_2726), .A3(net_2724), .A1(net_2711), .A2(net_1951) );
AND2_X4 inst_7841 ( .ZN(net_1400), .A2(net_785), .A1(net_640) );
CLKBUF_X2 inst_10088 ( .A(net_10049), .Z(net_10050) );
INV_X2 inst_5902 ( .A(net_7295), .ZN(net_2061) );
AOI22_X2 inst_7322 ( .ZN(net_3436), .A2(net_3435), .B2(net_3434), .A1(net_1309), .B1(net_1051) );
NAND2_X2 inst_3892 ( .A1(net_6978), .A2(net_1833), .ZN(net_1424) );
INV_X4 inst_4813 ( .ZN(net_4788), .A(net_1165) );
CLKBUF_X2 inst_8829 ( .A(net_8790), .Z(net_8791) );
NAND2_X2 inst_3930 ( .A1(net_6965), .A2(net_1833), .ZN(net_1368) );
NAND2_X4 inst_2867 ( .ZN(net_4284), .A1(net_4272), .A2(net_1655) );
CLKBUF_X2 inst_9725 ( .A(net_8697), .Z(net_9687) );
CLKBUF_X2 inst_9768 ( .A(net_9729), .Z(net_9730) );
NAND2_X2 inst_3398 ( .ZN(net_3540), .A2(net_3331), .A1(net_3239) );
SDFF_X2 inst_477 ( .Q(net_6871), .D(net_6871), .SE(net_3901), .SI(net_3894), .CK(net_11817) );
CLKBUF_X2 inst_7953 ( .A(net_7914), .Z(net_7915) );
CLKBUF_X2 inst_14235 ( .A(net_14196), .Z(net_14197) );
NAND2_X2 inst_3576 ( .ZN(net_2464), .A2(net_1976), .A1(net_1469) );
CLKBUF_X2 inst_10006 ( .A(net_9891), .Z(net_9968) );
SDFF_X2 inst_423 ( .D(net_6391), .SE(net_6052), .SI(net_316), .Q(net_316), .CK(net_13810) );
SDFF_X2 inst_835 ( .Q(net_7015), .D(net_7015), .SE(net_3899), .SI(net_3807), .CK(net_11895) );
NAND2_X2 inst_3305 ( .ZN(net_3636), .A1(net_3635), .A2(net_3229) );
NAND2_X2 inst_3082 ( .A1(net_6481), .A2(net_4927), .ZN(net_4921) );
NAND2_X2 inst_4137 ( .A2(net_1222), .ZN(net_1137), .A1(net_343) );
SDFF_X2 inst_1112 ( .SI(net_6667), .Q(net_6667), .D(net_3812), .SE(net_3465), .CK(net_9327) );
DFF_X1 inst_6852 ( .D(net_2553), .QN(net_217), .CK(net_9743) );
CLKBUF_X2 inst_10153 ( .A(net_10114), .Z(net_10115) );
CLKBUF_X2 inst_9678 ( .A(net_8607), .Z(net_9640) );
NAND2_X2 inst_4081 ( .A1(net_6521), .A2(net_1645), .ZN(net_971) );
SDFF_X2 inst_710 ( .SI(net_6782), .Q(net_6782), .SE(net_3816), .D(net_3779), .CK(net_8364) );
SDFF_X2 inst_941 ( .SI(net_7183), .Q(net_7183), .SE(net_3819), .D(net_3783), .CK(net_11563) );
NAND2_X2 inst_3350 ( .ZN(net_3547), .A1(net_3546), .A2(net_3226) );
CLKBUF_X2 inst_8869 ( .A(net_8830), .Z(net_8831) );
CLKBUF_X2 inst_8398 ( .A(net_8152), .Z(net_8360) );
CLKBUF_X2 inst_10375 ( .A(net_10336), .Z(net_10337) );
OAI21_X2 inst_1817 ( .ZN(net_5371), .B1(net_5343), .A(net_4338), .B2(net_3859) );
XNOR2_X2 inst_56 ( .ZN(net_2243), .A(net_2242), .B(net_2241) );
DFF_X1 inst_6835 ( .D(net_2620), .CK(net_10546), .Q(x138) );
SDFF_X2 inst_308 ( .SI(net_7524), .Q(net_7524), .D(net_5101), .SE(net_3988), .CK(net_9646) );
CLKBUF_X2 inst_11056 ( .A(net_11017), .Z(net_11018) );
OAI22_X2 inst_1546 ( .B2(net_3405), .A2(net_3360), .ZN(net_3359), .A1(net_3289), .B1(net_590) );
CLKBUF_X2 inst_11224 ( .A(net_11185), .Z(net_11186) );
CLKBUF_X2 inst_10081 ( .A(net_10042), .Z(net_10043) );
SDFF_X2 inst_455 ( .Q(net_6058), .SI(net_3919), .SE(net_3314), .D(net_3313), .CK(net_13169) );
CLKBUF_X2 inst_8449 ( .A(net_8410), .Z(net_8411) );
CLKBUF_X2 inst_10015 ( .A(net_9976), .Z(net_9977) );
NAND2_X4 inst_2871 ( .A1(net_5881), .ZN(net_4268), .A2(net_2579) );
OAI21_X2 inst_1694 ( .B2(net_5906), .ZN(net_5600), .A(net_5288), .B1(net_4105) );
NOR2_X2 inst_2540 ( .A2(net_7752), .A1(net_3208), .ZN(net_654) );
DFF_X1 inst_6833 ( .D(net_2586), .QN(net_190), .CK(net_12295) );
AOI222_X2 inst_7475 ( .C1(net_7528), .B1(net_7496), .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2155), .A1(net_2154) );
CLKBUF_X2 inst_13298 ( .A(net_8467), .Z(net_13260) );
NAND2_X2 inst_3629 ( .ZN(net_1954), .A1(net_1293), .A2(net_1116) );
CLKBUF_X2 inst_12593 ( .A(net_12554), .Z(net_12555) );
DFFR_X2 inst_7052 ( .QN(net_6021), .D(net_3132), .CK(net_8584), .RN(x1822) );
DFF_X1 inst_6602 ( .QN(net_7509), .D(net_5406), .CK(net_9245) );
CLKBUF_X2 inst_8114 ( .A(net_8075), .Z(net_8076) );
NAND2_X2 inst_3024 ( .A1(net_6882), .A2(net_5006), .ZN(net_4985) );
CLKBUF_X2 inst_13370 ( .A(net_13331), .Z(net_13332) );
CLKBUF_X2 inst_9946 ( .A(net_8270), .Z(net_9908) );
CLKBUF_X2 inst_8454 ( .A(net_8170), .Z(net_8416) );
NAND2_X1 inst_4414 ( .A2(net_5966), .A1(net_5965), .ZN(net_2878) );
DFFR_X1 inst_7129 ( .D(net_3369), .Q(net_297), .CK(net_13300), .RN(x1822) );
CLKBUF_X2 inst_11860 ( .A(net_11821), .Z(net_11822) );
CLKBUF_X2 inst_10052 ( .A(net_8995), .Z(net_10014) );
NAND2_X2 inst_3085 ( .A1(net_6450), .A2(net_4925), .ZN(net_4918) );
CLKBUF_X2 inst_8648 ( .A(net_8609), .Z(net_8610) );
AOI21_X4 inst_7620 ( .B2(net_5949), .B1(net_5948), .ZN(net_5608), .A(x1006) );
NAND2_X2 inst_3951 ( .A1(net_7118), .A2(net_1675), .ZN(net_1336) );
CLKBUF_X2 inst_8240 ( .A(net_7910), .Z(net_8202) );
NAND2_X1 inst_4282 ( .ZN(net_4585), .A2(net_3867), .A1(net_1856) );
INV_X4 inst_5428 ( .A(net_7257), .ZN(net_1997) );
NAND2_X2 inst_2943 ( .ZN(net_5503), .A1(net_4966), .A2(net_4965) );
OAI22_X2 inst_1593 ( .A1(net_3265), .B2(net_3200), .A2(net_3196), .ZN(net_3146), .B1(net_482) );
CLKBUF_X2 inst_13768 ( .A(net_13729), .Z(net_13730) );
INV_X4 inst_5661 ( .A(net_5989), .ZN(net_573) );
CLKBUF_X2 inst_9918 ( .A(net_9879), .Z(net_9880) );
CLKBUF_X2 inst_11541 ( .A(net_9134), .Z(net_11503) );
CLKBUF_X2 inst_14120 ( .A(net_14081), .Z(net_14082) );
SDFF_X2 inst_724 ( .Q(net_6840), .D(net_6840), .SE(net_3893), .SI(net_3813), .CK(net_11511) );
NAND2_X1 inst_4292 ( .ZN(net_4575), .A2(net_3867), .A1(net_1873) );
CLKBUF_X2 inst_12083 ( .A(net_9606), .Z(net_12045) );
NOR2_X2 inst_2449 ( .ZN(net_2862), .A1(net_2861), .A2(net_2860) );
DFF_X1 inst_6570 ( .QN(net_7506), .D(net_5092), .CK(net_9250) );
SDFF_X2 inst_975 ( .Q(net_6455), .D(net_6455), .SE(net_3820), .SI(net_3800), .CK(net_8069) );
CLKBUF_X2 inst_13683 ( .A(net_12169), .Z(net_13645) );
CLKBUF_X2 inst_13096 ( .A(net_13057), .Z(net_13058) );
NAND2_X2 inst_3191 ( .ZN(net_4735), .A2(net_3986), .A1(net_2129) );
NAND3_X2 inst_2789 ( .ZN(net_2311), .A1(net_1678), .A3(net_1601), .A2(net_1000) );
AND4_X2 inst_7792 ( .A4(net_2916), .ZN(net_2490), .A3(net_2489), .A2(net_2486), .A1(net_1656) );
CLKBUF_X2 inst_9504 ( .A(net_7844), .Z(net_9466) );
OAI22_X2 inst_1431 ( .B1(net_5859), .ZN(net_5798), .A2(net_5792), .B2(net_5791), .A1(net_5774) );
INV_X2 inst_5714 ( .ZN(net_4252), .A(net_4125) );
NAND2_X2 inst_3760 ( .A1(net_7033), .A2(net_1975), .ZN(net_1585) );
CLKBUF_X2 inst_12841 ( .A(net_9473), .Z(net_12803) );
CLKBUF_X2 inst_10110 ( .A(net_8015), .Z(net_10072) );
OR2_X4 inst_1398 ( .A2(net_7229), .A1(net_7228), .ZN(net_487) );
AOI21_X2 inst_7639 ( .ZN(net_3951), .B2(net_3757), .B1(net_2888), .A(net_927) );
CLKBUF_X2 inst_10783 ( .A(net_10744), .Z(net_10745) );
CLKBUF_X2 inst_8477 ( .A(net_7916), .Z(net_8439) );
DFFR_X1 inst_7122 ( .Q(net_6036), .D(net_4795), .CK(net_10037), .RN(x1822) );
NAND2_X4 inst_2849 ( .ZN(net_5474), .A1(net_4917), .A2(net_4916) );
OAI21_X2 inst_1804 ( .ZN(net_5386), .A(net_4712), .B2(net_3986), .B1(net_1094) );
CLKBUF_X2 inst_13808 ( .A(net_13769), .Z(net_13770) );
NOR2_X2 inst_2440 ( .A2(net_5975), .ZN(net_3164), .A1(net_3004) );
DFF_X1 inst_6418 ( .QN(net_6153), .D(net_5752), .CK(net_9046) );
CLKBUF_X2 inst_9261 ( .A(net_9222), .Z(net_9223) );
CLKBUF_X2 inst_11037 ( .A(net_10697), .Z(net_10999) );
NOR4_X2 inst_2183 ( .ZN(net_2300), .A2(net_2299), .A4(net_2275), .A1(net_1311), .A3(net_1052) );
CLKBUF_X2 inst_11981 ( .A(net_11898), .Z(net_11943) );
NAND2_X2 inst_3327 ( .ZN(net_3592), .A1(net_3591), .A2(net_3228) );
INV_X4 inst_5068 ( .A(net_785), .ZN(net_726) );
CLKBUF_X2 inst_10241 ( .A(net_10202), .Z(net_10203) );
NAND3_X2 inst_2659 ( .ZN(net_3941), .A1(net_3940), .A3(net_3858), .A2(net_1726) );
DFF_X1 inst_6545 ( .QN(net_7324), .D(net_5364), .CK(net_13013) );
OAI21_X2 inst_2134 ( .A(net_5922), .ZN(net_2852), .B1(net_2851), .B2(net_2850) );
OAI21_X2 inst_1744 ( .ZN(net_5528), .A(net_4823), .B2(net_4153), .B1(net_1259) );
CLKBUF_X2 inst_13878 ( .A(net_8141), .Z(net_13840) );
INV_X4 inst_4805 ( .ZN(net_4781), .A(net_1177) );
INV_X4 inst_5018 ( .ZN(net_1821), .A(net_1232) );
CLKBUF_X2 inst_11609 ( .A(net_11570), .Z(net_11571) );
INV_X4 inst_5628 ( .A(net_7695), .ZN(net_709) );
INV_X4 inst_5641 ( .A(net_7692), .ZN(net_838) );
CLKBUF_X2 inst_11958 ( .A(net_11919), .Z(net_11920) );
CLKBUF_X2 inst_11134 ( .A(net_11095), .Z(net_11096) );
SDFF_X2 inst_1155 ( .SI(net_6818), .Q(net_6818), .D(net_3788), .SE(net_3722), .CK(net_8331) );
NAND2_X2 inst_4117 ( .A2(net_1225), .ZN(net_1070), .A1(net_363) );
CLKBUF_X2 inst_11311 ( .A(net_9803), .Z(net_11273) );
SDFF_X2 inst_207 ( .Q(net_6307), .SI(net_6306), .D(net_3673), .SE(net_392), .CK(net_13562) );
CLKBUF_X2 inst_9329 ( .A(net_9290), .Z(net_9291) );
CLKBUF_X2 inst_8886 ( .A(net_8287), .Z(net_8848) );
CLKBUF_X2 inst_11198 ( .A(net_11159), .Z(net_11160) );
CLKBUF_X2 inst_10047 ( .A(net_8892), .Z(net_10009) );
CLKBUF_X2 inst_11639 ( .A(net_11600), .Z(net_11601) );
CLKBUF_X2 inst_11954 ( .A(net_11915), .Z(net_11916) );
CLKBUF_X2 inst_10490 ( .A(net_10451), .Z(net_10452) );
DFF_X1 inst_6940 ( .QN(net_6052), .D(net_2276), .CK(net_14366) );
CLKBUF_X2 inst_9615 ( .A(net_8869), .Z(net_9577) );
SDFF_X2 inst_712 ( .SI(net_6785), .Q(net_6785), .SE(net_3872), .D(net_3789), .CK(net_11325) );
CLKBUF_X2 inst_9912 ( .A(net_9714), .Z(net_9874) );
SDFF_X2 inst_1215 ( .SI(net_7205), .Q(net_7205), .D(net_3894), .SE(net_3750), .CK(net_10479) );
CLKBUF_X2 inst_9303 ( .A(net_7839), .Z(net_9265) );
SDFF_X2 inst_131 ( .QN(net_6219), .SI(net_6218), .SE(net_392), .D(net_153), .CK(net_14242) );
CLKBUF_X2 inst_14271 ( .A(net_14232), .Z(net_14233) );
CLKBUF_X2 inst_12436 ( .A(net_12397), .Z(net_12398) );
INV_X2 inst_6104 ( .A(net_7627), .ZN(net_1914) );
NAND2_X2 inst_3111 ( .A1(net_6618), .A2(net_4899), .ZN(net_4890) );
XNOR2_X2 inst_47 ( .B(net_6960), .ZN(net_2438), .A(net_1238) );
OAI21_X2 inst_2035 ( .B2(net_4476), .ZN(net_4468), .B1(net_4223), .A(net_3596) );
CLKBUF_X2 inst_12360 ( .A(net_12321), .Z(net_12322) );
CLKBUF_X2 inst_13530 ( .A(net_13491), .Z(net_13492) );
OAI21_X2 inst_1984 ( .B1(net_4851), .ZN(net_4845), .A(net_4582), .B2(net_3867) );
INV_X4 inst_5231 ( .A(net_460), .ZN(net_459) );
CLKBUF_X2 inst_11569 ( .A(net_11530), .Z(net_11531) );
CLKBUF_X2 inst_10442 ( .A(net_9287), .Z(net_10404) );
CLKBUF_X2 inst_11121 ( .A(net_11082), .Z(net_11083) );
CLKBUF_X2 inst_9458 ( .A(net_9419), .Z(net_9420) );
DFF_X1 inst_6520 ( .QN(net_7436), .D(net_5431), .CK(net_12483) );
CLKBUF_X2 inst_14356 ( .A(net_8768), .Z(net_14318) );
CLKBUF_X2 inst_12564 ( .A(net_12336), .Z(net_12526) );
CLKBUF_X2 inst_12397 ( .A(net_12358), .Z(net_12359) );
NAND2_X2 inst_4101 ( .A1(net_6940), .A2(net_1654), .ZN(net_951) );
DFF_X1 inst_6483 ( .QN(net_7414), .D(net_5569), .CK(net_9311) );
CLKBUF_X2 inst_10316 ( .A(net_10277), .Z(net_10278) );
CLKBUF_X2 inst_9469 ( .A(net_9430), .Z(net_9431) );
CLKBUF_X2 inst_12482 ( .A(net_12443), .Z(net_12444) );
INV_X4 inst_4792 ( .ZN(net_1269), .A(net_1268) );
AOI22_X2 inst_7381 ( .A2(net_5916), .B2(net_2957), .ZN(net_2940), .B1(net_2670), .A1(net_858) );
CLKBUF_X2 inst_14027 ( .A(net_7949), .Z(net_13989) );
SDFF_X2 inst_525 ( .SI(net_6644), .Q(net_6644), .SE(net_3850), .D(net_3836), .CK(net_9125) );
CLKBUF_X2 inst_12738 ( .A(net_9100), .Z(net_12700) );
SDFF_X2 inst_434 ( .Q(net_7386), .D(net_7386), .SE(net_3994), .SI(net_351), .CK(net_9751) );
CLKBUF_X2 inst_12196 ( .A(net_12157), .Z(net_12158) );
CLKBUF_X2 inst_11774 ( .A(net_11735), .Z(net_11736) );
NAND2_X2 inst_3455 ( .ZN(net_3068), .A1(net_2916), .A2(net_2907) );
CLKBUF_X2 inst_12424 ( .A(net_12385), .Z(net_12386) );
SDFF_X2 inst_1032 ( .Q(net_7548), .D(net_7548), .SE(net_3896), .SI(net_382), .CK(net_13115) );
CLKBUF_X2 inst_8985 ( .A(net_8946), .Z(net_8947) );
CLKBUF_X2 inst_14099 ( .A(net_14060), .Z(net_14061) );
CLKBUF_X2 inst_12638 ( .A(net_12599), .Z(net_12600) );
DFF_X1 inst_6711 ( .QN(net_7327), .D(net_5358), .CK(net_10152) );
OR2_X4 inst_1392 ( .A1(net_891), .ZN(net_811), .A2(net_399) );
INV_X2 inst_5932 ( .A(net_7333), .ZN(net_1749) );
AOI22_X2 inst_7376 ( .B1(net_7738), .A1(net_7709), .A2(net_5916), .B2(net_2957), .ZN(net_2945) );
CLKBUF_X2 inst_11816 ( .A(net_11705), .Z(net_11778) );
NAND2_X2 inst_4044 ( .A1(net_6925), .A2(net_1654), .ZN(net_1008) );
AOI222_X2 inst_7585 ( .A1(net_7396), .ZN(net_5444), .A2(net_1225), .B1(net_1224), .C1(net_1223), .B2(net_359), .C2(net_357) );
CLKBUF_X2 inst_11682 ( .A(net_11643), .Z(net_11644) );
OAI22_X2 inst_1476 ( .B1(net_4855), .A1(net_4228), .B2(net_4220), .ZN(net_4217), .A2(net_4216) );
CLKBUF_X2 inst_8265 ( .A(net_8226), .Z(net_8227) );
CLKBUF_X2 inst_11148 ( .A(net_8850), .Z(net_11110) );
NOR2_X4 inst_2249 ( .ZN(net_5637), .A1(net_5483), .A2(net_4449) );
CLKBUF_X2 inst_12339 ( .A(net_8199), .Z(net_12301) );
CLKBUF_X2 inst_11106 ( .A(net_9094), .Z(net_11068) );
CLKBUF_X2 inst_13773 ( .A(net_11291), .Z(net_13735) );
CLKBUF_X2 inst_8995 ( .A(net_8956), .Z(net_8957) );
INV_X4 inst_5404 ( .A(net_7696), .ZN(net_712) );
NOR2_X4 inst_2269 ( .ZN(net_5617), .A1(net_5462), .A2(net_4411) );
NOR2_X2 inst_2390 ( .ZN(net_4290), .A1(net_4138), .A2(net_4137) );
OAI21_X2 inst_1780 ( .ZN(net_5413), .B1(net_5412), .A(net_4692), .B2(net_3989) );
CLKBUF_X2 inst_11839 ( .A(net_9945), .Z(net_11801) );
OAI22_X2 inst_1436 ( .B1(net_5853), .ZN(net_5793), .A2(net_5782), .B2(net_5781), .A1(net_5769) );
INV_X2 inst_6033 ( .A(net_7584), .ZN(net_2127) );
CLKBUF_X2 inst_14305 ( .A(net_14266), .Z(net_14267) );
SDFF_X2 inst_852 ( .SI(net_7802), .Q(net_7005), .D(net_7005), .SE(net_3899), .CK(net_9025) );
CLKBUF_X2 inst_12792 ( .A(net_12753), .Z(net_12754) );
CLKBUF_X2 inst_8424 ( .A(net_8137), .Z(net_8386) );
NAND2_X2 inst_3871 ( .A1(net_6702), .A2(net_1497), .ZN(net_1457) );
CLKBUF_X2 inst_9268 ( .A(net_8655), .Z(net_9230) );
DFF_X1 inst_6663 ( .QN(net_7656), .D(net_5175), .CK(net_10552) );
NAND2_X1 inst_4306 ( .ZN(net_4560), .A2(net_3866), .A1(net_2100) );
CLKBUF_X2 inst_12528 ( .A(net_12489), .Z(net_12490) );
OAI22_X2 inst_1474 ( .B1(net_4855), .A1(net_4228), .B2(net_4225), .ZN(net_4221), .A2(net_4220) );
NAND2_X1 inst_4449 ( .A2(net_1256), .ZN(net_1132), .A1(net_1131) );
INV_X2 inst_6077 ( .A(net_7749), .ZN(net_5874) );
CLKBUF_X2 inst_11974 ( .A(net_7995), .Z(net_11936) );
AOI21_X2 inst_7637 ( .ZN(net_3953), .B2(net_3763), .B1(net_2890), .A(net_931) );
OAI21_X2 inst_2045 ( .B2(net_4457), .ZN(net_4455), .B1(net_4078), .A(net_3492) );
OAI21_X2 inst_1920 ( .B1(net_5335), .ZN(net_5143), .A(net_4745), .B2(net_3941) );
CLKBUF_X2 inst_11746 ( .A(net_11707), .Z(net_11708) );
CLKBUF_X2 inst_9022 ( .A(net_8983), .Z(net_8984) );
SDFF_X2 inst_1311 ( .D(net_6383), .SE(net_5799), .SI(net_368), .Q(net_368), .CK(net_13869) );
CLKBUF_X2 inst_9307 ( .A(net_9268), .Z(net_9269) );
NAND2_X2 inst_3415 ( .ZN(net_3442), .A2(net_3258), .A1(net_754) );
CLKBUF_X2 inst_13269 ( .A(net_13230), .Z(net_13231) );
CLKBUF_X2 inst_12787 ( .A(net_12748), .Z(net_12749) );
CLKBUF_X2 inst_9534 ( .A(net_9495), .Z(net_9496) );
CLKBUF_X2 inst_10780 ( .A(net_10741), .Z(net_10742) );
INV_X4 inst_4654 ( .ZN(net_4605), .A(net_4272) );
OAI221_X2 inst_1640 ( .ZN(net_5455), .B2(net_5383), .C2(net_5090), .A(net_5037), .C1(net_1151), .B1(net_721) );
CLKBUF_X2 inst_11359 ( .A(net_8264), .Z(net_11321) );
CLKBUF_X2 inst_11194 ( .A(net_11155), .Z(net_11156) );
NAND2_X2 inst_3234 ( .ZN(net_4283), .A2(net_4282), .A1(net_1635) );
NAND2_X2 inst_4143 ( .A1(net_1149), .ZN(net_912), .A2(net_702) );
CLKBUF_X2 inst_13928 ( .A(net_13889), .Z(net_13890) );
NAND3_X2 inst_2639 ( .ZN(net_5690), .A1(net_5667), .A2(net_5295), .A3(net_4241) );
INV_X4 inst_4747 ( .ZN(net_2754), .A(net_2630) );
AOI21_X2 inst_7682 ( .B1(net_7003), .ZN(net_4477), .A(net_2469), .B2(net_1100) );
CLKBUF_X2 inst_11122 ( .A(net_11083), .Z(net_11084) );
AOI222_X2 inst_7571 ( .A1(net_7551), .ZN(net_5225), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_383), .C2(net_381) );
INV_X4 inst_4630 ( .ZN(net_4192), .A(net_4044) );
NOR2_X2 inst_2509 ( .A2(net_3236), .ZN(net_1180), .A1(net_1179) );
INV_X2 inst_5971 ( .A(net_7437), .ZN(net_1507) );
INV_X2 inst_5897 ( .A(net_7433), .ZN(net_1459) );
NOR2_X2 inst_2542 ( .A2(net_5936), .ZN(net_2590), .A1(net_769) );
DFF_X1 inst_6632 ( .QN(net_7588), .D(net_5251), .CK(net_13161) );
NAND2_X2 inst_3091 ( .A1(net_6453), .A2(net_4925), .ZN(net_4912) );
NAND2_X2 inst_4197 ( .ZN(net_1215), .A1(net_650), .A2(net_307) );
CLKBUF_X2 inst_11791 ( .A(net_10839), .Z(net_11753) );
CLKBUF_X2 inst_9506 ( .A(net_9467), .Z(net_9468) );
DFF_X1 inst_6829 ( .D(net_2589), .QN(net_225), .CK(net_12303) );
AOI222_X2 inst_7567 ( .A1(net_7543), .ZN(net_5200), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_375), .C2(net_373) );
DFF_X1 inst_6590 ( .QN(net_7560), .D(net_5060), .CK(net_13165) );
SDFF_X2 inst_417 ( .D(net_6392), .SE(net_6052), .SI(net_317), .Q(net_317), .CK(net_13815) );
SDFF_X2 inst_671 ( .SI(net_7802), .Q(net_6703), .D(net_6703), .SE(net_3871), .CK(net_11101) );
AOI22_X2 inst_7400 ( .B1(net_5939), .ZN(net_2840), .A1(net_2839), .A2(net_2838), .B2(net_202) );
CLKBUF_X2 inst_13473 ( .A(net_13434), .Z(net_13435) );
CLKBUF_X2 inst_12733 ( .A(net_10835), .Z(net_12695) );
XNOR2_X2 inst_21 ( .ZN(net_2613), .A(net_2247), .B(net_1210) );
CLKBUF_X2 inst_9462 ( .A(net_8989), .Z(net_9424) );
CLKBUF_X2 inst_13745 ( .A(net_13706), .Z(net_13707) );
INV_X8 inst_4524 ( .ZN(net_3742), .A(net_3115) );
CLKBUF_X2 inst_11024 ( .A(net_10985), .Z(net_10986) );
INV_X4 inst_4871 ( .ZN(net_2855), .A(net_909) );
CLKBUF_X2 inst_10286 ( .A(net_8068), .Z(net_10248) );
INV_X4 inst_5520 ( .A(net_6689), .ZN(net_471) );
NAND2_X2 inst_3885 ( .A1(net_6427), .A2(net_1677), .ZN(net_1434) );
NOR2_X2 inst_2311 ( .A2(net_6203), .A1(net_5843), .ZN(net_5830) );
NAND2_X1 inst_4257 ( .ZN(net_4668), .A2(net_3993), .A1(net_1494) );
INV_X4 inst_4586 ( .ZN(net_4316), .A(net_4232) );
AOI21_X2 inst_7703 ( .B1(net_6880), .ZN(net_4087), .B2(net_2579), .A(net_2346) );
CLKBUF_X2 inst_13722 ( .A(net_12933), .Z(net_13684) );
SDFF_X2 inst_1317 ( .D(net_6381), .SE(net_5799), .SI(net_366), .Q(net_366), .CK(net_13864) );
DFF_X1 inst_6820 ( .QN(net_5964), .D(net_3012), .CK(net_12543) );
NAND2_X2 inst_3683 ( .A2(net_1798), .ZN(net_1767), .A1(net_1766) );
NAND2_X2 inst_2941 ( .ZN(net_5505), .A1(net_4970), .A2(net_4969) );
CLKBUF_X2 inst_13655 ( .A(net_11686), .Z(net_13617) );
CLKBUF_X2 inst_9623 ( .A(net_8482), .Z(net_9585) );
CLKBUF_X2 inst_12603 ( .A(net_12564), .Z(net_12565) );
CLKBUF_X2 inst_13528 ( .A(net_13489), .Z(net_13490) );
CLKBUF_X2 inst_12351 ( .A(net_8874), .Z(net_12313) );
CLKBUF_X2 inst_9861 ( .A(net_9822), .Z(net_9823) );
CLKBUF_X2 inst_9203 ( .A(net_9164), .Z(net_9165) );
SDFF_X2 inst_624 ( .SI(net_6634), .Q(net_6634), .SE(net_3851), .D(net_3813), .CK(net_9336) );
DFF_X2 inst_6284 ( .QN(net_6051), .D(net_2300), .CK(net_14347) );
INV_X2 inst_5728 ( .ZN(net_3968), .A(net_3967) );
CLKBUF_X2 inst_8442 ( .A(net_8403), .Z(net_8404) );
DFF_X1 inst_6404 ( .QN(net_6143), .D(net_5766), .CK(net_8164) );
CLKBUF_X2 inst_11930 ( .A(net_11891), .Z(net_11892) );
CLKBUF_X2 inst_10920 ( .A(net_10881), .Z(net_10882) );
DFF_X1 inst_6419 ( .QN(net_6174), .D(net_5751), .CK(net_11616) );
CLKBUF_X2 inst_9886 ( .A(net_9847), .Z(net_9848) );
CLKBUF_X2 inst_11247 ( .A(net_11208), .Z(net_11209) );
CLKBUF_X2 inst_9375 ( .A(net_9193), .Z(net_9337) );
NAND3_X2 inst_2637 ( .ZN(net_5692), .A1(net_5669), .A2(net_5299), .A3(net_4243) );
CLKBUF_X2 inst_9604 ( .A(net_9565), .Z(net_9566) );
NAND2_X2 inst_3624 ( .ZN(net_1959), .A1(net_1295), .A2(net_1130) );
CLKBUF_X2 inst_13207 ( .A(net_13062), .Z(net_13169) );
SDFF_X2 inst_236 ( .Q(net_6358), .SI(net_6357), .D(net_3597), .SE(net_392), .CK(net_13504) );
CLKBUF_X2 inst_11440 ( .A(net_11401), .Z(net_11402) );
INV_X8 inst_4539 ( .ZN(net_2970), .A(net_1819) );
CLKBUF_X2 inst_12389 ( .A(net_12350), .Z(net_12351) );
NAND2_X2 inst_3878 ( .A1(net_6436), .A2(net_1677), .ZN(net_1442) );
CLKBUF_X2 inst_13295 ( .A(net_10117), .Z(net_13257) );
CLKBUF_X2 inst_13262 ( .A(net_13223), .Z(net_13224) );
CLKBUF_X2 inst_9806 ( .A(net_9767), .Z(net_9768) );
NAND2_X2 inst_3172 ( .ZN(net_4761), .A2(net_3941), .A1(net_2055) );
SDFF_X2 inst_986 ( .Q(net_6472), .D(net_6472), .SE(net_3904), .SI(net_3809), .CK(net_8781) );
INV_X8 inst_4532 ( .ZN(net_5840), .A(net_392) );
INV_X4 inst_4983 ( .ZN(net_2652), .A(net_684) );
DFF_X2 inst_6277 ( .D(net_2613), .QN(net_192), .CK(net_12290) );
CLKBUF_X2 inst_12962 ( .A(net_9272), .Z(net_12924) );
OR2_X2 inst_1422 ( .ZN(net_2868), .A2(net_707), .A1(net_562) );
INV_X4 inst_5600 ( .A(net_5858), .ZN(net_603) );
CLKBUF_X2 inst_10263 ( .A(net_10224), .Z(net_10225) );
CLKBUF_X2 inst_8337 ( .A(net_8140), .Z(net_8299) );
NAND2_X2 inst_3508 ( .ZN(net_2559), .A2(net_2195), .A1(net_1382) );
INV_X4 inst_5132 ( .ZN(net_617), .A(net_582) );
DFF_X2 inst_6327 ( .QN(net_7817), .CK(net_11033), .D(x1398) );
CLKBUF_X2 inst_9702 ( .A(net_9663), .Z(net_9664) );
DFF_X1 inst_6893 ( .D(net_2517), .Q(net_170), .CK(net_10222) );
CLKBUF_X2 inst_10522 ( .A(net_10483), .Z(net_10484) );
SDFF_X2 inst_1221 ( .SI(net_7214), .Q(net_7214), .D(net_3807), .SE(net_3751), .CK(net_7831) );
CLKBUF_X2 inst_8675 ( .A(net_8636), .Z(net_8637) );
SDFF_X2 inst_1133 ( .SI(net_6657), .Q(net_6657), .D(net_3802), .SE(net_3471), .CK(net_10047) );
AOI21_X2 inst_7750 ( .B1(net_6876), .ZN(net_4095), .B2(net_2579), .A(net_2331) );
CLKBUF_X2 inst_12158 ( .A(net_8348), .Z(net_12120) );
INV_X4 inst_4580 ( .A(net_5089), .ZN(net_4332) );
CLKBUF_X2 inst_9990 ( .A(net_9951), .Z(net_9952) );
OAI21_X2 inst_2103 ( .ZN(net_3978), .A(net_3977), .B2(net_3877), .B1(net_1089) );
CLKBUF_X2 inst_7951 ( .A(net_7867), .Z(net_7913) );
CLKBUF_X2 inst_8710 ( .A(net_8671), .Z(net_8672) );
CLKBUF_X2 inst_14040 ( .A(net_8518), .Z(net_14002) );
INV_X4 inst_5139 ( .A(net_1224), .ZN(net_576) );
CLKBUF_X2 inst_10793 ( .A(net_10754), .Z(net_10755) );
NAND3_X2 inst_2664 ( .ZN(net_3932), .A3(net_3393), .A2(net_2930), .A1(net_2829) );
SDFF_X2 inst_339 ( .SI(net_7522), .Q(net_7522), .D(net_5094), .SE(net_3988), .CK(net_9757) );
INV_X4 inst_4750 ( .ZN(net_2630), .A(net_189) );
CLKBUF_X2 inst_13995 ( .A(net_10401), .Z(net_13957) );
SDFF_X2 inst_351 ( .SI(net_7669), .Q(net_7669), .D(net_4801), .SE(net_3866), .CK(net_8009) );
DFF_X1 inst_6615 ( .QN(net_7576), .D(net_5392), .CK(net_10312) );
CLKBUF_X2 inst_11615 ( .A(net_10750), .Z(net_11577) );
CLKBUF_X2 inst_10257 ( .A(net_10218), .Z(net_10219) );
CLKBUF_X2 inst_9557 ( .A(net_7933), .Z(net_9519) );
CLKBUF_X2 inst_8761 ( .A(net_7942), .Z(net_8723) );
AND2_X2 inst_7852 ( .ZN(net_3715), .A2(net_3327), .A1(net_394) );
DFF_X1 inst_6757 ( .QN(net_7283), .D(net_4869), .CK(net_12797) );
CLKBUF_X2 inst_12507 ( .A(net_12468), .Z(net_12469) );
CLKBUF_X2 inst_8170 ( .A(net_7945), .Z(net_8132) );
CLKBUF_X2 inst_7915 ( .A(net_7876), .Z(net_7877) );
INV_X2 inst_5862 ( .A(net_829), .ZN(net_585) );
AOI21_X2 inst_7651 ( .B2(net_3439), .ZN(net_3395), .A(net_3215), .B1(net_3082) );
CLKBUF_X2 inst_14007 ( .A(net_8036), .Z(net_13969) );
CLKBUF_X2 inst_10966 ( .A(net_10248), .Z(net_10928) );
OAI22_X2 inst_1560 ( .B2(net_3405), .A2(net_3360), .ZN(net_3345), .A1(net_3293), .B1(net_554) );
AOI21_X2 inst_7658 ( .B2(net_3439), .ZN(net_3379), .A(net_3213), .B1(net_1221) );
CLKBUF_X2 inst_11463 ( .A(net_9268), .Z(net_11425) );
CLKBUF_X2 inst_11381 ( .A(net_11342), .Z(net_11343) );
CLKBUF_X2 inst_12622 ( .A(net_11769), .Z(net_12584) );
CLKBUF_X2 inst_10868 ( .A(net_8838), .Z(net_10830) );
CLKBUF_X2 inst_10570 ( .A(net_10474), .Z(net_10532) );
CLKBUF_X2 inst_10994 ( .A(net_10955), .Z(net_10956) );
CLKBUF_X2 inst_8051 ( .A(net_8012), .Z(net_8013) );
CLKBUF_X2 inst_13915 ( .A(net_13876), .Z(net_13877) );
CLKBUF_X2 inst_8413 ( .A(net_8374), .Z(net_8375) );
NAND2_X2 inst_3932 ( .A2(net_1696), .ZN(net_1366), .A1(net_1365) );
CLKBUF_X2 inst_10203 ( .A(net_10164), .Z(net_10165) );
DFFR_X2 inst_7035 ( .QN(net_6002), .D(net_3199), .CK(net_13221), .RN(x1822) );
CLKBUF_X2 inst_13634 ( .A(net_13595), .Z(net_13596) );
CLKBUF_X2 inst_9224 ( .A(net_9185), .Z(net_9186) );
CLKBUF_X2 inst_11164 ( .A(net_11068), .Z(net_11126) );
CLKBUF_X2 inst_10161 ( .A(net_10122), .Z(net_10123) );
DFF_X2 inst_6295 ( .QN(net_5973), .D(net_1659), .CK(net_8555) );
SDFF_X2 inst_847 ( .Q(net_7027), .D(net_7027), .SE(net_3899), .SI(net_3800), .CK(net_10862) );
NAND3_X2 inst_2720 ( .ZN(net_2455), .A2(net_1803), .A3(net_1578), .A1(net_1347) );
DFF_X1 inst_6577 ( .QN(net_7566), .D(net_5073), .CK(net_13089) );
OAI21_X2 inst_1716 ( .ZN(net_5578), .B1(net_5548), .A(net_4688), .B2(net_3989) );
OAI21_X2 inst_1942 ( .B1(net_5240), .ZN(net_5083), .A(net_4735), .B2(net_3986) );
CLKBUF_X2 inst_11433 ( .A(net_11394), .Z(net_11395) );
CLKBUF_X2 inst_10857 ( .A(net_8936), .Z(net_10819) );
CLKBUF_X2 inst_9788 ( .A(net_8261), .Z(net_9750) );
INV_X2 inst_5950 ( .ZN(net_1113), .A(net_120) );
CLKBUF_X2 inst_13573 ( .A(net_13534), .Z(net_13535) );
CLKBUF_X2 inst_9136 ( .A(net_8810), .Z(net_9098) );
CLKBUF_X2 inst_11429 ( .A(net_11390), .Z(net_11391) );
NAND3_X2 inst_2648 ( .ZN(net_5955), .A3(net_3957), .A2(net_1484), .A1(net_783) );
DFFR_X2 inst_7055 ( .QN(net_5989), .D(net_3136), .CK(net_13220), .RN(x1822) );
CLKBUF_X2 inst_7919 ( .A(net_7880), .Z(net_7881) );
CLKBUF_X2 inst_8372 ( .A(net_8333), .Z(net_8334) );
SDFF_X2 inst_1146 ( .SI(net_6807), .Q(net_6807), .D(net_3808), .SE(net_3729), .CK(net_11301) );
CLKBUF_X2 inst_12947 ( .A(net_12908), .Z(net_12909) );
NAND2_X2 inst_3708 ( .A1(net_6496), .A2(net_1642), .ZN(net_1641) );
CLKBUF_X2 inst_13112 ( .A(net_13073), .Z(net_13074) );
INV_X4 inst_5512 ( .A(net_7265), .ZN(net_2055) );
CLKBUF_X2 inst_12265 ( .A(net_12226), .Z(net_12227) );
CLKBUF_X2 inst_11973 ( .A(net_11934), .Z(net_11935) );
NAND2_X2 inst_4023 ( .A1(net_6798), .A2(net_1651), .ZN(net_1029) );
NAND2_X2 inst_3781 ( .A1(net_6761), .A2(net_1635), .ZN(net_1564) );
NAND2_X2 inst_3673 ( .A1(net_7337), .A2(net_1798), .ZN(net_1784) );
NAND2_X2 inst_3105 ( .A1(net_6615), .A2(net_4899), .ZN(net_4896) );
INV_X4 inst_5162 ( .ZN(net_550), .A(net_549) );
INV_X8 inst_4519 ( .ZN(net_3722), .A(net_3117) );
INV_X4 inst_5349 ( .A(net_6010), .ZN(net_495) );
DFF_X2 inst_6210 ( .QN(net_7384), .D(net_4156), .CK(net_9518) );
CLKBUF_X2 inst_9899 ( .A(net_9860), .Z(net_9861) );
CLKBUF_X2 inst_9081 ( .A(net_8167), .Z(net_9043) );
NAND2_X2 inst_3539 ( .ZN(net_2528), .A2(net_2102), .A1(net_1187) );
NAND2_X2 inst_3552 ( .ZN(net_2515), .A2(net_2048), .A1(net_1782) );
NOR2_X2 inst_2457 ( .A2(net_5924), .ZN(net_3006), .A1(net_603) );
OAI21_X2 inst_1702 ( .B2(net_5908), .ZN(net_5592), .A(net_5215), .B1(net_4080) );
CLKBUF_X2 inst_8307 ( .A(net_8268), .Z(net_8269) );
CLKBUF_X2 inst_10188 ( .A(net_10149), .Z(net_10150) );
SDFF_X2 inst_274 ( .D(net_6399), .SE(net_5799), .SI(net_384), .Q(net_384), .CK(net_13908) );
SDFF_X2 inst_1277 ( .D(net_6388), .SE(net_6052), .SI(net_313), .Q(net_313), .CK(net_13726) );
AOI22_X2 inst_7329 ( .A2(net_3432), .B2(net_3431), .ZN(net_3417), .B1(net_2575), .A1(net_1252) );
NAND3_X2 inst_2817 ( .ZN(net_2281), .A3(net_1530), .A1(net_1323), .A2(net_945) );
CLKBUF_X2 inst_13135 ( .A(net_11160), .Z(net_13097) );
NAND2_X2 inst_4076 ( .A1(net_6937), .A2(net_1654), .ZN(net_976) );
OAI21_X2 inst_2092 ( .B2(net_4487), .ZN(net_4324), .B1(net_4105), .A(net_3668) );
CLKBUF_X2 inst_13436 ( .A(net_13397), .Z(net_13398) );
NAND2_X2 inst_3207 ( .ZN(net_4719), .A2(net_3986), .A1(net_1889) );
NAND2_X2 inst_3143 ( .ZN(net_4820), .A2(net_4153), .A1(net_2138) );
DFFR_X1 inst_7112 ( .QN(net_5859), .D(net_5798), .CK(net_10317), .RN(x1822) );
CLKBUF_X2 inst_11387 ( .A(net_11348), .Z(net_11349) );
NAND3_X2 inst_2696 ( .ZN(net_2696), .A3(net_2576), .A2(net_2436), .A1(net_2270) );
INV_X4 inst_5586 ( .A(net_7571), .ZN(net_1884) );
CLKBUF_X2 inst_14063 ( .A(net_14024), .Z(net_14025) );
CLKBUF_X2 inst_13784 ( .A(net_13745), .Z(net_13746) );
NAND2_X4 inst_2880 ( .ZN(net_3928), .A1(net_3847), .A2(net_574) );
OAI21_X2 inst_1771 ( .B1(net_5446), .ZN(net_5423), .A(net_4702), .B2(net_3989) );
CLKBUF_X2 inst_14402 ( .A(net_8318), .Z(net_14364) );
OAI22_X2 inst_1440 ( .B2(net_5894), .B1(net_4666), .ZN(net_4636), .A2(net_4634), .A1(net_4120) );
CLKBUF_X2 inst_13611 ( .A(net_13572), .Z(net_13573) );
CLKBUF_X2 inst_9415 ( .A(net_9376), .Z(net_9377) );
NAND3_X2 inst_2660 ( .ZN(net_3936), .A3(net_3391), .A2(net_2961), .A1(net_2841) );
CLKBUF_X2 inst_9854 ( .A(net_9172), .Z(net_9816) );
CLKBUF_X2 inst_13734 ( .A(net_9920), .Z(net_13696) );
AND2_X2 inst_7859 ( .ZN(net_1939), .A1(net_1938), .A2(net_1937) );
CLKBUF_X2 inst_13729 ( .A(net_13690), .Z(net_13691) );
NAND2_X2 inst_3355 ( .ZN(net_3535), .A1(net_3534), .A2(net_3226) );
NOR2_X2 inst_2389 ( .ZN(net_4291), .A1(net_4140), .A2(net_4139) );
INV_X2 inst_5912 ( .A(net_7587), .ZN(net_2132) );
CLKBUF_X2 inst_10802 ( .A(net_9130), .Z(net_10764) );
CLKBUF_X2 inst_12148 ( .A(net_11033), .Z(net_12110) );
DFF_X2 inst_6199 ( .QN(net_7533), .D(net_4529), .CK(net_12604) );
CLKBUF_X2 inst_8179 ( .A(net_7868), .Z(net_8141) );
INV_X4 inst_4946 ( .ZN(net_740), .A(net_739) );
OAI21_X2 inst_2148 ( .B1(net_5778), .ZN(net_2796), .A(net_2651), .B2(net_2649) );
DFF_X2 inst_6213 ( .QN(net_7383), .D(net_4158), .CK(net_9934) );
INV_X2 inst_5784 ( .ZN(net_2443), .A(net_2442) );
CLKBUF_X2 inst_13488 ( .A(net_13449), .Z(net_13450) );
CLKBUF_X2 inst_8354 ( .A(net_8128), .Z(net_8316) );
NAND2_X4 inst_2900 ( .A1(net_5891), .ZN(net_3400), .A2(net_538) );
OAI22_X2 inst_1591 ( .B2(net_3200), .A2(net_3196), .ZN(net_3171), .A1(net_3170), .B1(net_533) );
NAND2_X2 inst_3697 ( .ZN(net_1733), .A1(net_1281), .A2(net_1097) );
NAND2_X2 inst_3247 ( .ZN(net_3950), .A2(net_3733), .A1(net_1729) );
CLKBUF_X2 inst_13544 ( .A(net_13505), .Z(net_13506) );
SDFF_X2 inst_379 ( .SI(net_7674), .Q(net_7674), .D(net_4788), .SE(net_3866), .CK(net_13383) );
SDFF_X2 inst_926 ( .Q(net_7135), .D(net_7135), .SE(net_3903), .SI(net_3799), .CK(net_13351) );
CLKBUF_X2 inst_12348 ( .A(net_12309), .Z(net_12310) );
INV_X4 inst_5470 ( .A(net_7422), .ZN(net_1989) );
CLKBUF_X2 inst_10997 ( .A(net_8445), .Z(net_10959) );
CLKBUF_X2 inst_8312 ( .A(net_8257), .Z(net_8274) );
AND2_X4 inst_7827 ( .ZN(net_3113), .A2(net_3051), .A1(net_1243) );
CLKBUF_X2 inst_12856 ( .A(net_12817), .Z(net_12818) );
NAND3_X4 inst_2570 ( .A3(net_5889), .ZN(net_1819), .A2(net_1657), .A1(net_1656) );
NAND2_X2 inst_4153 ( .A2(net_1222), .ZN(net_1064), .A1(net_341) );
CLKBUF_X2 inst_13586 ( .A(net_11495), .Z(net_13548) );
CLKBUF_X2 inst_8684 ( .A(net_8645), .Z(net_8646) );
CLKBUF_X2 inst_10624 ( .A(net_10585), .Z(net_10586) );
INV_X4 inst_4960 ( .ZN(net_1172), .A(net_720) );
CLKBUF_X2 inst_14205 ( .A(net_13378), .Z(net_14167) );
CLKBUF_X2 inst_9098 ( .A(net_8426), .Z(net_9060) );
NAND2_X2 inst_3719 ( .A1(net_6771), .A2(net_1635), .ZN(net_1627) );
NAND2_X2 inst_3646 ( .A1(net_7067), .ZN(net_1817), .A2(net_791) );
SDFF_X2 inst_891 ( .Q(net_7122), .D(net_7122), .SE(net_3888), .SI(net_3803), .CK(net_11587) );
NAND2_X2 inst_4095 ( .A1(net_7199), .A2(net_1648), .ZN(net_957) );
CLKBUF_X2 inst_9479 ( .A(net_9440), .Z(net_9441) );
XNOR2_X2 inst_74 ( .ZN(net_1695), .B(net_1694), .A(net_768) );
CLKBUF_X2 inst_13357 ( .A(net_13318), .Z(net_13319) );
NOR2_X4 inst_2244 ( .ZN(net_5642), .A1(net_5488), .A2(net_4454) );
INV_X4 inst_5682 ( .A(net_6106), .ZN(net_3625) );
SDFF_X2 inst_288 ( .D(net_6396), .SE(net_6052), .SI(net_321), .Q(net_321), .CK(net_13826) );
CLKBUF_X2 inst_14414 ( .A(net_14375), .Z(net_14376) );
CLKBUF_X2 inst_11435 ( .A(net_11396), .Z(net_11397) );
NAND2_X2 inst_3284 ( .ZN(net_3678), .A1(net_3677), .A2(net_3231) );
CLKBUF_X2 inst_11729 ( .A(net_8447), .Z(net_11691) );
AOI22_X2 inst_7263 ( .B1(net_6954), .A1(net_6922), .A2(net_5298), .B2(net_5297), .ZN(net_5291) );
CLKBUF_X2 inst_14265 ( .A(net_14226), .Z(net_14227) );
SDFF_X2 inst_1298 ( .D(net_6387), .SE(net_6051), .SI(net_305), .Q(net_305), .CK(net_13723) );
INV_X8 inst_4512 ( .ZN(net_3891), .A(net_3163) );
INV_X4 inst_5648 ( .A(net_7381), .ZN(net_602) );
INV_X2 inst_5719 ( .ZN(net_4247), .A(net_4115) );
CLKBUF_X2 inst_9147 ( .A(net_8167), .Z(net_9109) );
CLKBUF_X2 inst_12032 ( .A(net_10030), .Z(net_11994) );
CLKBUF_X2 inst_8241 ( .A(net_8202), .Z(net_8203) );
DFF_X1 inst_6499 ( .QN(net_7421), .D(net_5534), .CK(net_12631) );
CLKBUF_X2 inst_8483 ( .A(net_8444), .Z(net_8445) );
SDFF_X2 inst_372 ( .SI(net_7644), .Q(net_7644), .D(net_4786), .SE(net_3867), .CK(net_7988) );
AOI22_X2 inst_7388 ( .A2(net_5916), .B2(net_2957), .ZN(net_2932), .B1(net_2931), .A1(net_712) );
CLKBUF_X2 inst_8031 ( .A(net_7990), .Z(net_7993) );
CLKBUF_X2 inst_13619 ( .A(net_13580), .Z(net_13581) );
CLKBUF_X2 inst_11234 ( .A(net_11195), .Z(net_11196) );
INV_X2 inst_5991 ( .A(net_6027), .ZN(net_2610) );
CLKBUF_X2 inst_9218 ( .A(net_9179), .Z(net_9180) );
CLKBUF_X2 inst_8512 ( .A(net_8188), .Z(net_8474) );
DFFS_X2 inst_6949 ( .QN(net_6407), .D(net_2722), .CK(net_14412), .SN(x1822) );
INV_X2 inst_5709 ( .ZN(net_4309), .A(net_4215) );
CLKBUF_X2 inst_11401 ( .A(net_11362), .Z(net_11363) );
INV_X2 inst_5835 ( .A(net_1149), .ZN(net_874) );
CLKBUF_X2 inst_11128 ( .A(net_11089), .Z(net_11090) );
NOR2_X2 inst_2397 ( .A1(net_5778), .ZN(net_3931), .A2(net_275) );
OAI21_X2 inst_1775 ( .B1(net_5438), .ZN(net_5419), .A(net_4698), .B2(net_3989) );
INV_X4 inst_5335 ( .A(net_6165), .ZN(net_3125) );
DFF_X2 inst_6223 ( .QN(net_7097), .D(net_3725), .CK(net_9714) );
CLKBUF_X2 inst_12802 ( .A(net_12763), .Z(net_12764) );
CLKBUF_X2 inst_13539 ( .A(net_13500), .Z(net_13501) );
SDFF_X2 inst_1172 ( .SI(net_6943), .Q(net_6943), .D(net_3831), .SE(net_3741), .CK(net_11693) );
CLKBUF_X2 inst_9709 ( .A(net_9670), .Z(net_9671) );
SDFF_X2 inst_1090 ( .SI(net_6929), .Q(net_6929), .D(net_3799), .SE(net_3741), .CK(net_8919) );
CLKBUF_X2 inst_9088 ( .A(net_8891), .Z(net_9050) );
NAND2_X2 inst_3903 ( .A1(net_6706), .A2(net_1497), .ZN(net_1407) );
NOR2_X2 inst_2372 ( .ZN(net_5213), .A2(net_4613), .A1(net_4444) );
AOI222_X2 inst_7467 ( .A2(net_2204), .B2(net_2202), .C2(net_2200), .ZN(net_2183), .A1(net_2182), .B1(net_2181), .C1(net_2180) );
CLKBUF_X2 inst_13454 ( .A(net_13415), .Z(net_13416) );
NAND3_X2 inst_2575 ( .ZN(net_5764), .A1(net_5659), .A2(net_5283), .A3(net_4233) );
INV_X4 inst_5007 ( .A(net_7816), .ZN(net_3780) );
CLKBUF_X2 inst_10923 ( .A(net_10884), .Z(net_10885) );
SDFF_X2 inst_1239 ( .SI(net_6533), .Q(net_6533), .D(net_3811), .SE(net_3755), .CK(net_8613) );
CLKBUF_X2 inst_13521 ( .A(net_12306), .Z(net_13483) );
CLKBUF_X2 inst_12496 ( .A(net_12457), .Z(net_12458) );
INV_X4 inst_5655 ( .A(net_6028), .ZN(net_462) );
CLKBUF_X2 inst_11874 ( .A(net_10744), .Z(net_11836) );
CLKBUF_X2 inst_8991 ( .A(net_8952), .Z(net_8953) );
INV_X2 inst_5874 ( .ZN(net_413), .A(x1034) );
CLKBUF_X2 inst_13832 ( .A(net_13793), .Z(net_13794) );
CLKBUF_X2 inst_14068 ( .A(net_14029), .Z(net_14030) );
NAND2_X2 inst_3126 ( .ZN(net_4837), .A2(net_4153), .A1(net_2198) );
DFFR_X2 inst_7094 ( .QN(net_6421), .D(net_2738), .CK(net_10236), .RN(x1822) );
CLKBUF_X2 inst_12547 ( .A(net_12508), .Z(net_12509) );
CLKBUF_X2 inst_11319 ( .A(net_10412), .Z(net_11281) );
SDFF_X2 inst_503 ( .Q(net_7109), .D(net_7109), .SI(net_3894), .SE(net_3888), .CK(net_10503) );
CLKBUF_X2 inst_8028 ( .A(net_7989), .Z(net_7990) );
CLKBUF_X2 inst_12107 ( .A(net_12068), .Z(net_12069) );
CLKBUF_X2 inst_8770 ( .A(net_8731), .Z(net_8732) );
CLKBUF_X2 inst_8556 ( .A(net_8366), .Z(net_8518) );
CLKBUF_X2 inst_14445 ( .A(net_14406), .Z(net_14407) );
CLKBUF_X2 inst_8724 ( .A(net_8685), .Z(net_8686) );
INV_X4 inst_5340 ( .A(net_7565), .ZN(net_1902) );
CLKBUF_X2 inst_8300 ( .A(net_8261), .Z(net_8262) );
CLKBUF_X2 inst_13235 ( .A(net_13196), .Z(net_13197) );
CLKBUF_X2 inst_10580 ( .A(net_10541), .Z(net_10542) );
CLKBUF_X2 inst_8907 ( .A(net_8844), .Z(net_8869) );
NAND2_X2 inst_3193 ( .ZN(net_4733), .A2(net_3986), .A1(net_1913) );
OAI21_X2 inst_1936 ( .B1(net_5551), .ZN(net_5109), .A(net_4741), .B2(net_3988) );
DFF_X1 inst_6458 ( .QN(net_6111), .D(net_5601), .CK(net_11173) );
INV_X4 inst_5088 ( .A(net_3150), .ZN(net_733) );
OAI21_X2 inst_2099 ( .B2(net_4403), .ZN(net_4317), .B1(net_4030), .A(net_3494) );
NAND2_X2 inst_4193 ( .ZN(net_1828), .A1(net_652), .A2(net_309) );
NAND2_X2 inst_4069 ( .A1(net_7200), .A2(net_1648), .ZN(net_983) );
CLKBUF_X2 inst_13316 ( .A(net_13277), .Z(net_13278) );
DFFR_X2 inst_7074 ( .D(net_2812), .QN(net_287), .CK(net_12330), .RN(x1822) );
CLKBUF_X2 inst_14200 ( .A(net_10893), .Z(net_14162) );
CLKBUF_X2 inst_12858 ( .A(net_9491), .Z(net_12820) );
SDFF_X2 inst_686 ( .Q(net_6752), .D(net_6752), .SE(net_3815), .SI(net_3790), .CK(net_10914) );
SDFF_X2 inst_1097 ( .SI(net_6795), .Q(net_6795), .D(net_3798), .SE(net_3722), .CK(net_11084) );
INV_X4 inst_5433 ( .A(net_7748), .ZN(net_2650) );
CLKBUF_X2 inst_9871 ( .A(net_8131), .Z(net_9833) );
CLKBUF_X2 inst_11079 ( .A(net_11040), .Z(net_11041) );
INV_X4 inst_4892 ( .A(net_1683), .ZN(net_1045) );
NAND2_X4 inst_2888 ( .ZN(net_4105), .A2(net_3330), .A1(net_2843) );
CLKBUF_X2 inst_9382 ( .A(net_9279), .Z(net_9344) );
DFF_X1 inst_6804 ( .D(net_3749), .CK(net_10424), .Q(x361) );
CLKBUF_X2 inst_12683 ( .A(net_12644), .Z(net_12645) );
CLKBUF_X2 inst_12633 ( .A(net_9488), .Z(net_12595) );
NAND2_X2 inst_3643 ( .ZN(net_2228), .A2(net_1918), .A1(net_1692) );
CLKBUF_X2 inst_12330 ( .A(net_12291), .Z(net_12292) );
CLKBUF_X2 inst_9235 ( .A(net_9196), .Z(net_9197) );
SDFF_X2 inst_967 ( .Q(net_6446), .D(net_6446), .SE(net_3820), .SI(net_3804), .CK(net_8417) );
CLKBUF_X2 inst_13117 ( .A(net_8014), .Z(net_13079) );
CLKBUF_X2 inst_10635 ( .A(net_8279), .Z(net_10597) );
CLKBUF_X2 inst_9075 ( .A(net_9036), .Z(net_9037) );
OAI21_X2 inst_2119 ( .B2(net_3297), .ZN(net_3294), .B1(net_3293), .A(net_3076) );
OAI21_X2 inst_1929 ( .ZN(net_5116), .A(net_4774), .B2(net_3941), .B1(net_1066) );
CLKBUF_X2 inst_12665 ( .A(net_12626), .Z(net_12627) );
NAND2_X2 inst_3391 ( .ZN(net_3766), .A2(net_3366), .A1(net_2883) );
CLKBUF_X2 inst_9422 ( .A(net_8234), .Z(net_9384) );
CLKBUF_X2 inst_8519 ( .A(net_8480), .Z(net_8481) );
CLKBUF_X2 inst_11495 ( .A(net_10673), .Z(net_11457) );
CLKBUF_X2 inst_7863 ( .A(x821), .Z(net_7825) );
CLKBUF_X2 inst_12200 ( .A(net_12161), .Z(net_12162) );
CLKBUF_X2 inst_9025 ( .A(net_8283), .Z(net_8987) );
CLKBUF_X2 inst_12472 ( .A(net_9587), .Z(net_12434) );
OAI21_X2 inst_1794 ( .ZN(net_5396), .A(net_4723), .B2(net_3986), .B1(net_1081) );
CLKBUF_X2 inst_12029 ( .A(net_11990), .Z(net_11991) );
SDFF_X2 inst_1227 ( .SI(net_7221), .Q(net_7221), .D(net_3795), .SE(net_3751), .CK(net_10616) );
NOR2_X2 inst_2324 ( .A2(net_6294), .A1(net_5840), .ZN(net_5817) );
CLKBUF_X2 inst_9443 ( .A(net_8744), .Z(net_9405) );
INV_X2 inst_5856 ( .ZN(net_642), .A(net_641) );
INV_X2 inst_5732 ( .ZN(net_3960), .A(net_3959) );
CLKBUF_X2 inst_8126 ( .A(net_8087), .Z(net_8088) );
NAND2_X2 inst_3047 ( .A1(net_7016), .A2(net_4979), .ZN(net_4960) );
INV_X2 inst_5957 ( .A(net_7665), .ZN(net_1844) );
NAND2_X2 inst_3847 ( .A1(net_6564), .A2(net_1705), .ZN(net_1490) );
NAND2_X4 inst_2897 ( .A1(net_5890), .ZN(net_3404), .A2(net_582) );
NOR2_X2 inst_2529 ( .ZN(net_1652), .A2(net_772), .A1(net_564) );
CLKBUF_X2 inst_11807 ( .A(net_11768), .Z(net_11769) );
OAI21_X2 inst_1787 ( .B1(net_5438), .ZN(net_5404), .A(net_4678), .B2(net_3988) );
INV_X2 inst_5756 ( .A(net_3400), .ZN(net_3326) );
CLKBUF_X2 inst_12581 ( .A(net_12542), .Z(net_12543) );
AOI22_X2 inst_7274 ( .B1(net_7088), .A1(net_7056), .A2(net_5280), .B2(net_5279), .ZN(net_5274) );
CLKBUF_X2 inst_11376 ( .A(net_11337), .Z(net_11338) );
CLKBUF_X2 inst_14290 ( .A(net_14251), .Z(net_14252) );
CLKBUF_X2 inst_9741 ( .A(net_8800), .Z(net_9703) );
CLKBUF_X2 inst_14369 ( .A(net_14330), .Z(net_14331) );
INV_X2 inst_5943 ( .A(net_7321), .ZN(net_1799) );
CLKBUF_X2 inst_9891 ( .A(net_9852), .Z(net_9853) );
OAI22_X2 inst_1540 ( .B1(net_4637), .A1(net_4030), .B2(net_4018), .ZN(net_4015), .A2(net_4014) );
DFF_X2 inst_6310 ( .QN(net_7795), .CK(net_11826), .D(x1580) );
CLKBUF_X2 inst_9493 ( .A(net_9454), .Z(net_9455) );
CLKBUF_X2 inst_9748 ( .A(net_9709), .Z(net_9710) );
NAND2_X2 inst_3536 ( .ZN(net_2531), .A2(net_2167), .A1(net_1477) );
NAND3_X2 inst_2742 ( .ZN(net_2359), .A3(net_1535), .A1(net_1458), .A2(net_947) );
OAI221_X2 inst_1660 ( .C2(net_5894), .ZN(net_4669), .B1(net_4666), .B2(net_4508), .C1(net_4132), .A(net_3626) );
CLKBUF_X2 inst_10113 ( .A(net_10074), .Z(net_10075) );
AOI222_X2 inst_7515 ( .B1(net_7375), .C1(net_7311), .A2(net_2211), .B2(net_2209), .C2(net_2207), .ZN(net_2024), .A1(net_2023) );
NAND2_X1 inst_4375 ( .ZN(net_4352), .A2(net_3859), .A1(net_2019) );
INV_X4 inst_5243 ( .ZN(net_1146), .A(net_447) );
CLKBUF_X2 inst_13416 ( .A(net_13377), .Z(net_13378) );
CLKBUF_X2 inst_12355 ( .A(net_11831), .Z(net_12317) );
SDFF_X2 inst_517 ( .Q(net_6719), .D(net_6719), .SI(net_3898), .SE(net_3871), .CK(net_8379) );
NOR2_X2 inst_2346 ( .ZN(net_5658), .A1(net_5510), .A2(net_4480) );
SDFF_X2 inst_1261 ( .D(net_6389), .SE(net_5799), .SI(net_374), .Q(net_374), .CK(net_13887) );
INV_X4 inst_5368 ( .A(net_7720), .ZN(net_916) );
CLKBUF_X2 inst_8967 ( .A(net_8928), .Z(net_8929) );
CLKBUF_X2 inst_12486 ( .A(net_12447), .Z(net_12448) );
CLKBUF_X2 inst_12123 ( .A(net_9910), .Z(net_12085) );
CLKBUF_X2 inst_10220 ( .A(net_10181), .Z(net_10182) );
INV_X16 inst_6130 ( .ZN(net_4436), .A(net_3840) );
INV_X4 inst_5382 ( .A(net_6001), .ZN(net_452) );
CLKBUF_X2 inst_13653 ( .A(net_13614), .Z(net_13615) );
SDFF_X2 inst_310 ( .D(net_6393), .SE(net_5801), .SI(net_338), .Q(net_338), .CK(net_13903) );
CLKBUF_X2 inst_8900 ( .A(net_8861), .Z(net_8862) );
CLKBUF_X2 inst_12291 ( .A(net_12252), .Z(net_12253) );
AOI22_X2 inst_7250 ( .B1(net_6818), .A1(net_6786), .A2(net_5316), .B2(net_5315), .ZN(net_5310) );
CLKBUF_X2 inst_9746 ( .A(net_8613), .Z(net_9708) );
AOI22_X2 inst_7363 ( .A2(net_2991), .B2(net_2990), .ZN(net_2975), .A1(net_1202), .B1(net_1201) );
SDFF_X2 inst_1005 ( .SI(net_7802), .Q(net_6465), .D(net_6465), .SE(net_3904), .CK(net_11249) );
DFFR_X2 inst_6979 ( .D(net_3744), .QN(net_288), .CK(net_12348), .RN(x1822) );
OAI22_X2 inst_1580 ( .ZN(net_3202), .A1(net_3201), .B2(net_3200), .A2(net_3193), .B1(net_605) );
NAND3_X2 inst_2688 ( .ZN(net_3157), .A2(net_2939), .A3(net_2845), .A1(net_2778) );
OAI21_X2 inst_1842 ( .B1(net_5357), .ZN(net_5330), .A(net_4370), .B2(net_3853) );
HA_X1 inst_6172 ( .S(net_1691), .CO(net_887), .A(net_886), .B(net_797) );
INV_X4 inst_5592 ( .A(net_7554), .ZN(net_2148) );
NOR2_X2 inst_2351 ( .ZN(net_5653), .A1(net_5505), .A2(net_4472) );
CLKBUF_X2 inst_8067 ( .A(net_8028), .Z(net_8029) );
CLKBUF_X2 inst_12302 ( .A(net_11776), .Z(net_12264) );
INV_X4 inst_5125 ( .A(net_2968), .ZN(net_591) );
OAI21_X2 inst_1853 ( .B1(net_5335), .ZN(net_5319), .A(net_4360), .B2(net_3853) );
AOI222_X2 inst_7534 ( .B2(net_2135), .C2(net_2133), .A2(net_1910), .ZN(net_1900), .A1(net_1899), .B1(net_1898), .C1(net_1897) );
AOI222_X2 inst_7576 ( .A1(net_7539), .ZN(net_5208), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_371), .C2(net_369) );
CLKBUF_X2 inst_11101 ( .A(net_8813), .Z(net_11063) );
SDFF_X2 inst_264 ( .Q(net_6370), .SI(net_6369), .D(net_3568), .SE(net_392), .CK(net_14078) );
NAND2_X2 inst_3703 ( .A1(net_7105), .ZN(net_1676), .A2(net_1675) );
DFF_X1 inst_6737 ( .QN(net_7348), .D(net_4858), .CK(net_12695) );
SDFFR_X2 inst_1333 ( .SI(net_7740), .Q(net_7740), .D(net_4596), .SE(net_3931), .CK(net_13199), .RN(x1822) );
NAND2_X2 inst_3710 ( .A1(net_7167), .ZN(net_1638), .A2(net_1637) );
CLKBUF_X2 inst_12613 ( .A(net_12574), .Z(net_12575) );
NAND2_X2 inst_3953 ( .A1(net_6570), .A2(net_1705), .ZN(net_1332) );
AOI22_X2 inst_7315 ( .B1(net_6676), .A1(net_6644), .A2(net_5139), .B2(net_5138), .ZN(net_5124) );
OAI22_X2 inst_1551 ( .B2(net_3405), .A2(net_3360), .ZN(net_3354), .A1(net_717), .B1(net_444) );
SDFF_X2 inst_1260 ( .D(net_6389), .SE(net_5800), .SI(net_354), .Q(net_354), .CK(net_13809) );
CLKBUF_X2 inst_9579 ( .A(net_9540), .Z(net_9541) );
SDFF_X2 inst_1088 ( .SI(net_7071), .Q(net_7071), .D(net_3813), .SE(net_3742), .CK(net_10830) );
DFF_X1 inst_6490 ( .QN(net_7402), .D(net_5560), .CK(net_12506) );
CLKBUF_X2 inst_13200 ( .A(net_10121), .Z(net_13162) );
CLKBUF_X2 inst_10190 ( .A(net_10151), .Z(net_10152) );
CLKBUF_X2 inst_8692 ( .A(net_8653), .Z(net_8654) );
CLKBUF_X2 inst_11672 ( .A(net_9797), .Z(net_11634) );
NAND2_X2 inst_3332 ( .ZN(net_3582), .A1(net_3581), .A2(net_3228) );
CLKBUF_X2 inst_7885 ( .A(net_7829), .Z(net_7847) );
CLKBUF_X2 inst_13165 ( .A(net_13126), .Z(net_13127) );
INV_X4 inst_4898 ( .A(net_3805), .ZN(net_3133) );
NAND3_X2 inst_2717 ( .ZN(net_2459), .A2(net_1809), .A3(net_1585), .A1(net_1394) );
INV_X2 inst_5844 ( .A(net_1150), .ZN(net_741) );
CLKBUF_X2 inst_13142 ( .A(net_13103), .Z(net_13104) );
CLKBUF_X2 inst_8781 ( .A(net_8159), .Z(net_8743) );
DFF_X1 inst_6433 ( .QN(net_6076), .D(net_5737), .CK(net_8446) );
CLKBUF_X2 inst_13836 ( .A(net_8943), .Z(net_13798) );
NAND2_X2 inst_4176 ( .A2(net_7093), .ZN(net_915), .A1(net_569) );
SDFF_X2 inst_129 ( .Q(net_6192), .SI(net_6191), .D(net_3918), .SE(net_392), .CK(net_13746) );
NAND3_X2 inst_2740 ( .ZN(net_2361), .A3(net_1629), .A1(net_1473), .A2(net_1035) );
OAI21_X2 inst_1754 ( .ZN(net_5449), .B1(net_5448), .A(net_4671), .B2(net_3993) );
CLKBUF_X2 inst_12941 ( .A(net_12902), .Z(net_12903) );
CLKBUF_X2 inst_9922 ( .A(net_9883), .Z(net_9884) );
DFFR_X2 inst_6974 ( .QN(net_7788), .D(net_3995), .CK(net_10194), .RN(x1822) );
CLKBUF_X2 inst_12955 ( .A(net_12916), .Z(net_12917) );
NAND2_X2 inst_2931 ( .ZN(net_5520), .A1(net_4993), .A2(net_4992) );
INV_X4 inst_4768 ( .ZN(net_2431), .A(net_1933) );
AOI211_X2 inst_7789 ( .ZN(net_2621), .C2(net_2616), .C1(net_1973), .B(net_1040), .A(x149) );
NAND3_X2 inst_2727 ( .ZN(net_2374), .A3(net_1633), .A1(net_1457), .A2(net_1029) );
NOR2_X2 inst_2530 ( .ZN(net_3982), .A1(net_772), .A2(net_409) );
CLKBUF_X2 inst_7974 ( .A(net_7854), .Z(net_7936) );
OAI22_X2 inst_1503 ( .B1(net_4660), .A1(net_4105), .B2(net_4095), .ZN(net_4092), .A2(net_4091) );
CLKBUF_X2 inst_12234 ( .A(net_10508), .Z(net_12196) );
CLKBUF_X2 inst_8848 ( .A(net_8718), .Z(net_8810) );
INV_X4 inst_5656 ( .A(net_6082), .ZN(net_3542) );
DFF_X2 inst_6305 ( .Q(net_6381), .D(net_6380), .CK(net_13839) );
CLKBUF_X2 inst_7874 ( .A(net_7835), .Z(net_7836) );
SDFF_X2 inst_777 ( .SI(net_6905), .Q(net_6905), .D(net_3812), .SE(net_3781), .CK(net_11460) );
CLKBUF_X2 inst_8317 ( .A(net_8278), .Z(net_8279) );
NAND2_X2 inst_3802 ( .A1(net_6629), .A2(net_1624), .ZN(net_1543) );
HA_X1 inst_6164 ( .S(net_1712), .CO(net_1711), .B(net_1225), .A(net_905) );
CLKBUF_X2 inst_14175 ( .A(net_14136), .Z(net_14137) );
CLKBUF_X2 inst_12926 ( .A(net_12887), .Z(net_12888) );
INV_X4 inst_5016 ( .A(net_7800), .ZN(net_3883) );
CLKBUF_X2 inst_10276 ( .A(net_10237), .Z(net_10238) );
CLKBUF_X2 inst_11094 ( .A(net_11055), .Z(net_11056) );
CLKBUF_X2 inst_10718 ( .A(net_10679), .Z(net_10680) );
SDFF_X2 inst_933 ( .SI(net_7175), .Q(net_7175), .SE(net_3819), .D(net_3812), .CK(net_12152) );
DFFR_X2 inst_7000 ( .QN(net_7717), .D(net_3352), .CK(net_10747), .RN(x1822) );
CLKBUF_X2 inst_9983 ( .A(net_9944), .Z(net_9945) );
NAND2_X2 inst_3724 ( .A1(net_7030), .A2(net_1975), .ZN(net_1621) );
CLKBUF_X2 inst_14393 ( .A(net_14354), .Z(net_14355) );
CLKBUF_X2 inst_14138 ( .A(net_14099), .Z(net_14100) );
CLKBUF_X2 inst_13902 ( .A(net_13863), .Z(net_13864) );
CLKBUF_X2 inst_14362 ( .A(net_14323), .Z(net_14324) );
CLKBUF_X2 inst_10509 ( .A(net_10470), .Z(net_10471) );
SDFF_X2 inst_1013 ( .SI(net_6507), .Q(net_6507), .SE(net_3889), .D(net_3784), .CK(net_8767) );
INV_X16 inst_6146 ( .ZN(net_1705), .A(net_698) );
CLKBUF_X2 inst_13978 ( .A(net_13939), .Z(net_13940) );
CLKBUF_X2 inst_11909 ( .A(net_11870), .Z(net_11871) );
NAND2_X2 inst_3613 ( .ZN(net_2269), .A2(net_1934), .A1(net_1302) );
INV_X4 inst_4965 ( .ZN(net_905), .A(net_715) );
CLKBUF_X2 inst_13039 ( .A(net_9980), .Z(net_13001) );
CLKBUF_X2 inst_9439 ( .A(net_9400), .Z(net_9401) );
CLKBUF_X2 inst_11158 ( .A(net_11119), .Z(net_11120) );
NOR2_X2 inst_2354 ( .ZN(net_5650), .A1(net_5502), .A2(net_4469) );
CLKBUF_X2 inst_9447 ( .A(net_9408), .Z(net_9409) );
CLKBUF_X2 inst_8735 ( .A(net_8163), .Z(net_8697) );
AND4_X4 inst_7790 ( .ZN(net_2385), .A1(net_2384), .A4(net_1835), .A2(net_1668), .A3(net_1045) );
CLKBUF_X2 inst_14054 ( .A(net_14015), .Z(net_14016) );
CLKBUF_X2 inst_12870 ( .A(net_12831), .Z(net_12832) );
CLKBUF_X2 inst_8481 ( .A(net_8314), .Z(net_8443) );
CLKBUF_X2 inst_10729 ( .A(net_8698), .Z(net_10691) );
NAND2_X2 inst_3515 ( .ZN(net_2552), .A2(net_2145), .A1(net_1369) );
SDFF_X2 inst_124 ( .Q(net_6198), .SI(net_6197), .D(net_3372), .SE(net_392), .CK(net_14246) );
CLKBUF_X2 inst_13315 ( .A(net_13276), .Z(net_13277) );
CLKBUF_X2 inst_12316 ( .A(net_12277), .Z(net_12278) );
CLKBUF_X2 inst_10883 ( .A(net_10844), .Z(net_10845) );
CLKBUF_X2 inst_10982 ( .A(net_10943), .Z(net_10944) );
NAND2_X2 inst_3869 ( .A2(net_1696), .ZN(net_1460), .A1(net_1459) );
NAND2_X2 inst_3488 ( .ZN(net_2656), .A1(net_2655), .A2(net_2654) );
CLKBUF_X2 inst_13849 ( .A(net_12274), .Z(net_13811) );
CLKBUF_X2 inst_12531 ( .A(net_12492), .Z(net_12493) );
CLKBUF_X2 inst_11593 ( .A(net_11554), .Z(net_11555) );
SDFF_X2 inst_1270 ( .D(net_7802), .SI(net_6529), .Q(net_6529), .SE(net_3755), .CK(net_11209) );
DFF_X2 inst_6332 ( .QN(net_7823), .CK(net_8238), .D(x1351) );
NAND2_X2 inst_3448 ( .A1(net_7761), .ZN(net_2974), .A2(net_2973) );
CLKBUF_X2 inst_8001 ( .A(net_7946), .Z(net_7963) );
INV_X2 inst_6088 ( .A(net_7619), .ZN(net_1188) );
CLKBUF_X2 inst_12689 ( .A(net_11168), .Z(net_12651) );
INV_X8 inst_4563 ( .ZN(net_1654), .A(net_478) );
CLKBUF_X2 inst_10123 ( .A(net_10084), .Z(net_10085) );
CLKBUF_X2 inst_13032 ( .A(net_12993), .Z(net_12994) );
INV_X4 inst_5504 ( .A(net_7404), .ZN(net_2125) );
INV_X4 inst_5361 ( .A(net_5997), .ZN(net_469) );
CLKBUF_X2 inst_12489 ( .A(net_12450), .Z(net_12451) );
CLKBUF_X2 inst_13049 ( .A(net_13010), .Z(net_13011) );
AOI22_X2 inst_7453 ( .A2(net_2934), .B2(net_2664), .ZN(net_711), .A1(net_710), .B1(net_709) );
OAI22_X2 inst_1519 ( .B1(net_4650), .B2(net_4458), .A1(net_4080), .A2(net_4078), .ZN(net_4059) );
CLKBUF_X1 inst_7243 ( .A(x130657), .Z(x145) );
OAI21_X2 inst_2156 ( .ZN(net_2688), .B1(net_2687), .A(net_2619), .B2(net_2422) );
CLKBUF_X2 inst_13389 ( .A(net_13350), .Z(net_13351) );
CLKBUF_X2 inst_9936 ( .A(net_9897), .Z(net_9898) );
CLKBUF_X2 inst_8461 ( .A(net_8422), .Z(net_8423) );
INV_X4 inst_4989 ( .A(net_7093), .ZN(net_1152) );
CLKBUF_X2 inst_12142 ( .A(net_12103), .Z(net_12104) );
NAND2_X1 inst_4324 ( .ZN(net_4540), .A2(net_3870), .A1(net_1344) );
INV_X2 inst_5746 ( .ZN(net_3718), .A(net_3415) );
INV_X4 inst_5417 ( .ZN(net_505), .A(net_298) );
INV_X4 inst_5597 ( .A(net_6960), .ZN(net_829) );
DFFR_X2 inst_7009 ( .D(net_3279), .QN(net_267), .CK(net_12342), .RN(x1822) );
CLKBUF_X2 inst_12705 ( .A(net_12666), .Z(net_12667) );
NOR2_X2 inst_2515 ( .A2(net_3238), .ZN(net_1139), .A1(net_1138) );
CLKBUF_X2 inst_8531 ( .A(net_8492), .Z(net_8493) );
CLKBUF_X2 inst_12244 ( .A(net_12056), .Z(net_12206) );
OAI22_X2 inst_1491 ( .B1(net_4666), .A1(net_4132), .B2(net_4122), .ZN(net_4119), .A2(net_4118) );
CLKBUF_X2 inst_8070 ( .A(net_8031), .Z(net_8032) );
CLKBUF_X2 inst_12747 ( .A(net_12708), .Z(net_12709) );
CLKBUF_X2 inst_8703 ( .A(net_8664), .Z(net_8665) );
CLKBUF_X2 inst_12900 ( .A(net_7966), .Z(net_12862) );
XNOR2_X2 inst_117 ( .ZN(net_5863), .A(net_816), .B(net_791) );
NAND3_X2 inst_2676 ( .ZN(net_3460), .A3(net_3306), .A1(net_2966), .A2(net_2946) );
INV_X4 inst_5172 ( .A(net_820), .ZN(net_535) );
CLKBUF_X2 inst_8566 ( .A(net_8527), .Z(net_8528) );
SDFF_X2 inst_154 ( .Q(net_6224), .SI(net_6223), .SE(net_392), .D(net_130), .CK(net_14088) );
CLKBUF_X2 inst_13104 ( .A(net_13065), .Z(net_13066) );
NAND2_X2 inst_4106 ( .A1(net_7208), .A2(net_1648), .ZN(net_946) );
CLKBUF_X2 inst_9794 ( .A(net_9755), .Z(net_9756) );
SDFF_X2 inst_465 ( .Q(net_6879), .D(net_6879), .SE(net_3901), .SI(net_3897), .CK(net_11758) );
INV_X2 inst_6057 ( .ZN(net_1115), .A(net_122) );
CLKBUF_X2 inst_11367 ( .A(net_11328), .Z(net_11329) );
NOR2_X2 inst_2304 ( .A2(net_6210), .A1(net_5843), .ZN(net_5837) );
CLKBUF_X2 inst_12325 ( .A(net_8021), .Z(net_12287) );
CLKBUF_X2 inst_10078 ( .A(net_8387), .Z(net_10040) );
CLKBUF_X2 inst_13427 ( .A(net_13388), .Z(net_13389) );
CLKBUF_X2 inst_10368 ( .A(net_10152), .Z(net_10330) );
NAND2_X1 inst_4240 ( .ZN(net_4687), .A2(net_3989), .A1(net_2110) );
CLKBUF_X2 inst_11701 ( .A(net_11662), .Z(net_11663) );
CLKBUF_X2 inst_10813 ( .A(net_10774), .Z(net_10775) );
NOR4_X2 inst_2173 ( .ZN(net_3248), .A4(net_3124), .A1(net_2642), .A3(net_2482), .A2(net_824) );
CLKBUF_X2 inst_12570 ( .A(net_12531), .Z(net_12532) );
OAI21_X2 inst_1790 ( .B1(net_5432), .ZN(net_5401), .A(net_4675), .B2(net_3988) );
DFF_X1 inst_6621 ( .QN(net_7582), .D(net_5386), .CK(net_10302) );
DFFR_X2 inst_7048 ( .QN(net_6017), .D(net_3126), .CK(net_8592), .RN(x1822) );
NAND2_X2 inst_3214 ( .ZN(net_4712), .A2(net_3986), .A1(net_1875) );
CLKBUF_X2 inst_10989 ( .A(net_10552), .Z(net_10951) );
CLKBUF_X2 inst_12940 ( .A(net_8711), .Z(net_12902) );
OAI21_X2 inst_1905 ( .B1(net_5359), .ZN(net_5164), .A(net_4764), .B2(net_3941) );
DFF_X1 inst_6355 ( .QN(net_6203), .D(net_5829), .CK(net_13700) );
CLKBUF_X2 inst_11917 ( .A(net_11878), .Z(net_11879) );
CLKBUF_X2 inst_13982 ( .A(net_13943), .Z(net_13944) );
NOR2_X4 inst_2264 ( .ZN(net_5622), .A1(net_5467), .A2(net_4419) );
SDFF_X2 inst_243 ( .Q(net_6351), .SI(net_6350), .D(net_3611), .SE(net_392), .CK(net_13941) );
OR2_X4 inst_1378 ( .ZN(net_3443), .A2(net_3246), .A1(net_2605) );
CLKBUF_X2 inst_14156 ( .A(net_14117), .Z(net_14118) );
CLKBUF_X2 inst_14049 ( .A(net_14010), .Z(net_14011) );
NAND3_X2 inst_2697 ( .ZN(net_2695), .A3(net_2574), .A2(net_2434), .A1(net_2269) );
CLKBUF_X2 inst_10196 ( .A(net_9991), .Z(net_10158) );
XNOR2_X2 inst_15 ( .ZN(net_2639), .B(net_2638), .A(net_2485) );
NAND2_X2 inst_3747 ( .A1(net_6904), .A2(net_1639), .ZN(net_1598) );
CLKBUF_X2 inst_8189 ( .A(net_8150), .Z(net_8151) );
CLKBUF_X2 inst_11902 ( .A(net_11863), .Z(net_11864) );
AOI22_X2 inst_7281 ( .B1(net_7218), .A1(net_7186), .ZN(net_5245), .A2(net_5244), .B2(net_5243) );
NAND2_X2 inst_3496 ( .A2(net_2644), .ZN(net_2623), .A1(net_412) );
DFF_X1 inst_6704 ( .QN(net_7287), .D(net_5371), .CK(net_10163) );
CLKBUF_X2 inst_9501 ( .A(net_9462), .Z(net_9463) );
CLKBUF_X2 inst_13082 ( .A(net_13043), .Z(net_13044) );
CLKBUF_X2 inst_9830 ( .A(net_9791), .Z(net_9792) );
CLKBUF_X2 inst_13642 ( .A(net_13603), .Z(net_13604) );
CLKBUF_X2 inst_12020 ( .A(net_11981), .Z(net_11982) );
CLKBUF_X2 inst_8799 ( .A(net_8760), .Z(net_8761) );
OAI21_X2 inst_2123 ( .B1(net_3268), .B2(net_3087), .ZN(net_3064), .A(net_2912) );
NAND2_X2 inst_3229 ( .ZN(net_4526), .A2(net_4293), .A1(net_1733) );
INV_X4 inst_4918 ( .A(net_3794), .ZN(net_3201) );
CLKBUF_X2 inst_8615 ( .A(net_8000), .Z(net_8577) );
NAND2_X2 inst_4135 ( .A1(net_1150), .ZN(net_935), .A2(net_866) );
OR2_X4 inst_1369 ( .ZN(net_3975), .A2(net_3738), .A1(net_3230) );
NAND2_X2 inst_3988 ( .A1(net_6713), .A2(net_1497), .ZN(net_1276) );
SDFF_X2 inst_349 ( .SI(net_7677), .Q(net_7677), .D(net_4802), .SE(net_3866), .CK(net_10281) );
CLKBUF_X2 inst_14145 ( .A(net_14106), .Z(net_14107) );
CLKBUF_X2 inst_10690 ( .A(net_10651), .Z(net_10652) );
DFF_X1 inst_6548 ( .Q(net_7773), .D(net_5609), .CK(net_12416) );
CLKBUF_X2 inst_14381 ( .A(net_14096), .Z(net_14343) );
NAND2_X1 inst_4249 ( .ZN(net_4677), .A2(net_3988), .A1(net_2176) );
NAND2_X1 inst_4235 ( .ZN(net_4692), .A2(net_3989), .A1(net_2181) );
CLKBUF_X2 inst_13940 ( .A(net_13901), .Z(net_13902) );
NAND4_X2 inst_2561 ( .A1(net_2299), .ZN(net_1825), .A3(net_1824), .A4(net_1823), .A2(net_1820) );
AOI21_X2 inst_7767 ( .B1(net_7135), .ZN(net_5908), .B2(net_2582), .A(net_2294) );
CLKBUF_X2 inst_13629 ( .A(net_10561), .Z(net_13591) );
CLKBUF_X2 inst_11507 ( .A(net_11468), .Z(net_11469) );
CLKBUF_X2 inst_9570 ( .A(net_9531), .Z(net_9532) );
INV_X2 inst_6024 ( .A(net_7663), .ZN(net_1897) );
CLKBUF_X2 inst_8495 ( .A(net_8456), .Z(net_8457) );
CLKBUF_X2 inst_8974 ( .A(net_8312), .Z(net_8936) );
CLKBUF_X2 inst_8163 ( .A(net_8039), .Z(net_8125) );
CLKBUF_X2 inst_13669 ( .A(net_13630), .Z(net_13631) );
CLKBUF_X2 inst_13257 ( .A(net_13218), .Z(net_13219) );
CLKBUF_X2 inst_9583 ( .A(net_9544), .Z(net_9545) );
NAND2_X1 inst_4226 ( .ZN(net_4701), .A2(net_3989), .A1(net_2203) );
NOR2_X4 inst_2252 ( .ZN(net_5634), .A1(net_5479), .A2(net_4440) );
CLKBUF_X2 inst_12289 ( .A(net_9748), .Z(net_12251) );
CLKBUF_X2 inst_12514 ( .A(net_12475), .Z(net_12476) );
CLKBUF_X2 inst_9222 ( .A(net_9183), .Z(net_9184) );
NAND2_X1 inst_4229 ( .ZN(net_4698), .A2(net_3989), .A1(net_2185) );
CLKBUF_X2 inst_12843 ( .A(net_11881), .Z(net_12805) );
INV_X2 inst_5795 ( .ZN(net_2231), .A(net_2230) );
CLKBUF_X2 inst_12112 ( .A(net_10259), .Z(net_12074) );
CLKBUF_X2 inst_12065 ( .A(net_12026), .Z(net_12027) );
NOR2_X4 inst_2238 ( .ZN(net_5660), .A1(net_5513), .A2(net_4482) );
NAND3_X2 inst_2763 ( .ZN(net_2338), .A3(net_1623), .A1(net_1425), .A2(net_966) );
INV_X4 inst_5207 ( .ZN(net_3001), .A(net_491) );
INV_X8 inst_4543 ( .ZN(net_2581), .A(net_1279) );
INV_X4 inst_5072 ( .A(net_3109), .ZN(net_799) );
CLKBUF_X2 inst_14334 ( .A(net_14295), .Z(net_14296) );
CLKBUF_X2 inst_10301 ( .A(net_8346), .Z(net_10263) );
CLKBUF_X2 inst_14347 ( .A(net_14308), .Z(net_14309) );
NAND2_X2 inst_3151 ( .ZN(net_4812), .A2(net_4153), .A1(net_2121) );
CLKBUF_X2 inst_10554 ( .A(net_10515), .Z(net_10516) );
DFF_X1 inst_6798 ( .D(net_3939), .CK(net_12832), .Q(x620) );
SDFF_X2 inst_761 ( .Q(net_6884), .D(net_6884), .SE(net_3901), .SI(net_3803), .CK(net_11727) );
CLKBUF_X2 inst_13073 ( .A(net_12297), .Z(net_13035) );
CLKBUF_X2 inst_10764 ( .A(net_10725), .Z(net_10726) );
INV_X4 inst_4867 ( .A(net_2705), .ZN(net_1101) );
CLKBUF_X2 inst_13342 ( .A(net_10929), .Z(net_13304) );
NAND2_X1 inst_4436 ( .A1(net_7604), .A2(net_2131), .ZN(net_1378) );
NAND3_X2 inst_2803 ( .ZN(net_2295), .A1(net_1706), .A3(net_1544), .A2(net_950) );
CLKBUF_X2 inst_8180 ( .A(net_8141), .Z(net_8142) );
CLKBUF_X2 inst_13042 ( .A(net_13003), .Z(net_13004) );
NAND2_X2 inst_4120 ( .A2(net_1228), .ZN(net_1108), .A1(net_383) );
INV_X2 inst_5801 ( .ZN(net_1923), .A(net_265) );
CLKBUF_X2 inst_9363 ( .A(net_9324), .Z(net_9325) );
CLKBUF_X2 inst_9211 ( .A(net_9172), .Z(net_9173) );
INV_X4 inst_5525 ( .A(net_6136), .ZN(net_3661) );
DFF_X1 inst_6674 ( .QN(net_7251), .D(net_5155), .CK(net_12802) );
CLKBUF_X2 inst_10003 ( .A(net_8045), .Z(net_9965) );
NOR2_X4 inst_2259 ( .ZN(net_5627), .A1(net_5472), .A2(net_4430) );
INV_X4 inst_5097 ( .A(net_7801), .ZN(net_3814) );
CLKBUF_X2 inst_12935 ( .A(net_12896), .Z(net_12897) );
NAND3_X2 inst_2641 ( .ZN(net_5688), .A1(net_5665), .A2(net_5293), .A3(net_4239) );
DFF_X2 inst_6196 ( .QN(net_6555), .D(net_5042), .CK(net_8815) );
CLKBUF_X2 inst_14314 ( .A(net_10151), .Z(net_14276) );
OAI222_X2 inst_1638 ( .C2(net_4157), .ZN(net_4156), .A2(net_4155), .B2(net_4154), .A1(net_2437), .B1(net_1647), .C1(net_536) );
DFF_X1 inst_6462 ( .QN(net_6131), .D(net_5597), .CK(net_10954) );
CLKBUF_X2 inst_11450 ( .A(net_8072), .Z(net_11412) );
INV_X2 inst_5771 ( .ZN(net_2983), .A(net_2982) );
CLKBUF_X2 inst_9812 ( .A(net_8019), .Z(net_9774) );
NAND2_X2 inst_3220 ( .ZN(net_4706), .A2(net_3986), .A1(net_1872) );
CLKBUF_X2 inst_14101 ( .A(net_13305), .Z(net_14063) );
CLKBUF_X2 inst_12824 ( .A(net_12785), .Z(net_12786) );
CLKBUF_X2 inst_11915 ( .A(net_8003), .Z(net_11877) );
CLKBUF_X2 inst_8177 ( .A(net_8138), .Z(net_8139) );
CLKBUF_X2 inst_12280 ( .A(net_12241), .Z(net_12242) );
CLKBUF_X2 inst_11072 ( .A(net_10794), .Z(net_11034) );
CLKBUF_X2 inst_11983 ( .A(net_11944), .Z(net_11945) );
INV_X4 inst_5354 ( .A(net_6093), .ZN(net_3475) );
DFF_X1 inst_6428 ( .QN(net_6183), .D(net_5742), .CK(net_10673) );
CLKBUF_X2 inst_14221 ( .A(net_14182), .Z(net_14183) );
AOI22_X2 inst_7312 ( .B1(net_6685), .A1(net_6653), .A2(net_5139), .B2(net_5138), .ZN(net_5131) );
INV_X4 inst_5373 ( .A(net_6078), .ZN(net_3575) );
AOI222_X2 inst_7560 ( .A1(net_7548), .ZN(net_5232), .A2(net_1228), .B1(net_1227), .C1(net_1226), .B2(net_380), .C2(net_378) );
INV_X4 inst_4783 ( .ZN(net_2642), .A(net_1660) );
CLKBUF_X2 inst_9047 ( .A(net_9008), .Z(net_9009) );
NAND2_X2 inst_3862 ( .A1(net_7462), .A2(net_1696), .ZN(net_1470) );
DFF_X1 inst_6556 ( .QN(net_7264), .D(net_5162), .CK(net_13009) );
DFF_X1 inst_6532 ( .QN(net_7479), .D(net_5419), .CK(net_9270) );
CLKBUF_X2 inst_10749 ( .A(net_10710), .Z(net_10711) );
CLKBUF_X2 inst_10847 ( .A(net_10808), .Z(net_10809) );
INV_X4 inst_5304 ( .A(net_7428), .ZN(net_1983) );
CLKBUF_X2 inst_14326 ( .A(net_12085), .Z(net_14288) );
CLKBUF_X2 inst_12737 ( .A(net_12698), .Z(net_12699) );
CLKBUF_X2 inst_10482 ( .A(net_9106), .Z(net_10444) );
SDFF_X2 inst_633 ( .SI(net_6645), .Q(net_6645), .SE(net_3851), .D(net_3775), .CK(net_9112) );
CLKBUF_X2 inst_12837 ( .A(net_12641), .Z(net_12799) );
SDFF_X2 inst_524 ( .SI(net_6648), .Q(net_6648), .D(net_3902), .SE(net_3850), .CK(net_12049) );
CLKBUF_X2 inst_13027 ( .A(net_12988), .Z(net_12989) );
NAND2_X2 inst_4060 ( .A1(net_6522), .A2(net_1645), .ZN(net_992) );
XNOR2_X2 inst_104 ( .ZN(net_2253), .A(net_1152), .B(net_1140) );
NOR2_X4 inst_2285 ( .ZN(net_5914), .A2(net_5871), .A1(net_3020) );
CLKBUF_X2 inst_10500 ( .A(net_10461), .Z(net_10462) );
NOR2_X2 inst_2331 ( .A2(net_6287), .A1(net_5843), .ZN(net_5810) );
NAND2_X2 inst_3344 ( .ZN(net_3559), .A1(net_3558), .A2(net_3226) );
INV_X8 inst_4478 ( .ZN(net_4927), .A(net_4263) );
INV_X2 inst_6096 ( .A(net_7632), .ZN(net_1856) );
CLKBUF_X2 inst_11878 ( .A(net_11839), .Z(net_11840) );
CLKBUF_X2 inst_9752 ( .A(net_9446), .Z(net_9714) );
NAND2_X2 inst_3447 ( .A1(net_7765), .ZN(net_3007), .A2(net_3006) );
NOR2_X2 inst_2377 ( .ZN(net_5152), .A2(net_4626), .A1(net_4422) );
NOR2_X2 inst_2522 ( .ZN(net_3862), .A1(net_1728), .A2(net_449) );
CLKBUF_X2 inst_13793 ( .A(net_9269), .Z(net_13755) );
INV_X4 inst_4862 ( .A(net_7799), .ZN(net_3293) );
CLKBUF_X2 inst_11910 ( .A(net_11871), .Z(net_11872) );
INV_X4 inst_4663 ( .ZN(net_5884), .A(net_3923) );
CLKBUF_X2 inst_10360 ( .A(net_10321), .Z(net_10322) );
SDFF_X2 inst_882 ( .Q(net_7112), .D(net_7112), .SE(net_3888), .SI(net_3811), .CK(net_12158) );
CLKBUF_X2 inst_10673 ( .A(net_10504), .Z(net_10635) );
CLKBUF_X2 inst_13935 ( .A(net_13896), .Z(net_13897) );
CLKBUF_X2 inst_7967 ( .A(net_7928), .Z(net_7929) );
CLKBUF_X2 inst_9848 ( .A(net_9809), .Z(net_9810) );
INV_X4 inst_5216 ( .ZN(net_480), .A(net_479) );
CLKBUF_X2 inst_13700 ( .A(net_13661), .Z(net_13662) );
NAND2_X2 inst_2938 ( .ZN(net_5508), .A1(net_4976), .A2(net_4975) );
INV_X4 inst_5257 ( .A(net_842), .ZN(net_434) );
CLKBUF_X2 inst_8011 ( .A(net_7864), .Z(net_7973) );
CLKBUF_X2 inst_9116 ( .A(net_9077), .Z(net_9078) );
CLKBUF_X2 inst_11226 ( .A(net_11187), .Z(net_11188) );
INV_X4 inst_5083 ( .A(net_7809), .ZN(net_3785) );
DFF_X1 inst_6931 ( .D(net_2387), .Q(net_248), .CK(net_8022) );
SDFF_X2 inst_708 ( .SI(net_6780), .Q(net_6780), .SE(net_3816), .D(net_3804), .CK(net_11142) );
SDFFR_X2 inst_1346 ( .D(net_3897), .SE(net_3256), .SI(net_148), .Q(net_148), .CK(net_8550), .RN(x1822) );
NAND2_X2 inst_3523 ( .ZN(net_2544), .A2(net_2112), .A1(net_1410) );
OR2_X4 inst_1374 ( .ZN(net_3447), .A2(net_3248), .A1(net_2595) );
INV_X4 inst_4855 ( .A(net_1240), .ZN(net_1060) );
INV_X2 inst_5811 ( .ZN(net_1106), .A(net_1105) );
CLKBUF_X2 inst_9046 ( .A(net_8458), .Z(net_9008) );
NAND2_X2 inst_3510 ( .ZN(net_2557), .A2(net_2179), .A1(net_1464) );
NOR2_X2 inst_2510 ( .A2(net_3234), .ZN(net_1173), .A1(net_1172) );
INV_X4 inst_5108 ( .A(net_2889), .ZN(net_700) );
DFF_X1 inst_6723 ( .QN(net_7356), .D(net_5333), .CK(net_12982) );
SDFF_X2 inst_1071 ( .SI(net_6532), .Q(net_6532), .D(net_3812), .SE(net_3755), .CK(net_8629) );
NAND2_X1 inst_4277 ( .ZN(net_4591), .A2(net_3867), .A1(net_1914) );
DFF_X1 inst_6421 ( .QN(net_6176), .D(net_5749), .CK(net_8745) );
DFF_X2 inst_6316 ( .QN(net_7793), .CK(net_11822), .D(x1595) );
INV_X4 inst_5291 ( .A(net_7687), .ZN(net_411) );
CLKBUF_X2 inst_11352 ( .A(net_11313), .Z(net_11314) );
CLKBUF_X2 inst_13211 ( .A(net_13172), .Z(net_13173) );
CLKBUF_X2 inst_11548 ( .A(net_11509), .Z(net_11510) );
CLKBUF_X2 inst_14199 ( .A(net_14160), .Z(net_14161) );
OAI21_X2 inst_1994 ( .ZN(net_4522), .B1(net_4521), .B2(net_4518), .A(net_3702) );
CLKBUF_X2 inst_13132 ( .A(net_13093), .Z(net_13094) );
CLKBUF_X2 inst_9192 ( .A(net_9153), .Z(net_9154) );
INV_X4 inst_5298 ( .A(net_7423), .ZN(net_2156) );
CLKBUF_X2 inst_14436 ( .A(net_9512), .Z(net_14398) );
CLKBUF_X2 inst_10108 ( .A(net_10069), .Z(net_10070) );
CLKBUF_X2 inst_13191 ( .A(net_13152), .Z(net_13153) );
CLKBUF_X2 inst_8940 ( .A(net_8901), .Z(net_8902) );
OAI21_X2 inst_2162 ( .ZN(net_2898), .A(net_303), .B2(net_301), .B1(net_279) );
SDFF_X2 inst_392 ( .SI(net_7313), .Q(net_7313), .D(net_4776), .SE(net_3859), .CK(net_12761) );
XNOR2_X2 inst_120 ( .ZN(net_5866), .B(net_1651), .A(net_818) );
DFF_X1 inst_6780 ( .QN(net_6164), .D(net_4322), .CK(net_7945) );
AOI21_X2 inst_7747 ( .B1(net_6606), .ZN(net_4020), .B2(net_2583), .A(net_2288) );
CLKBUF_X2 inst_10917 ( .A(net_8480), .Z(net_10879) );
NAND2_X2 inst_4165 ( .ZN(net_2222), .A1(net_871), .A2(net_459) );
NAND2_X1 inst_4398 ( .A2(net_3297), .ZN(net_3083), .A1(net_3082) );
OAI22_X2 inst_1514 ( .B1(net_4650), .A1(net_4080), .B2(net_4072), .ZN(net_4069), .A2(net_4068) );
NOR2_X4 inst_2272 ( .ZN(net_5614), .A1(net_5459), .A2(net_4408) );
CLKBUF_X2 inst_8361 ( .A(net_7883), .Z(net_8323) );
SDFF_X2 inst_567 ( .D(net_7807), .SI(net_6772), .Q(net_6772), .SE(net_3816), .CK(net_11167) );
OAI22_X2 inst_1608 ( .B2(net_3200), .A2(net_3187), .ZN(net_3112), .A1(net_3111), .B1(net_494) );
NAND2_X2 inst_3200 ( .ZN(net_4726), .A2(net_3986), .A1(net_1861) );
CLKBUF_X2 inst_11631 ( .A(net_7933), .Z(net_11593) );
CLKBUF_X2 inst_9134 ( .A(net_9095), .Z(net_9096) );
OAI22_X2 inst_1484 ( .B1(net_4666), .ZN(net_4136), .A2(net_4135), .B2(net_4134), .A1(net_4132) );
OAI22_X2 inst_1601 ( .B2(net_3200), .A2(net_3193), .ZN(net_3135), .A1(net_827), .B1(net_796) );
NAND2_X2 inst_3526 ( .ZN(net_2541), .A2(net_2094), .A1(net_1384) );
CLKBUF_X2 inst_9010 ( .A(net_8059), .Z(net_8972) );
SDFF_X2 inst_856 ( .SI(net_7041), .Q(net_7041), .SE(net_3818), .D(net_3811), .CK(net_9021) );
INV_X4 inst_5677 ( .A(net_6167), .ZN(net_3562) );

endmodule
