module c1355 (
n43gat,
n190gat,
n99gat,
n78gat,
n85gat,
n232gat,
n211gat,
n226gat,
n155gat,
n176gat,
n162gat,
n64gat,
n230gat,
n92gat,
n228gat,
n127gat,
n22gat,
n1gat,
n113gat,
n183gat,
n148gat,
n29gat,
n197gat,
n134gat,
n204gat,
n218gat,
n227gat,
n8gat,
n169gat,
n225gat,
n36gat,
n57gat,
n231gat,
n106gat,
n233gat,
n50gat,
n15gat,
n71gat,
n120gat,
n229gat,
n141gat,
n1328gat,
n1348gat,
n1338gat,
n1331gat,
n1339gat,
n1344gat,
n1346gat,
n1353gat,
n1337gat,
n1333gat,
n1347gat,
n1340gat,
n1354gat,
n1351gat,
n1355gat,
n1352gat,
n1343gat,
n1329gat,
n1332gat,
n1336gat,
n1324gat,
n1335gat,
n1334gat,
n1349gat,
n1330gat,
n1327gat,
n1341gat,
n1326gat,
n1345gat,
n1342gat,
n1350gat,
n1325gat);

// Start PIs
input n43gat;
input n190gat;
input n99gat;
input n78gat;
input n85gat;
input n232gat;
input n211gat;
input n226gat;
input n155gat;
input n176gat;
input n162gat;
input n64gat;
input n230gat;
input n92gat;
input n228gat;
input n127gat;
input n22gat;
input n1gat;
input n113gat;
input n183gat;
input n148gat;
input n29gat;
input n197gat;
input n134gat;
input n204gat;
input n218gat;
input n227gat;
input n8gat;
input n169gat;
input n225gat;
input n36gat;
input n57gat;
input n231gat;
input n106gat;
input n233gat;
input n50gat;
input n15gat;
input n71gat;
input n120gat;
input n229gat;
input n141gat;

// Start POs
output n1328gat;
output n1348gat;
output n1338gat;
output n1331gat;
output n1339gat;
output n1344gat;
output n1346gat;
output n1353gat;
output n1337gat;
output n1333gat;
output n1347gat;
output n1340gat;
output n1354gat;
output n1351gat;
output n1355gat;
output n1352gat;
output n1343gat;
output n1329gat;
output n1332gat;
output n1336gat;
output n1324gat;
output n1335gat;
output n1334gat;
output n1349gat;
output n1330gat;
output n1327gat;
output n1341gat;
output n1326gat;
output n1345gat;
output n1342gat;
output n1350gat;
output n1325gat;

// Start wires
wire n43gat;
wire net_107;
wire net_47;
wire n190gat;
wire n1328gat;
wire n99gat;
wire net_61;
wire net_137;
wire n1338gat;
wire net_132;
wire net_54;
wire net_105;
wire net_62;
wire net_6;
wire n176gat;
wire net_129;
wire net_119;
wire net_98;
wire net_23;
wire net_117;
wire net_12;
wire net_74;
wire net_53;
wire net_93;
wire n1353gat;
wire net_135;
wire net_130;
wire n1347gat;
wire net_147;
wire net_127;
wire net_14;
wire n1351gat;
wire net_113;
wire net_26;
wire n204gat;
wire net_76;
wire net_101;
wire net_32;
wire net_111;
wire n1332gat;
wire n1329gat;
wire net_90;
wire net_40;
wire net_100;
wire n8gat;
wire net_85;
wire net_69;
wire n225gat;
wire net_124;
wire n57gat;
wire net_141;
wire n1330gat;
wire net_83;
wire net_115;
wire n1345gat;
wire n120gat;
wire net_4;
wire net_95;
wire net_17;
wire net_78;
wire net_27;
wire net_56;
wire net_87;
wire net_0;
wire n232gat;
wire net_35;
wire n211gat;
wire net_22;
wire net_16;
wire n64gat;
wire net_39;
wire n228gat;
wire n92gat;
wire net_144;
wire net_102;
wire net_2;
wire net_59;
wire net_9;
wire net_42;
wire n22gat;
wire net_120;
wire n1337gat;
wire net_109;
wire net_80;
wire net_65;
wire net_50;
wire n183gat;
wire n1354gat;
wire n1340gat;
wire net_96;
wire net_66;
wire net_38;
wire net_44;
wire n197gat;
wire net_136;
wire net_134;
wire net_19;
wire n1352gat;
wire net_89;
wire net_45;
wire net_126;
wire n1336gat;
wire n1324gat;
wire net_34;
wire net_108;
wire n1334gat;
wire n50gat;
wire n15gat;
wire net_63;
wire n1342gat;
wire n229gat;
wire n141gat;
wire n1348gat;
wire net_116;
wire net_30;
wire n78gat;
wire n1331gat;
wire net_91;
wire net_106;
wire net_99;
wire net_24;
wire net_55;
wire net_46;
wire net_140;
wire net_118;
wire net_104;
wire net_146;
wire net_72;
wire net_122;
wire net_25;
wire net_70;
wire net_7;
wire n1333gat;
wire n113gat;
wire net_5;
wire net_52;
wire n148gat;
wire net_128;
wire n1355gat;
wire net_138;
wire net_13;
wire n218gat;
wire net_94;
wire net_11;
wire n169gat;
wire net_18;
wire net_123;
wire n36gat;
wire n1335gat;
wire net_131;
wire net_114;
wire n1349gat;
wire n1327gat;
wire net_29;
wire n231gat;
wire net_68;
wire n1341gat;
wire net_142;
wire net_77;
wire n71gat;
wire net_20;
wire net_31;
wire n1350gat;
wire net_36;
wire net_49;
wire net_15;
wire net_57;
wire net_41;
wire net_71;
wire n85gat;
wire n226gat;
wire n155gat;
wire net_3;
wire net_84;
wire n162gat;
wire net_112;
wire net_92;
wire net_1;
wire net_103;
wire n1339gat;
wire net_139;
wire n230gat;
wire n127gat;
wire net_43;
wire n1344gat;
wire net_10;
wire n1346gat;
wire net_28;
wire net_21;
wire net_51;
wire net_79;
wire n1gat;
wire net_143;
wire net_97;
wire net_88;
wire n29gat;
wire net_145;
wire net_60;
wire n134gat;
wire net_81;
wire net_58;
wire n227gat;
wire n1343gat;
wire net_82;
wire net_67;
wire net_64;
wire net_37;
wire net_110;
wire net_121;
wire net_73;
wire net_33;
wire net_48;
wire net_86;
wire net_75;
wire net_8;
wire n1326gat;
wire n106gat;
wire n233gat;
wire net_133;
wire net_125;
wire n1325gat;

// Start cells
NAND2_X1 inst_145 ( .A1(net_112), .ZN(net_104), .A2(net_103) );
XNOR2_X1 inst_103 ( .B(net_147), .ZN(n1324gat), .A(n1gat) );
NAND3_X1 inst_125 ( .A2(net_105), .ZN(net_99), .A3(net_91), .A1(net_86) );
NAND2_X1 inst_138 ( .ZN(net_92), .A2(net_90), .A1(net_77) );
NAND2_X1 inst_159 ( .A1(net_138), .ZN(net_128), .A2(net_127) );
XOR2_X1 inst_15 ( .Z(net_28), .A(n120gat), .B(n113gat) );
NAND2_X1 inst_134 ( .A1(net_116), .ZN(net_100), .A2(net_73) );
AND2_X4 inst_179 ( .A2(net_94), .A1(net_93), .ZN(net_76) );
XNOR2_X1 inst_24 ( .ZN(net_13), .A(n92gat), .B(n85gat) );
NOR2_X1 inst_114 ( .ZN(net_103), .A2(net_95), .A1(net_94) );
XOR2_X1 inst_6 ( .Z(net_15), .A(n99gat), .B(n71gat) );
NAND2_X1 inst_131 ( .ZN(net_5), .A2(n233gat), .A1(n228gat) );
XNOR2_X1 inst_76 ( .B(net_122), .ZN(n1351gat), .A(n190gat) );
NAND2_X1 inst_160 ( .A1(net_136), .A2(net_134), .ZN(net_129) );
NAND2_X1 inst_150 ( .A2(net_115), .ZN(net_114), .A1(net_112) );
XNOR2_X1 inst_33 ( .ZN(net_40), .A(net_32), .B(net_20) );
INV_X1 inst_172 ( .A(net_145), .ZN(net_75) );
XNOR2_X1 inst_83 ( .B(net_98), .ZN(n1344gat), .A(n141gat) );
XNOR2_X1 inst_47 ( .ZN(net_47), .B(net_22), .A(net_12) );
XOR2_X1 inst_19 ( .Z(net_35), .A(n50gat), .B(n43gat) );
NAND3_X1 inst_123 ( .A1(net_118), .ZN(net_87), .A2(net_86), .A3(net_82) );
NAND3_X1 inst_121 ( .A2(net_112), .ZN(net_83), .A3(net_82), .A1(net_73) );
XOR2_X1 inst_2 ( .Z(net_10), .A(n85gat), .B(n57gat) );
XOR2_X1 inst_8 ( .Z(net_17), .A(n29gat), .B(n1gat) );
NOR2_X1 inst_118 ( .ZN(net_134), .A1(net_111), .A2(net_99) );
XNOR2_X1 inst_86 ( .B(net_104), .ZN(n1341gat), .A(n120gat) );
NAND2_X1 inst_153 ( .ZN(net_121), .A2(net_120), .A1(net_116) );
XOR2_X1 inst_20 ( .Z(net_36), .A(n204gat), .B(n176gat) );
XNOR2_X1 inst_27 ( .ZN(net_22), .A(n162gat), .B(n134gat) );
XNOR2_X1 inst_38 ( .ZN(net_60), .A(net_34), .B(net_19) );
XNOR2_X1 inst_100 ( .B(net_132), .ZN(n1327gat), .A(n22gat) );
XNOR2_X1 inst_52 ( .ZN(net_59), .B(net_58), .A(net_52) );
XNOR2_X1 inst_90 ( .B(net_128), .ZN(n1337gat), .A(n92gat) );
NAND2_X1 inst_140 ( .A2(net_115), .A1(net_105), .ZN(net_96) );
XNOR2_X1 inst_40 ( .ZN(net_44), .A(net_39), .B(net_9) );
NAND2_X1 inst_162 ( .A2(net_142), .ZN(net_132), .A1(net_131) );
NAND2_X1 inst_167 ( .ZN(net_141), .A2(net_140), .A1(net_138) );
XNOR2_X1 inst_93 ( .B(net_137), .ZN(n1334gat), .A(n71gat) );
XNOR2_X1 inst_81 ( .B(net_108), .ZN(n1346gat), .A(n155gat) );
XNOR2_X1 inst_95 ( .B(net_146), .ZN(n1332gat), .A(n57gat) );
XOR2_X1 inst_1 ( .Z(net_9), .A(n92gat), .B(n64gat) );
XNOR2_X1 inst_72 ( .B(net_119), .ZN(n1355gat), .A(n218gat) );
NAND2_X1 inst_139 ( .ZN(net_95), .A2(net_90), .A1(net_78) );
NAND2_X1 inst_155 ( .ZN(net_123), .A2(net_120), .A1(net_105) );
XNOR2_X1 inst_59 ( .ZN(net_67), .A(net_57), .B(net_3) );
NAND2_X1 inst_135 ( .A1(net_118), .ZN(net_111), .A2(net_74) );
XNOR2_X1 inst_44 ( .ZN(net_58), .B(net_21), .A(net_8) );
XNOR2_X1 inst_55 ( .ZN(net_63), .B(net_56), .A(net_54) );
INV_X1 inst_174 ( .A(net_131), .ZN(net_72) );
NOR2_X1 inst_115 ( .ZN(net_142), .A1(net_100), .A2(net_99) );
XNOR2_X1 inst_37 ( .ZN(net_43), .A(net_37), .B(net_30) );
NAND2_X1 inst_148 ( .A1(net_112), .ZN(net_109), .A2(net_107) );
NAND2_X1 inst_164 ( .A1(net_138), .ZN(net_135), .A2(net_134) );
XOR2_X1 inst_5 ( .Z(net_14), .A(n99gat), .B(n106gat) );
NAND2_X1 inst_157 ( .A1(net_136), .A2(net_127), .ZN(net_125) );
XNOR2_X1 inst_84 ( .B(net_101), .ZN(n1343gat), .A(n134gat) );
XNOR2_X1 inst_51 ( .ZN(net_57), .B(net_56), .A(net_49) );
NAND2_X1 inst_142 ( .A2(net_107), .A1(net_105), .ZN(net_98) );
XNOR2_X1 inst_80 ( .B(net_97), .ZN(n1347gat), .A(n162gat) );
INV_X1 inst_173 ( .ZN(net_112), .A(net_86) );
OR3_X4 inst_105 ( .A2(net_136), .A1(net_131), .ZN(net_89), .A3(net_79) );
XNOR2_X1 inst_68 ( .ZN(net_74), .B(net_71), .A(net_41) );
XNOR2_X1 inst_78 ( .B(net_114), .ZN(n1349gat), .A(n176gat) );
XNOR2_X1 inst_42 ( .ZN(net_54), .B(net_38), .A(net_28) );
INV_X1 inst_175 ( .ZN(net_116), .A(net_74) );
XNOR2_X1 inst_53 ( .ZN(net_61), .A(net_60), .B(net_51) );
INV_X1 inst_177 ( .ZN(net_105), .A(net_84) );
NAND2_X1 inst_133 ( .ZN(net_7), .A2(n233gat), .A1(n231gat) );
XNOR2_X1 inst_26 ( .ZN(net_21), .A(n22gat), .B(n15gat) );
NAND2_X1 inst_151 ( .ZN(net_117), .A1(net_116), .A2(net_115) );
NOR2_X1 inst_112 ( .ZN(net_115), .A1(net_94), .A2(net_92) );
XNOR2_X1 inst_64 ( .ZN(net_145), .B(net_69), .A(net_42) );
NOR2_X1 inst_107 ( .A1(net_116), .A2(net_105), .ZN(net_82) );
XNOR2_X1 inst_67 ( .ZN(net_131), .B(net_64), .A(net_40) );
NAND2_X1 inst_127 ( .ZN(net_1), .A2(n233gat), .A1(n229gat) );
XNOR2_X1 inst_70 ( .ZN(net_138), .B(net_67), .A(net_44) );
NAND2_X1 inst_129 ( .ZN(net_3), .A2(n233gat), .A1(n226gat) );
XNOR2_X1 inst_92 ( .B(net_133), .ZN(n1335gat), .A(n78gat) );
XNOR2_X1 inst_29 ( .ZN(net_30), .A(n197gat), .B(n169gat) );
XOR2_X1 inst_17 ( .Z(net_32), .A(n50gat), .B(n22gat) );
XOR2_X1 inst_11 ( .Z(net_24), .A(n218gat), .B(n211gat) );
NAND2_X1 inst_146 ( .ZN(net_106), .A1(net_105), .A2(net_103) );
XOR2_X1 inst_14 ( .Z(net_27), .A(n155gat), .B(n127gat) );
NAND3_X1 inst_122 ( .A2(net_116), .ZN(net_85), .A1(net_84), .A3(net_80) );
XNOR2_X1 inst_31 ( .ZN(net_33), .A(n176gat), .B(n169gat) );
XNOR2_X1 inst_25 ( .ZN(net_18), .A(n211gat), .B(n183gat) );
NAND2_X1 inst_126 ( .ZN(net_0), .A2(n233gat), .A1(n225gat) );
NAND2_X1 inst_158 ( .A2(net_134), .A1(net_131), .ZN(net_126) );
NAND2_X1 inst_141 ( .A1(net_118), .A2(net_107), .ZN(net_97) );
XNOR2_X1 inst_62 ( .ZN(net_70), .A(net_63), .B(net_6) );
NOR2_X1 inst_110 ( .ZN(net_79), .A1(net_78), .A2(net_77) );
XNOR2_X1 inst_74 ( .B(net_113), .ZN(n1353gat), .A(n204gat) );
XNOR2_X1 inst_57 ( .ZN(net_65), .A(net_53), .B(net_4) );
XNOR2_X1 inst_35 ( .ZN(net_42), .A(net_17), .B(net_10) );
XNOR2_X1 inst_99 ( .B(net_144), .ZN(n1328gat), .A(n29gat) );
XNOR2_X1 inst_48 ( .ZN(net_50), .A(net_49), .B(net_48) );
XNOR2_X1 inst_69 ( .ZN(net_73), .B(net_65), .A(net_47) );
XNOR2_X1 inst_46 ( .ZN(net_48), .B(net_31), .A(net_26) );
XNOR2_X1 inst_82 ( .B(net_109), .ZN(n1345gat), .A(n148gat) );
NAND2_X1 inst_136 ( .A1(net_136), .ZN(net_94), .A2(net_72) );
XNOR2_X1 inst_30 ( .ZN(net_31), .A(n148gat), .B(n141gat) );
XNOR2_X1 inst_102 ( .B(net_139), .ZN(n1325gat), .A(n8gat) );
NOR2_X1 inst_108 ( .A2(net_118), .A1(net_112), .ZN(net_80) );
NAND2_X1 inst_165 ( .A2(net_140), .ZN(net_137), .A1(net_136) );
XNOR2_X1 inst_32 ( .ZN(net_52), .A(net_35), .B(net_29) );
XOR2_X1 inst_22 ( .Z(net_38), .A(n134gat), .B(n127gat) );
NAND2_X1 inst_144 ( .A1(net_116), .A2(net_103), .ZN(net_102) );
XNOR2_X1 inst_34 ( .ZN(net_41), .A(net_27), .B(net_18) );
XOR2_X1 inst_12 ( .Z(net_25), .A(n204gat), .B(n197gat) );
XNOR2_X1 inst_56 ( .ZN(net_64), .A(net_50), .B(net_5) );
XNOR2_X1 inst_71 ( .ZN(net_84), .B(net_68), .A(net_43) );
XOR2_X1 inst_21 ( .Z(net_37), .A(n141gat), .B(n113gat) );
OR3_X4 inst_104 ( .A2(net_145), .A1(net_138), .ZN(net_88), .A3(net_76) );
XNOR2_X1 inst_60 ( .ZN(net_68), .A(net_59), .B(net_1) );
NAND2_X1 inst_169 ( .A1(net_145), .ZN(net_144), .A2(net_134) );
NAND2_X1 inst_168 ( .ZN(net_143), .A2(net_142), .A1(net_136) );
XNOR2_X1 inst_97 ( .B(net_129), .ZN(n1330gat), .A(n43gat) );
NAND2_X1 inst_161 ( .A1(net_145), .ZN(net_130), .A2(net_127) );
NAND3_X1 inst_124 ( .A1(net_112), .ZN(net_110), .A3(net_91), .A2(net_84) );
XOR2_X1 inst_18 ( .Z(net_34), .A(n64gat), .B(n57gat) );
XOR2_X1 inst_16 ( .Z(net_29), .A(n36gat), .B(n29gat) );
XNOR2_X1 inst_88 ( .B(net_124), .ZN(n1339gat), .A(n106gat) );
XOR2_X1 inst_3 ( .Z(net_11), .A(n190gat), .B(n183gat) );
NAND2_X1 inst_156 ( .A1(net_131), .A2(net_127), .ZN(net_124) );
XOR2_X1 inst_9 ( .Z(net_19), .A(n78gat), .B(n71gat) );
NOR2_X1 inst_113 ( .ZN(net_107), .A2(net_95), .A1(net_93) );
NAND2_X1 inst_170 ( .ZN(net_146), .A1(net_145), .A2(net_140) );
XNOR2_X1 inst_50 ( .ZN(net_55), .A(net_54), .B(net_48) );
NAND2_X1 inst_137 ( .ZN(net_91), .A2(net_89), .A1(net_88) );
XNOR2_X1 inst_41 ( .ZN(net_51), .A(net_14), .B(net_13) );
NAND2_X1 inst_130 ( .ZN(net_4), .A2(n233gat), .A1(n232gat) );
XNOR2_X1 inst_91 ( .B(net_130), .ZN(n1336gat), .A(n85gat) );
NAND2_X1 inst_132 ( .ZN(net_6), .A2(n233gat), .A1(n227gat) );
NAND2_X1 inst_143 ( .A1(net_118), .A2(net_103), .ZN(net_101) );
INV_X1 inst_176 ( .ZN(net_118), .A(net_73) );
NAND2_X1 inst_152 ( .A2(net_120), .ZN(net_119), .A1(net_118) );
XNOR2_X1 inst_58 ( .ZN(net_66), .A(net_61), .B(net_2) );
XNOR2_X1 inst_36 ( .ZN(net_49), .A(net_25), .B(net_24) );
NAND2_X1 inst_147 ( .A1(net_116), .ZN(net_108), .A2(net_107) );
XNOR2_X1 inst_87 ( .B(net_106), .ZN(n1340gat), .A(n113gat) );
XNOR2_X1 inst_61 ( .ZN(net_69), .A(net_55), .B(net_0) );
XNOR2_X1 inst_45 ( .ZN(net_46), .B(net_16), .A(net_15) );
XNOR2_X1 inst_96 ( .B(net_126), .ZN(n1331gat), .A(n50gat) );
XNOR2_X1 inst_101 ( .B(net_143), .ZN(n1326gat), .A(n15gat) );
XOR2_X1 inst_0 ( .Z(net_8), .A(n8gat), .B(n1gat) );
XOR2_X1 inst_10 ( .Z(net_20), .A(n78gat), .B(n106gat) );
XOR2_X1 inst_4 ( .Z(net_12), .A(n218gat), .B(n190gat) );
XNOR2_X1 inst_65 ( .ZN(net_86), .B(net_66), .A(net_45) );
AND2_X4 inst_178 ( .A1(net_138), .ZN(net_77), .A2(net_75) );
XNOR2_X1 inst_89 ( .B(net_125), .ZN(n1338gat), .A(n99gat) );
XNOR2_X1 inst_28 ( .ZN(net_23), .A(n148gat), .B(n120gat) );
NOR2_X1 inst_111 ( .ZN(net_120), .A1(net_93), .A2(net_92) );
XNOR2_X1 inst_66 ( .ZN(net_136), .B(net_70), .A(net_46) );
NOR2_X1 inst_117 ( .ZN(net_140), .A2(net_110), .A1(net_100) );
XNOR2_X1 inst_98 ( .B(net_135), .ZN(n1329gat), .A(n36gat) );
XNOR2_X1 inst_63 ( .ZN(net_71), .A(net_62), .B(net_7) );
XOR2_X1 inst_7 ( .Z(net_16), .A(n43gat), .B(n15gat) );
XNOR2_X1 inst_49 ( .ZN(net_53), .A(net_52), .B(net_51) );
NAND3_X1 inst_120 ( .A1(net_105), .ZN(net_81), .A3(net_80), .A2(net_74) );
NAND2_X1 inst_154 ( .ZN(net_122), .A1(net_118), .A2(net_115) );
XOR2_X1 inst_13 ( .Z(net_26), .A(n162gat), .B(n155gat) );
NAND4_X1 inst_119 ( .ZN(net_90), .A2(net_87), .A1(net_85), .A3(net_83), .A4(net_81) );
XNOR2_X1 inst_75 ( .B(net_123), .ZN(n1352gat), .A(n197gat) );
NAND2_X1 inst_166 ( .A2(net_142), .ZN(net_139), .A1(net_138) );
NOR2_X1 inst_116 ( .ZN(net_127), .A1(net_111), .A2(net_110) );
NAND2_X1 inst_163 ( .A2(net_140), .ZN(net_133), .A1(net_131) );
XNOR2_X1 inst_85 ( .B(net_102), .ZN(n1342gat), .A(n127gat) );
XNOR2_X1 inst_54 ( .ZN(net_62), .A(net_60), .B(net_58) );
XNOR2_X1 inst_79 ( .B(net_96), .ZN(n1348gat), .A(n169gat) );
NOR2_X1 inst_109 ( .A2(net_138), .ZN(net_78), .A1(net_75) );
OR2_X4 inst_106 ( .A2(net_136), .ZN(net_93), .A1(net_72) );
NAND2_X1 inst_149 ( .A2(net_120), .ZN(net_113), .A1(net_112) );
XNOR2_X1 inst_43 ( .ZN(net_45), .A(net_36), .B(net_23) );
XNOR2_X1 inst_39 ( .ZN(net_56), .B(net_33), .A(net_11) );
NAND2_X1 inst_128 ( .ZN(net_2), .A2(n233gat), .A1(n230gat) );
XNOR2_X1 inst_73 ( .B(net_121), .ZN(n1354gat), .A(n211gat) );
XOR2_X1 inst_23 ( .Z(net_39), .A(n8gat), .B(n36gat) );
NAND2_X1 inst_171 ( .ZN(net_147), .A1(net_145), .A2(net_142) );
XNOR2_X1 inst_77 ( .B(net_117), .ZN(n1350gat), .A(n183gat) );
XNOR2_X1 inst_94 ( .B(net_141), .ZN(n1333gat), .A(n64gat) );

endmodule
