module usb_phy_ispd (
phy_tx_mode,
DataOut_i_3_,
tau_clk,
DataOut_i_1_,
DataOut_i_7_,
DataOut_i_5_,
rxd,
rst,
TxValid_i,
rxdp,
rxdn,
DataOut_i_2_,
DataOut_i_0_,
DataOut_i_4_,
DataOut_i_6_,
DataIn_o_2_,
txdn,
txdp,
LineState_o_0_,
RxValid_o,
txoe,
LineState_o_1_,
DataIn_o_7_,
DataIn_o_4_,
usb_rst,
DataIn_o_5_,
DataIn_o_3_,
RxError_o,
g1897_u0_o,
DataIn_o_1_,
TxReady_o,
DataIn_o_0_,
RxActive_o,
DataIn_o_6_);

// Start PIs
input phy_tx_mode;
input DataOut_i_3_;
input tau_clk;
input DataOut_i_1_;
input DataOut_i_7_;
input DataOut_i_5_;
input rxd;
input rst;
input TxValid_i;
input rxdp;
input rxdn;
input DataOut_i_2_;
input DataOut_i_0_;
input DataOut_i_4_;
input DataOut_i_6_;

// Start POs
output DataIn_o_2_;
output txdn;
output txdp;
output LineState_o_0_;
output RxValid_o;
output txoe;
output LineState_o_1_;
output DataIn_o_7_;
output DataIn_o_4_;
output usb_rst;
output DataIn_o_5_;
output DataIn_o_3_;
output RxError_o;
output g1897_u0_o;
output DataIn_o_1_;
output TxReady_o;
output DataIn_o_0_;
output RxActive_o;
output DataIn_o_6_;

// Start wires
wire newNet_120;
wire newNet_199;
wire n_707;
wire newNet_235;
wire newNet_110;
wire n_479;
wire g1778_db;
wire newNet_10;
wire n_990;
wire n_960;
wire i_tx_phy_bit_cnt_2_;
wire newNet_166;
wire newNet_130;
wire n_959;
wire n_980;
wire newNet_24;
wire i_tx_phy_sd_raw_o;
wire n_297;
wire newNet_79;
wire n_192;
wire i_tx_phy_hold_reg_d_11;
wire n_210;
wire newNet_117;
wire newNet_73;
wire newNet_63;
wire n_184;
wire n_61;
wire g2068_p;
wire n_232;
wire n_362;
wire newNet_193;
wire i_tx_phy_txoe_r1;
wire newNet_2;
wire newNet_25;
wire newNet_247;
wire n_331;
wire n_341;
wire n_509;
wire g1980_p;
wire i_rx_phy_bit_cnt_2_;
wire n_484;
wire g1741_p;
wire newNet_38;
wire n_353;
wire n_737;
wire newNet_292;
wire n_157;
wire g2050_p;
wire n_701;
wire n_749;
wire newNet_124;
wire i_rx_phy_dpll_state_1_;
wire newNet_149;
wire newNet_101;
wire n_125;
wire newNet_83;
wire i_tx_phy_one_cnt_2_;
wire n_323;
wire n_410;
wire newNet_189;
wire newNet_160;
wire newNet_113;
wire newNet_53;
wire n_274;
wire g1965_p;
wire n_256;
wire n_977;
wire g2108_p;
wire newNet_272;
wire n_373;
wire n_395;
wire n_318;
wire newNet_92;
wire newNet_19;
wire i_rx_phy_bit_stuff_err_reg_Q;
wire n_763;
wire n_233;
wire newNet_26;
wire FE_RN_0_0;
wire n_53;
wire newNet_297;
wire n_426;
wire newNet_46;
wire n_227;
wire n_404;
wire n_507;
wire n_629;
wire newNet_214;
wire newNet_279;
wire newNet_183;
wire newNet_201;
wire n_223;
wire newNet_157;
wire newNet_286;
wire newNet_139;
wire newNet_140;
wire newNet_256;
wire newNet_174;
wire n_231;
wire newNet_277;
wire n_332;
wire n_391;
wire newNet_99;
wire n_165;
wire n_947;
wire newNet_237;
wire i_rx_phy_one_cnt_0_;
wire n_435;
wire newNet_108;
wire g1778_da;
wire newNet_150;
wire n_937;
wire newNet_309;
wire newNet_220;
wire newNet_269;
wire newNet_268;
wire n_974;
wire newNet_226;
wire n_511;
wire RxActive_o;
wire i_rx_phy_rxd_s0;
wire g1742_p;
wire n_37;
wire n_290;
wire n_154;
wire n_300;
wire n_97;
wire rxd;
wire newNet_119;
wire g1757_p;
wire newNet_3;
wire n_958;
wire newNet_158;
wire i_rx_phy_bit_cnt_0_;
wire n_324;
wire newNet_244;
wire g1777_db;
wire n_486;
wire n_127;
wire n_141;
wire n_800;
wire newNet_234;
wire newNet_313;
wire newNet_261;
wire n_361;
wire n_748;
wire TxReady_o;
wire n_115;
wire n_70;
wire n_126;
wire newNet_188;
wire n_183;
wire n_665;
wire newNet_8;
wire newNet_29;
wire n_246;
wire n_170;
wire newNet_257;
wire newNet_116;
wire g2413_p;
wire newNet_51;
wire newNet_5;
wire n_427;
wire i_rx_phy_shift_en;
wire g1780_db;
wire n_360;
wire n_366;
wire n_447;
wire n_359;
wire newNet_74;
wire newNet_23;
wire newNet_260;
wire g2113_p;
wire n_485;
wire n_450;
wire newNet_47;
wire n_884;
wire n_222;
wire newNet_228;
wire n_796;
wire newNet_41;
wire n_991;
wire n_434;
wire n_506;
wire n_52;
wire n_166;
wire n_195;
wire n_405;
wire g1782_sb;
wire n_424;
wire newNet_271;
wire newNet_66;
wire n_273;
wire newNet_207;
wire newNet_121;
wire n_258;
wire newNet_109;
wire n_77;
wire newNet_255;
wire newNet_0;
wire n_944;
wire g2506_p;
wire newNet_50;
wire n_920;
wire g1975_p;
wire newNet_56;
wire newNet_112;
wire n_152;
wire newNet_169;
wire newNet_138;
wire i_tx_phy_hold_reg_10;
wire newNet_293;
wire n_894;
wire n_919;
wire newNet_137;
wire g2067_p;
wire n_406;
wire newNet_204;
wire n_727;
wire n_266;
wire n_976;
wire n_325;
wire n_312;
wire n_459;
wire newNet_285;
wire n_389;
wire n_69;
wire newNet_177;
wire newNet_39;
wire n_794;
wire n_296;
wire newNet_94;
wire i_rx_phy_rxdn_s_r;
wire newNet_236;
wire n_317;
wire newNet_122;
wire DataOut_i_2_;
wire newNet_267;
wire n_364;
wire n_935;
wire newNet_312;
wire newNet_181;
wire n_461;
wire g1779_db;
wire newNet_274;
wire txoe;
wire newNet_280;
wire n_161;
wire newNet_241;
wire g15_p;
wire DataIn_o_4_;
wire newNet_216;
wire newNet_197;
wire newNet_245;
wire n_299;
wire n_334;
wire newNet_65;
wire n_257;
wire newNet_48;
wire newNet_42;
wire n_58;
wire n_35;
wire n_742;
wire newNet_36;
wire n_310;
wire newNet_143;
wire g1738_p;
wire newNet_294;
wire newNet_107;
wire n_631;
wire newNet_221;
wire n_735;
wire n_878;
wire i_tx_phy_hold_reg_d_17;
wire g1777_da;
wire n_529;
wire n_764;
wire n_453;
wire newNet_52;
wire newNet_288;
wire LineState_o_1_;
wire n_431;
wire newNet_89;
wire n_972;
wire n_167;
wire n_235;
wire n_175;
wire n_351;
wire n_182;
wire g1739_p;
wire n_916;
wire n_369;
wire n_51;
wire n_225;
wire n_982;
wire newNet_258;
wire newNet_75;
wire g1776_da;
wire newNet_17;
wire newNet_205;
wire newNet_299;
wire i_rx_phy_se0_r_reg_Q;
wire g2063_sb;
wire newNet_164;
wire n_85;
wire newNet_192;
wire rst_cnt_4_;
wire rst_cnt_3_;
wire n_124;
wire g2651_p;
wire n_885;
wire n_425;
wire newNet_303;
wire newNet_93;
wire n_138;
wire n_505;
wire i_rx_phy_rxdn_s_r_reg_Q;
wire newNet_296;
wire i_tx_phy_append_eop_sync4;
wire n_490;
wire newNet_82;
wire n_759;
wire i_tx_phy_state_2_;
wire n_132;
wire n_269;
wire n_914;
wire n_708;
wire n_590;
wire g2385_p;
wire n_9;
wire i_rx_phy_rxdp_s;
wire DataIn_o_3_;
wire newNet_118;
wire newNet_106;
wire n_15;
wire n_632;
wire n_217;
wire n_130;
wire newNet_308;
wire n_330;
wire newNet_176;
wire newNet_152;
wire n_413;
wire newNet_239;
wire newNet_142;
wire n_57;
wire n_743;
wire txdp;
wire n_354;
wire newNet_167;
wire n_934;
wire n_255;
wire n_168;
wire g1881_p;
wire DataOut_i_3_;
wire newNet_198;
wire i_tx_phy_sft_done;
wire n_263;
wire n_460;
wire g11_p;
wire newNet_35;
wire n_921;
wire n_452;
wire newNet_304;
wire i_tx_phy_ld_data_reg_Q;
wire n_539;
wire g2494_p;
wire rxdp;
wire g1855_sb;
wire n_407;
wire newNet_100;
wire n_915;
wire n_758;
wire newNet_232;
wire n_176;
wire newNet_287;
wire n_888;
wire n_209;
wire n_244;
wire n_436;
wire n_191;
wire n_968;
wire newNet_128;
wire n_116;
wire newNet_240;
wire newNet_186;
wire n_322;
wire n_277;
wire n_105;
wire n_342;
wire newNet_301;
wire n_840;
wire newNet_54;
wire n_306;
wire newNet_49;
wire newNet_180;
wire n_12;
wire g1897_u0_o;
wire newNet_254;
wire n_21;
wire n_28;
wire DataOut_i_0_;
wire n_169;
wire DataIn_o_6_;
wire i_tx_phy_one_cnt_1_;
wire g1923_p;
wire newNet_295;
wire n_499;
wire n_388;
wire n_27;
wire g1779_sb;
wire n_245;
wire newNet_96;
wire i_tx_phy_tx_ip;
wire newNet_208;
wire newNet_307;
wire n_333;
wire n_788;
wire g2069_p;
wire n_567;
wire n_852;
wire newNet_22;
wire n_924;
wire newNet_141;
wire n_559;
wire g1781_db;
wire n_930;
wire n_709;
wire n_411;
wire n_540;
wire n_925;
wire n_967;
wire n_472;
wire newNet_311;
wire newNet_227;
wire n_864;
wire newNet_156;
wire newNet_87;
wire n_666;
wire newNet_59;
wire n_756;
wire i_rx_phy_sync_err;
wire i_tx_phy_sft_done_r;
wire n_700;
wire g1776_db;
wire newNet_202;
wire n_133;
wire n_446;
wire n_598;
wire newNet_187;
wire newNet_310;
wire n_224;
wire newNet_215;
wire newNet_273;
wire newNet_259;
wire n_50;
wire newNet_68;
wire n_64;
wire newNet_151;
wire n_131;
wire newNet_134;
wire n_340;
wire n_482;
wire newNet_305;
wire newNet_238;
wire n_804;
wire newNet_191;
wire n_722;
wire newNet_7;
wire n_415;
wire newNet_170;
wire DataIn_o_7_;
wire n_338;
wire newNet_178;
wire n_259;
wire n_604;
wire n_969;
wire newNet_243;
wire i_tx_phy_hold_reg_d_15;
wire n_574;
wire newNet_80;
wire newNet_223;
wire newNet_16;
wire n_444;
wire n_782;
wire g1778_sb;
wire DataOut_i_4_;
wire i_tx_phy_sd_bs_o;
wire newNet_281;
wire newNet_264;
wire g1780_sb;
wire newNet_145;
wire g2128_p;
wire rst;
wire n_948;
wire newNet_211;
wire n_292;
wire newNet_61;
wire n_952;
wire newNet_162;
wire n_951;
wire n_228;
wire n_33;
wire n_538;
wire g2674_p;
wire newNet_155;
wire n_268;
wire n_922;
wire n_471;
wire n_754;
wire n_873;
wire n_710;
wire n_941;
wire newNet_88;
wire n_439;
wire n_237;
wire i_rx_phy_byte_err;
wire n_11;
wire i_tx_phy_one_cnt_0_;
wire n_163;
wire n_400;
wire newNet_230;
wire n_573;
wire n_7;
wire n_74;
wire n_22;
wire i_rx_phy_rx_valid_r;
wire newNet_57;
wire n_120;
wire newNet_200;
wire newNet_76;
wire n_971;
wire newNet_276;
wire newNet_95;
wire n_455;
wire RxError_o;
wire i_rx_phy_rxd_s1_reg_Q;
wire n_841;
wire g1781_da;
wire n_316;
wire newNet_62;
wire n_741;
wire i_tx_phy_hold_reg_d_reg_1__Q;
wire n_420;
wire newNet_30;
wire n_699;
wire newNet_263;
wire newNet_21;
wire n_704;
wire n_368;
wire n_785;
wire n_352;
wire LineState_o_0_;
wire newNet_13;
wire n_193;
wire i_tx_phy_hold_reg_4;
wire newNet_253;
wire rxdn;
wire i_rx_phy_sd_nrzi;
wire i_rx_phy_rx_valid1;
wire n_56;
wire n_989;
wire i_tx_phy_hold_reg_6;
wire n_933;
wire n_201;
wire phy_tx_mode;
wire newNet_11;
wire i_rx_phy_se0_s;
wire n_377;
wire newNet_195;
wire n_480;
wire n_423;
wire g1884_p;
wire n_88;
wire n_71;
wire newNet_123;
wire newNet_67;
wire newNet_252;
wire g1781_sb;
wire n_387;
wire newNet_249;
wire n_926;
wire n_394;
wire newNet_222;
wire n_462;
wire i_rx_phy_rxdp_s0;
wire n_103;
wire newNet_219;
wire n_386;
wire n_293;
wire i_tx_phy_hold_reg_d_reg_5__Q;
wire g2412_p;
wire newNet_171;
wire newNet_196;
wire n_923;
wire newNet_265;
wire n_755;
wire newNet_282;
wire newNet_28;
wire n_963;
wire n_339;
wire newNet_70;
wire newNet_289;
wire newNet_144;
wire n_443;
wire newNet_185;
wire n_940;
wire g2057_p;
wire n_63;
wire newNet_270;
wire i_tx_phy_hold_reg;
wire n_304;
wire n_966;
wire i_rx_phy_one_cnt_2_;
wire n_100;
wire n_414;
wire n_283;
wire n_697;
wire i_rx_phy_dpll_state_0_;
wire n_55;
wire newNet_154;
wire n_347;
wire rst_cnt_0_;
wire newNet_251;
wire newNet_190;
wire newNet_18;
wire n_734;
wire n_949;
wire n_409;
wire g1942_p;
wire g2028_p;
wire n_783;
wire n_252;
wire newNet_15;
wire n_320;
wire newNet_77;
wire n_243;
wire newNet_210;
wire newNet_248;
wire newNet_34;
wire txdn;
wire n_970;
wire n_291;
wire newNet_90;
wire n_275;
wire newNet_12;
wire n_401;
wire n_301;
wire n_278;
wire i_tx_phy_bit_cnt_1_;
wire newNet_126;
wire newNet_14;
wire i_tx_phy_hold_reg_7;
wire newNet_242;
wire newNet_115;
wire newNet_146;
wire tau_clk;
wire n_988;
wire n_421;
wire i_tx_phy_append_eop_sync2;
wire newNet_275;
wire DataOut_i_5_;
wire newNet_233;
wire newNet_133;
wire i_rx_phy_rxd_r;
wire n_593;
wire newNet_290;
wire newNet_163;
wire n_375;
wire newNet_98;
wire newNet_302;
wire n_454;
wire newNet_206;
wire n_108;
wire newNet_165;
wire newNet_27;
wire rst_cnt_1_;
wire n_433;
wire n_932;
wire g1780_da;
wire n_267;
wire newNet_184;
wire n_913;
wire n_984;
wire n_111;
wire n_142;
wire i_rx_phy_rxdp_s_r;
wire g2063_db;
wire n_139;
wire n_121;
wire n_583;
wire n_280;
wire newNet_105;
wire newNet_31;
wire n_118;
wire n_48;
wire n_927;
wire newNet_153;
wire n_786;
wire DataOut_i_1_;
wire i_tx_phy_hold_reg_5;
wire n_767;
wire newNet_40;
wire i_tx_phy_hold_reg_d_reg_3__Q;
wire n_367;
wire n_489;
wire newNet_85;
wire n_523;
wire n_440;
wire n_957;
wire n_122;
wire n_204;
wire newNet_6;
wire newNet_262;
wire n_726;
wire n_457;
wire n_481;
wire n_198;
wire newNet_129;
wire newNet_71;
wire n_226;
wire n_962;
wire usb_rst;
wire n_385;
wire i_rx_phy_rx_en;
wire i_tx_phy_data_done;
wire n_487;
wire DataIn_o_5_;
wire g2116_p;
wire newNet_103;
wire TxValid_i;
wire newNet_225;
wire newNet_182;
wire newNet_161;
wire newNet_4;
wire newNet_32;
wire i_rx_phy_se0_r;
wire n_230;
wire newNet_172;
wire n_449;
wire i_tx_phy_hold_reg_d_reg_6__Q;
wire newNet_69;
wire g1855_db;
wire n_203;
wire n_456;
wire i_tx_phy_bit_cnt_0_;
wire n_66;
wire n_90;
wire i_rx_phy_rxd_s;
wire n_661;
wire newNet_81;
wire i_rx_phy_fs_ce_r1;
wire n_992;
wire i_rx_phy_fs_state_0_;
wire n_185;
wire newNet_1;
wire i_tx_phy_sd_nrzi_o;
wire i_tx_phy_hold_reg_d_13;
wire newNet_213;
wire g1782_db;
wire g1901_p;
wire i_rx_phy_rxd_s1;
wire n_155;
wire newNet_266;
wire n_311;
wire newNet_9;
wire n_153;
wire n_965;
wire newNet_159;
wire newNet_283;
wire newNet_250;
wire n_294;
wire DataIn_o_0_;
wire n_417;
wire newNet_55;
wire newNet_229;
wire newNet_217;
wire i_tx_phy_append_eop;
wire n_308;
wire newNet_147;
wire n_355;
wire n_428;
wire newNet_300;
wire n_265;
wire n_213;
wire FE_RN_2_0;
wire n_350;
wire n_229;
wire g1776_sb;
wire n_458;
wire n_943;
wire i_tx_phy_hold_reg_d;
wire n_254;
wire newNet_136;
wire n_392;
wire newNet_284;
wire i_tx_phy_state_1_;
wire i_tx_phy_append_eop_sync1;
wire n_288;
wire newNet_102;
wire newNet_168;
wire n_238;
wire newNet_125;
wire i_rx_phy_rxdn_s0;
wire newNet_203;
wire n_112;
wire RxValid_o;
wire n_910;
wire n_928;
wire g1779_da;
wire g1782_da;
wire newNet_127;
wire g1737_p;
wire n_706;
wire n_344;
wire newNet_246;
wire newNet_132;
wire newNet_33;
wire n_240;
wire n_882;
wire newNet_291;
wire n_276;
wire g2035_p;
wire FE_RN_1_0;
wire n_10;
wire i_tx_phy_hold_reg_8;
wire n_432;
wire n_752;
wire i_rx_phy_one_cnt_1_;
wire DataIn_o_1_;
wire newNet_20;
wire newNet_111;
wire newNet_114;
wire newNet_104;
wire n_942;
wire g2141_p;
wire n_18;
wire newNet_212;
wire g2066_p;
wire n_981;
wire n_753;
wire n_239;
wire newNet_179;
wire n_49;
wire n_660;
wire g1857_p;
wire n_483;
wire n_319;
wire newNet_135;
wire i_tx_phy_txoe_r2;
wire g2103_p;
wire n_309;
wire i_rx_phy_byte_err_reg_Q;
wire n_337;
wire newNet_86;
wire i_tx_phy_ld_data;
wire newNet_209;
wire n_251;
wire newNet_60;
wire newNet_131;
wire i_tx_phy_hold_reg_d_12;
wire i_rx_phy_rxdn_s;
wire newNet_44;
wire newNet_306;
wire n_60;
wire i_rx_phy_bit_stuff_err;
wire n_492;
wire newNet_72;
wire n_106;
wire n_164;
wire n_81;
wire newNet_97;
wire g41_p;
wire n_186;
wire n_197;
wire newNet_45;
wire newNet_37;
wire n_248;
wire n_961;
wire newNet_173;
wire n_416;
wire newNet_64;
wire n_289;
wire n_123;
wire newNet_78;
wire i_rx_phy_sync_err_reg_Q;
wire n_588;
wire g1740_p;
wire i_tx_phy_hold_reg_d_14;
wire n_370;
wire i_rx_phy_sd_r;
wire g2063_da;
wire newNet_224;
wire newNet_43;
wire n_343;
wire n_54;
wire n_307;
wire newNet_58;
wire n_945;
wire n_384;
wire newNet_91;
wire g1855_da;
wire newNet_148;
wire g1743_p;
wire n_91;
wire n_172;
wire n_703;
wire n_8;
wire DataOut_i_7_;
wire n_911;
wire n_365;
wire n_313;
wire g2130_p;
wire n_390;
wire n_150;
wire i_rx_phy_fs_state_2_;
wire newNet_84;
wire DataIn_o_2_;
wire n_493;
wire n_380;
wire newNet_194;
wire g2091_p;
wire newNet_175;
wire i_tx_phy_hold_reg_9;
wire n_929;
wire newNet_278;
wire newNet_231;
wire n_628;
wire DataOut_i_6_;
wire n_467;
wire n_378;
wire n_938;
wire i_rx_phy_fs_ce_r2;
wire g1777_sb;
wire n_241;
wire newNet_298;
wire i_rx_phy_rxdp_s_r_reg_Q;
wire newNet_218;

// Start cells
in01f80 newInst_312 ( .a(newNet_96), .o(newNet_312) );
no02f80 g2096_u0 ( .a(n_984), .b(usb_rst), .o(n_103) );
no02f80 g1950_u0 ( .a(n_210), .b(n_882), .o(n_296) );
in01f80 newInst_252 ( .a(newNet_251), .o(newNet_252) );
in01f80 g2511_u0 ( .a(n_763), .o(n_764) );
ao12f80 g1845_u0 ( .a(n_961), .b(n_157), .c(n_352), .o(n_406) );
na02f80 g2512_u0 ( .a(n_759), .b(n_885), .o(n_763) );
na02f80 g2027_u0 ( .a(n_55), .b(n_50), .o(n_182) );
in01f80 g2003_u0 ( .a(n_982), .o(n_217) );
na02f80 g2111_u0 ( .a(i_tx_phy_bit_cnt_1_), .b(n_56), .o(n_804) );
in01f80 newInst_224 ( .a(newNet_223), .o(newNet_224) );
in01f80 newInst_54 ( .a(newNet_53), .o(newNet_54) );
na02f80 g1916_u0 ( .a(n_37), .b(n_764), .o(n_331) );
in01f80 g27_u0 ( .a(n_224), .o(n_559) );
no02f80 g1896_u0 ( .a(n_132), .b(n_70), .o(n_197) );
in01f80 newInst_211 ( .a(newNet_210), .o(newNet_211) );
in01f80 newInst_305 ( .a(newNet_304), .o(newNet_305) );
ms00f80 i_tx_phy_one_cnt_reg_0__u0 ( .ck(newNet_71), .d(n_378), .o(i_tx_phy_one_cnt_0_) );
na02f80 g2000_u0 ( .a(i_rx_phy_rxd_s0), .b(n_130), .o(n_131) );
no02f80 g2057_u0 ( .a(i_rx_phy_sd_r), .b(n_243), .o(g2057_p) );
oa12f80 g1977_u0 ( .a(n_183), .b(n_185), .c(n_224), .o(n_225) );
na03f80 g1649_u0 ( .a(i_rx_phy_byte_err), .b(i_rx_phy_sync_err), .c(i_rx_phy_bit_stuff_err), .o(RxError_o) );
in01f80 newInst_3 ( .a(newNet_1), .o(newNet_3) );
ms00f80 i_rx_phy_se0_s_reg_u0 ( .ck(newNet_166), .d(n_471), .o(i_rx_phy_se0_s) );
in01f80 g2190_u0 ( .a(RxActive_o), .o(n_509) );
in01f80 newInst_217 ( .a(newNet_216), .o(newNet_217) );
in01f80 newInst_268 ( .a(newNet_267), .o(newNet_268) );
in01f80 newInst_74 ( .a(newNet_54), .o(newNet_74) );
ms00f80 i_rx_phy_rxdp_s_reg_u0 ( .ck(newNet_181), .d(n_309), .o(i_rx_phy_rxdp_s) );
in01f80 newInst_68 ( .a(newNet_42), .o(newNet_68) );
no02f80 g1961_u0 ( .a(n_233), .b(n_318), .o(n_320) );
na02f80 g2087_u0 ( .a(i_tx_phy_one_cnt_2_), .b(n_873), .o(n_163) );
in01f80 g2491_u0 ( .a(n_735), .o(n_737) );
na02f80 g2461_u0 ( .a(n_257), .b(n_929), .o(n_701) );
in01f80 newInst_204 ( .a(newNet_203), .o(newNet_204) );
na04m80 g1936_u0 ( .a(n_182), .b(n_15), .c(i_tx_phy_bit_cnt_2_), .d(n_77), .o(n_263) );
in01f80 g2092_u0 ( .a(n_111), .o(n_112) );
na02f80 g1739_u0 ( .a(n_456), .b(n_974), .o(g1739_p) );
in01f80 newInst_143 ( .a(newNet_93), .o(newNet_143) );
ms00f80 i_tx_phy_append_eop_sync2_reg_u0 ( .ck(newNet_142), .d(n_316), .o(i_tx_phy_append_eop_sync2) );
in01f80 g2152_u0 ( .a(i_rx_phy_bit_cnt_0_), .o(n_37) );
no02f80 g2626_u0 ( .a(n_224), .b(n_888), .o(n_928) );
in01f80 newInst_2 ( .a(newNet_1), .o(newNet_2) );
in01f80 i_rx_phy_bit_stuff_err_reg_u1 ( .a(i_rx_phy_bit_stuff_err_reg_Q), .o(i_rx_phy_bit_stuff_err) );
ms00f80 rst_cnt_reg_4__u0 ( .ck(newNet_5), .d(n_423), .o(rst_cnt_4_) );
no02f80 g2640_u0 ( .a(n_980), .b(n_947), .o(n_948) );
in01f80 g2440_u0 ( .a(i_rx_phy_rxdp_s), .o(n_666) );
in01f80 g2182_u0 ( .a(i_tx_phy_bit_cnt_0_), .o(n_56) );
in01f80 g2026_u0 ( .a(n_182), .o(n_210) );
in01f80 newInst_36 ( .a(newNet_26), .o(newNet_36) );
oa12f80 g2502_u0 ( .a(n_754), .b(n_944), .c(n_752), .o(n_755) );
in01f80 newInst_294 ( .a(newNet_293), .o(newNet_294) );
na03f80 g1926_u0 ( .a(n_259), .b(n_50), .c(g2674_p), .o(n_299) );
no02f80 g2068_u0 ( .a(n_353), .b(i_rx_phy_bit_cnt_0_), .o(g2068_p) );
in01f80 newInst_156 ( .a(newNet_63), .o(newNet_156) );
in01f80 g2219_u0 ( .a(i_tx_phy_one_cnt_1_), .o(n_49) );
in01f80 g2173_u0 ( .a(rst_cnt_1_), .o(n_22) );
in01f80 newInst_7 ( .a(newNet_1), .o(newNet_7) );
oa12f80 g1928_u0 ( .a(n_131), .b(n_127), .c(i_rx_phy_rxd_s1), .o(n_229) );
ms00f80 i_rx_phy_se0_r_reg_u0 ( .ck(newNet_171), .d(n_446), .o(i_rx_phy_se0_r_reg_Q) );
no02f80 g2639_u0 ( .a(n_794), .b(n_111), .o(n_945) );
ms00f80 i_tx_phy_hold_reg_reg_3__u0 ( .ck(newNet_90), .d(n_485), .o(i_tx_phy_hold_reg_6) );
in01f80 newInst_173 ( .a(newNet_172), .o(newNet_173) );
na02f80 g2627_u0 ( .a(n_930), .b(n_933), .o(n_934) );
in01f80 g2599_u0 ( .a(n_885), .o(n_882) );
na02f80 g2048_u0 ( .a(n_277), .b(i_tx_phy_sd_bs_o), .o(n_278) );
in01f80 newInst_108 ( .a(newNet_107), .o(newNet_108) );
na02f80 g1931_u0 ( .a(n_169), .b(n_296), .o(n_294) );
ao12f80 g1859_u0 ( .a(n_391), .b(n_88), .c(n_390), .o(n_421) );
no02f80 g1725_u0 ( .a(n_385), .b(n_416), .o(n_428) );
in01f80 g2149_u0 ( .a(n_306), .o(n_70) );
in01f80 i_rx_phy_rxd_s1_reg_u1 ( .a(i_rx_phy_rxd_s1_reg_Q), .o(i_rx_phy_rxd_s1) );
na02f80 g1782_u3 ( .a(g1782_da), .b(g1782_db), .o(n_452) );
na02f80 g1778_u3 ( .a(g1778_da), .b(g1778_db), .o(n_456) );
in01f80 newInst_73 ( .a(newNet_72), .o(newNet_73) );
in01f80 i_tx_phy_hold_reg_d_reg_5__u1 ( .a(i_tx_phy_hold_reg_d_reg_5__Q), .o(i_tx_phy_hold_reg_d_15) );
na02f80 g1907_u0 ( .a(n_106), .b(n_103), .o(n_268) );
na02f80 g2015_u0 ( .a(n_277), .b(n_48), .o(n_280) );
ao12f80 g1846_u0 ( .a(n_961), .b(n_354), .c(n_334), .o(n_405) );
in01f80 g2035_u1 ( .a(g2035_p), .o(n_126) );
in01f80 g1742_u1 ( .a(g1742_p), .o(n_483) );
in01f80 newInst_65 ( .a(newNet_37), .o(newNet_65) );
na02f80 g1813_u0 ( .a(n_434), .b(DataOut_i_7_), .o(n_462) );
in01f80 g1964_u0 ( .a(n_289), .o(n_290) );
in01f80 newInst_150 ( .a(newNet_149), .o(newNet_150) );
no02f80 g2130_u0 ( .a(n_884), .b(n_509), .o(g2130_p) );
in01f80 newInst_142 ( .a(newNet_141), .o(newNet_142) );
ms00f80 i_rx_phy_fs_ce_reg_u0 ( .ck(newNet_284), .d(i_rx_phy_fs_ce_r2), .o(n_885) );
ao22s80 g1879_u0 ( .a(n_225), .b(i_tx_phy_sd_nrzi_o), .c(n_873), .d(txdp), .o(n_308) );
ms00f80 i_rx_phy_hold_reg_reg_1__u0 ( .ck(newNet_272), .d(DataIn_o_2_), .o(DataIn_o_1_) );
na02f80 g2053_u0 ( .a(n_804), .b(n_168), .o(n_169) );
in01f80 g1857_u1 ( .a(g1857_p), .o(n_433) );
in01f80 g1738_u1 ( .a(g1738_p), .o(n_487) );
in01f80 newInst_12 ( .a(newNet_11), .o(newNet_12) );
na02f80 g23_u0 ( .a(n_604), .b(n_926), .o(n_938) );
in01f80 newInst_88 ( .a(newNet_87), .o(newNet_88) );
na02f80 g1958_u0 ( .a(n_574), .b(n_841), .o(n_257) );
in01f80 newInst_134 ( .a(newNet_125), .o(newNet_134) );
in01f80 newInst_287 ( .a(newNet_286), .o(newNet_287) );
in01f80 newInst_226 ( .a(newNet_225), .o(newNet_226) );
ms00f80 i_rx_phy_rx_en_reg_u0 ( .ck(newNet_233), .d(txoe), .o(i_rx_phy_rx_en) );
in01f80 newInst_17 ( .a(newNet_16), .o(newNet_17) );
no02f80 g2506_u0 ( .a(n_910), .b(n_460), .o(g2506_p) );
in01f80 newInst_232 ( .a(newNet_231), .o(newNet_232) );
in01f80 newInst_21 ( .a(newNet_20), .o(newNet_21) );
ms00f80 i_tx_phy_hold_reg_reg_2__u0 ( .ck(newNet_95), .d(n_486), .o(i_tx_phy_hold_reg_5) );
in01f80 g2050_u1 ( .a(g2050_p), .o(n_172) );
in01f80 newInst_260 ( .a(newNet_259), .o(newNet_260) );
in01f80 newInst_111 ( .a(newNet_110), .o(newNet_111) );
in01f80 newInst_49 ( .a(newNet_48), .o(newNet_49) );
in01f80 newInst_149 ( .a(newNet_148), .o(newNet_149) );
no02f80 FE_RC_1_0 ( .a(FE_RN_2_0), .b(FE_RN_1_0), .o(FE_RN_0_0) );
in01f80 newInst_231 ( .a(newNet_230), .o(newNet_231) );
in01f80 newInst_181 ( .a(newNet_180), .o(newNet_181) );
in01f80 g2637_u0 ( .a(n_794), .o(n_940) );
na02f80 g1873_u0 ( .a(n_280), .b(n_273), .o(n_338) );
in01f80 newInst_300 ( .a(newNet_105), .o(newNet_300) );
na02f80 g2030_u0 ( .a(i_tx_phy_hold_reg_d_12), .b(n_124), .o(n_97) );
ao12f80 g1986_u0 ( .a(n_241), .b(n_384), .c(n_240), .o(n_313) );
in01f80 newInst_80 ( .a(newNet_79), .o(newNet_80) );
ms00f80 i_rx_phy_one_cnt_reg_1__u0 ( .ck(newNet_242), .d(n_427), .o(i_rx_phy_one_cnt_1_) );
na02f80 g1741_u0 ( .a(n_454), .b(n_974), .o(g1741_p) );
ao12f80 g2069_u1 ( .a(g2069_p), .b(n_115), .c(i_tx_phy_one_cnt_0_), .o(n_116) );
in01f80 g1740_u1 ( .a(g1740_p), .o(n_485) );
in01f80 newInst_242 ( .a(newNet_241), .o(newNet_242) );
in01f80 newInst_214 ( .a(newNet_24), .o(newNet_214) );
in01f80 g22_u0 ( .a(n_852), .o(n_988) );
in01f80 newInst_20 ( .a(newNet_19), .o(newNet_20) );
ms00f80 i_tx_phy_TxReady_o_reg_u0 ( .ck(newNet_155), .d(n_392), .o(TxReady_o) );
oa12f80 g1745_u0 ( .a(n_252), .b(n_311), .c(n_384), .o(n_380) );
in01f80 newInst_97 ( .a(newNet_96), .o(newNet_97) );
ms00f80 i_rx_phy_rx_valid1_reg_u0 ( .ck(newNet_232), .d(n_431), .o(i_rx_phy_rx_valid1) );
na02f80 g1897_u0 ( .a(n_764), .b(i_rx_phy_shift_en), .o(g1897_u0_o) );
na03f80 g42_u0 ( .a(n_737), .b(n_593), .c(n_590), .o(n_968) );
in01f80 newInst_306 ( .a(newNet_305), .o(newNet_306) );
in01f80 newInst_165 ( .a(newNet_164), .o(newNet_165) );
in01f80 newInst_29 ( .a(newNet_28), .o(newNet_29) );
in01f80 newInst_225 ( .a(newNet_13), .o(newNet_225) );
no02f80 g11_u0 ( .a(n_980), .b(n_947), .o(g11_p) );
in01f80 g2195_u0 ( .a(rst), .o(n_318) );
na02f80 g1951_u0 ( .a(n_182), .b(n_885), .o(n_343) );
no02f80 g2465_u0 ( .a(n_318), .b(n_540), .o(n_706) );
na03f80 g1924_u0 ( .a(n_325), .b(n_53), .c(g2674_p), .o(n_352) );
ms00f80 i_rx_phy_rx_valid_r_reg_u0 ( .ck(newNet_228), .d(n_433), .o(i_rx_phy_rx_valid_r) );
ao22s80 g2062_u0 ( .a(i_tx_phy_append_eop_sync4), .b(n_852), .c(n_48), .d(g2674_p), .o(n_204) );
in01f80 g1954_u0 ( .a(n_258), .o(n_259) );
na02f80 g2063_u3 ( .a(g2063_da), .b(g2063_db), .o(n_203) );
in01f80 newInst_210 ( .a(newNet_209), .o(newNet_210) );
no02f80 g2392_u0 ( .a(n_932), .b(n_952), .o(n_590) );
in01f80 newInst_298 ( .a(newNet_297), .o(newNet_298) );
ms00f80 i_tx_phy_append_eop_sync1_reg_u0 ( .ck(newNet_145), .d(n_317), .o(i_tx_phy_append_eop_sync1) );
in01f80 g2257_u0 ( .a(rst_cnt_3_), .o(n_69) );
na02f80 g2108_u0 ( .a(i_rx_phy_rx_valid_r), .b(n_882), .o(g2108_p) );
na02f80 g2459_u0 ( .a(n_910), .b(n_980), .o(n_697) );
ms00f80 i_rx_phy_fs_ce_r2_reg_u0 ( .ck(newNet_287), .d(i_rx_phy_fs_ce_r1), .o(i_rx_phy_fs_ce_r2) );
na02f80 g1742_u0 ( .a(n_453), .b(n_974), .o(g1742_p) );
in01f80 newInst_59 ( .a(newNet_58), .o(newNet_59) );
in01f80 newInst_69 ( .a(newNet_68), .o(newNet_69) );
ms00f80 i_tx_phy_append_eop_sync3_reg_u0 ( .ck(newNet_139), .d(n_338), .o(n_224) );
na02f80 g1975_u0 ( .a(i_rx_phy_rxdp_s0), .b(LineState_o_0_), .o(g1975_p) );
in01f80 newInst_10 ( .a(newNet_9), .o(newNet_10) );
in01f80 g1776_u0 ( .a(i_tx_phy_ld_data), .o(g1776_sb) );
in01f80 newInst_255 ( .a(newNet_254), .o(newNet_255) );
in01f80 newInst_216 ( .a(newNet_215), .o(newNet_216) );
in01f80 newInst_168 ( .a(newNet_167), .o(newNet_168) );
na02f80 g2063_u2 ( .a(i_rx_phy_sd_r), .b(n_852), .o(g2063_db) );
in01f80 g1998_u0 ( .a(n_949), .o(n_782) );
in01f80 newInst_129 ( .a(newNet_53), .o(newNet_129) );
in01f80 newInst_28 ( .a(newNet_22), .o(newNet_28) );
in01f80 newInst_263 ( .a(newNet_70), .o(newNet_263) );
na02f80 g1776_u3 ( .a(g1776_da), .b(g1776_db), .o(n_458) );
ms00f80 i_rx_phy_rxd_s1_reg_u0 ( .ck(newNet_213), .d(i_rx_phy_rxd_s0), .o(i_rx_phy_rxd_s1_reg_Q) );
ao12f80 g2057_u1 ( .a(g2057_p), .b(i_rx_phy_sd_r), .c(n_243), .o(n_122) );
ms00f80 i_tx_phy_tx_ip_sync_reg_u0 ( .ck(newNet_41), .d(n_319), .o(n_238) );
ms00f80 i_rx_phy_hold_reg_reg_0__u0 ( .ck(newNet_274), .d(DataIn_o_1_), .o(DataIn_o_0_) );
in01f80 newInst_53 ( .a(newNet_52), .o(newNet_53) );
in01f80 newInst_33 ( .a(newNet_32), .o(newNet_33) );
in01f80 g2095_u0 ( .a(n_103), .o(n_384) );
in01f80 g1923_u1 ( .a(g1923_p), .o(n_390) );
na02f80 g1780_u3 ( .a(g1780_da), .b(g1780_db), .o(n_454) );
in01f80 newInst_114 ( .a(newNet_113), .o(newNet_114) );
in01f80 newInst_19 ( .a(newNet_3), .o(newNet_19) );
in01f80 g2270_u0 ( .a(n_353), .o(n_18) );
in01f80 newInst_282 ( .a(newNet_281), .o(newNet_282) );
oa12f80 g1854_u0 ( .a(n_133), .b(n_231), .c(i_tx_phy_hold_reg_d_13), .o(n_232) );
no02f80 g2122_u0 ( .a(n_52), .b(n_28), .o(n_58) );
na02f80 g2043_u0 ( .a(n_948), .b(n_794), .o(n_175) );
na02f80 g2632_u0 ( .a(n_64), .b(i_tx_phy_sft_done), .o(n_932) );
no02f80 g1981_u0 ( .a(LineState_o_0_), .b(LineState_o_1_), .o(n_191) );
ms00f80 i_rx_phy_hold_reg_reg_6__u0 ( .ck(newNet_253), .d(DataIn_o_7_), .o(DataIn_o_6_) );
na03f80 g1982_u0 ( .a(n_125), .b(i_tx_phy_hold_reg_d_17), .c(i_tx_phy_bit_cnt_2_), .o(n_133) );
na02f80 g35_u0 ( .a(n_722), .b(n_926), .o(n_741) );
na02f80 g2109_u0 ( .a(n_115), .b(n_873), .o(n_154) );
in01f80 g1975_u1 ( .a(g1975_p), .o(n_226) );
in01f80 newInst_274 ( .a(newNet_273), .o(newNet_274) );
in01f80 newInst_157 ( .a(newNet_156), .o(newNet_157) );
in01f80 newInst_197 ( .a(newNet_182), .o(newNet_197) );
na03f80 g1927_u0 ( .a(n_296), .b(i_tx_phy_sd_raw_o), .c(n_85), .o(n_297) );
in01f80 g2648_u0 ( .a(i_tx_phy_state_1_), .o(n_735) );
in01f80 g2227_u0 ( .a(n_980), .o(n_91) );
ms00f80 i_tx_phy_txdp_reg_u0 ( .ck(newNet_35), .d(n_366), .o(txdp) );
no02f80 g2069_u0 ( .a(n_115), .b(i_tx_phy_one_cnt_0_), .o(g2069_p) );
ao22s80 g1937_u0 ( .a(n_100), .b(n_885), .c(i_tx_phy_sd_nrzi_o), .d(n_873), .o(n_195) );
in01f80 newInst_122 ( .a(newNet_45), .o(newNet_122) );
in01f80 newInst_295 ( .a(newNet_294), .o(newNet_295) );
in01f80 g2604_u0 ( .a(n_929), .o(n_888) );
in01f80 g2413_u1 ( .a(g2413_p), .o(n_628) );
oa12f80 g2655_u0 ( .a(n_965), .b(n_734), .c(n_937), .o(n_966) );
ms00f80 i_tx_phy_hold_reg_d_reg_5__u0 ( .ck(newNet_106), .d(i_tx_phy_hold_reg_8), .o(i_tx_phy_hold_reg_d_reg_5__Q) );
in01f80 newInst_176 ( .a(newNet_175), .o(newNet_176) );
in01f80 newInst_109 ( .a(newNet_108), .o(newNet_109) );
ao12f80 g1726_u0 ( .a(n_384), .b(n_292), .c(n_256), .o(n_370) );
na02f80 g1697_u0 ( .a(n_490), .b(n_786), .o(n_506) );
na02f80 g2622_u0 ( .a(n_920), .b(n_921), .o(n_922) );
in01f80 newInst_125 ( .a(newNet_124), .o(newNet_125) );
ms00f80 i_rx_phy_rxdn_s0_reg_u0 ( .ck(newNet_206), .d(rxdn), .o(i_rx_phy_rxdn_s0) );
na02f80 g2431_u0 ( .a(n_749), .b(n_754), .o(n_660) );
in01f80 g2117_u0 ( .a(n_164), .o(n_108) );
ao12f80 g1983_u0 ( .a(n_167), .b(n_192), .c(i_tx_phy_hold_reg_d), .o(n_255) );
no02f80 g2024_u0 ( .a(i_rx_phy_rxd_s0), .b(n_130), .o(n_127) );
in01f80 g2272_u0 ( .a(i_tx_phy_one_cnt_2_), .o(n_33) );
in01f80 newInst_42 ( .a(newNet_25), .o(newNet_42) );
na02f80 g2635_u0 ( .a(n_938), .b(n_943), .o(n_944) );
in01f80 newInst_135 ( .a(newNet_134), .o(newNet_135) );
in01f80 newInst_4 ( .a(newNet_3), .o(newNet_4) );
ms00f80 i_tx_phy_tx_ip_reg_u0 ( .ck(newNet_45), .d(n_976), .o(i_tx_phy_tx_ip) );
in01f80 g2610_u0 ( .a(n_929), .o(n_894) );
no02f80 g1806_u0 ( .a(n_232), .b(n_300), .o(n_369) );
in01f80 g1734_u0 ( .a(n_753), .o(n_460) );
in01f80 g2091_u1 ( .a(g2091_p), .o(n_183) );
in01f80 newInst_243 ( .a(newNet_31), .o(newNet_243) );
in01f80 newInst_64 ( .a(newNet_63), .o(newNet_64) );
no02f80 g1923_u0 ( .a(n_312), .b(n_540), .o(g1923_p) );
na02f80 g1855_u1 ( .a(rst_cnt_4_), .b(g1855_sb), .o(g1855_da) );
na02f80 g1780_u2 ( .a(i_tx_phy_hold_reg_7), .b(i_tx_phy_ld_data), .o(g1780_db) );
in01f80 newInst_102 ( .a(newNet_64), .o(newNet_102) );
ao22s80 g2059_u0 ( .a(i_tx_phy_tx_ip), .b(n_885), .c(n_238), .d(n_984), .o(n_239) );
na02f80 g1914_u0 ( .a(n_296), .b(n_56), .o(n_301) );
in01f80 g1746_u0 ( .a(n_479), .o(n_505) );
na02f80 g2653_u0 ( .a(i_rx_phy_shift_en), .b(rst), .o(n_961) );
in01f80 newInst_288 ( .a(newNet_120), .o(newNet_288) );
na03f80 g26_u0 ( .a(n_443), .b(RxActive_o), .c(rst), .o(n_708) );
ms00f80 i_rx_phy_fs_state_reg_2__u0 ( .ck(newNet_276), .d(n_758), .o(i_rx_phy_fs_state_2_) );
in01f80 g2112_u0 ( .a(n_389), .o(n_81) );
in01f80 i_tx_phy_hold_reg_d_reg_3__u1 ( .a(i_tx_phy_hold_reg_d_reg_3__Q), .o(i_tx_phy_hold_reg_d_13) );
ms00f80 i_tx_phy_sd_bs_o_reg_u0 ( .ck(newNet_64), .d(n_361), .o(i_tx_phy_sd_bs_o) );
na02f80 g1868_u0 ( .a(n_116), .b(n_340), .o(n_341) );
no02f80 g1962_u0 ( .a(n_239), .b(n_318), .o(n_319) );
no02f80 g1718_u0 ( .a(n_916), .b(n_467), .o(n_783) );
in01f80 newInst_233 ( .a(newNet_7), .o(newNet_233) );
no02f80 g1967_u0 ( .a(n_235), .b(FE_RN_2_0), .o(n_316) );
na02f80 g1855_u2 ( .a(n_11), .b(n_274), .o(g1855_db) );
in01f80 newInst_81 ( .a(newNet_80), .o(newNet_81) );
ms00f80 i_rx_phy_sd_nrzi_reg_u0 ( .ck(newNet_178), .d(n_365), .o(i_rx_phy_sd_nrzi) );
in01f80 g24_u0 ( .a(n_941), .o(n_942) );
in01f80 g2103_u1 ( .a(g2103_p), .o(n_277) );
in01f80 newInst_18 ( .a(newNet_17), .o(newNet_18) );
ao12f80 g1775_u0 ( .a(n_368), .b(n_384), .c(n_306), .o(n_385) );
na02f80 g1955_u0 ( .a(n_182), .b(i_tx_phy_sd_raw_o), .o(n_258) );
na02m80 FE_RC_0_0 ( .a(FE_RN_0_0), .b(n_629), .o(n_632) );
in01f80 g1952_u0 ( .a(n_324), .o(n_325) );
na03f80 g1774_u0 ( .a(n_425), .b(n_175), .c(n_949), .o(n_440) );
ao12f80 g1870_u0 ( .a(n_343), .b(n_126), .c(n_231), .o(n_339) );
in01f80 newInst_63 ( .a(newNet_31), .o(newNet_63) );
in01f80 newInst_241 ( .a(newNet_240), .o(newNet_241) );
ao12f80 g2056_u0 ( .a(n_164), .b(n_888), .c(n_737), .o(n_165) );
na02f80 g2104_u0 ( .a(i_rx_phy_one_cnt_0_), .b(n_873), .o(n_157) );
ms00f80 i_tx_phy_hold_reg_reg_5__u0 ( .ck(newNet_81), .d(n_483), .o(i_tx_phy_hold_reg_8) );
ao22s80 g1933_u0 ( .a(n_122), .b(n_266), .c(n_150), .d(i_rx_phy_sd_nrzi), .o(n_267) );
in01f80 newInst_303 ( .a(newNet_280), .o(newNet_303) );
in01f80 newInst_50 ( .a(newNet_49), .o(newNet_50) );
in01f80 newInst_297 ( .a(newNet_296), .o(newNet_297) );
na02f80 g1762_u0 ( .a(i_rx_phy_rx_valid_r), .b(n_446), .o(n_443) );
in01f80 newInst_167 ( .a(newNet_132), .o(newNet_167) );
ms00f80 i_rx_phy_dpll_state_reg_0__u0 ( .ck(newNet_299), .d(n_449), .o(i_rx_phy_dpll_state_0_) );
in01f80 g1828_u0 ( .a(i_tx_phy_ld_data), .o(n_434) );
in01f80 g2527_u0 ( .a(n_788), .o(n_786) );
no02f80 g1811_u0 ( .a(n_377), .b(n_400), .o(n_415) );
ao12f80 g1838_u0 ( .a(n_416), .b(n_251), .c(n_268), .o(n_367) );
na02f80 g1810_u0 ( .a(n_197), .b(n_69), .o(n_256) );
in01f80 newInst_307 ( .a(newNet_72), .o(newNet_307) );
in01f80 newInst_23 ( .a(newNet_15), .o(newNet_23) );
in01f80 g2273_u0 ( .a(n_243), .o(n_130) );
na03f80 g2482_u0 ( .a(n_439), .b(n_794), .c(n_90), .o(n_726) );
in01f80 newInst_281 ( .a(newNet_119), .o(newNet_281) );
in01f80 newInst_257 ( .a(newNet_256), .o(newNet_257) );
in01f80 newInst_202 ( .a(newNet_189), .o(newNet_202) );
in01f80 g2161_u0 ( .a(i_tx_phy_append_eop_sync2), .o(n_12) );
ao12f80 g1695_u0 ( .a(FE_RN_2_0), .b(n_704), .c(n_935), .o(n_459) );
na02f80 g2088_u0 ( .a(i_tx_phy_one_cnt_0_), .b(n_873), .o(n_161) );
no02f80 g1865_u0 ( .a(n_274), .b(n_11), .o(n_275) );
na02f80 g1872_u0 ( .a(n_227), .b(i_rx_phy_rxdp_s_r), .o(n_309) );
no02f80 g2652_u0 ( .a(n_984), .b(n_324), .o(n_958) );
in01f80 newInst_121 ( .a(newNet_7), .o(newNet_121) );
na02f80 g1778_u2 ( .a(i_tx_phy_hold_reg_5), .b(i_tx_phy_ld_data), .o(g1778_db) );
in01f80 newInst_30 ( .a(newNet_29), .o(newNet_30) );
na02f80 g2114_u0 ( .a(n_852), .b(txdn), .o(n_153) );
ao22s80 g2623_u0 ( .a(n_919), .b(n_945), .c(n_722), .d(n_916), .o(n_920) );
in01f80 newInst_254 ( .a(newNet_112), .o(newNet_254) );
na02f80 g1776_u2 ( .a(i_tx_phy_hold_reg), .b(i_tx_phy_ld_data), .o(g1776_db) );
na02f80 g1922_u0 ( .a(n_71), .b(n_66), .o(n_274) );
na02f80 g2656_u0 ( .a(n_583), .b(n_737), .o(n_967) );
no02f80 g2124_u0 ( .a(i_rx_phy_dpll_state_1_), .b(i_rx_phy_dpll_state_0_), .o(n_88) );
no02f80 g2479_u0 ( .a(n_788), .b(n_697), .o(n_722) );
in01f80 g2084_u0 ( .a(i_rx_phy_rxd_r), .o(n_244) );
ms00f80 i_tx_phy_sd_nrzi_o_reg_u0 ( .ck(newNet_62), .d(n_276), .o(i_tx_phy_sd_nrzi_o) );
in01f80 newInst_71 ( .a(newNet_66), .o(newNet_71) );
in01f80 i_rx_phy_rxdn_s_r_reg_u1 ( .a(i_rx_phy_rxdn_s_r_reg_Q), .o(i_rx_phy_rxdn_s_r) );
na02f80 g2090_u0 ( .a(i_tx_phy_append_eop), .b(n_12), .o(n_63) );
na03f80 g1925_u0 ( .a(n_350), .b(n_583), .c(n_800), .o(n_351) );
ms00f80 i_tx_phy_append_eop_reg_u0 ( .ck(newNet_150), .d(n_409), .o(i_tx_phy_append_eop) );
na03f80 g58_u0 ( .a(n_788), .b(n_112), .c(n_919), .o(n_921) );
na02f80 g1777_u2 ( .a(i_tx_phy_hold_reg_4), .b(i_tx_phy_ld_data), .o(g1777_db) );
in01f80 g41_u1 ( .a(g41_p), .o(n_700) );
in01f80 newInst_248 ( .a(newNet_247), .o(newNet_248) );
ao12f80 g2501_u0 ( .a(n_318), .b(n_755), .c(n_756), .o(n_758) );
in01f80 newInst_153 ( .a(newNet_152), .o(newNet_153) );
in01f80 newInst_209 ( .a(newNet_208), .o(newNet_209) );
ms00f80 i_rx_phy_byte_err_reg_u0 ( .ck(newNet_301), .d(n_499), .o(i_rx_phy_byte_err_reg_Q) );
ao12f80 g1851_u0 ( .a(FE_RN_2_0), .b(n_267), .c(RxActive_o), .o(n_365) );
in01f80 newInst_179 ( .a(newNet_157), .o(newNet_179) );
in01f80 newInst_101 ( .a(newNet_14), .o(newNet_101) );
in01f80 newInst_62 ( .a(newNet_53), .o(newNet_62) );
in01f80 g1819_u0 ( .a(n_426), .o(n_446) );
no02f80 g2035_u0 ( .a(n_125), .b(n_124), .o(g2035_p) );
na02f80 g1724_u0 ( .a(n_919), .b(n_914), .o(n_492) );
in01f80 newInst_106 ( .a(newNet_20), .o(newNet_106) );
ao12f80 g1853_u0 ( .a(FE_RN_2_0), .b(n_153), .c(n_265), .o(n_364) );
ms00f80 i_rx_phy_rxdn_s1_reg_u0 ( .ck(newNet_201), .d(i_rx_phy_rxdn_s0), .o(LineState_o_1_) );
in01f80 newInst_1 ( .a(newNet_0), .o(newNet_1) );
ms00f80 i_tx_phy_append_eop_sync4_reg_u0 ( .ck(newNet_138), .d(n_288), .o(i_tx_phy_append_eop_sync4) );
ms00f80 i_rx_phy_rxdn_s_reg_u0 ( .ck(newNet_196), .d(n_310), .o(i_rx_phy_rxdn_s) );
in01f80 newInst_140 ( .a(newNet_66), .o(newNet_140) );
ms00f80 rst_cnt_reg_0__u0 ( .ck(newNet_18), .d(n_362), .o(rst_cnt_0_) );
in01f80 g2157_u0 ( .a(i_rx_phy_dpll_state_0_), .o(n_60) );
ao12f80 g2066_u1 ( .a(g2066_p), .b(n_105), .c(n_240), .o(n_106) );
in01f80 newInst_89 ( .a(newNet_88), .o(newNet_89) );
na02f80 g1782_u1 ( .a(DataOut_i_6_), .b(g1782_sb), .o(g1782_da) );
oa12f80 g2058_u0 ( .a(n_35), .b(i_tx_phy_sd_bs_o), .c(i_tx_phy_sd_nrzi_o), .o(n_100) );
in01f80 newInst_273 ( .a(newNet_78), .o(newNet_273) );
na02f80 g1942_u0 ( .a(i_tx_phy_data_done), .b(n_937), .o(g1942_p) );
ms00f80 i_tx_phy_sft_done_r_reg_u0 ( .ck(newNet_60), .d(i_tx_phy_sft_done), .o(i_tx_phy_sft_done_r) );
in01f80 g2385_u1 ( .a(g2385_p), .o(n_567) );
ms00f80 i_tx_phy_hold_reg_reg_4__u0 ( .ck(newNet_86), .d(n_484), .o(i_tx_phy_hold_reg_7) );
na02f80 g1681_u0 ( .a(n_493), .b(n_440), .o(n_511) );
in01f80 newInst_234 ( .a(newNet_33), .o(newNet_234) );
na02f80 g2495_u0 ( .a(n_467), .b(n_914), .o(n_742) );
no02f80 g1808_u0 ( .a(n_307), .b(n_384), .o(n_368) );
in01f80 g2020_u0 ( .a(n_759), .o(n_248) );
in01f80 newInst_272 ( .a(newNet_271), .o(newNet_272) );
ms00f80 i_rx_phy_hold_reg_reg_3__u0 ( .ck(newNet_264), .d(DataIn_o_4_), .o(DataIn_o_3_) );
in01f80 newInst_266 ( .a(newNet_265), .o(newNet_266) );
no02f80 g2139_u0 ( .a(n_50), .b(n_49), .o(n_51) );
in01f80 newInst_201 ( .a(newNet_45), .o(newNet_201) );
in01f80 newInst_51 ( .a(newNet_50), .o(newNet_51) );
in01f80 newInst_188 ( .a(newNet_158), .o(newNet_188) );
in01f80 g1830_u0 ( .a(i_rx_phy_rxdn_s), .o(n_424) );
ao12f80 g1821_u0 ( .a(FE_RN_2_0), .b(n_435), .c(n_389), .o(n_436) );
in01f80 newInst_112 ( .a(newNet_111), .o(newNet_112) );
in01f80 newInst_107 ( .a(newNet_49), .o(newNet_107) );
in01f80 g2119_u0 ( .a(n_697), .o(n_90) );
in01f80 newInst_236 ( .a(newNet_235), .o(newNet_236) );
in01f80 newInst_183 ( .a(newNet_182), .o(newNet_183) );
in01f80 newInst_139 ( .a(newNet_68), .o(newNet_139) );
in01f80 newInst_240 ( .a(newNet_51), .o(newNet_240) );
na02f80 g1778_u1 ( .a(DataOut_i_2_), .b(g1778_sb), .o(g1778_da) );
in01f80 newInst_148 ( .a(newNet_147), .o(newNet_148) );
na03f80 g2508_u0 ( .a(n_763), .b(i_rx_phy_rx_valid1), .c(rst), .o(n_767) );
in01f80 g2438_u0 ( .a(n_666), .o(n_665) );
in01f80 newInst_256 ( .a(newNet_255), .o(newNet_256) );
in01f80 newInst_22 ( .a(newNet_21), .o(newNet_22) );
in01f80 g2183_u0 ( .a(n_57), .o(n_15) );
in01f80 i_tx_phy_hold_reg_d_reg_1__u1 ( .a(i_tx_phy_hold_reg_d_reg_1__Q), .o(i_tx_phy_hold_reg_d_11) );
in01f80 g1979_u0 ( .a(n_222), .o(n_223) );
in01f80 g1935_u0 ( .a(n_263), .o(n_293) );
in01f80 newInst_133 ( .a(newNet_125), .o(newNet_133) );
in01f80 newInst_269 ( .a(newNet_268), .o(newNet_269) );
in01f80 newInst_308 ( .a(newNet_307), .o(newNet_308) );
in01f80 g1779_u0 ( .a(i_tx_phy_ld_data), .o(g1779_sb) );
in01f80 g2667_u0 ( .a(n_796), .o(n_794) );
in01f80 newInst_144 ( .a(newNet_143), .o(newNet_144) );
na02f80 g1781_u2 ( .a(i_tx_phy_hold_reg_8), .b(i_tx_phy_ld_data), .o(g1781_db) );
ms00f80 i_tx_phy_hold_reg_d_reg_4__u0 ( .ck(newNet_109), .d(i_tx_phy_hold_reg_7), .o(i_tx_phy_hold_reg_d_14) );
oa12f80 g1744_u0 ( .a(i_rx_phy_se0_r), .b(n_353), .c(i_rx_phy_bit_cnt_2_), .o(n_472) );
in01f80 newInst_195 ( .a(newNet_194), .o(newNet_195) );
in01f80 g12_u0 ( .a(i_rx_phy_rx_en), .o(n_540) );
no02f80 g2054_u0 ( .a(n_168), .b(i_tx_phy_hold_reg_d_11), .o(n_167) );
in01f80 g2258_u0 ( .a(i_rx_phy_se0_s), .o(n_9) );
ao12f80 g1837_u0 ( .a(FE_RN_2_0), .b(n_63), .c(n_968), .o(n_409) );
na03f80 g25_u0 ( .a(n_735), .b(n_952), .c(n_894), .o(n_841) );
in01f80 g2155_u0 ( .a(i_tx_phy_one_cnt_0_), .o(n_50) );
in01f80 newInst_190 ( .a(newNet_189), .o(newNet_190) );
in01f80 newInst_94 ( .a(newNet_93), .o(newNet_94) );
in01f80 newInst_203 ( .a(newNet_202), .o(newNet_203) );
no02f80 g1963_u0 ( .a(n_201), .b(n_318), .o(n_291) );
in01f80 newInst_119 ( .a(newNet_93), .o(newNet_119) );
in01f80 g61_u0 ( .a(n_942), .o(n_919) );
na03f80 g2505_u0 ( .a(n_61), .b(n_426), .c(n_9), .o(n_753) );
in01f80 g2412_u1 ( .a(g2412_p), .o(n_629) );
na02f80 g1900_u0 ( .a(n_118), .b(n_764), .o(n_334) );
na02f80 g2115_u0 ( .a(n_120), .b(n_873), .o(n_152) );
in01f80 g1767_u0 ( .a(n_941), .o(n_467) );
in01f80 newInst_35 ( .a(newNet_34), .o(newNet_35) );
in01f80 g2669_u0 ( .a(i_rx_phy_fs_state_0_), .o(n_980) );
ms00f80 i_tx_phy_hold_reg_d_reg_0__u0 ( .ck(newNet_121), .d(i_tx_phy_hold_reg), .o(i_tx_phy_hold_reg_d) );
na03f80 g1816_u0 ( .a(n_421), .b(n_435), .c(rst), .o(n_449) );
in01f80 newInst_155 ( .a(newNet_154), .o(newNet_155) );
in01f80 newInst_46 ( .a(newNet_14), .o(newNet_46) );
no02f80 g2665_u0 ( .a(n_913), .b(n_981), .o(n_982) );
in01f80 newInst_219 ( .a(newNet_218), .o(newNet_219) );
in01f80 newInst_154 ( .a(newNet_153), .o(newNet_154) );
in01f80 newInst_198 ( .a(newNet_197), .o(newNet_198) );
na02f80 g1980_u0 ( .a(i_rx_phy_rxdn_s0), .b(LineState_o_1_), .o(g1980_p) );
in01f80 newInst_200 ( .a(newNet_199), .o(newNet_200) );
in01f80 newInst_292 ( .a(newNet_291), .o(newNet_292) );
in01f80 newInst_72 ( .a(newNet_7), .o(newNet_72) );
in01f80 g2145_u0 ( .a(n_559), .o(n_48) );
in01f80 newInst_126 ( .a(newNet_125), .o(newNet_126) );
in01f80 g2127_u0 ( .a(n_400), .o(n_85) );
na02f80 g2672_u0 ( .a(n_988), .b(n_989), .o(n_990) );
no02f80 g2050_u0 ( .a(n_804), .b(n_785), .o(g2050_p) );
ao12f80 g1840_u0 ( .a(n_322), .b(n_330), .c(n_952), .o(n_538) );
na02f80 g1906_u0 ( .a(n_191), .b(rst), .o(n_416) );
na02f80 g2385_u0 ( .a(n_885), .b(n_559), .o(g2385_p) );
oa12f80 g1934_u0 ( .a(n_184), .b(n_186), .c(n_48), .o(n_265) );
in01f80 newInst_249 ( .a(newNet_129), .o(newNet_249) );
in01f80 newInst_130 ( .a(newNet_129), .o(newNet_130) );
oa12f80 g1932_u0 ( .a(n_193), .b(n_97), .c(n_804), .o(n_228) );
in01f80 newInst_100 ( .a(newNet_99), .o(newNet_100) );
in01f80 g1741_u1 ( .a(g1741_p), .o(n_484) );
in01f80 newInst_141 ( .a(newNet_140), .o(newNet_141) );
in01f80 newInst_92 ( .a(newNet_91), .o(newNet_92) );
in01f80 newInst_57 ( .a(newNet_56), .o(newNet_57) );
ao12f80 g2657_u0 ( .a(n_318), .b(n_970), .c(n_974), .o(n_976) );
in01f80 g2645_u0 ( .a(n_951), .o(n_952) );
in01f80 FE_RC_2_0 ( .a(n_631), .o(FE_RN_1_0) );
no02f80 g2413_u0 ( .a(n_753), .b(n_727), .o(g2413_p) );
in01f80 newInst_235 ( .a(newNet_234), .o(newNet_235) );
in01f80 newInst_174 ( .a(newNet_38), .o(newNet_174) );
no02f80 g2091_u0 ( .a(phy_tx_mode), .b(n_984), .o(g2091_p) );
na02f80 g1782_u2 ( .a(i_tx_phy_hold_reg_9), .b(i_tx_phy_ld_data), .o(g1782_db) );
na02f80 g2390_u0 ( .a(n_972), .b(n_894), .o(n_574) );
in01f80 newInst_261 ( .a(newNet_260), .o(newNet_261) );
ms00f80 i_rx_phy_rxdp_s_r_reg_u0 ( .ck(newNet_184), .d(n_226), .o(i_rx_phy_rxdp_s_r_reg_Q) );
ao12f80 g1882_u0 ( .a(n_230), .b(n_132), .c(n_306), .o(n_307) );
in01f80 newInst_304 ( .a(newNet_303), .o(newNet_304) );
in01f80 g56_u0 ( .a(n_916), .o(n_926) );
in01f80 g2601_u0 ( .a(n_885), .o(n_884) );
in01f80 newInst_40 ( .a(newNet_16), .o(newNet_40) );
ms00f80 i_rx_phy_rxd_s0_reg_u0 ( .ck(newNet_217), .d(rxd), .o(i_rx_phy_rxd_s0) );
no02f80 g2140_u0 ( .a(n_49), .b(n_33), .o(n_55) );
ao12f80 g1881_u1 ( .a(g1881_p), .b(i_rx_phy_bit_cnt_2_), .c(n_141), .o(n_142) );
na02f80 g1871_u0 ( .a(n_223), .b(i_rx_phy_rxdn_s_r), .o(n_310) );
in01f80 newInst_271 ( .a(newNet_270), .o(newNet_271) );
in01f80 newInst_123 ( .a(newNet_122), .o(newNet_123) );
in01f80 newInst_99 ( .a(newNet_98), .o(newNet_99) );
in01f80 g2573_u0 ( .a(g2674_p), .o(n_852) );
na02f80 g1852_u0 ( .a(n_304), .b(n_360), .o(n_392) );
in01f80 newInst_82 ( .a(newNet_22), .o(newNet_82) );
na02f80 g2513_u0 ( .a(n_58), .b(n_53), .o(n_759) );
ao12f80 g1856_u0 ( .a(n_339), .b(n_343), .c(i_tx_phy_bit_cnt_2_), .o(n_377) );
in01f80 newInst_284 ( .a(newNet_176), .o(newNet_284) );
in01f80 newInst_227 ( .a(newNet_226), .o(newNet_227) );
in01f80 newInst_91 ( .a(newNet_11), .o(newNet_91) );
in01f80 g1942_u1 ( .a(g1942_p), .o(n_350) );
in01f80 newInst_118 ( .a(newNet_117), .o(newNet_118) );
in01f80 newInst_15 ( .a(newNet_14), .o(newNet_15) );
na02f80 g64_u0 ( .a(n_754), .b(n_509), .o(n_924) );
in01f80 g2253_u0 ( .a(n_21), .o(n_240) );
in01f80 newInst_279 ( .a(newNet_278), .o(newNet_279) );
ms00f80 i_rx_phy_dpll_state_reg_1__u0 ( .ck(newNet_295), .d(n_436), .o(i_rx_phy_dpll_state_1_) );
in01f80 g2130_u1 ( .a(g2130_p), .o(n_150) );
in01f80 newInst_160 ( .a(newNet_159), .o(newNet_160) );
ms00f80 i_tx_phy_hold_reg_d_reg_7__u0 ( .ck(newNet_104), .d(i_tx_phy_hold_reg_10), .o(i_tx_phy_hold_reg_d_17) );
na02f80 g2103_u0 ( .a(rst), .b(n_882), .o(g2103_p) );
in01f80 newInst_189 ( .a(newNet_188), .o(newNet_189) );
in01f80 newInst_182 ( .a(newNet_36), .o(newNet_182) );
na03f80 g54_u0 ( .a(n_492), .b(n_217), .c(n_209), .o(n_915) );
na02f80 g2099_u0 ( .a(n_57), .b(i_tx_phy_bit_cnt_0_), .o(n_168) );
na03f80 g2660_u0 ( .a(n_972), .b(n_894), .c(TxValid_i), .o(n_974) );
na02f80 g1918_u0 ( .a(n_353), .b(n_763), .o(n_354) );
na02f80 g2138_u0 ( .a(i_tx_phy_sd_bs_o), .b(i_tx_phy_sd_nrzi_o), .o(n_35) );
in01f80 newInst_246 ( .a(newNet_245), .o(newNet_246) );
ms00f80 i_rx_phy_hold_reg_reg_7__u0 ( .ck(newNet_248), .d(i_rx_phy_sd_nrzi), .o(DataIn_o_7_) );
na02f80 g2477_u0 ( .a(n_741), .b(n_726), .o(n_727) );
in01f80 newInst_138 ( .a(newNet_137), .o(newNet_138) );
in01f80 g2028_u1 ( .a(g2028_p), .o(n_246) );
na03f80 g2464_u0 ( .a(n_706), .b(n_461), .c(n_511), .o(n_707) );
in01f80 i_rx_phy_byte_err_reg_u1 ( .a(i_rx_phy_byte_err_reg_Q), .o(i_rx_phy_byte_err) );
ms00f80 i_rx_phy_fs_state_reg_0__u0 ( .ck(newNet_283), .d(n_529), .o(i_rx_phy_fs_state_0_) );
in01f80 g1777_u0 ( .a(i_tx_phy_ld_data), .o(g1777_sb) );
no02f80 g2066_u0 ( .a(n_105), .b(n_240), .o(g2066_p) );
ms00f80 i_rx_phy_one_cnt_reg_2__u0 ( .ck(newNet_239), .d(n_962), .o(i_rx_phy_one_cnt_2_) );
in01f80 g2643_u0 ( .a(n_796), .o(n_788) );
ao12f80 g1815_u0 ( .a(n_400), .b(n_154), .c(n_341), .o(n_401) );
na04m80 g1880_u0 ( .a(n_323), .b(n_350), .c(n_737), .d(n_108), .o(n_360) );
in01f80 g2174_u0 ( .a(i_tx_phy_append_eop_sync4), .o(n_7) );
in01f80 newInst_187 ( .a(newNet_186), .o(newNet_187) );
in01f80 newInst_245 ( .a(newNet_204), .o(newNet_245) );
in01f80 newInst_32 ( .a(newNet_0), .o(newNet_32) );
in01f80 newInst_79 ( .a(newNet_60), .o(newNet_79) );
na02f80 g1719_u0 ( .a(n_926), .b(n_982), .o(n_480) );
ms00f80 rst_cnt_reg_3__u0 ( .ck(newNet_6), .d(n_417), .o(rst_cnt_3_) );
no02f80 g10_u0 ( .a(n_911), .b(n_913), .o(n_914) );
in01f80 newInst_85 ( .a(newNet_84), .o(newNet_85) );
na03f80 g32_u0 ( .a(n_743), .b(n_938), .c(n_748), .o(n_749) );
in01f80 newInst_270 ( .a(newNet_0), .o(newNet_270) );
in01f80 FE_RC_3_0 ( .a(rst), .o(FE_RN_2_0) );
ao22s80 g2061_u0 ( .a(i_tx_phy_append_eop_sync1), .b(n_885), .c(i_tx_phy_append_eop_sync2), .d(n_864), .o(n_235) );
ao12f80 g1985_u0 ( .a(n_213), .b(n_852), .c(txoe), .o(n_283) );
in01f80 newInst_116 ( .a(newNet_115), .o(newNet_116) );
in01f80 i_rx_phy_sync_err_reg_u1 ( .a(i_rx_phy_sync_err_reg_Q), .o(i_rx_phy_sync_err) );
in01f80 g2278_u0 ( .a(i_rx_phy_one_cnt_0_), .o(n_53) );
in01f80 g1780_u0 ( .a(i_tx_phy_ld_data), .o(g1780_sb) );
in01f80 newInst_60 ( .a(newNet_59), .o(newNet_60) );
in01f80 g2072_u0 ( .a(i_tx_phy_sft_done_r), .o(n_64) );
na02f80 g2389_u0 ( .a(n_840), .b(n_567), .o(n_573) );
na02f80 g2638_u0 ( .a(n_413), .b(n_424), .o(n_941) );
oa12f80 g1978_u0 ( .a(n_927), .b(n_952), .c(n_224), .o(n_539) );
in01f80 g1980_u1 ( .a(g1980_p), .o(n_222) );
in01f80 newInst_196 ( .a(newNet_195), .o(newNet_196) );
in01f80 g2159_u0 ( .a(n_52), .o(n_120) );
in01f80 newInst_186 ( .a(newNet_185), .o(newNet_186) );
in01f80 g2642_u0 ( .a(i_rx_phy_fs_state_2_), .o(n_947) );
in01f80 newInst_103 ( .a(newNet_102), .o(newNet_103) );
in01f80 newInst_218 ( .a(newNet_82), .o(newNet_218) );
in01f80 newInst_159 ( .a(newNet_129), .o(newNet_159) );
ao12f80 g1709_u0 ( .a(n_370), .b(n_384), .c(rst_cnt_3_), .o(n_386) );
no02f80 g2625_u0 ( .a(n_888), .b(n_661), .o(n_927) );
ms00f80 i_tx_phy_ld_data_reg_u0 ( .ck(newNet_73), .d(n_387), .o(i_tx_phy_ld_data_reg_Q) );
in01f80 newInst_58 ( .a(newNet_57), .o(newNet_58) );
in01f80 newInst_43 ( .a(newNet_42), .o(newNet_43) );
in01f80 newInst_26 ( .a(newNet_25), .o(newNet_26) );
ao12f80 g2068_u1 ( .a(g2068_p), .b(n_353), .c(i_rx_phy_bit_cnt_0_), .o(n_118) );
in01f80 g2042_u0 ( .a(n_175), .o(n_176) );
in01f80 newInst_16 ( .a(newNet_15), .o(newNet_16) );
na02f80 g1814_u0 ( .a(i_tx_phy_hold_reg_10), .b(i_tx_phy_ld_data), .o(n_450) );
no02f80 g2113_u0 ( .a(i_rx_phy_dpll_state_1_), .b(n_60), .o(g2113_p) );
no02f80 g1817_u0 ( .a(n_666), .b(n_540), .o(n_413) );
na03f80 g1973_u0 ( .a(i_tx_phy_hold_reg_d_14), .b(n_192), .c(i_tx_phy_bit_cnt_2_), .o(n_193) );
in01f80 g2487_u0 ( .a(n_735), .o(n_734) );
in01f80 newInst_278 ( .a(newNet_277), .o(newNet_278) );
in01f80 newInst_221 ( .a(newNet_220), .o(newNet_221) );
no02f80 g2412_u0 ( .a(n_481), .b(n_628), .o(g2412_p) );
in01f80 newInst_169 ( .a(newNet_168), .o(newNet_169) );
in01f80 newInst_131 ( .a(newNet_130), .o(newNet_131) );
ms00f80 i_tx_phy_bit_cnt_reg_1__u0 ( .ck(newNet_132), .d(n_394), .o(i_tx_phy_bit_cnt_1_) );
in01f80 newInst_13 ( .a(newNet_12), .o(newNet_13) );
in01f80 newInst_37 ( .a(newNet_36), .o(newNet_37) );
in01f80 g1739_u1 ( .a(g1739_p), .o(n_486) );
no02f80 g2040_u0 ( .a(n_384), .b(n_240), .o(n_241) );
in01f80 newInst_146 ( .a(newNet_104), .o(newNet_146) );
no02f80 g2010_u0 ( .a(n_185), .b(i_tx_phy_sd_nrzi_o), .o(n_186) );
in01f80 newInst_296 ( .a(newNet_91), .o(newNet_296) );
in01f80 g13_u0 ( .a(n_794), .o(n_913) );
in01f80 g2128_u1 ( .a(g2128_p), .o(n_400) );
in01f80 g2504_u0 ( .a(n_753), .o(n_754) );
in01f80 g1653_u0 ( .a(n_632), .o(n_529) );
no02f80 g2137_u0 ( .a(n_53), .b(n_52), .o(n_54) );
in01f80 g2676_u0 ( .a(n_885), .o(n_984) );
in01f80 g51_u0 ( .a(n_583), .o(n_588) );
ms00f80 i_tx_phy_bit_cnt_reg_2__u0 ( .ck(newNet_128), .d(n_415), .o(i_tx_phy_bit_cnt_2_) );
na02f80 g2011_u0 ( .a(n_384), .b(rst_cnt_4_), .o(n_252) );
na02f80 g2677_u0 ( .a(n_710), .b(n_509), .o(n_989) );
na02f80 g2658_u0 ( .a(n_559), .b(i_tx_phy_tx_ip), .o(n_970) );
in01f80 newInst_104 ( .a(newNet_103), .o(newNet_104) );
ms00f80 i_tx_phy_one_cnt_reg_1__u0 ( .ck(newNet_2), .d(n_401), .o(i_tx_phy_one_cnt_1_) );
no02f80 g1707_u0 ( .a(n_472), .b(n_444), .o(n_499) );
no02f80 g1968_u0 ( .a(n_204), .b(FE_RN_2_0), .o(n_288) );
na02f80 g2630_u0 ( .a(n_965), .b(n_932), .o(n_933) );
in01f80 g2661_u0 ( .a(n_971), .o(n_972) );
in01f80 newInst_207 ( .a(newNet_180), .o(newNet_207) );
in01f80 newInst_283 ( .a(newNet_282), .o(newNet_283) );
in01f80 newInst_177 ( .a(newNet_176), .o(newNet_177) );
no02f80 g2651_u0 ( .a(n_139), .b(n_54), .o(g2651_p) );
na02f80 g2668_u0 ( .a(n_980), .b(i_rx_phy_fs_state_2_), .o(n_981) );
in01f80 g1974_u0 ( .a(n_226), .o(n_227) );
in01f80 g1733_u0 ( .a(n_753), .o(n_461) );
in01f80 newInst_83 ( .a(newNet_82), .o(newNet_83) );
no02f80 g2397_u0 ( .a(n_952), .b(n_735), .o(n_598) );
ms00f80 i_tx_phy_hold_reg_reg_0__u0 ( .ck(newNet_101), .d(n_489), .o(i_tx_phy_hold_reg) );
na02f80 g2503_u0 ( .a(n_480), .b(n_742), .o(n_752) );
no02f80 g1884_u0 ( .a(i_tx_phy_one_cnt_2_), .b(n_51), .o(g1884_p) );
na02f80 g2116_u0 ( .a(n_57), .b(n_56), .o(g2116_p) );
ms00f80 i_tx_phy_sft_done_reg_u0 ( .ck(newNet_55), .d(n_293), .o(i_tx_phy_sft_done) );
na02f80 g1760_u0 ( .a(n_446), .b(RxActive_o), .o(n_444) );
na02f80 g1965_u0 ( .a(n_965), .b(n_937), .o(g1965_p) );
in01f80 newInst_124 ( .a(newNet_121), .o(newNet_124) );
no02f80 g2028_u0 ( .a(n_244), .b(n_243), .o(g2028_p) );
in01f80 newInst_259 ( .a(newNet_258), .o(newNet_259) );
na02f80 g2671_u0 ( .a(n_990), .b(n_991), .o(n_992) );
in01f80 newInst_313 ( .a(newNet_312), .o(newNet_313) );
na02f80 g2012_u0 ( .a(n_224), .b(n_183), .o(n_184) );
na02f80 g2093_u0 ( .a(n_910), .b(n_91), .o(n_111) );
ms00f80 i_tx_phy_hold_reg_reg_6__u0 ( .ck(newNet_78), .d(n_482), .o(i_tx_phy_hold_reg_9) );
ms00f80 i_rx_phy_sync_err_reg_u0 ( .ck(newNet_158), .d(n_925), .o(i_rx_phy_sync_err_reg_Q) );
in01f80 g2664_u0 ( .a(n_974), .o(n_977) );
in01f80 g1959_u0 ( .a(n_573), .o(n_322) );
ms00f80 i_tx_phy_hold_reg_d_reg_3__u0 ( .ck(newNet_114), .d(i_tx_phy_hold_reg_6), .o(i_tx_phy_hold_reg_d_reg_3__Q) );
in01f80 newInst_110 ( .a(newNet_71), .o(newNet_110) );
ms00f80 i_tx_phy_hold_reg_reg_1__u0 ( .ck(newNet_100), .d(n_487), .o(i_tx_phy_hold_reg_4) );
in01f80 g2218_u0 ( .a(n_49), .o(n_115) );
in01f80 g1965_u1 ( .a(g1965_p), .o(n_289) );
in01f80 i_tx_phy_hold_reg_d_reg_6__u1 ( .a(i_tx_phy_hold_reg_d_reg_6__Q), .o(n_785) );
na02f80 g2463_u0 ( .a(n_707), .b(n_708), .o(n_709) );
in01f80 newInst_237 ( .a(newNet_236), .o(newNet_237) );
in01f80 newInst_137 ( .a(newNet_136), .o(newNet_137) );
no02f80 g33_u0 ( .a(i_tx_phy_data_done), .b(n_929), .o(n_593) );
no02f80 g41_u0 ( .a(n_588), .b(n_888), .o(g41_p) );
na02f80 g15_u0 ( .a(n_948), .b(n_796), .o(g15_p) );
in01f80 newInst_24 ( .a(newNet_23), .o(newNet_24) );
ms00f80 i_rx_phy_hold_reg_reg_2__u0 ( .ck(newNet_269), .d(DataIn_o_3_), .o(DataIn_o_2_) );
na02f80 g1876_u0 ( .a(n_278), .b(n_297), .o(n_361) );
in01f80 newInst_291 ( .a(newNet_224), .o(newNet_291) );
in01f80 newInst_277 ( .a(newNet_271), .o(newNet_277) );
in01f80 newInst_86 ( .a(newNet_85), .o(newNet_86) );
in01f80 newInst_117 ( .a(newNet_116), .o(newNet_117) );
na02f80 g2016_u0 ( .a(n_384), .b(n_105), .o(n_251) );
in01f80 g2634_u0 ( .a(n_932), .o(n_937) );
ms00f80 i_rx_phy_bit_cnt_reg_1__u0 ( .ck(newNet_311), .d(n_405), .o(n_353) );
no02f80 g2131_u0 ( .a(n_70), .b(n_69), .o(n_71) );
na02f80 g1913_u0 ( .a(n_343), .b(i_tx_phy_bit_cnt_0_), .o(n_332) );
in01f80 newInst_48 ( .a(newNet_24), .o(newNet_48) );
na02f80 g1743_u0 ( .a(n_452), .b(n_974), .o(g1743_p) );
in01f80 g2141_u1 ( .a(g2141_p), .o(n_185) );
in01f80 newInst_171 ( .a(newNet_170), .o(newNet_171) );
ao22s80 g2624_u0 ( .a(n_927), .b(n_928), .c(n_934), .d(n_929), .o(n_935) );
no02f80 g1680_u0 ( .a(n_386), .b(n_416), .o(n_417) );
ms00f80 i_rx_phy_bit_cnt_reg_2__u0 ( .ck(newNet_306), .d(n_414), .o(i_rx_phy_bit_cnt_2_) );
in01f80 g1702_u0 ( .a(n_404), .o(n_423) );
na03f80 g40_u0 ( .a(n_559), .b(n_734), .c(n_927), .o(n_963) );
na02f80 g1902_u0 ( .a(i_rx_phy_bit_cnt_2_), .b(n_763), .o(n_359) );
in01f80 newInst_301 ( .a(newNet_300), .o(newNet_301) );
in01f80 newInst_55 ( .a(newNet_54), .o(newNet_55) );
oa12f80 g1878_u0 ( .a(n_351), .b(n_290), .c(n_583), .o(n_387) );
in01f80 newInst_213 ( .a(newNet_212), .o(newNet_213) );
in01f80 newInst_6 ( .a(newNet_2), .o(newNet_6) );
na02f80 g34_u0 ( .a(n_873), .b(n_139), .o(n_960) );
in01f80 newInst_170 ( .a(newNet_169), .o(newNet_170) );
ms00f80 i_tx_phy_data_done_reg_u0 ( .ck(newNet_123), .d(n_166), .o(i_tx_phy_data_done) );
oa12f80 g1748_u0 ( .a(n_447), .b(n_9), .c(n_885), .o(n_471) );
no02f80 g14_u0 ( .a(n_788), .b(n_981), .o(n_604) );
in01f80 newInst_162 ( .a(newNet_161), .o(newNet_162) );
in01f80 g1737_u1 ( .a(g1737_p), .o(n_489) );
ms00f80 i_rx_phy_rx_active_reg_u0 ( .ck(newNet_238), .d(n_709), .o(RxActive_o) );
ms00f80 i_tx_phy_txoe_r2_reg_u0 ( .ck(newNet_27), .d(n_291), .o(i_tx_phy_txoe_r2) );
in01f80 newInst_267 ( .a(newNet_266), .o(newNet_267) );
in01f80 g2113_u1 ( .a(g2113_p), .o(n_389) );
in01f80 newInst_96 ( .a(newNet_73), .o(newNet_96) );
ao12f80 g1843_u0 ( .a(n_400), .b(n_332), .c(n_301), .o(n_395) );
no03m80 g2644_u0 ( .a(n_929), .b(n_952), .c(n_735), .o(n_583) );
no03m80 g2014_u0 ( .a(i_tx_phy_txoe_r2), .b(i_tx_phy_txoe_r1), .c(n_864), .o(n_213) );
na02f80 g1903_u0 ( .a(n_289), .b(n_165), .o(n_304) );
ms00f80 i_rx_phy_rxd_s_reg_u0 ( .ck(newNet_211), .d(n_229), .o(i_rx_phy_rxd_s) );
ao12f80 g1884_u1 ( .a(g1884_p), .b(i_tx_phy_one_cnt_2_), .c(n_51), .o(n_138) );
no02f80 g1956_u0 ( .a(n_929), .b(n_965), .o(n_323) );
ms00f80 i_tx_phy_one_cnt_reg_2__u0 ( .ck(newNet_67), .d(n_388), .o(i_tx_phy_one_cnt_2_) );
na02f80 g1781_u3 ( .a(g1781_da), .b(g1781_db), .o(n_453) );
in01f80 newInst_132 ( .a(newNet_131), .o(newNet_132) );
in01f80 g1743_u1 ( .a(g1743_p), .o(n_482) );
no02f80 g2123_u0 ( .a(n_57), .b(n_56), .o(n_125) );
in01f80 newInst_145 ( .a(newNet_144), .o(newNet_145) );
in01f80 newInst_93 ( .a(newNet_92), .o(newNet_93) );
in01f80 newInst_289 ( .a(newNet_288), .o(newNet_289) );
in01f80 g1731_u0 ( .a(n_754), .o(n_490) );
in01f80 newInst_84 ( .a(newNet_83), .o(newNet_84) );
in01f80 g2568_u0 ( .a(n_841), .o(n_840) );
ms00f80 i_tx_phy_txdn_reg_u0 ( .ck(newNet_39), .d(n_364), .o(txdn) );
na02f80 g2118_u0 ( .a(TxValid_i), .b(rst), .o(n_164) );
na02f80 g1776_u1 ( .a(DataOut_i_0_), .b(g1776_sb), .o(g1776_da) );
ms00f80 i_rx_phy_rx_valid_reg_u0 ( .ck(newNet_224), .d(n_373), .o(RxValid_o) );
no02f80 g2100_u0 ( .a(n_878), .b(RxActive_o), .o(n_61) );
in01f80 newInst_128 ( .a(newNet_127), .o(newNet_128) );
in01f80 i_tx_phy_ld_data_reg_u1 ( .a(i_tx_phy_ld_data_reg_Q), .o(i_tx_phy_ld_data) );
in01f80 newInst_25 ( .a(newNet_24), .o(newNet_25) );
ao12f80 g1729_u0 ( .a(n_961), .b(n_359), .c(n_347), .o(n_414) );
ao22s80 g2060_u0 ( .a(i_tx_phy_append_eop), .b(g2674_p), .c(i_tx_phy_append_eop_sync1), .d(n_984), .o(n_237) );
na02f80 g1779_u1 ( .a(DataOut_i_3_), .b(g1779_sb), .o(g1779_da) );
ao12f80 g1877_u0 ( .a(n_228), .b(n_254), .c(i_tx_phy_bit_cnt_2_), .o(n_337) );
in01f80 g2108_u1 ( .a(g2108_p), .o(n_155) );
in01f80 g2106_u0 ( .a(n_598), .o(n_661) );
in01f80 newInst_208 ( .a(newNet_207), .o(newNet_208) );
in01f80 newInst_52 ( .a(newNet_38), .o(newNet_52) );
in01f80 g2116_u1 ( .a(g2116_p), .o(n_192) );
na02f80 g1757_u0 ( .a(n_969), .b(rst), .o(g1757_p) );
in01f80 g1781_u0 ( .a(i_tx_phy_ld_data), .o(g1781_sb) );
in01f80 g1782_u0 ( .a(i_tx_phy_ld_data), .o(g1782_sb) );
in01f80 newInst_105 ( .a(newNet_3), .o(newNet_105) );
in01f80 newInst_0 ( .a(tau_clk), .o(newNet_0) );
ms00f80 i_tx_phy_state_reg_0__u0 ( .ck(newNet_51), .d(n_459), .o(n_929) );
no02f80 g1921_u0 ( .a(n_255), .b(i_tx_phy_bit_cnt_2_), .o(n_300) );
in01f80 g2460_u0 ( .a(n_703), .o(n_704) );
na02f80 g1807_u0 ( .a(n_142), .b(n_764), .o(n_347) );
in01f80 newInst_70 ( .a(newNet_69), .o(newNet_70) );
na03f80 g1894_u0 ( .a(g2674_p), .b(n_170), .c(rst), .o(n_273) );
na03f80 g57_u0 ( .a(n_666), .b(i_rx_phy_rxdn_s), .c(i_rx_phy_rx_en), .o(n_916) );
na03f80 g2636_u0 ( .a(n_112), .b(n_940), .c(n_942), .o(n_943) );
ms00f80 i_rx_phy_rxdn_s_r_reg_u0 ( .ck(newNet_200), .d(n_222), .o(i_rx_phy_rxdn_s_r_reg_Q) );
in01f80 g2226_u0 ( .a(n_91), .o(n_74) );
ao12f80 g1661_u0 ( .a(FE_RN_2_0), .b(n_506), .c(n_660), .o(n_523) );
ao12f80 g1758_u0 ( .a(n_318), .b(n_538), .c(n_539), .o(n_432) );
ms00f80 i_rx_phy_hold_reg_reg_5__u0 ( .ck(newNet_257), .d(DataIn_o_6_), .o(DataIn_o_5_) );
in01f80 newInst_247 ( .a(newNet_246), .o(newNet_247) );
in01f80 g1905_u0 ( .a(n_416), .o(n_269) );
no02f80 g2128_u0 ( .a(n_27), .b(n_318), .o(g2128_p) );
in01f80 g2178_u0 ( .a(n_56), .o(n_77) );
no02f80 g2136_u0 ( .a(n_21), .b(n_22), .o(n_66) );
na02f80 g31_u0 ( .a(n_957), .b(n_958), .o(n_959) );
ms00f80 i_rx_phy_bit_cnt_reg_0__u0 ( .ck(newNet_313), .d(n_407), .o(i_rx_phy_bit_cnt_0_) );
in01f80 newInst_87 ( .a(newNet_33), .o(newNet_87) );
na02f80 g1703_u0 ( .a(n_380), .b(n_269), .o(n_404) );
na04m80 g2628_u0 ( .a(n_735), .b(n_984), .c(n_952), .d(n_929), .o(n_930) );
in01f80 newInst_76 ( .a(newNet_75), .o(newNet_76) );
ao22s80 g2065_u0 ( .a(n_238), .b(g2674_p), .c(i_tx_phy_txoe_r1), .d(n_984), .o(n_233) );
in01f80 newInst_14 ( .a(newNet_0), .o(newNet_14) );
ms00f80 i_tx_phy_hold_reg_d_reg_6__u0 ( .ck(newNet_105), .d(i_tx_phy_hold_reg_9), .o(i_tx_phy_hold_reg_d_reg_6__Q) );
in01f80 g11_u1 ( .a(g11_p), .o(n_911) );
in01f80 newInst_222 ( .a(newNet_221), .o(newNet_222) );
in01f80 newInst_265 ( .a(newNet_4), .o(newNet_265) );
in01f80 newInst_11 ( .a(newNet_0), .o(newNet_11) );
in01f80 newInst_193 ( .a(newNet_192), .o(newNet_193) );
in01f80 newInst_175 ( .a(newNet_174), .o(newNet_175) );
in01f80 newInst_45 ( .a(newNet_44), .o(newNet_45) );
in01f80 newInst_238 ( .a(newNet_237), .o(newNet_238) );
in01f80 newInst_311 ( .a(newNet_310), .o(newNet_311) );
na02f80 g1696_u0 ( .a(n_938), .b(n_480), .o(n_481) );
in01f80 newInst_215 ( .a(newNet_214), .o(newNet_215) );
na02f80 g1717_u0 ( .a(n_916), .b(n_74), .o(n_439) );
in01f80 newInst_180 ( .a(newNet_179), .o(newNet_180) );
in01f80 newInst_178 ( .a(newNet_177), .o(newNet_178) );
no02f80 g2135_u0 ( .a(n_37), .b(n_18), .o(n_141) );
na02f80 g1867_u0 ( .a(n_121), .b(n_958), .o(n_375) );
in01f80 g2162_u0 ( .a(rst_cnt_4_), .o(n_11) );
in01f80 newInst_164 ( .a(newNet_107), .o(newNet_164) );
no02f80 g1857_u0 ( .a(n_155), .b(RxValid_o), .o(g1857_p) );
in01f80 g2595_u0 ( .a(n_885), .o(n_878) );
in01f80 newInst_206 ( .a(newNet_205), .o(newNet_206) );
in01f80 newInst_172 ( .a(newNet_48), .o(newNet_172) );
ms00f80 i_tx_phy_hold_reg_d_reg_2__u0 ( .ck(newNet_118), .d(i_tx_phy_hold_reg_5), .o(i_tx_phy_hold_reg_d_12) );
no02f80 g1899_u0 ( .a(n_258), .b(n_984), .o(n_340) );
ao12f80 g39_u0 ( .a(n_977), .b(n_840), .c(n_567), .o(n_699) );
na02f80 g1915_u0 ( .a(n_343), .b(n_15), .o(n_344) );
na02f80 g1764_u0 ( .a(n_767), .b(n_410), .o(n_431) );
in01f80 g2172_u0 ( .a(n_22), .o(n_105) );
in01f80 newInst_67 ( .a(newNet_66), .o(newNet_67) );
in01f80 newInst_262 ( .a(newNet_261), .o(newNet_262) );
in01f80 newInst_290 ( .a(newNet_289), .o(newNet_290) );
ms00f80 usb_rst_reg_u0 ( .ck(newNet_70), .d(n_275), .o(usb_rst) );
na04m80 g1858_u0 ( .a(n_195), .b(n_238), .c(rst), .d(i_tx_phy_txoe_r1), .o(n_276) );
in01f80 newInst_34 ( .a(newNet_33), .o(newNet_34) );
in01f80 newInst_77 ( .a(newNet_76), .o(newNet_77) );
in01f80 g2275_u0 ( .a(i_rx_phy_rxd_s), .o(n_243) );
ms00f80 i_tx_phy_state_reg_1__u0 ( .ck(newNet_47), .d(n_420), .o(i_tx_phy_state_1_) );
in01f80 g1860_u0 ( .a(n_197), .o(n_198) );
na02f80 g1919_u0 ( .a(i_rx_phy_bit_cnt_0_), .b(n_763), .o(n_355) );
in01f80 g2593_u0 ( .a(n_885), .o(n_873) );
in01f80 newInst_285 ( .a(newNet_230), .o(newNet_285) );
ao12f80 g2052_u0 ( .a(i_tx_phy_append_eop_sync2), .b(n_7), .c(n_48), .o(n_123) );
in01f80 newInst_302 ( .a(newNet_140), .o(newNet_302) );
in01f80 newInst_276 ( .a(newNet_275), .o(newNet_276) );
in01f80 newInst_98 ( .a(newNet_97), .o(newNet_98) );
in01f80 g2584_u0 ( .a(n_885), .o(n_864) );
in01f80 newInst_27 ( .a(newNet_26), .o(newNet_27) );
in01f80 newInst_212 ( .a(newNet_147), .o(newNet_212) );
in01f80 g1991_u0 ( .a(n_66), .o(n_132) );
in01f80 newInst_113 ( .a(newNet_112), .o(newNet_113) );
no02f80 g1822_u0 ( .a(n_424), .b(n_665), .o(n_425) );
in01f80 newInst_56 ( .a(newNet_15), .o(newNet_56) );
ms00f80 i_tx_phy_hold_reg_reg_7__u0 ( .ck(newNet_74), .d(n_507), .o(i_tx_phy_hold_reg_10) );
na02f80 g1781_u1 ( .a(DataOut_i_5_), .b(g1781_sb), .o(g1781_da) );
in01f80 newInst_136 ( .a(newNet_135), .o(newNet_136) );
in01f80 newInst_39 ( .a(newNet_38), .o(newNet_39) );
na04m80 g1824_u0 ( .a(n_764), .b(i_rx_phy_bit_cnt_2_), .c(rst), .d(n_141), .o(n_410) );
na02f80 g2029_u0 ( .a(n_244), .b(n_243), .o(n_245) );
na02f80 g2662_u0 ( .a(n_735), .b(n_951), .o(n_971) );
in01f80 i_rx_phy_rxdp_s_r_reg_u1 ( .a(i_rx_phy_rxdp_s_r_reg_Q), .o(i_rx_phy_rxdp_s_r) );
no02f80 g1869_u0 ( .a(n_313), .b(n_416), .o(n_362) );
in01f80 newInst_158 ( .a(newNet_157), .o(newNet_158) );
in01f80 newInst_184 ( .a(newNet_183), .o(newNet_184) );
in01f80 newInst_90 ( .a(newNet_89), .o(newNet_90) );
in01f80 newInst_205 ( .a(newNet_204), .o(newNet_205) );
in01f80 g2224_u0 ( .a(n_28), .o(n_139) );
no02f80 g2141_u0 ( .a(n_8), .b(n_984), .o(g2141_p) );
in01f80 newInst_5 ( .a(newNet_4), .o(newNet_5) );
na02f80 g2466_u0 ( .a(n_461), .b(n_511), .o(n_710) );
na03f80 g2497_u0 ( .a(n_112), .b(n_788), .c(n_942), .o(n_748) );
in01f80 newInst_8 ( .a(newNet_7), .o(newNet_8) );
in01f80 g2160_u0 ( .a(i_rx_phy_one_cnt_1_), .o(n_52) );
na02f80 g1987_u0 ( .a(n_246), .b(n_245), .o(n_312) );
na02f80 g2036_u0 ( .a(n_125), .b(n_124), .o(n_231) );
na04m80 g1747_u0 ( .a(n_248), .b(n_266), .c(n_426), .d(i_rx_phy_sd_nrzi), .o(n_479) );
na02f80 g1780_u1 ( .a(DataOut_i_4_), .b(g1780_sb), .o(g1780_da) );
na02f80 g1820_u0 ( .a(n_424), .b(n_666), .o(n_426) );
na02f80 g20_u0 ( .a(n_852), .b(i_rx_phy_shift_en), .o(n_991) );
in01f80 newInst_151 ( .a(newNet_113), .o(newNet_151) );
no02f80 g1966_u0 ( .a(n_237), .b(n_318), .o(n_317) );
ao12f80 g1763_u0 ( .a(n_400), .b(n_163), .c(n_342), .o(n_388) );
in01f80 newInst_229 ( .a(newNet_68), .o(newNet_229) );
in01f80 g1901_u1 ( .a(g1901_p), .o(n_373) );
in01f80 newInst_163 ( .a(newNet_162), .o(newNet_163) );
in01f80 newInst_192 ( .a(newNet_118), .o(newNet_192) );
in01f80 g1855_u0 ( .a(n_274), .o(g1855_sb) );
in01f80 g2251_u0 ( .a(i_tx_phy_data_done), .o(n_10) );
in01f80 g2646_u0 ( .a(i_tx_phy_state_2_), .o(n_951) );
na02f80 g1842_u0 ( .a(n_308), .b(rst), .o(n_366) );
na02f80 g1779_u2 ( .a(i_tx_phy_hold_reg_6), .b(i_tx_phy_ld_data), .o(g1779_db) );
ms00f80 i_rx_phy_one_cnt_reg_0__u0 ( .ck(newNet_244), .d(n_406), .o(i_rx_phy_one_cnt_0_) );
in01f80 newInst_258 ( .a(newNet_163), .o(newNet_258) );
ms00f80 i_tx_phy_sd_raw_o_reg_u0 ( .ck(newNet_61), .d(n_411), .o(i_tx_phy_sd_raw_o) );
na03f80 g1875_u0 ( .a(n_390), .b(i_rx_phy_dpll_state_1_), .c(n_60), .o(n_435) );
in01f80 g2670_u0 ( .a(i_rx_phy_fs_state_2_), .o(n_910) );
in01f80 newInst_250 ( .a(newNet_249), .o(newNet_250) );
in01f80 newInst_75 ( .a(newNet_61), .o(newNet_75) );
ms00f80 i_rx_phy_rxdp_s0_reg_u0 ( .ck(newNet_191), .d(rxdp), .o(i_rx_phy_rxdp_s0) );
in01f80 g2063_u0 ( .a(n_852), .o(g2063_sb) );
in01f80 g1757_u1 ( .a(g1757_p), .o(n_420) );
in01f80 newInst_251 ( .a(newNet_250), .o(newNet_251) );
ao12f80 g1844_u0 ( .a(n_400), .b(n_344), .c(n_294), .o(n_394) );
in01f80 newInst_194 ( .a(newNet_193), .o(newNet_194) );
na04m80 g36_u0 ( .a(n_699), .b(n_700), .c(n_701), .d(n_968), .o(n_703) );
in01f80 newInst_310 ( .a(newNet_309), .o(newNet_310) );
in01f80 newInst_280 ( .a(newNet_279), .o(newNet_280) );
in01f80 newInst_286 ( .a(newNet_285), .o(newNet_286) );
in01f80 newInst_161 ( .a(newNet_160), .o(newNet_161) );
in01f80 newInst_115 ( .a(newNet_48), .o(newNet_115) );
in01f80 newInst_120 ( .a(newNet_119), .o(newNet_120) );
ms00f80 rst_cnt_reg_1__u0 ( .ck(newNet_13), .d(n_367), .o(rst_cnt_1_) );
oa12f80 g1984_u0 ( .a(n_172), .b(i_tx_phy_hold_reg_d_15), .c(n_168), .o(n_254) );
na02f80 g2063_u1 ( .a(n_130), .b(g2063_sb), .o(g2063_da) );
in01f80 g2537_u0 ( .a(n_965), .o(n_800) );
na03f80 g1711_u0 ( .a(n_782), .b(n_176), .c(n_783), .o(n_493) );
na03f80 g1728_u0 ( .a(n_974), .b(n_462), .c(n_450), .o(n_507) );
in01f80 g2186_u0 ( .a(i_tx_phy_bit_cnt_1_), .o(n_57) );
in01f80 g2254_u0 ( .a(rst_cnt_0_), .o(n_21) );
ms00f80 rst_cnt_reg_2__u0 ( .ck(newNet_10), .d(n_428), .o(n_306) );
ms00f80 i_tx_phy_txoe_r1_reg_u0 ( .ck(newNet_31), .d(n_320), .o(i_tx_phy_txoe_r1) );
ms00f80 i_rx_phy_rxd_r_reg_u0 ( .ck(newNet_222), .d(n_130), .o(i_rx_phy_rxd_r) );
ao12f80 g2067_u1 ( .a(g2067_p), .b(n_120), .c(i_rx_phy_one_cnt_0_), .o(n_121) );
ao12f80 g2651_u1 ( .a(g2651_p), .b(n_139), .c(n_54), .o(n_957) );
in01f80 newInst_223 ( .a(newNet_88), .o(newNet_223) );
in01f80 newInst_61 ( .a(newNet_2), .o(newNet_61) );
na04m80 g2654_u0 ( .a(n_963), .b(n_966), .c(n_967), .d(n_968), .o(n_969) );
na02f80 g1904_u0 ( .a(n_283), .b(rst), .o(n_333) );
in01f80 newInst_95 ( .a(newNet_94), .o(newNet_95) );
in01f80 g2225_u0 ( .a(i_rx_phy_one_cnt_2_), .o(n_28) );
in01f80 newInst_244 ( .a(newNet_243), .o(newNet_244) );
in01f80 g2194_u0 ( .a(i_tx_phy_bit_cnt_2_), .o(n_124) );
in01f80 newInst_127 ( .a(newNet_126), .o(newNet_127) );
in01f80 g2158_u0 ( .a(phy_tx_mode), .o(n_8) );
in01f80 g2506_u1 ( .a(g2506_p), .o(n_756) );
in01f80 newInst_41 ( .a(newNet_40), .o(newNet_41) );
ao22s80 g2064_u0 ( .a(i_tx_phy_txoe_r2), .b(n_852), .c(i_tx_phy_txoe_r1), .d(g2674_p), .o(n_201) );
in01f80 newInst_38 ( .a(newNet_37), .o(newNet_38) );
ms00f80 i_rx_phy_hold_reg_reg_4__u0 ( .ck(newNet_262), .d(DataIn_o_5_), .o(DataIn_o_4_) );
ms00f80 i_tx_phy_bit_cnt_reg_0__u0 ( .ck(newNet_133), .d(n_395), .o(i_tx_phy_bit_cnt_0_) );
na02f80 g2494_u0 ( .a(n_741), .b(n_742), .o(g2494_p) );
in01f80 newInst_264 ( .a(newNet_263), .o(newNet_264) );
in01f80 newInst_239 ( .a(newNet_204), .o(newNet_239) );
na02f80 g1759_u0 ( .a(n_446), .b(g2674_p), .o(n_447) );
na02f80 g1809_u0 ( .a(n_198), .b(rst_cnt_3_), .o(n_292) );
in01f80 newInst_275 ( .a(newNet_266), .o(newNet_275) );
ao12f80 g1841_u0 ( .a(n_961), .b(n_355), .c(n_331), .o(n_407) );
in01f80 i_rx_phy_se0_r_reg_u1 ( .a(i_rx_phy_se0_r_reg_Q), .o(i_rx_phy_se0_r) );
ms00f80 i_rx_phy_sd_r_reg_u0 ( .ck(newNet_173), .d(n_203), .o(i_rx_phy_sd_r) );
na02f80 g1849_u0 ( .a(n_138), .b(n_340), .o(n_342) );
ms00f80 i_tx_phy_hold_reg_d_reg_1__u0 ( .ck(newNet_120), .d(i_tx_phy_hold_reg_4), .o(i_tx_phy_hold_reg_d_reg_1__Q) );
ao12f80 g2650_u0 ( .a(n_961), .b(n_959), .c(n_960), .o(n_962) );
ms00f80 i_rx_phy_fs_state_reg_1__u0 ( .ck(newNet_280), .d(n_523), .o(n_796) );
na02f80 g1917_u0 ( .a(n_930), .b(n_841), .o(n_330) );
no02f80 g1881_u0 ( .a(i_rx_phy_bit_cnt_2_), .b(n_141), .o(g1881_p) );
in01f80 g2051_u0 ( .a(n_123), .o(n_170) );
ms00f80 i_rx_phy_rxdp_s1_reg_u0 ( .ck(newNet_187), .d(i_rx_phy_rxdp_s0), .o(LineState_o_0_) );
in01f80 g2129_u0 ( .a(n_150), .o(n_266) );
in01f80 newInst_309 ( .a(newNet_308), .o(newNet_309) );
no02f80 g1874_u0 ( .a(n_390), .b(n_389), .o(n_391) );
no02f80 g2620_u0 ( .a(n_923), .b(n_924), .o(n_925) );
in01f80 newInst_31 ( .a(newNet_30), .o(newNet_31) );
na02f80 g1737_u0 ( .a(n_458), .b(n_974), .o(g1737_p) );
ms00f80 i_rx_phy_fs_ce_r1_reg_u0 ( .ck(newNet_290), .d(n_81), .o(i_rx_phy_fs_ce_r1) );
in01f80 newInst_228 ( .a(newNet_227), .o(newNet_228) );
ms00f80 i_tx_phy_state_reg_2__u0 ( .ck(newNet_46), .d(n_432), .o(i_tx_phy_state_2_) );
in01f80 g2494_u1 ( .a(g2494_p), .o(n_743) );
in01f80 newInst_293 ( .a(newNet_292), .o(newNet_293) );
no02f80 g1908_u0 ( .a(n_132), .b(n_306), .o(n_230) );
ao12f80 g1848_u0 ( .a(n_400), .b(n_161), .c(n_299), .o(n_378) );
in01f80 newInst_166 ( .a(newNet_165), .o(newNet_166) );
in01f80 newInst_47 ( .a(newNet_21), .o(newNet_47) );
in01f80 newInst_147 ( .a(newNet_146), .o(newNet_147) );
ao12f80 g1812_u0 ( .a(n_961), .b(n_152), .c(n_375), .o(n_427) );
no02f80 g44_u0 ( .a(n_971), .b(n_894), .o(n_965) );
ao12f80 g2621_u0 ( .a(n_922), .b(n_915), .c(n_916), .o(n_923) );
in01f80 newInst_199 ( .a(newNet_198), .o(newNet_199) );
in01f80 newInst_44 ( .a(newNet_43), .o(newNet_44) );
ao12f80 g2055_u0 ( .a(n_164), .b(n_10), .c(i_tx_phy_tx_ip), .o(n_166) );
in01f80 g2674_u0 ( .a(n_984), .o(g2674_p) );
ms00f80 i_rx_phy_bit_stuff_err_reg_u0 ( .ck(newNet_302), .d(n_505), .o(i_rx_phy_bit_stuff_err_reg_Q) );
in01f80 newInst_191 ( .a(newNet_190), .o(newNet_191) );
in01f80 newInst_299 ( .a(newNet_298), .o(newNet_299) );
in01f80 newInst_253 ( .a(newNet_252), .o(newNet_253) );
in01f80 newInst_66 ( .a(newNet_65), .o(newNet_66) );
na02f80 g1953_u0 ( .a(n_759), .b(i_rx_phy_sd_nrzi), .o(n_324) );
no02f80 g2067_u0 ( .a(n_120), .b(i_rx_phy_one_cnt_0_), .o(g2067_p) );
in01f80 g15_u1 ( .a(g15_p), .o(n_949) );
na02f80 g1777_u1 ( .a(DataOut_i_1_), .b(g1777_sb), .o(g1777_da) );
in01f80 newInst_152 ( .a(newNet_151), .o(newNet_152) );
in01f80 newInst_78 ( .a(newNet_77), .o(newNet_78) );
na02f80 g2415_u0 ( .a(n_753), .b(n_74), .o(n_631) );
in01f80 g1778_u0 ( .a(i_tx_phy_ld_data), .o(g1778_sb) );
in01f80 newInst_9 ( .a(newNet_8), .o(newNet_9) );
na02f80 g1740_u0 ( .a(n_455), .b(n_974), .o(g1740_p) );
na02f80 g1855_u3 ( .a(g1855_da), .b(g1855_db), .o(n_311) );
in01f80 g2038_u0 ( .a(n_604), .o(n_209) );
in01f80 newInst_185 ( .a(newNet_87), .o(newNet_185) );
na02f80 g1777_u3 ( .a(g1777_da), .b(g1777_db), .o(n_457) );
in01f80 newInst_230 ( .a(newNet_229), .o(newNet_230) );
na02f80 g1901_u0 ( .a(n_764), .b(i_rx_phy_rx_valid1), .o(g1901_p) );
ao12f80 g1736_u0 ( .a(n_27), .b(n_369), .c(n_337), .o(n_411) );
na02f80 g1738_u0 ( .a(n_457), .b(n_974), .o(g1738_p) );
in01f80 g2164_u0 ( .a(n_238), .o(n_27) );
in01f80 newInst_220 ( .a(newNet_219), .o(newNet_220) );
ms00f80 i_rx_phy_shift_en_reg_u0 ( .ck(newNet_163), .d(n_992), .o(i_rx_phy_shift_en) );
ms00f80 i_tx_phy_txoe_reg_u0 ( .ck(newNet_22), .d(n_333), .o(txoe) );
na02f80 g1779_u3 ( .a(g1779_da), .b(g1779_db), .o(n_455) );

endmodule
