module s386 (
v4,
v3,
v5,
v1,
v0,
blif_clk_net,
v2,
v6,
blif_reset_net,
v13_D_11,
v13_D_6,
v13_D_10,
v13_D_12,
v13_D_7,
v13_D_8,
v13_D_9);

// Start PIs
input v4;
input v3;
input v5;
input v1;
input v0;
input blif_clk_net;
input v2;
input v6;
input blif_reset_net;

// Start POs
output v13_D_11;
output v13_D_6;
output v13_D_10;
output v13_D_12;
output v13_D_7;
output v13_D_8;
output v13_D_9;

// Start wires
wire net_166;
wire net_107;
wire net_47;
wire net_159;
wire v13_D_7;
wire net_61;
wire net_137;
wire net_132;
wire net_54;
wire net_105;
wire net_62;
wire net_6;
wire net_129;
wire net_119;
wire net_98;
wire net_23;
wire net_117;
wire net_12;
wire net_151;
wire net_74;
wire v13_D_12;
wire net_53;
wire net_93;
wire net_168;
wire net_135;
wire net_130;
wire net_147;
wire net_127;
wire net_14;
wire net_113;
wire net_26;
wire net_76;
wire blif_clk_net;
wire net_101;
wire net_32;
wire net_111;
wire net_90;
wire net_40;
wire net_100;
wire net_85;
wire net_69;
wire net_124;
wire net_161;
wire net_141;
wire net_160;
wire v1;
wire net_83;
wire net_115;
wire v2;
wire net_4;
wire net_95;
wire net_17;
wire net_78;
wire net_27;
wire net_164;
wire net_56;
wire net_87;
wire v13_D_11;
wire net_0;
wire net_155;
wire net_35;
wire v6;
wire net_16;
wire net_22;
wire net_39;
wire net_157;
wire net_144;
wire net_102;
wire v3;
wire net_2;
wire net_59;
wire net_9;
wire net_42;
wire net_120;
wire net_109;
wire net_80;
wire net_65;
wire blif_reset_net;
wire net_50;
wire net_162;
wire net_96;
wire net_66;
wire net_38;
wire net_44;
wire net_167;
wire net_136;
wire net_134;
wire net_19;
wire net_89;
wire net_45;
wire net_126;
wire net_34;
wire net_108;
wire v13_D_6;
wire net_150;
wire net_63;
wire net_152;
wire net_116;
wire net_30;
wire net_91;
wire net_24;
wire net_55;
wire net_99;
wire net_106;
wire net_46;
wire net_140;
wire net_118;
wire net_148;
wire net_104;
wire net_146;
wire v13_D_8;
wire net_72;
wire net_122;
wire net_25;
wire v0;
wire net_7;
wire net_70;
wire net_5;
wire net_52;
wire net_165;
wire net_128;
wire v5;
wire net_138;
wire net_13;
wire net_94;
wire net_11;
wire net_18;
wire net_123;
wire net_131;
wire net_114;
wire net_29;
wire net_68;
wire net_149;
wire net_142;
wire v13_D_10;
wire net_77;
wire net_20;
wire net_31;
wire net_36;
wire net_49;
wire net_158;
wire v4;
wire net_15;
wire net_41;
wire net_57;
wire net_71;
wire net_153;
wire net_156;
wire net_3;
wire net_84;
wire net_154;
wire net_1;
wire net_92;
wire net_112;
wire net_103;
wire net_139;
wire net_43;
wire net_10;
wire net_28;
wire net_169;
wire net_21;
wire net_51;
wire net_79;
wire net_143;
wire net_97;
wire net_88;
wire net_145;
wire net_60;
wire net_81;
wire net_163;
wire net_58;
wire v13_D_9;
wire net_67;
wire net_82;
wire net_64;
wire net_37;
wire net_110;
wire net_121;
wire net_73;
wire net_33;
wire net_48;
wire net_8;
wire net_75;
wire net_86;
wire net_133;
wire net_125;

// Start cells
DFFR_X2 inst_145 ( .QN(net_146), .RN(net_97), .D(net_90), .CK(net_165) );
INV_X4 inst_103 ( .ZN(net_43), .A(v1) );
INV_X4 inst_125 ( .ZN(net_24), .A(net_19) );
INV_X2 inst_138 ( .A(net_133), .ZN(net_132) );
CLKBUF_X2 inst_159 ( .A(net_151), .Z(net_152) );
NOR2_X2 inst_15 ( .A2(net_139), .ZN(net_13), .A1(net_12) );
INV_X4 inst_134 ( .ZN(net_94), .A(net_87) );
NAND4_X2 inst_24 ( .A3(net_74), .ZN(net_64), .A2(net_63), .A4(net_62), .A1(net_2) );
INV_X4 inst_114 ( .A(net_143), .ZN(net_14) );
NOR4_X2 inst_6 ( .A3(net_75), .A4(net_73), .A2(net_40), .A1(net_17), .ZN(v13_D_9) );
INV_X4 inst_131 ( .A(net_46), .ZN(net_32) );
NAND2_X2 inst_76 ( .A2(net_142), .ZN(net_122), .A1(net_51) );
CLKBUF_X2 inst_160 ( .A(net_152), .Z(net_153) );
AND4_X2 inst_150 ( .A3(net_146), .A4(net_129), .ZN(net_44), .A2(net_43), .A1(v4) );
NAND3_X2 inst_33 ( .ZN(net_102), .A2(net_74), .A1(net_68), .A3(net_65) );
CLKBUF_X2 inst_172 ( .A(net_164), .Z(net_165) );
NAND2_X2 inst_83 ( .A1(net_111), .ZN(net_78), .A2(net_31) );
NAND2_X4 inst_47 ( .ZN(net_85), .A2(net_31), .A1(net_24) );
NOR2_X2 inst_19 ( .ZN(net_49), .A1(net_23), .A2(net_14) );
INV_X4 inst_123 ( .ZN(net_25), .A(net_18) );
INV_X4 inst_121 ( .ZN(net_15), .A(net_14) );
OR2_X2 inst_2 ( .A2(net_147), .A1(net_143), .ZN(net_9) );
NOR3_X2 inst_8 ( .ZN(net_119), .A3(net_116), .A2(net_114), .A1(net_49) );
INV_X4 inst_118 ( .ZN(net_77), .A(net_75) );
NAND2_X2 inst_86 ( .ZN(net_110), .A2(net_72), .A1(net_52) );
AND2_X4 inst_153 ( .A2(net_148), .A1(net_147), .ZN(net_6) );
NOR2_X2 inst_20 ( .A1(net_132), .ZN(net_59), .A2(net_41) );
NAND3_X4 inst_27 ( .ZN(net_90), .A2(net_88), .A1(net_82), .A3(net_66) );
NAND3_X2 inst_38 ( .ZN(net_130), .A1(net_67), .A3(net_37), .A2(net_33) );
INV_X4 inst_100 ( .A(net_134), .ZN(net_133) );
NAND2_X4 inst_52 ( .A1(net_112), .ZN(net_106), .A2(net_68) );
NAND2_X2 inst_90 ( .A2(net_121), .A1(net_120), .ZN(net_112) );
INV_X2 inst_140 ( .ZN(net_0), .A(v2) );
NAND3_X2 inst_40 ( .ZN(net_81), .A3(net_48), .A2(net_39), .A1(net_30) );
CLKBUF_X2 inst_162 ( .A(net_154), .Z(net_155) );
CLKBUF_X2 inst_167 ( .A(blif_clk_net), .Z(net_160) );
NAND2_X2 inst_93 ( .A2(net_100), .A1(net_80), .ZN(v13_D_11) );
NAND2_X2 inst_81 ( .ZN(net_72), .A1(net_71), .A2(net_57) );
INV_X4 inst_95 ( .A(net_144), .ZN(net_138) );
OR2_X4 inst_1 ( .ZN(net_28), .A1(net_27), .A2(net_26) );
NAND2_X2 inst_72 ( .ZN(net_55), .A1(net_54), .A2(net_53) );
INV_X2 inst_139 ( .A(net_117), .ZN(net_116) );
AND2_X2 inst_155 ( .ZN(net_124), .A2(net_31), .A1(v1) );
NAND2_X2 inst_59 ( .ZN(net_141), .A1(net_19), .A2(net_7) );
INV_X4 inst_135 ( .ZN(net_95), .A(net_93) );
NAND3_X2 inst_44 ( .A1(net_103), .ZN(net_96), .A3(net_92), .A2(net_91) );
NAND2_X2 inst_55 ( .ZN(net_140), .A1(net_131), .A2(v2) );
CLKBUF_X2 inst_174 ( .A(net_166), .Z(net_167) );
INV_X4 inst_115 ( .A(net_146), .ZN(net_16) );
NAND3_X2 inst_37 ( .A2(net_147), .A1(net_105), .ZN(net_67), .A3(v4) );
DFFR_X2 inst_148 ( .QN(net_147), .RN(net_97), .D(net_95), .CK(net_156) );
CLKBUF_X2 inst_164 ( .A(net_154), .Z(net_157) );
NOR4_X2 inst_5 ( .A2(net_77), .A1(net_76), .A3(net_63), .ZN(v13_D_12), .A4(v0) );
CLKBUF_X2 inst_157 ( .A(net_149), .Z(net_150) );
NAND2_X2 inst_84 ( .A1(net_122), .ZN(net_109), .A2(net_71) );
NAND2_X4 inst_51 ( .A1(net_126), .ZN(net_120), .A2(net_31) );
INV_X2 inst_142 ( .ZN(net_40), .A(net_39) );
NAND2_X2 inst_80 ( .ZN(net_88), .A1(net_74), .A2(net_56) );
CLKBUF_X2 inst_173 ( .A(net_155), .Z(net_166) );
INV_X4 inst_105 ( .A(net_148), .ZN(net_34) );
NAND2_X2 inst_68 ( .ZN(net_121), .A2(net_65), .A1(v1) );
NAND2_X2 inst_78 ( .A1(net_134), .ZN(net_70), .A2(net_42) );
NAND3_X2 inst_42 ( .A1(net_110), .A3(net_92), .A2(net_91), .ZN(net_87) );
CLKBUF_X2 inst_175 ( .A(net_167), .Z(net_168) );
NAND2_X2 inst_53 ( .A2(net_145), .ZN(net_3), .A1(v1) );
INV_X4 inst_133 ( .A(net_85), .ZN(net_56) );
NAND4_X2 inst_26 ( .A4(net_102), .A1(net_101), .ZN(net_89), .A3(net_88), .A2(net_64) );
AND4_X2 inst_151 ( .A1(net_75), .A4(net_62), .A3(net_47), .ZN(v13_D_10), .A2(v1) );
INV_X4 inst_112 ( .ZN(net_75), .A(net_5) );
NAND2_X2 inst_64 ( .A2(net_143), .A1(net_140), .ZN(net_105) );
INV_X4 inst_107 ( .ZN(net_12), .A(v3) );
NAND2_X2 inst_67 ( .ZN(net_45), .A2(net_25), .A1(net_16) );
INV_X4 inst_127 ( .ZN(net_65), .A(net_36) );
NAND2_X2 inst_70 ( .A2(net_129), .ZN(net_48), .A1(net_28) );
INV_X4 inst_129 ( .ZN(net_38), .A(net_24) );
NAND2_X2 inst_92 ( .ZN(net_100), .A2(net_99), .A1(net_77) );
NAND3_X2 inst_29 ( .A2(net_136), .ZN(net_21), .A3(net_6), .A1(net_1) );
NOR2_X2 inst_17 ( .A1(net_147), .ZN(net_54), .A2(net_31) );
NOR2_X4 inst_11 ( .A1(net_131), .ZN(net_129), .A2(v3) );
DFFR_X2 inst_146 ( .QN(net_145), .RN(net_97), .D(net_89), .CK(net_161) );
NOR2_X2 inst_14 ( .A2(net_143), .ZN(net_125), .A1(net_63) );
INV_X4 inst_122 ( .ZN(net_68), .A(net_16) );
NAND3_X2 inst_31 ( .ZN(net_37), .A1(net_13), .A3(net_10), .A2(net_9) );
NAND4_X2 inst_25 ( .A2(net_115), .ZN(net_107), .A1(net_65), .A4(net_31), .A3(v0) );
INV_X4 inst_126 ( .A(net_147), .ZN(net_22) );
CLKBUF_X2 inst_158 ( .A(net_150), .Z(net_151) );
INV_X2 inst_141 ( .A(net_71), .ZN(net_17) );
NAND2_X2 inst_62 ( .A2(net_125), .A1(net_114), .ZN(net_33) );
INV_X4 inst_110 ( .ZN(net_5), .A(net_2) );
NAND2_X2 inst_74 ( .ZN(net_57), .A1(net_35), .A2(net_21) );
NAND2_X2 inst_57 ( .ZN(net_11), .A2(net_3), .A1(v0) );
NAND3_X2 inst_35 ( .A3(net_65), .ZN(net_60), .A2(net_54), .A1(v5) );
INV_X4 inst_99 ( .A(net_135), .ZN(net_134) );
NAND2_X4 inst_48 ( .A1(net_118), .ZN(net_113), .A2(net_85) );
NAND2_X2 inst_69 ( .ZN(net_47), .A1(net_46), .A2(net_4) );
NAND2_X4 inst_46 ( .A2(net_143), .A1(net_139), .ZN(net_36) );
NAND2_X2 inst_82 ( .ZN(net_126), .A2(net_70), .A1(net_43) );
INV_X4 inst_136 ( .ZN(net_98), .A(net_96) );
NAND3_X2 inst_30 ( .A1(net_147), .A2(net_129), .ZN(net_117), .A3(net_26) );
INV_X4 inst_102 ( .ZN(net_63), .A(v5) );
INV_X4 inst_108 ( .A(net_145), .ZN(net_2) );
CLKBUF_X2 inst_165 ( .A(net_157), .Z(net_158) );
NAND3_X2 inst_32 ( .A1(net_147), .ZN(net_142), .A2(net_135), .A3(net_34) );
NOR2_X2 inst_22 ( .A2(net_116), .ZN(net_79), .A1(net_59) );
DFFR_X2 inst_144 ( .QN(net_143), .RN(net_97), .D(net_86), .CK(net_169) );
NAND3_X2 inst_34 ( .A1(net_133), .ZN(net_50), .A3(net_18), .A2(v2) );
NOR2_X4 inst_12 ( .A2(net_146), .ZN(net_115), .A1(net_22) );
NAND2_X2 inst_56 ( .A2(net_143), .ZN(net_10), .A1(v2) );
NAND2_X2 inst_71 ( .ZN(net_76), .A2(net_62), .A1(net_46) );
NOR2_X2 inst_21 ( .ZN(net_73), .A1(net_69), .A2(net_44) );
INV_X4 inst_104 ( .ZN(net_74), .A(v0) );
NAND2_X2 inst_60 ( .A1(net_31), .ZN(net_29), .A2(net_5) );
CLKBUF_X2 inst_169 ( .A(net_155), .Z(net_162) );
CLKBUF_X2 inst_168 ( .A(net_160), .Z(net_161) );
INV_X4 inst_97 ( .A(net_138), .ZN(net_137) );
CLKBUF_X2 inst_161 ( .A(net_153), .Z(net_154) );
INV_X4 inst_124 ( .A(net_68), .ZN(net_46) );
NOR2_X2 inst_18 ( .ZN(net_62), .A2(net_36), .A1(net_8) );
NOR2_X2 inst_16 ( .ZN(net_53), .A1(net_36), .A2(v5) );
NAND2_X2 inst_88 ( .A1(net_130), .ZN(net_108), .A2(net_31) );
OR2_X2 inst_3 ( .ZN(net_52), .A2(net_51), .A1(net_15) );
CLKBUF_X2 inst_156 ( .A(blif_clk_net), .Z(net_149) );
NOR3_X2 inst_9 ( .A1(net_119), .ZN(net_86), .A3(net_85), .A2(net_84) );
INV_X4 inst_113 ( .ZN(net_8), .A(net_6) );
CLKBUF_X2 inst_170 ( .A(net_162), .Z(net_163) );
NAND2_X4 inst_50 ( .A2(net_124), .A1(net_123), .ZN(net_82) );
INV_X2 inst_137 ( .A(net_137), .ZN(net_136) );
NAND3_X2 inst_41 ( .ZN(net_104), .A1(net_78), .A3(net_55), .A2(net_50) );
INV_X4 inst_130 ( .ZN(net_39), .A(net_25) );
NAND2_X2 inst_91 ( .A2(net_107), .A1(net_106), .ZN(net_99) );
INV_X4 inst_132 ( .ZN(net_92), .A(net_38) );
INV_X1 inst_143 ( .ZN(net_97), .A(blif_reset_net) );
CLKBUF_X2 inst_176 ( .A(net_168), .Z(net_169) );
AND3_X1 inst_152 ( .A1(net_92), .A2(net_91), .A3(net_83), .ZN(v13_D_6) );
NAND2_X2 inst_58 ( .A2(net_146), .A1(net_145), .ZN(net_19) );
NAND3_X2 inst_36 ( .ZN(net_66), .A2(net_65), .A1(net_45), .A3(net_11) );
DFFR_X2 inst_147 ( .QN(net_148), .RN(net_97), .D(net_94), .CK(net_151) );
NAND2_X2 inst_87 ( .ZN(net_83), .A2(net_81), .A1(net_60) );
NAND2_X2 inst_61 ( .A1(net_71), .ZN(net_30), .A2(net_0) );
NAND2_X4 inst_45 ( .ZN(net_7), .A1(net_6), .A2(v0) );
INV_X4 inst_96 ( .ZN(net_139), .A(net_138) );
INV_X4 inst_101 ( .A(net_138), .ZN(net_131) );
OR2_X4 inst_0 ( .A1(net_147), .A2(net_143), .ZN(net_41) );
NOR3_X2 inst_10 ( .A1(net_85), .A2(net_84), .A3(net_79), .ZN(v13_D_7) );
NOR4_X2 inst_4 ( .A1(net_76), .A2(net_75), .A3(net_74), .ZN(v13_D_8), .A4(v6) );
NAND2_X2 inst_65 ( .A2(net_114), .ZN(net_35), .A1(net_34) );
NAND2_X2 inst_89 ( .A2(net_109), .A1(net_108), .ZN(net_103) );
NAND3_X2 inst_28 ( .A3(net_147), .A1(net_26), .ZN(net_20), .A2(net_12) );
INV_X4 inst_111 ( .A(net_34), .ZN(net_31) );
NAND2_X2 inst_66 ( .ZN(net_42), .A1(net_41), .A2(net_20) );
INV_X4 inst_117 ( .ZN(net_27), .A(net_14) );
INV_X4 inst_98 ( .A(net_136), .ZN(net_135) );
NAND2_X2 inst_63 ( .A2(net_128), .A1(net_127), .ZN(net_51) );
NOR3_X2 inst_7 ( .A1(net_132), .A2(net_74), .ZN(net_69), .A3(net_68) );
NAND2_X4 inst_49 ( .A1(net_113), .ZN(net_101), .A2(v1) );
INV_X4 inst_120 ( .ZN(net_91), .A(net_84) );
AND2_X2 inst_154 ( .ZN(net_1), .A2(v2), .A1(v3) );
NOR2_X2 inst_13 ( .A1(net_147), .A2(net_138), .ZN(net_114) );
INV_X4 inst_119 ( .ZN(net_71), .A(net_14) );
NAND2_X2 inst_75 ( .ZN(net_58), .A1(net_36), .A2(net_29) );
CLKBUF_X2 inst_166 ( .A(net_158), .Z(net_159) );
INV_X4 inst_116 ( .ZN(net_18), .A(net_8) );
CLKBUF_X2 inst_163 ( .A(net_155), .Z(net_156) );
NAND2_X2 inst_85 ( .ZN(net_123), .A2(net_61), .A1(net_38) );
NAND2_X2 inst_54 ( .ZN(net_84), .A2(net_43), .A1(v0) );
NAND2_X2 inst_79 ( .A1(net_117), .ZN(net_111), .A2(net_27) );
INV_X4 inst_109 ( .ZN(net_128), .A(net_34) );
INV_X4 inst_106 ( .ZN(net_26), .A(v4) );
DFFR_X2 inst_149 ( .QN(net_144), .D(net_98), .RN(net_97), .CK(net_159) );
NAND3_X2 inst_43 ( .A1(net_104), .ZN(net_93), .A3(net_92), .A2(net_91) );
NAND3_X2 inst_39 ( .ZN(net_80), .A2(net_74), .A3(net_58), .A1(net_32) );
INV_X4 inst_128 ( .ZN(net_23), .A(net_22) );
NAND2_X2 inst_73 ( .A1(net_141), .ZN(net_118), .A2(net_65) );
NOR2_X1 inst_23 ( .A2(net_147), .A1(net_137), .ZN(net_127) );
CLKBUF_X2 inst_171 ( .A(net_163), .Z(net_164) );
NAND2_X2 inst_77 ( .A1(net_115), .ZN(net_61), .A2(net_53) );
NAND2_X1 inst_94 ( .ZN(net_4), .A2(v0), .A1(v5) );

endmodule
