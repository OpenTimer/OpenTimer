module s1196 (
G1,
G11,
G8,
G5,
G9,
G3,
G13,
G4,
G12,
G2,
blif_clk_net,
G7,
blif_reset_net,
G10,
G0,
G6,
G549,
G542,
G530,
G552,
G45,
G547,
G548,
G537,
G551,
G532,
G539,
G546,
G535,
G550);

// Start PIs
input G1;
input G11;
input G8;
input G5;
input G9;
input G3;
input G13;
input G4;
input G12;
input G2;
input blif_clk_net;
input G7;
input blif_reset_net;
input G10;
input G0;
input G6;

// Start POs
output G549;
output G542;
output G530;
output G552;
output G45;
output G547;
output G548;
output G537;
output G551;
output G532;
output G539;
output G546;
output G535;
output G550;

// Start wires
wire net_568;
wire net_47;
wire net_416;
wire net_215;
wire net_54;
wire net_526;
wire G546;
wire net_429;
wire net_557;
wire net_129;
wire net_373;
wire net_119;
wire net_98;
wire net_151;
wire net_356;
wire net_53;
wire net_452;
wire net_210;
wire net_545;
wire net_284;
wire net_168;
wire net_560;
wire G6;
wire net_477;
wire net_439;
wire net_385;
wire net_259;
wire net_269;
wire net_548;
wire net_469;
wire net_501;
wire net_187;
wire net_111;
wire net_264;
wire net_90;
wire net_225;
wire net_283;
wire net_85;
wire net_263;
wire net_252;
wire net_124;
wire net_343;
wire net_404;
wire net_240;
wire net_160;
wire net_322;
wire net_511;
wire net_4;
wire net_420;
wire net_447;
wire net_295;
wire net_410;
wire net_508;
wire net_390;
wire net_307;
wire net_35;
wire net_586;
wire net_344;
wire net_16;
wire net_239;
wire net_193;
wire net_257;
wire net_310;
wire net_233;
wire net_474;
wire net_120;
wire net_292;
wire net_201;
wire net_472;
wire net_109;
wire net_80;
wire net_65;
wire net_96;
wire net_484;
wire net_167;
wire net_207;
wire net_136;
wire net_280;
wire net_126;
wire net_495;
wire net_278;
wire net_34;
wire net_458;
wire net_108;
wire net_598;
wire net_571;
wire net_63;
wire net_593;
wire net_617;
wire net_601;
wire net_274;
wire net_554;
wire net_425;
wire net_321;
wire net_287;
wire net_189;
wire net_490;
wire G551;
wire G539;
wire net_99;
wire net_46;
wire net_480;
wire net_216;
wire net_433;
wire net_584;
wire net_544;
wire net_368;
wire net_224;
wire net_52;
wire net_538;
wire net_165;
wire net_608;
wire net_510;
wire net_370;
wire net_464;
wire net_366;
wire net_13;
wire net_413;
wire net_446;
wire net_114;
wire G13;
wire net_248;
wire net_384;
wire net_36;
wire net_198;
wire net_253;
wire net_311;
wire net_276;
wire G45;
wire net_494;
wire net_209;
wire net_3;
wire net_547;
wire net_294;
wire net_154;
wire net_507;
wire net_616;
wire net_371;
wire net_238;
wire net_529;
wire net_28;
wire G532;
wire net_587;
wire net_485;
wire net_97;
wire net_192;
wire G9;
wire net_503;
wire net_256;
wire net_460;
wire net_82;
wire net_64;
wire net_457;
wire net_291;
wire net_121;
wire net_597;
wire net_200;
wire net_308;
wire net_75;
wire net_515;
wire net_600;
wire net_396;
wire net_206;
wire net_195;
wire net_125;
wire net_397;
wire net_107;
wire net_166;
wire net_223;
wire net_235;
wire net_530;
wire net_606;
wire net_623;
wire net_603;
wire net_594;
wire net_320;
wire net_271;
wire net_23;
wire net_117;
wire net_74;
wire net_579;
wire net_401;
wire net_250;
wire net_205;
wire net_242;
wire net_312;
wire net_130;
wire net_572;
wire net_359;
wire net_440;
wire net_286;
wire G11;
wire net_147;
wire net_481;
wire net_369;
wire net_470;
wire net_26;
wire net_403;
wire net_334;
wire blif_clk_net;
wire net_32;
wire net_430;
wire net_365;
wire net_282;
wire net_426;
wire net_380;
wire net_141;
wire net_467;
wire net_83;
wire net_609;
wire net_541;
wire net_414;
wire net_372;
wire net_437;
wire net_528;
wire net_56;
wire net_566;
wire net_456;
wire net_155;
wire net_335;
wire net_506;
wire net_181;
wire net_336;
wire net_624;
wire net_349;
wire net_39;
wire net_555;
wire net_245;
wire net_2;
wire net_9;
wire net_395;
wire net_331;
wire net_298;
wire net_493;
wire net_475;
wire G549;
wire G8;
wire net_563;
wire net_386;
wire net_605;
wire net_277;
wire net_199;
wire net_502;
wire net_431;
wire net_89;
wire net_290;
wire net_338;
wire net_243;
wire net_400;
wire net_222;
wire net_602;
wire net_313;
wire net_152;
wire net_489;
wire net_175;
wire net_106;
wire net_607;
wire net_258;
wire net_140;
wire net_247;
wire net_329;
wire net_279;
wire net_148;
wire net_419;
wire net_25;
wire net_70;
wire net_251;
wire net_194;
wire net_615;
wire net_478;
wire net_244;
wire net_585;
wire net_441;
wire net_128;
wire net_596;
wire net_138;
wire net_333;
wire net_549;
wire net_374;
wire net_411;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_77;
wire net_214;
wire net_249;
wire net_20;
wire net_49;
wire net_518;
wire G1;
wire net_15;
wire net_57;
wire net_71;
wire net_156;
wire net_394;
wire net_92;
wire net_1;
wire net_112;
wire net_139;
wire net_551;
wire net_537;
wire net_332;
wire net_180;
wire net_409;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire G550;
wire net_492;
wire net_463;
wire net_432;
wire net_88;
wire net_197;
wire net_513;
wire net_204;
wire net_81;
wire net_232;
wire net_604;
wire net_163;
wire net_402;
wire net_67;
wire net_202;
wire net_268;
wire net_110;
wire net_379;
wire net_459;
wire net_483;
wire net_48;
wire net_33;
wire net_8;
wire net_203;
wire net_450;
wire net_289;
wire net_505;
wire net_621;
wire net_435;
wire net_176;
wire net_137;
wire net_296;
wire net_132;
wire net_613;
wire net_237;
wire net_105;
wire net_614;
wire net_532;
wire net_12;
wire net_93;
wire net_578;
wire net_302;
wire net_569;
wire net_127;
wire net_327;
wire net_357;
wire net_348;
wire net_76;
wire net_626;
wire net_101;
wire net_388;
wire net_326;
wire net_353;
wire net_589;
wire net_519;
wire net_100;
wire net_412;
wire net_536;
wire net_455;
wire net_221;
wire net_115;
wire net_393;
wire net_442;
wire net_17;
wire net_319;
wire net_542;
wire net_453;
wire net_575;
wire net_595;
wire net_581;
wire net_378;
wire net_164;
wire net_408;
wire net_377;
wire net_87;
wire net_0;
wire net_288;
wire net_423;
wire net_328;
wire net_157;
wire net_540;
wire net_512;
wire net_42;
wire blif_reset_net;
wire net_50;
wire net_234;
wire net_38;
wire net_66;
wire net_466;
wire net_342;
wire net_612;
wire net_19;
wire net_443;
wire net_504;
wire net_522;
wire net_270;
wire net_183;
wire net_618;
wire net_150;
wire G0;
wire net_303;
wire net_304;
wire net_352;
wire net_491;
wire net_30;
wire net_436;
wire net_24;
wire net_392;
wire net_622;
wire net_186;
wire net_118;
wire net_421;
wire net_146;
wire net_550;
wire net_122;
wire net_417;
wire net_7;
wire net_172;
wire net_428;
wire net_94;
wire net_246;
wire net_461;
wire net_219;
wire net_18;
wire G542;
wire net_309;
wire net_482;
wire net_131;
wire net_196;
wire net_29;
wire net_358;
wire net_142;
wire net_149;
wire net_516;
wire net_31;
wire net_387;
wire net_330;
wire net_535;
wire net_498;
wire net_158;
wire net_41;
wire G3;
wire net_577;
wire net_360;
wire net_570;
wire net_525;
wire net_444;
wire net_213;
wire net_325;
wire net_301;
wire net_260;
wire G547;
wire net_299;
wire net_438;
wire net_580;
wire net_314;
wire net_182;
wire net_521;
wire net_60;
wire net_590;
wire net_337;
wire net_341;
wire net_267;
wire net_273;
wire net_424;
wire net_468;
wire net_58;
wire net_576;
wire net_488;
wire net_73;
wire G5;
wire net_465;
wire net_86;
wire net_177;
wire net_523;
wire G12;
wire net_407;
wire net_476;
wire net_564;
wire net_382;
wire net_179;
wire net_159;
wire G552;
wire net_61;
wire net_583;
wire net_449;
wire net_383;
wire net_62;
wire net_6;
wire net_553;
wire net_534;
wire net_217;
wire net_351;
wire net_427;
wire net_486;
wire net_135;
wire net_340;
wire net_265;
wire net_517;
wire net_434;
wire net_406;
wire net_473;
wire net_220;
wire net_14;
wire net_293;
wire net_324;
wire net_113;
wire net_497;
wire net_454;
wire net_418;
wire net_462;
wire net_40;
wire net_69;
wire net_543;
wire net_161;
wire net_625;
wire net_300;
wire net_339;
wire net_95;
wire net_173;
wire net_361;
wire net_78;
wire net_27;
wire net_317;
wire net_305;
wire G2;
wire net_514;
wire net_191;
wire net_261;
wire net_22;
wire net_376;
wire net_558;
wire net_354;
wire net_524;
wire net_144;
wire net_102;
wire net_227;
wire net_59;
wire G548;
wire net_363;
wire net_445;
wire net_573;
wire net_162;
wire net_44;
wire net_230;
wire net_520;
wire net_422;
wire net_134;
wire net_546;
wire net_561;
wire net_567;
wire net_45;
wire net_381;
wire net_591;
wire net_185;
wire net_588;
wire net_272;
wire G4;
wire net_178;
wire net_208;
wire net_236;
wire G535;
wire net_487;
wire net_212;
wire G10;
wire net_315;
wire net_552;
wire net_415;
wire net_116;
wire net_556;
wire net_347;
wire G537;
wire net_91;
wire net_297;
wire net_346;
wire G7;
wire net_55;
wire net_559;
wire net_255;
wire net_266;
wire net_345;
wire net_104;
wire net_620;
wire net_448;
wire net_619;
wire net_72;
wire net_350;
wire net_229;
wire net_398;
wire net_306;
wire net_241;
wire net_5;
wire net_405;
wire net_500;
wire net_355;
wire net_184;
wire net_599;
wire net_11;
wire net_610;
wire net_123;
wire net_527;
wire net_262;
wire net_362;
wire net_389;
wire net_68;
wire net_318;
wire net_451;
wire net_323;
wire net_275;
wire net_539;
wire net_399;
wire net_153;
wire net_316;
wire net_218;
wire net_84;
wire net_174;
wire net_611;
wire net_231;
wire net_562;
wire net_103;
wire net_375;
wire net_226;
wire net_364;
wire net_43;
wire net_10;
wire net_228;
wire net_592;
wire net_21;
wire net_79;
wire net_143;
wire net_190;
wire net_391;
wire net_533;
wire net_145;
wire net_285;
wire net_281;
wire net_254;
wire net_37;
wire net_582;
wire net_188;
wire net_496;
wire G530;
wire net_509;
wire net_574;
wire net_479;
wire net_211;
wire net_133;

// Start cells
INV_X2 inst_537 ( .ZN(net_245), .A(net_244) );
INV_X4 inst_481 ( .A(net_195), .ZN(net_162) );
DFFR_X1 inst_551 ( .RN(net_464), .D(net_264), .Q(net_8), .CK(net_623) );
NAND2_X2 inst_228 ( .ZN(net_141), .A2(net_50), .A1(net_22) );
NAND4_X2 inst_125 ( .ZN(net_568), .A3(net_480), .A1(net_479), .A4(net_438), .A2(net_429) );
INV_X4 inst_486 ( .A(net_227), .ZN(net_220) );
INV_X2 inst_506 ( .A(net_536), .ZN(net_535) );
INV_X4 inst_495 ( .ZN(net_381), .A(net_374) );
INV_X4 inst_353 ( .A(net_562), .ZN(net_561) );
NAND2_X4 inst_207 ( .A2(net_563), .A1(net_487), .ZN(net_190) );
NAND3_X2 inst_159 ( .A2(net_527), .A3(net_522), .ZN(net_481), .A1(net_151) );
INV_X4 inst_395 ( .ZN(net_478), .A(G7) );
NAND3_X2 inst_134 ( .A3(net_519), .ZN(net_144), .A2(net_133), .A1(net_53) );
NAND2_X2 inst_244 ( .ZN(net_173), .A2(net_148), .A1(net_99) );
NAND2_X2 inst_333 ( .A2(net_440), .A1(net_403), .ZN(G547) );
INV_X4 inst_452 ( .ZN(net_77), .A(net_76) );
INV_X4 inst_430 ( .A(net_334), .ZN(net_169) );
NAND3_X4 inst_131 ( .ZN(net_551), .A2(net_544), .A1(net_543), .A3(net_469) );
INV_X4 inst_406 ( .A(net_72), .ZN(net_26) );
NAND2_X4 inst_214 ( .A2(net_538), .ZN(net_430), .A1(net_415) );
INV_X4 inst_462 ( .ZN(net_145), .A(net_99) );
NAND3_X2 inst_160 ( .ZN(net_531), .A1(net_371), .A2(net_312), .A3(net_77) );
NAND2_X2 inst_328 ( .A1(net_531), .ZN(net_444), .A2(net_442) );
NOR2_X2 inst_47 ( .A1(net_520), .ZN(net_66), .A2(G4) );
OR2_X2 inst_19 ( .ZN(net_537), .A1(net_381), .A2(net_2) );
DFFR_X2 inst_548 ( .QN(net_527), .RN(net_464), .D(net_236), .CK(net_622) );
INV_X2 inst_515 ( .ZN(net_507), .A(G6) );
OR2_X4 inst_8 ( .ZN(net_230), .A2(net_213), .A1(net_158) );
INV_X4 inst_370 ( .ZN(net_502), .A(net_501) );
AND2_X4 inst_573 ( .ZN(net_355), .A2(net_354), .A1(net_206) );
NOR2_X2 inst_100 ( .ZN(net_336), .A1(net_335), .A2(net_321) );
INV_X4 inst_459 ( .ZN(net_262), .A(net_180) );
NAND2_X2 inst_279 ( .ZN(net_291), .A2(net_225), .A1(net_166) );
INV_X4 inst_445 ( .A(net_206), .ZN(net_96) );
NOR2_X2 inst_93 ( .ZN(net_288), .A2(net_287), .A1(net_63) );
NOR2_X2 inst_81 ( .ZN(net_235), .A2(net_160), .A1(net_59) );
CLKBUF_X2 inst_612 ( .A(net_597), .Z(net_598) );
CLKBUF_X2 inst_606 ( .A(net_591), .Z(net_592) );
INV_X4 inst_367 ( .ZN(net_548), .A(G6) );
INV_X2 inst_525 ( .A(net_42), .ZN(net_33) );
NAND3_X2 inst_139 ( .ZN(net_241), .A1(net_238), .A3(net_217), .A2(net_169) );
DFFR_X1 inst_559 ( .RN(net_464), .D(net_377), .QN(net_9), .CK(net_586) );
CLKBUF_X2 inst_584 ( .A(blif_clk_net), .Z(net_570) );
INV_X2 inst_521 ( .A(net_496), .ZN(net_495) );
INV_X4 inst_434 ( .ZN(net_80), .A(net_49) );
INV_X4 inst_470 ( .ZN(net_160), .A(net_124) );
INV_X2 inst_535 ( .ZN(net_242), .A(net_164) );
INV_X4 inst_450 ( .ZN(net_270), .A(net_68) );
INV_X2 inst_520 ( .A(net_498), .ZN(net_497) );
NAND2_X2 inst_237 ( .A1(net_559), .A2(net_169), .ZN(net_106) );
NAND3_X2 inst_148 ( .ZN(net_300), .A3(net_275), .A2(net_229), .A1(net_110) );
DFFR_X1 inst_554 ( .RN(net_464), .D(net_330), .Q(net_5), .CK(net_603) );
INV_X4 inst_377 ( .ZN(net_14), .A(G8) );
NAND3_X1 inst_191 ( .A2(net_513), .A3(net_492), .ZN(net_472), .A1(net_191) );
NOR2_X2 inst_51 ( .A1(net_562), .ZN(net_213), .A2(net_15) );
NAND3_X2 inst_142 ( .ZN(net_475), .A3(net_254), .A2(net_212), .A1(net_115) );
NAND2_X2 inst_315 ( .ZN(net_407), .A2(net_392), .A1(net_386) );
NOR2_X2 inst_80 ( .ZN(net_189), .A2(net_188), .A1(net_107) );
NAND2_X4 inst_216 ( .ZN(net_488), .A2(net_486), .A1(net_432) );
NOR2_X2 inst_78 ( .ZN(net_179), .A2(net_178), .A1(net_136) );
NAND2_X2 inst_241 ( .A2(net_493), .ZN(net_116), .A1(net_115) );
NAND3_X2 inst_177 ( .A3(net_492), .ZN(net_450), .A1(net_449), .A2(net_347) );
NAND3_X2 inst_183 ( .ZN(net_458), .A3(net_454), .A2(net_436), .A1(net_395) );
NAND3_X2 inst_151 ( .ZN(net_333), .A2(net_332), .A3(net_291), .A1(net_241) );
NOR2_X2 inst_64 ( .A1(net_148), .ZN(net_129), .A2(net_128) );
INV_X4 inst_415 ( .ZN(net_49), .A(net_37) );
CLKBUF_X2 inst_615 ( .A(net_596), .Z(net_601) );
INV_X4 inst_393 ( .ZN(net_37), .A(G4) );
NOR2_X2 inst_107 ( .ZN(net_359), .A2(net_351), .A1(net_186) );
NOR2_X2 inst_92 ( .ZN(net_273), .A1(net_272), .A2(net_202) );
MUX2_X2 inst_345 ( .B(net_120), .Z(net_102), .A(net_101), .S(net_18) );
NAND2_X2 inst_223 ( .ZN(net_70), .A2(net_13), .A1(G3) );
INV_X4 inst_402 ( .A(net_28), .ZN(net_25) );
NAND2_X2 inst_340 ( .A2(net_466), .A1(net_452), .ZN(G532) );
INV_X4 inst_494 ( .ZN(net_378), .A(net_363) );
INV_X4 inst_487 ( .ZN(net_239), .A(net_187) );
NAND2_X2 inst_329 ( .ZN(net_445), .A2(net_426), .A1(net_333) );
AND2_X4 inst_574 ( .A1(net_420), .ZN(net_393), .A2(net_383) );
INV_X4 inst_386 ( .A(net_19), .ZN(net_15) );
NAND3_X2 inst_158 ( .ZN(net_544), .A1(net_485), .A2(net_74), .A3(net_72) );
NAND3_X2 inst_141 ( .A2(net_334), .ZN(net_243), .A3(net_242), .A1(net_149) );
NAND2_X4 inst_200 ( .A2(net_521), .ZN(net_90), .A1(net_54) );
INV_X2 inst_507 ( .A(net_535), .ZN(net_533) );
AND2_X4 inst_571 ( .A2(net_493), .ZN(net_212), .A1(G11) );
NOR2_X2 inst_57 ( .A1(net_133), .ZN(net_86), .A2(net_85) );
NAND2_X2 inst_338 ( .ZN(net_465), .A1(net_462), .A2(net_455) );
DFFR_X1 inst_552 ( .RN(net_464), .D(net_305), .Q(net_12), .CK(net_612) );
CLKBUF_X2 inst_599 ( .A(net_584), .Z(net_585) );
INV_X4 inst_417 ( .ZN(net_115), .A(net_42) );
AND2_X2 inst_579 ( .ZN(net_142), .A2(net_141), .A1(net_79) );
OR2_X2 inst_21 ( .ZN(net_437), .A2(net_436), .A1(net_378) );
INV_X4 inst_469 ( .ZN(net_215), .A(net_178) );
NAND2_X2 inst_281 ( .A1(net_500), .ZN(net_299), .A2(net_237) );
CLKBUF_X2 inst_585 ( .A(net_570), .Z(net_571) );
OR2_X2 inst_18 ( .A1(net_538), .ZN(net_375), .A2(net_332) );
INV_X2 inst_541 ( .A(net_365), .ZN(net_358) );
INV_X4 inst_410 ( .ZN(net_312), .A(net_29) );
NAND2_X4 inst_208 ( .ZN(net_522), .A1(net_474), .A2(net_75) );
NOR2_X2 inst_88 ( .A1(net_416), .ZN(net_234), .A2(net_129) );
NAND2_X2 inst_316 ( .ZN(net_412), .A2(net_411), .A1(net_366) );
NAND2_X2 inst_220 ( .ZN(net_520), .A2(G3), .A1(G1) );
OR2_X4 inst_9 ( .ZN(net_539), .A1(net_527), .A2(net_14) );
NOR2_X2 inst_113 ( .ZN(net_390), .A2(net_384), .A1(net_383) );
INV_X2 inst_505 ( .A(net_555), .ZN(net_554) );
INV_X4 inst_356 ( .A(net_555), .ZN(net_553) );
INV_X4 inst_383 ( .A(net_44), .ZN(net_22) );
INV_X4 inst_360 ( .A(net_529), .ZN(net_528) );
NAND2_X4 inst_198 ( .A2(net_494), .ZN(net_117), .A1(net_37) );
NOR2_X2 inst_50 ( .ZN(net_526), .A1(net_42), .A2(net_34) );
NAND2_X2 inst_245 ( .ZN(net_195), .A2(net_123), .A1(net_50) );
AND2_X4 inst_569 ( .ZN(net_35), .A2(G11), .A1(G9) );
CLKBUF_X2 inst_624 ( .A(net_609), .Z(net_610) );
NAND2_X2 inst_260 ( .ZN(net_194), .A1(net_173), .A2(net_61) );
NAND3_X2 inst_147 ( .ZN(net_545), .A3(net_540), .A1(net_536), .A2(net_182) );
NAND2_X2 inst_313 ( .ZN(net_486), .A1(net_98), .A2(net_4) );
NAND2_X2 inst_293 ( .ZN(net_329), .A2(net_314), .A1(net_245) );
CLKBUF_X2 inst_636 ( .A(net_621), .Z(net_622) );
CLKBUF_X2 inst_632 ( .A(net_595), .Z(net_618) );
DFFR_X2 inst_549 ( .RN(net_464), .D(net_290), .QN(net_1), .CK(net_619) );
NAND2_X2 inst_234 ( .A1(net_508), .ZN(net_84), .A2(net_45) );
XNOR2_X2 inst_0 ( .ZN(net_264), .A(net_263), .B(net_262) );
INV_X2 inst_522 ( .ZN(net_13), .A(G2) );
NAND3_X2 inst_184 ( .ZN(net_461), .A1(net_460), .A2(net_311), .A3(net_7) );
NAND2_X2 inst_236 ( .A2(net_200), .ZN(net_168), .A1(G6) );
INV_X4 inst_433 ( .ZN(net_200), .A(net_70) );
DFFR_X1 inst_553 ( .Q(net_547), .RN(net_464), .D(net_303), .CK(net_607) );
INV_X4 inst_478 ( .ZN(net_187), .A(net_159) );
NOR2_X2 inst_65 ( .A2(net_525), .A1(net_507), .ZN(net_130) );
INV_X2 inst_536 ( .ZN(net_219), .A(net_218) );
NAND2_X2 inst_242 ( .ZN(net_118), .A1(net_117), .A2(net_69) );
INV_X2 inst_516 ( .A(net_507), .ZN(net_506) );
NOR2_X2 inst_98 ( .ZN(net_310), .A2(net_288), .A1(net_159) );
NAND2_X2 inst_263 ( .ZN(net_211), .A2(net_209), .A1(net_178) );
NAND3_X1 inst_190 ( .A1(net_557), .ZN(net_429), .A3(net_425), .A2(net_252) );
NAND3_X2 inst_185 ( .A2(net_451), .A3(net_423), .A1(net_417), .ZN(G551) );
OR2_X2 inst_13 ( .ZN(net_170), .A1(net_169), .A2(net_168) );
NOR2_X2 inst_75 ( .ZN(net_171), .A2(net_132), .A1(net_96) );
NAND2_X2 inst_332 ( .ZN(net_479), .A2(net_435), .A1(net_337) );
NAND3_X2 inst_166 ( .A2(net_420), .ZN(net_402), .A3(net_396), .A1(net_318) );
NOR2_X1 inst_116 ( .A2(net_495), .ZN(net_175), .A1(net_140) );
CLKBUF_X2 inst_598 ( .A(net_583), .Z(net_584) );
INV_X4 inst_416 ( .A(net_72), .ZN(net_36) );
NAND3_X2 inst_163 ( .A3(net_387), .ZN(net_386), .A2(net_384), .A1(net_204) );
INV_X4 inst_471 ( .ZN(net_192), .A(net_134) );
INV_X4 inst_394 ( .A(net_35), .ZN(net_31) );
NOR2_X2 inst_79 ( .ZN(net_186), .A1(net_185), .A2(net_154) );
NOR2_X2 inst_106 ( .ZN(net_357), .A2(net_343), .A1(net_272) );
INV_X4 inst_422 ( .ZN(net_57), .A(net_39) );
NAND2_X2 inst_219 ( .ZN(net_24), .A2(G5), .A1(G3) );
NAND2_X4 inst_201 ( .A1(net_553), .ZN(net_88), .A2(net_19) );
CLKBUF_X2 inst_605 ( .A(net_576), .Z(net_591) );
NAND2_X2 inst_304 ( .ZN(net_541), .A2(net_378), .A1(net_319) );
INV_X2 inst_542 ( .ZN(net_406), .A(net_405) );
NAND2_X2 inst_255 ( .A1(net_497), .A2(net_203), .ZN(net_191) );
INV_X4 inst_453 ( .ZN(net_335), .A(net_79) );
NAND3_X4 inst_128 ( .ZN(net_93), .A2(net_92), .A3(net_91), .A1(net_52) );
NOR2_X2 inst_73 ( .A2(net_334), .ZN(net_317), .A1(net_145) );
INV_X4 inst_493 ( .ZN(net_350), .A(net_340) );
INV_X4 inst_378 ( .ZN(net_19), .A(G1) );
NOR4_X2 inst_23 ( .A3(net_496), .ZN(net_307), .A4(net_306), .A1(net_221), .A2(net_94) );
NAND2_X2 inst_339 ( .A1(net_568), .ZN(net_466), .A2(net_456) );
INV_X8 inst_351 ( .ZN(net_75), .A(net_32) );
INV_X4 inst_361 ( .A(net_526), .ZN(net_525) );
INV_X4 inst_408 ( .A(net_210), .ZN(net_148) );
NAND2_X2 inst_325 ( .ZN(net_567), .A2(net_428), .A1(net_375) );
INV_X4 inst_461 ( .A(net_335), .ZN(net_95) );
INV_X4 inst_385 ( .ZN(net_41), .A(net_14) );
NAND2_X4 inst_197 ( .ZN(net_45), .A2(net_41), .A1(net_35) );
NAND2_X2 inst_250 ( .ZN(net_157), .A2(net_89), .A1(G6) );
NAND3_X2 inst_179 ( .A3(net_492), .ZN(net_452), .A1(net_368), .A2(net_308) );
NOR4_X2 inst_24 ( .ZN(net_377), .A4(net_367), .A2(net_345), .A3(net_307), .A1(net_207) );
NOR2_X2 inst_114 ( .A2(net_537), .ZN(net_400), .A1(G12) );
CLKBUF_X2 inst_617 ( .A(net_602), .Z(net_603) );
NOR2_X2 inst_76 ( .A1(net_200), .ZN(net_172), .A2(net_164) );
INV_X4 inst_397 ( .ZN(net_48), .A(net_21) );
INV_X2 inst_504 ( .A(net_558), .ZN(net_557) );
NAND3_X2 inst_150 ( .ZN(net_331), .A1(net_280), .A3(net_276), .A2(net_184) );
NAND3_X2 inst_172 ( .ZN(net_417), .A1(net_416), .A3(net_411), .A2(net_8) );
INV_X4 inst_362 ( .A(net_526), .ZN(net_523) );
NAND2_X2 inst_277 ( .ZN(net_289), .A2(net_283), .A1(net_119) );
NOR2_X2 inst_83 ( .ZN(net_198), .A1(net_192), .A2(net_141) );
NAND4_X2 inst_121 ( .ZN(net_294), .A1(net_177), .A3(net_168), .A4(net_157), .A2(net_106) );
INV_X2 inst_534 ( .ZN(net_136), .A(net_135) );
INV_X4 inst_440 ( .ZN(net_58), .A(net_57) );
NAND2_X2 inst_306 ( .ZN(net_484), .A2(net_379), .A1(net_50) );
OR3_X4 inst_2 ( .ZN(net_339), .A2(net_338), .A3(net_337), .A1(net_310) );
CLKBUF_X2 inst_596 ( .A(net_581), .Z(net_582) );
AND2_X2 inst_578 ( .ZN(net_138), .A2(net_137), .A1(net_91) );
NOR2_X2 inst_52 ( .ZN(net_137), .A2(net_56), .A1(G3) );
NOR2_X2 inst_90 ( .ZN(net_249), .A2(net_215), .A1(net_171) );
NAND2_X2 inst_267 ( .ZN(net_229), .A1(net_222), .A2(net_60) );
NAND3_X2 inst_140 ( .ZN(net_267), .A3(net_199), .A1(net_50), .A2(net_29) );
NAND2_X2 inst_221 ( .ZN(net_521), .A1(net_19), .A2(G5) );
DFFR_X1 inst_556 ( .RN(net_464), .D(net_352), .QN(net_11), .CK(net_599) );
CLKBUF_X2 inst_637 ( .A(net_581), .Z(net_623) );
NAND2_X2 inst_289 ( .ZN(net_319), .A2(net_277), .A1(net_155) );
DFFR_X2 inst_547 ( .RN(net_464), .D(net_248), .QN(net_6), .CK(net_624) );
INV_X2 inst_530 ( .A(net_335), .ZN(net_104) );
INV_X4 inst_432 ( .ZN(net_133), .A(net_47) );
INV_X4 inst_420 ( .ZN(net_542), .A(net_50) );
NAND2_X2 inst_282 ( .A1(net_554), .A2(net_534), .ZN(net_332) );
INV_X4 inst_368 ( .A(net_505), .ZN(net_504) );
INV_X2 inst_513 ( .A(net_511), .ZN(net_510) );
NOR2_X4 inst_44 ( .A2(net_551), .A1(net_550), .ZN(net_413) );
NAND2_X2 inst_274 ( .A1(net_511), .ZN(net_279), .A2(net_208) );
NAND3_X2 inst_174 ( .A2(net_517), .A1(net_456), .ZN(net_422), .A3(net_406) );
INV_X4 inst_371 ( .A(net_499), .ZN(net_496) );
NAND2_X2 inst_314 ( .ZN(net_399), .A1(net_326), .A2(net_4) );
INV_X4 inst_435 ( .A(net_148), .ZN(net_64) );
NAND3_X2 inst_164 ( .ZN(net_480), .A3(net_387), .A2(net_11), .A1(G13) );
OR3_X2 inst_5 ( .ZN(net_318), .A2(net_317), .A3(net_246), .A1(net_234) );
CLKBUF_X2 inst_597 ( .A(blif_clk_net), .Z(net_583) );
NAND3_X2 inst_157 ( .ZN(net_371), .A1(net_362), .A2(net_286), .A3(net_271) );
CLKBUF_X2 inst_621 ( .A(net_606), .Z(net_607) );
NOR2_X2 inst_68 ( .A2(net_384), .ZN(net_297), .A1(net_58) );
NAND2_X4 inst_213 ( .A1(net_517), .ZN(net_415), .A2(net_405) );
CLKBUF_X2 inst_604 ( .A(net_589), .Z(net_590) );
NOR2_X2 inst_53 ( .A1(net_507), .ZN(net_247), .A2(net_101) );
CLKBUF_X2 inst_628 ( .A(net_613), .Z(net_614) );
NAND2_X4 inst_205 ( .ZN(net_209), .A1(net_131), .A2(net_43) );
INV_X4 inst_472 ( .ZN(net_159), .A(net_140) );
INV_X4 inst_447 ( .A(net_117), .ZN(net_65) );
INV_X4 inst_380 ( .ZN(net_20), .A(net_14) );
INV_X4 inst_457 ( .ZN(net_275), .A(net_90) );
NAND2_X2 inst_292 ( .ZN(net_327), .A2(net_299), .A1(net_194) );
INV_X4 inst_379 ( .ZN(net_50), .A(net_13) );
NAND4_X2 inst_127 ( .A2(net_468), .A1(net_443), .A4(net_421), .A3(net_410), .ZN(G550) );
NAND3_X2 inst_186 ( .A3(net_532), .A2(net_448), .A1(net_404), .ZN(G542) );
OR2_X2 inst_17 ( .ZN(net_286), .A2(net_285), .A1(net_44) );
INV_X4 inst_413 ( .ZN(net_46), .A(net_31) );
NAND3_X2 inst_146 ( .ZN(net_276), .A3(net_275), .A2(net_255), .A1(net_230) );
NAND2_X2 inst_249 ( .ZN(net_153), .A1(net_152), .A2(net_135) );
NAND2_X2 inst_334 ( .A2(net_447), .A1(net_399), .ZN(G548) );
NAND3_X2 inst_187 ( .A1(net_532), .A3(net_472), .ZN(net_463), .A2(net_398) );
NAND2_X4 inst_206 ( .ZN(net_536), .A2(net_116), .A1(net_93) );
NAND4_X2 inst_122 ( .A4(net_476), .A1(net_475), .ZN(net_309), .A2(net_257), .A3(net_214) );
NOR4_X2 inst_25 ( .A1(net_549), .ZN(net_453), .A2(net_416), .A4(net_388), .A3(net_57) );
INV_X4 inst_354 ( .ZN(net_560), .A(G3) );
INV_X4 inst_405 ( .ZN(net_40), .A(net_25) );
INV_X4 inst_492 ( .ZN(net_268), .A(net_267) );
NAND2_X2 inst_240 ( .A1(net_506), .A2(net_493), .ZN(net_114) );
NAND2_X2 inst_326 ( .ZN(net_441), .A2(net_431), .A1(net_380) );
NOR2_X2 inst_110 ( .ZN(net_373), .A2(net_361), .A1(net_349) );
INV_X2 inst_518 ( .ZN(net_503), .A(net_501) );
NOR2_X2 inst_74 ( .ZN(net_165), .A1(net_87), .A2(net_82) );
NAND2_X2 inst_288 ( .A1(net_558), .ZN(net_316), .A2(net_268) );
INV_X4 inst_396 ( .ZN(net_210), .A(net_56) );
NAND2_X2 inst_229 ( .ZN(net_67), .A2(net_66), .A1(G6) );
NOR2_X2 inst_99 ( .ZN(net_313), .A2(net_295), .A1(net_203) );
NOR2_X2 inst_69 ( .A2(net_493), .ZN(net_185), .A1(net_43) );
INV_X4 inst_373 ( .ZN(net_427), .A(G13) );
NOR2_X2 inst_82 ( .A2(net_514), .A1(net_504), .ZN(net_238) );
NOR2_X2 inst_108 ( .A2(net_522), .ZN(net_367), .A1(net_344) );
CLKBUF_X2 inst_595 ( .A(net_577), .Z(net_581) );
NAND2_X2 inst_283 ( .A2(net_533), .A1(net_500), .ZN(net_301) );
NOR4_X2 inst_22 ( .A2(net_497), .ZN(net_205), .A1(net_204), .A3(net_203), .A4(net_143) );
NAND2_X2 inst_311 ( .ZN(net_397), .A2(net_396), .A1(net_243) );
INV_X4 inst_460 ( .ZN(net_272), .A(net_94) );
INV_X4 inst_372 ( .ZN(net_494), .A(G6) );
NAND3_X2 inst_169 ( .ZN(net_408), .A1(net_397), .A3(net_391), .A2(net_389) );
NAND2_X4 inst_215 ( .A2(net_499), .A1(net_492), .ZN(net_432) );
NAND2_X2 inst_307 ( .ZN(net_391), .A2(net_390), .A1(net_200) );
CLKBUF_X2 inst_638 ( .A(net_615), .Z(net_624) );
INV_X4 inst_421 ( .ZN(net_60), .A(net_38) );
NAND3_X2 inst_161 ( .ZN(net_379), .A3(net_364), .A2(net_285), .A1(net_278) );
DFFR_X1 inst_560 ( .RN(net_464), .D(net_382), .Q(net_4), .CK(net_582) );
CLKBUF_X2 inst_586 ( .A(net_571), .Z(net_572) );
DFFR_X1 inst_555 ( .RN(net_464), .D(net_348), .QN(net_0), .CK(net_600) );
OR2_X2 inst_16 ( .ZN(net_253), .A1(net_197), .A2(net_176) );
NAND2_X2 inst_276 ( .A2(net_334), .ZN(net_282), .A1(net_281) );
INV_X4 inst_431 ( .ZN(net_231), .A(net_46) );
INV_X8 inst_348 ( .A(net_507), .ZN(net_499) );
OR3_X2 inst_3 ( .A2(net_317), .ZN(net_274), .A1(net_201), .A3(net_174) );
NAND3_X2 inst_156 ( .ZN(net_362), .A3(net_342), .A2(net_270), .A1(net_216) );
AND2_X4 inst_577 ( .A1(net_427), .ZN(net_411), .A2(net_400) );
AND3_X4 inst_566 ( .A2(net_495), .A3(net_217), .ZN(net_207), .A1(net_206) );
NAND2_X2 inst_296 ( .ZN(net_341), .A2(net_324), .A1(net_242) );
NOR2_X2 inst_91 ( .ZN(net_261), .A1(net_260), .A2(net_259) );
NAND3_X2 inst_132 ( .A3(net_554), .ZN(net_154), .A1(net_120), .A2(net_119) );
NAND2_X2 inst_342 ( .A2(net_467), .A1(net_445), .ZN(G537) );
INV_X2 inst_526 ( .A(net_148), .ZN(net_51) );
NOR3_X2 inst_36 ( .ZN(net_349), .A3(net_2), .A1(G13), .A2(G12) );
INV_X4 inst_463 ( .A(net_335), .ZN(net_100) );
INV_X2 inst_503 ( .A(net_559), .ZN(net_558) );
NOR2_X2 inst_96 ( .ZN(net_296), .A2(net_258), .A1(net_231) );
NOR2_X4 inst_45 ( .ZN(net_460), .A1(net_454), .A2(net_85) );
INV_X4 inst_451 ( .ZN(net_103), .A(net_74) );
NOR2_X2 inst_101 ( .A2(net_529), .ZN(net_340), .A1(net_1) );
NAND2_X2 inst_319 ( .A1(net_554), .A2(net_425), .ZN(net_424) );
NAND2_X2 inst_269 ( .ZN(net_240), .A1(net_239), .A2(net_238) );
INV_X4 inst_458 ( .A(net_203), .ZN(net_140) );
INV_X4 inst_444 ( .A(net_206), .ZN(net_63) );
INV_X4 inst_400 ( .A(net_92), .ZN(net_23) );
CLKBUF_X2 inst_614 ( .A(net_586), .Z(net_600) );
NAND2_X2 inst_261 ( .A1(net_498), .ZN(net_196), .A2(net_195) );
INV_X2 inst_514 ( .A(net_515), .ZN(net_509) );
INV_X2 inst_500 ( .A(net_564), .ZN(net_563) );
INV_X2 inst_510 ( .A(net_520), .ZN(net_518) );
NAND2_X2 inst_268 ( .ZN(net_237), .A2(net_193), .A1(net_180) );
INV_X4 inst_369 ( .ZN(net_501), .A(net_499) );
DFFR_X2 inst_550 ( .RN(net_464), .D(net_274), .QN(net_2), .CK(net_617) );
NOR2_X2 inst_63 ( .ZN(net_565), .A1(net_123), .A2(net_56) );
NAND4_X2 inst_119 ( .A4(net_554), .ZN(net_476), .A3(net_217), .A1(net_125), .A2(net_25) );
CLKBUF_X2 inst_603 ( .A(net_588), .Z(net_589) );
NAND2_X2 inst_327 ( .A2(net_492), .ZN(net_443), .A1(net_376) );
NOR2_X2 inst_85 ( .ZN(net_224), .A1(net_223), .A2(net_156) );
NAND2_X2 inst_291 ( .ZN(net_325), .A2(net_304), .A1(net_240) );
NAND2_X2 inst_266 ( .ZN(net_226), .A2(net_187), .A1(net_121) );
INV_X4 inst_473 ( .ZN(net_255), .A(net_145) );
NAND2_X4 inst_217 ( .A2(net_530), .ZN(net_454), .A1(net_442) );
AND2_X4 inst_572 ( .A1(net_507), .ZN(net_354), .A2(net_1) );
NOR2_X2 inst_77 ( .A2(net_554), .ZN(net_174), .A1(net_173) );
NAND3_X2 inst_171 ( .A1(net_411), .ZN(net_410), .A3(net_262), .A2(net_195) );
DFFR_X1 inst_558 ( .Q(net_469), .RN(net_464), .D(net_372), .CK(net_590) );
INV_X4 inst_427 ( .ZN(net_76), .A(net_50) );
NAND2_X2 inst_257 ( .ZN(net_306), .A2(net_101), .A1(net_98) );
CLKBUF_X2 inst_594 ( .A(net_579), .Z(net_580) );
NAND3_X2 inst_145 ( .A2(net_505), .A3(net_493), .ZN(net_266), .A1(net_219) );
NAND2_X2 inst_290 ( .A1(net_504), .ZN(net_324), .A2(net_282) );
INV_X4 inst_374 ( .ZN(net_17), .A(G9) );
NAND2_X2 inst_272 ( .A2(net_535), .ZN(net_277), .A1(net_126) );
INV_X2 inst_502 ( .ZN(net_559), .A(G3) );
NOR2_X2 inst_103 ( .ZN(net_343), .A2(net_313), .A1(net_233) );
INV_X4 inst_485 ( .ZN(net_416), .A(net_223) );
AND4_X2 inst_565 ( .ZN(net_352), .A2(net_316), .A4(net_265), .A1(net_147), .A3(net_144) );
NAND2_X2 inst_248 ( .A2(net_166), .A1(net_152), .ZN(net_143) );
CLKBUF_X2 inst_622 ( .A(net_582), .Z(net_608) );
NAND3_X2 inst_138 ( .ZN(net_285), .A3(net_216), .A1(net_215), .A2(net_47) );
INV_X4 inst_389 ( .ZN(net_477), .A(net_17) );
INV_X4 inst_357 ( .ZN(net_552), .A(net_463) );
INV_X4 inst_409 ( .A(net_167), .ZN(net_101) );
NAND3_X2 inst_180 ( .A3(net_439), .A1(net_412), .A2(net_385), .ZN(G552) );
NOR3_X2 inst_33 ( .A3(net_335), .ZN(net_322), .A1(net_293), .A2(net_263) );
NAND2_X2 inst_312 ( .ZN(net_398), .A1(net_338), .A2(net_4) );
CLKBUF_X2 inst_609 ( .A(net_594), .Z(net_595) );
INV_X2 inst_517 ( .A(net_506), .ZN(net_505) );
NAND2_X2 inst_309 ( .ZN(net_394), .A1(net_393), .A2(net_358) );
NAND2_X2 inst_232 ( .ZN(net_108), .A1(net_75), .A2(net_43) );
MUX2_X2 inst_347 ( .Z(net_347), .B(net_335), .S(net_320), .A(net_300) );
NAND2_X2 inst_301 ( .ZN(net_366), .A2(net_353), .A1(net_170) );
INV_X4 inst_363 ( .A(net_514), .ZN(net_513) );
NOR3_X2 inst_27 ( .A2(net_512), .A1(net_505), .ZN(net_232), .A3(net_231) );
NAND2_X2 inst_247 ( .A1(net_499), .A2(net_334), .ZN(net_127) );
NAND2_X2 inst_297 ( .ZN(net_485), .A2(net_346), .A1(net_73) );
INV_X4 inst_403 ( .ZN(net_32), .A(G7) );
NAND2_X2 inst_302 ( .ZN(net_369), .A1(net_368), .A2(net_0) );
NAND2_X2 inst_310 ( .ZN(net_395), .A1(net_393), .A2(net_365) );
NAND2_X2 inst_322 ( .A1(net_538), .ZN(net_435), .A2(net_424) );
NAND2_X2 inst_253 ( .ZN(net_181), .A1(net_180), .A2(net_114) );
NAND2_X4 inst_211 ( .ZN(net_383), .A2(net_374), .A1(net_360) );
CLKBUF_X2 inst_619 ( .A(net_604), .Z(net_605) );
NAND3_X2 inst_162 ( .A2(net_420), .A1(net_387), .ZN(net_385), .A3(net_327) );
CLKBUF_X2 inst_589 ( .A(net_574), .Z(net_575) );
DFFR_X1 inst_561 ( .RN(net_464), .D(net_458), .Q(G45), .CK(net_580) );
INV_X4 inst_412 ( .A(net_210), .ZN(net_30) );
INV_X4 inst_449 ( .ZN(net_166), .A(net_107) );
CLKBUF_X2 inst_639 ( .A(net_614), .Z(net_625) );
NAND3_X2 inst_155 ( .A2(net_562), .A3(net_548), .A1(net_547), .ZN(net_546) );
INV_X4 inst_464 ( .ZN(net_134), .A(net_123) );
CLKBUF_X2 inst_602 ( .A(net_587), .Z(net_588) );
NOR2_X2 inst_59 ( .A1(net_148), .ZN(net_135), .A2(net_117) );
NAND3_X2 inst_135 ( .ZN(net_482), .A2(net_167), .A3(net_166), .A1(net_36) );
NAND2_X2 inst_341 ( .ZN(net_467), .A2(net_465), .A1(net_449) );
NAND2_X4 inst_196 ( .ZN(net_112), .A1(net_34), .A2(G7) );
INV_X2 inst_532 ( .A(net_272), .ZN(net_121) );
NOR2_X2 inst_55 ( .A2(net_561), .ZN(net_540), .A1(net_72) );
NOR3_X2 inst_37 ( .ZN(net_372), .A2(net_355), .A3(net_336), .A1(net_331) );
INV_X4 inst_498 ( .ZN(net_419), .A(net_418) );
NAND2_X2 inst_264 ( .ZN(net_281), .A2(net_222), .A1(net_148) );
NOR2_X2 inst_84 ( .ZN(net_202), .A2(net_163), .A1(net_139) );
NAND3_X2 inst_173 ( .A1(net_449), .ZN(net_421), .A2(net_420), .A3(net_407) );
NAND2_X2 inst_298 ( .A1(net_449), .ZN(net_353), .A2(net_341) );
NAND2_X2 inst_303 ( .ZN(net_376), .A2(net_369), .A1(net_298) );
CLKBUF_X2 inst_611 ( .A(net_596), .Z(net_597) );
NAND2_X2 inst_224 ( .ZN(net_529), .A2(net_41), .A1(net_32) );
NOR2_X4 inst_42 ( .ZN(net_125), .A1(net_103), .A2(net_83) );
NAND2_X2 inst_287 ( .ZN(net_490), .A1(net_312), .A2(net_294) );
NAND2_X2 inst_323 ( .A2(net_492), .ZN(net_439), .A1(net_9) );
CLKBUF_X2 inst_618 ( .A(net_579), .Z(net_604) );
INV_X4 inst_426 ( .A(net_75), .ZN(net_74) );
CLKBUF_X2 inst_588 ( .A(net_573), .Z(net_574) );
INV_X8 inst_350 ( .ZN(net_42), .A(net_20) );
NAND2_X2 inst_231 ( .A1(net_92), .A2(net_91), .ZN(net_73) );
NAND2_X2 inst_270 ( .ZN(net_252), .A2(net_183), .A1(net_117) );
INV_X4 inst_474 ( .ZN(net_302), .A(net_146) );
NOR3_X2 inst_26 ( .ZN(net_156), .A2(net_137), .A1(net_109), .A3(net_78) );
INV_X4 inst_437 ( .A(net_64), .ZN(net_53) );
INV_X4 inst_490 ( .ZN(net_221), .A(net_220) );
CLKBUF_X2 inst_626 ( .A(net_611), .Z(net_612) );
NOR2_X2 inst_70 ( .A1(net_569), .ZN(net_151), .A2(net_150) );
NAND3_X4 inst_129 ( .ZN(net_374), .A3(net_350), .A2(net_108), .A1(net_84) );
NAND3_X2 inst_189 ( .A2(net_556), .ZN(net_468), .A1(net_427), .A3(net_3) );
OR2_X2 inst_11 ( .A2(net_168), .ZN(net_147), .A1(net_100) );
CLKBUF_X2 inst_631 ( .A(net_616), .Z(net_617) );
NAND3_X2 inst_188 ( .A2(net_461), .A3(net_457), .A1(net_434), .ZN(G535) );
OR2_X2 inst_14 ( .ZN(net_236), .A1(net_235), .A2(net_165) );
INV_X4 inst_475 ( .ZN(net_155), .A(net_154) );
INV_X4 inst_441 ( .ZN(net_94), .A(net_59) );
NOR3_X2 inst_31 ( .ZN(net_305), .A2(net_205), .A3(net_189), .A1(net_179) );
INV_X2 inst_528 ( .ZN(net_128), .A(net_81) );
NAND2_X2 inst_252 ( .ZN(net_177), .A2(net_118), .A1(net_30) );
NOR2_X2 inst_62 ( .ZN(net_113), .A1(net_112), .A2(net_68) );
DFFR_X1 inst_557 ( .RN(net_464), .D(net_370), .QN(net_10), .CK(net_572) );
NAND2_X2 inst_251 ( .A1(net_210), .ZN(net_199), .A2(net_111) );
INV_X4 inst_352 ( .ZN(net_562), .A(G3) );
AND2_X4 inst_575 ( .A1(net_537), .ZN(net_517), .A2(net_427) );
INV_X4 inst_398 ( .ZN(net_320), .A(net_22) );
NAND2_X2 inst_286 ( .ZN(net_473), .A2(net_289), .A1(net_122) );
INV_X4 inst_436 ( .A(net_75), .ZN(net_52) );
INV_X4 inst_484 ( .A(net_344), .ZN(net_218) );
CLKBUF_X2 inst_627 ( .A(net_600), .Z(net_613) );
NAND2_X2 inst_300 ( .A2(net_546), .A1(net_545), .ZN(net_363) );
NOR2_X2 inst_102 ( .ZN(net_474), .A1(net_1), .A2(G6) );
NOR3_X2 inst_32 ( .ZN(net_321), .A2(net_320), .A1(net_284), .A3(net_71) );
NAND2_X1 inst_344 ( .ZN(net_431), .A2(net_430), .A1(net_315) );
INV_X4 inst_428 ( .A(net_120), .ZN(net_59) );
INV_X4 inst_446 ( .ZN(net_204), .A(net_64) );
INV_X4 inst_364 ( .A(net_514), .ZN(net_512) );
NAND3_X2 inst_144 ( .A2(net_519), .ZN(net_265), .A3(net_196), .A1(net_127) );
CLKBUF_X2 inst_629 ( .A(net_614), .Z(net_615) );
NAND2_X4 inst_195 ( .ZN(net_54), .A1(net_24), .A2(G4) );
INV_X4 inst_407 ( .A(net_320), .ZN(net_39) );
CLKBUF_X2 inst_623 ( .A(net_608), .Z(net_609) );
INV_X4 inst_411 ( .A(net_216), .ZN(net_38) );
NOR2_X2 inst_97 ( .ZN(net_303), .A1(net_302), .A2(net_249) );
CLKBUF_X2 inst_616 ( .A(net_601), .Z(net_602) );
NAND4_X2 inst_124 ( .ZN(net_543), .A2(net_539), .A1(net_522), .A4(net_167), .A3(net_152) );
INV_X2 inst_533 ( .ZN(net_132), .A(net_131) );
CLKBUF_X2 inst_620 ( .A(net_605), .Z(net_606) );
NAND3_X2 inst_137 ( .A1(net_507), .ZN(net_491), .A3(net_260), .A2(net_50) );
INV_X4 inst_425 ( .A(net_312), .ZN(net_79) );
INV_X1 inst_545 ( .ZN(net_433), .A(net_432) );
NAND3_X4 inst_130 ( .ZN(net_550), .A3(net_482), .A1(net_481), .A2(net_356) );
NAND2_X2 inst_227 ( .A2(net_216), .ZN(net_85), .A1(net_83) );
INV_X4 inst_399 ( .ZN(net_167), .A(net_92) );
INV_X2 inst_527 ( .A(net_133), .ZN(net_61) );
NAND2_X2 inst_226 ( .A2(net_560), .ZN(net_81), .A1(net_50) );
NAND3_X2 inst_176 ( .A1(net_492), .ZN(net_446), .A3(net_260), .A2(net_259) );
NOR2_X2 inst_58 ( .A1(net_169), .ZN(net_105), .A2(net_70) );
INV_X4 inst_414 ( .ZN(net_120), .A(net_72) );
NOR2_X2 inst_87 ( .ZN(net_228), .A1(net_227), .A2(net_55) );
NOR2_X2 inst_61 ( .ZN(net_569), .A2(net_526), .A1(net_23) );
DFFR_X1 inst_562 ( .RN(net_464), .D(net_459), .QN(net_3), .CK(net_577) );
INV_X2 inst_531 ( .ZN(net_489), .A(net_108) );
NAND2_X4 inst_203 ( .ZN(net_487), .A1(net_90), .A2(net_50) );
NAND2_X4 inst_212 ( .A2(net_484), .A1(net_483), .ZN(net_405) );
INV_X2 inst_499 ( .ZN(net_564), .A(net_562) );
NAND2_X2 inst_335 ( .A1(net_567), .A2(net_456), .ZN(net_455) );
INV_X4 inst_466 ( .A(net_384), .ZN(net_260) );
OR2_X4 inst_10 ( .ZN(net_326), .A1(net_296), .A2(net_273) );
OR3_X2 inst_4 ( .ZN(net_308), .A1(net_256), .A3(net_224), .A2(net_66) );
INV_X4 inst_456 ( .A(net_96), .ZN(net_87) );
AND2_X2 inst_581 ( .A1(net_334), .ZN(net_284), .A2(net_283) );
CLKBUF_X2 inst_600 ( .A(net_585), .Z(net_586) );
NOR3_X2 inst_28 ( .A2(net_499), .ZN(net_233), .A1(net_227), .A3(net_43) );
NAND2_X2 inst_275 ( .A1(net_501), .ZN(net_280), .A2(net_250) );
NOR2_X1 inst_117 ( .ZN(net_197), .A1(net_98), .A2(net_31) );
INV_X4 inst_438 ( .ZN(net_368), .A(net_57) );
INV_X2 inst_501 ( .ZN(net_566), .A(net_562) );
NOR2_X2 inst_49 ( .ZN(net_152), .A1(net_28), .A2(G11) );
NAND2_X4 inst_204 ( .ZN(net_254), .A1(net_88), .A2(net_67) );
CLKBUF_X2 inst_587 ( .A(net_570), .Z(net_573) );
NAND3_X2 inst_154 ( .A3(net_491), .A1(net_490), .ZN(net_360), .A2(net_267) );
CLKBUF_X2 inst_592 ( .A(net_572), .Z(net_578) );
DFFR_X2 inst_546 ( .RN(net_464), .D(net_113), .Q(net_7), .CK(net_626) );
NAND2_X2 inst_324 ( .A2(net_492), .ZN(net_440), .A1(net_325) );
INV_X4 inst_465 ( .ZN(net_124), .A(net_103) );
NOR2_X2 inst_109 ( .ZN(net_370), .A2(net_357), .A1(net_232) );
NOR2_X2 inst_54 ( .A1(net_334), .ZN(net_71), .A2(net_70) );
AND2_X4 inst_570 ( .ZN(net_337), .A2(net_91), .A1(net_35) );
INV_X4 inst_390 ( .A(net_83), .ZN(net_29) );
CLKBUF_X2 inst_640 ( .A(net_625), .Z(net_626) );
NOR2_X4 inst_43 ( .ZN(net_244), .A2(net_210), .A1(net_209) );
INV_X4 inst_359 ( .A(net_531), .ZN(net_530) );
NAND2_X2 inst_256 ( .A1(net_558), .ZN(net_292), .A2(net_192) );
NOR2_X2 inst_94 ( .A2(net_523), .ZN(net_338), .A1(net_228) );
INV_X4 inst_454 ( .ZN(net_123), .A(net_80) );
CLKBUF_X2 inst_630 ( .A(net_615), .Z(net_616) );
INV_X4 inst_375 ( .ZN(net_456), .A(G12) );
INV_X4 inst_401 ( .ZN(net_216), .A(net_24) );
NAND2_X2 inst_262 ( .A1(net_247), .ZN(net_208), .A2(net_7) );
INV_X2 inst_512 ( .A(net_515), .ZN(net_514) );
INV_X4 inst_355 ( .A(net_557), .ZN(net_556) );
NAND2_X2 inst_243 ( .A1(net_558), .A2(net_270), .ZN(net_122) );
NAND2_X2 inst_285 ( .A1(net_503), .ZN(net_304), .A2(net_253) );
CLKBUF_X2 inst_591 ( .A(net_576), .Z(net_577) );
INV_X4 inst_424 ( .ZN(net_206), .A(net_40) );
INV_X4 inst_497 ( .ZN(net_425), .A(net_415) );
NAND2_X4 inst_218 ( .ZN(net_532), .A2(net_489), .A1(net_488) );
OR2_X2 inst_15 ( .ZN(net_248), .A1(net_247), .A2(net_175) );
NAND2_X1 inst_343 ( .A1(net_564), .ZN(net_69), .A2(net_48) );
OR3_X2 inst_6 ( .ZN(net_328), .A2(net_297), .A3(net_269), .A1(net_261) );
NAND2_X4 inst_194 ( .ZN(net_555), .A2(net_21), .A1(G3) );
INV_X2 inst_543 ( .A(net_436), .ZN(net_426) );
NAND2_X2 inst_337 ( .ZN(net_462), .A2(net_460), .A1(net_279) );
NAND4_X2 inst_123 ( .A3(net_566), .A1(net_565), .ZN(net_364), .A2(net_120), .A4(net_5) );
INV_X2 inst_509 ( .A(net_520), .ZN(net_519) );
NAND2_X2 inst_299 ( .ZN(net_356), .A2(net_354), .A1(net_26) );
INV_X4 inst_418 ( .A(net_48), .ZN(net_47) );
INV_X4 inst_476 ( .ZN(net_344), .A(net_98) );
NAND4_X2 inst_118 ( .ZN(net_214), .A2(net_213), .A1(net_212), .A3(net_65), .A4(net_62) );
NOR2_X2 inst_86 ( .ZN(net_287), .A1(net_227), .A2(net_98) );
NAND3_X2 inst_153 ( .A1(net_527), .ZN(net_346), .A3(net_92), .A2(net_41) );
OR2_X2 inst_20 ( .A2(net_436), .ZN(net_434), .A1(net_359) );
INV_X4 inst_442 ( .ZN(net_180), .A(net_60) );
CLKBUF_X2 inst_613 ( .A(net_598), .Z(net_599) );
NOR2_X4 inst_38 ( .ZN(net_91), .A1(net_34), .A2(net_20) );
INV_X4 inst_381 ( .ZN(net_92), .A(net_17) );
NAND2_X2 inst_295 ( .A1(net_473), .ZN(net_414), .A2(net_334) );
INV_X8 inst_349 ( .A(net_499), .ZN(net_498) );
INV_X4 inst_483 ( .ZN(net_263), .A(net_255) );
AND2_X4 inst_576 ( .ZN(net_401), .A2(net_400), .A1(net_317) );
NAND2_X4 inst_209 ( .A2(net_471), .A1(net_470), .ZN(net_365) );
NAND2_X2 inst_259 ( .A2(net_384), .A1(net_255), .ZN(net_193) );
NOR2_X4 inst_40 ( .ZN(net_493), .A2(net_477), .A1(net_112) );
NAND2_X2 inst_320 ( .A1(net_456), .ZN(net_436), .A2(net_425) );
NAND3_X2 inst_167 ( .ZN(net_403), .A2(net_323), .A1(net_239), .A3(net_4) );
CLKBUF_X2 inst_607 ( .A(net_592), .Z(net_593) );
NAND2_X2 inst_246 ( .A2(net_528), .ZN(net_126), .A1(net_43) );
CLKBUF_X2 inst_635 ( .A(net_620), .Z(net_621) );
NOR2_X2 inst_95 ( .ZN(net_295), .A1(net_287), .A2(net_130) );
XNOR2_X2 inst_1 ( .B(net_524), .ZN(net_323), .A(net_251) );
NOR2_X2 inst_72 ( .A2(net_529), .ZN(net_163), .A1(net_43) );
INV_X2 inst_519 ( .A(net_501), .ZN(net_500) );
INV_X4 inst_439 ( .ZN(net_203), .A(net_55) );
NAND2_X2 inst_331 ( .ZN(net_448), .A2(net_433), .A1(net_339) );
AND2_X2 inst_582 ( .ZN(net_293), .A1(net_292), .A2(net_281) );
NOR2_X2 inst_115 ( .ZN(net_459), .A2(net_453), .A1(net_401) );
NAND2_X2 inst_235 ( .ZN(net_89), .A1(net_81), .A2(net_54) );
NAND2_X4 inst_210 ( .ZN(net_538), .A1(net_365), .A2(G13) );
NAND2_X2 inst_317 ( .ZN(net_418), .A1(net_414), .A2(net_413) );
NAND2_X2 inst_278 ( .ZN(net_290), .A2(net_226), .A1(net_97) );
INV_X4 inst_467 ( .ZN(net_388), .A(net_335) );
NAND2_X2 inst_239 ( .ZN(net_111), .A2(net_80), .A1(G6) );
NOR2_X2 inst_105 ( .A1(net_558), .ZN(net_351), .A2(net_12) );
INV_X4 inst_488 ( .ZN(net_449), .A(net_263) );
INV_X4 inst_387 ( .A(net_34), .ZN(net_16) );
CLKBUF_X2 inst_593 ( .A(net_578), .Z(net_579) );
NAND3_X2 inst_175 ( .A1(net_430), .ZN(net_428), .A2(net_218), .A3(net_181) );
NAND2_X2 inst_254 ( .A2(net_212), .ZN(net_183), .A1(net_182) );
CLKBUF_X2 inst_625 ( .A(net_610), .Z(net_611) );
NAND2_X2 inst_225 ( .ZN(net_68), .A1(net_44), .A2(net_37) );
CLKBUF_X2 inst_601 ( .A(net_586), .Z(net_587) );
NAND3_X2 inst_133 ( .ZN(net_188), .A3(net_182), .A2(net_46), .A1(net_40) );
INV_X2 inst_508 ( .A(net_526), .ZN(net_524) );
AND2_X4 inst_568 ( .ZN(net_21), .A2(G6), .A1(G4) );
NOR2_X2 inst_112 ( .ZN(net_396), .A2(net_383), .A1(net_95) );
INV_X2 inst_523 ( .ZN(net_44), .A(G0) );
INV_X4 inst_365 ( .A(net_512), .ZN(net_511) );
NOR2_X2 inst_67 ( .A2(net_509), .A1(net_203), .ZN(net_139) );
NAND3_X2 inst_181 ( .A3(net_444), .A1(net_422), .A2(net_394), .ZN(G539) );
NAND2_X2 inst_305 ( .A2(net_542), .A1(net_541), .ZN(net_483) );
INV_X4 inst_479 ( .ZN(net_227), .A(net_160) );
NOR3_X2 inst_29 ( .A1(net_558), .ZN(net_256), .A3(net_255), .A2(net_104) );
INV_X4 inst_391 ( .ZN(net_119), .A(net_56) );
CLKBUF_X2 inst_590 ( .A(net_575), .Z(net_576) );
NAND2_X4 inst_202 ( .A1(net_515), .A2(net_217), .ZN(net_178) );
NAND4_X2 inst_126 ( .A2(net_468), .A1(net_446), .A3(net_409), .A4(net_402), .ZN(G549) );
INV_X4 inst_480 ( .A(net_173), .ZN(net_161) );
CLKBUF_X2 inst_634 ( .A(net_616), .Z(net_620) );
INV_X4 inst_419 ( .A(net_101), .ZN(net_55) );
INV_X4 inst_477 ( .ZN(net_223), .A(net_192) );
AND4_X4 inst_564 ( .ZN(net_492), .A3(net_427), .A1(net_414), .A4(net_413), .A2(G12) );
INV_X2 inst_538 ( .ZN(net_251), .A(net_250) );
INV_X4 inst_423 ( .A(net_115), .ZN(net_62) );
NOR3_X2 inst_35 ( .A3(net_527), .A2(net_505), .ZN(net_345), .A1(net_344) );
INV_X4 inst_382 ( .ZN(net_83), .A(net_19) );
NOR2_X2 inst_48 ( .ZN(net_43), .A1(net_17), .A2(net_16) );
INV_X4 inst_358 ( .A(net_535), .ZN(net_534) );
NOR2_X2 inst_46 ( .A1(net_427), .ZN(net_420), .A2(G12) );
NAND3_X2 inst_136 ( .A1(net_368), .A3(net_275), .ZN(net_184), .A2(net_128) );
NOR3_X2 inst_30 ( .A2(net_558), .ZN(net_269), .A3(net_198), .A1(net_142) );
NAND2_X2 inst_330 ( .A2(net_492), .ZN(net_447), .A1(net_10) );
CLKBUF_X2 inst_610 ( .A(net_584), .Z(net_596) );
NAND2_X2 inst_233 ( .ZN(net_384), .A1(net_83), .A2(net_49) );
NAND3_X2 inst_165 ( .ZN(net_389), .A1(net_388), .A3(net_387), .A2(net_162) );
NAND2_X2 inst_271 ( .A2(net_524), .ZN(net_258), .A1(net_220) );
INV_X4 inst_443 ( .ZN(net_98), .A(net_62) );
CLKBUF_X2 inst_633 ( .A(net_618), .Z(net_619) );
NOR3_X2 inst_34 ( .ZN(net_342), .A1(net_150), .A2(net_112), .A3(net_6) );
OR2_X2 inst_12 ( .A2(net_168), .ZN(net_149), .A1(net_148) );
INV_X2 inst_529 ( .ZN(net_97), .A(net_96) );
INV_X2 inst_524 ( .ZN(net_27), .A(G5) );
NOR2_X2 inst_56 ( .ZN(net_78), .A1(net_50), .A2(net_38) );
NOR2_X2 inst_71 ( .A1(net_320), .ZN(net_158), .A2(net_134) );
NAND2_X2 inst_308 ( .ZN(net_392), .A2(net_390), .A1(net_146) );
NOR2_X2 inst_104 ( .ZN(net_348), .A2(net_322), .A1(net_105) );
INV_X4 inst_448 ( .ZN(net_99), .A(net_76) );
NOR2_X2 inst_60 ( .A2(net_518), .ZN(net_109), .A1(net_76) );
INV_X4 inst_455 ( .A(net_231), .ZN(net_82) );
NAND3_X2 inst_168 ( .A2(net_510), .ZN(net_404), .A1(net_306), .A3(net_4) );
INV_X4 inst_384 ( .ZN(net_56), .A(net_27) );
NAND2_X2 inst_321 ( .ZN(net_549), .A2(net_419), .A1(G12) );
INV_X4 inst_496 ( .ZN(net_387), .A(net_383) );
CLKBUF_X2 inst_608 ( .A(net_593), .Z(net_594) );
NAND2_X2 inst_336 ( .A1(net_450), .A2(net_437), .ZN(G530) );
DFFR_X1 inst_563 ( .D(net_552), .RN(net_464), .QN(G546), .CK(net_595) );
AND2_X2 inst_583 ( .A1(net_420), .ZN(net_361), .A2(net_360) );
AND2_X2 inst_580 ( .ZN(net_201), .A1(net_200), .A2(net_199) );
NAND3_X2 inst_170 ( .A1(net_411), .ZN(net_409), .A2(net_292), .A3(net_161) );
NAND2_X2 inst_258 ( .A2(net_558), .ZN(net_259), .A1(net_39) );
INV_X4 inst_376 ( .ZN(net_34), .A(G10) );
NAND2_X4 inst_199 ( .A2(net_478), .ZN(net_107), .A1(net_42) );
NOR2_X4 inst_41 ( .ZN(net_131), .A1(net_107), .A2(G11) );
INV_X2 inst_511 ( .A(net_516), .ZN(net_515) );
NAND3_X2 inst_143 ( .A2(net_337), .ZN(net_257), .A1(net_254), .A3(net_124) );
NAND3_X2 inst_152 ( .ZN(net_470), .A1(net_309), .A3(net_210), .A2(net_50) );
NAND2_X2 inst_265 ( .ZN(net_225), .A2(net_188), .A1(net_153) );
INV_X4 inst_482 ( .ZN(net_222), .A(net_192) );
INV_X4 inst_468 ( .A(net_204), .ZN(net_146) );
INV_X1 inst_544 ( .ZN(net_464), .A(blif_reset_net) );
NAND2_X2 inst_238 ( .A2(net_519), .ZN(net_110), .A1(net_51) );
INV_X2 inst_540 ( .ZN(net_315), .A(net_314) );
INV_X2 inst_539 ( .ZN(net_311), .A(net_6) );
INV_X4 inst_429 ( .ZN(net_217), .A(net_45) );
INV_X4 inst_404 ( .ZN(net_72), .A(G11) );
NAND3_X2 inst_178 ( .A3(net_492), .ZN(net_451), .A2(net_328), .A1(net_302) );
NOR2_X2 inst_89 ( .ZN(net_246), .A2(net_172), .A1(net_64) );
NOR2_X2 inst_111 ( .ZN(net_382), .A1(net_381), .A2(net_373) );
NOR2_X2 inst_66 ( .A1(net_558), .ZN(net_164), .A2(net_133) );
INV_X4 inst_388 ( .A(net_34), .ZN(net_28) );
OR3_X2 inst_7 ( .A3(net_538), .ZN(net_380), .A2(net_334), .A1(net_185) );
NAND3_X2 inst_182 ( .A2(net_503), .ZN(net_457), .A1(net_456), .A3(net_441) );
INV_X4 inst_392 ( .A(net_28), .ZN(net_18) );
NAND4_X2 inst_120 ( .ZN(net_271), .A4(net_270), .A3(net_247), .A1(net_235), .A2(net_138) );
NAND2_X2 inst_273 ( .A1(net_554), .ZN(net_278), .A2(net_244) );
NAND2_X2 inst_294 ( .ZN(net_330), .A2(net_301), .A1(net_266) );
NAND2_X2 inst_222 ( .ZN(net_516), .A1(net_28), .A2(G7) );
NAND2_X2 inst_284 ( .A2(net_533), .ZN(net_314), .A1(net_223) );
INV_X4 inst_489 ( .ZN(net_250), .A(net_220) );
NAND3_X1 inst_192 ( .A2(net_502), .ZN(net_438), .A3(net_430), .A1(net_329) );
NAND2_X2 inst_280 ( .A1(net_556), .ZN(net_298), .A2(net_297) );
INV_X4 inst_366 ( .A(net_516), .ZN(net_508) );
MUX2_X2 inst_346 ( .S(net_529), .Z(net_176), .A(net_102), .B(net_43) );
INV_X4 inst_491 ( .ZN(net_283), .A(net_190) );
AND3_X4 inst_567 ( .ZN(net_442), .A3(net_427), .A1(net_418), .A2(G12) );
NAND2_X4 inst_193 ( .ZN(net_334), .A1(net_27), .A2(G4) );
NAND3_X2 inst_149 ( .ZN(net_471), .A3(net_211), .A1(net_86), .A2(net_50) );
NAND2_X2 inst_318 ( .ZN(net_423), .A1(net_420), .A2(net_408) );
NOR2_X4 inst_39 ( .ZN(net_182), .A1(net_48), .A2(net_27) );
NAND2_X2 inst_230 ( .ZN(net_150), .A1(net_33), .A2(G11) );

endmodule
