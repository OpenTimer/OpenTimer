module c880 (
n201gat,
n189gat,
n17gat,
n72gat,
n152gat,
n255gat,
n159gat,
n85gat,
n267gat,
n87gat,
n116gat,
n74gat,
n55gat,
n90gat,
n210gat,
n96gat,
n228gat,
n260gat,
n143gat,
n80gat,
n207gat,
n153gat,
n268gat,
n171gat,
n1gat,
n135gat,
n111gat,
n237gat,
n183gat,
n130gat,
n29gat,
n261gat,
n101gat,
n59gat,
n138gat,
n149gat,
n195gat,
n86gat,
n177gat,
n219gat,
n42gat,
n121gat,
n146gat,
n91gat,
n26gat,
n156gat,
n68gat,
n13gat,
n246gat,
n8gat,
n75gat,
n73gat,
n36gat,
n88gat,
n126gat,
n106gat,
n165gat,
n259gat,
n89gat,
n51gat,
n420gat,
n389gat,
n879gat,
n865gat,
n850gat,
n446gat,
n767gat,
n390gat,
n874gat,
n864gat,
n768gat,
n421gat,
n863gat,
n419gat,
n388gat,
n449gat,
n450gat,
n880gat,
n423gat,
n866gat,
n447gat,
n391gat,
n448gat,
n878gat,
n418gat,
n422gat);

// Start PIs
input n201gat;
input n189gat;
input n17gat;
input n72gat;
input n152gat;
input n255gat;
input n159gat;
input n85gat;
input n267gat;
input n87gat;
input n116gat;
input n74gat;
input n55gat;
input n90gat;
input n210gat;
input n96gat;
input n228gat;
input n260gat;
input n143gat;
input n80gat;
input n207gat;
input n153gat;
input n268gat;
input n171gat;
input n1gat;
input n135gat;
input n111gat;
input n237gat;
input n183gat;
input n130gat;
input n29gat;
input n261gat;
input n101gat;
input n59gat;
input n138gat;
input n149gat;
input n195gat;
input n86gat;
input n177gat;
input n219gat;
input n42gat;
input n121gat;
input n146gat;
input n91gat;
input n26gat;
input n156gat;
input n68gat;
input n13gat;
input n246gat;
input n8gat;
input n75gat;
input n73gat;
input n36gat;
input n88gat;
input n126gat;
input n106gat;
input n165gat;
input n259gat;
input n89gat;
input n51gat;

// Start POs
output n420gat;
output n389gat;
output n879gat;
output n865gat;
output n850gat;
output n446gat;
output n767gat;
output n390gat;
output n874gat;
output n864gat;
output n768gat;
output n421gat;
output n863gat;
output n419gat;
output n388gat;
output n449gat;
output n450gat;
output n880gat;
output n423gat;
output n866gat;
output n447gat;
output n391gat;
output n448gat;
output n878gat;
output n418gat;
output n422gat;

// Start wires
wire net_47;
wire net_176;
wire net_137;
wire n159gat;
wire net_132;
wire net_54;
wire n768gat;
wire net_105;
wire n419gat;
wire net_129;
wire net_119;
wire net_98;
wire net_12;
wire net_151;
wire net_53;
wire net_93;
wire net_168;
wire net_127;
wire net_76;
wire net_101;
wire net_187;
wire net_111;
wire net_90;
wire n26gat;
wire net_100;
wire net_85;
wire net_124;
wire net_160;
wire net_115;
wire n878gat;
wire net_4;
wire net_17;
wire n51gat;
wire n865gat;
wire n17gat;
wire net_164;
wire net_87;
wire net_0;
wire net_35;
wire n87gat;
wire net_16;
wire n74gat;
wire net_193;
wire net_157;
wire n260gat;
wire net_42;
wire net_120;
wire net_109;
wire net_80;
wire net_65;
wire net_50;
wire n183gat;
wire n130gat;
wire net_96;
wire net_66;
wire net_38;
wire n446gat;
wire net_167;
wire net_136;
wire net_19;
wire n177gat;
wire net_126;
wire n91gat;
wire net_34;
wire net_108;
wire net_183;
wire n88gat;
wire net_150;
wire net_63;
wire n879gat;
wire n255gat;
wire net_30;
wire net_189;
wire net_99;
wire net_24;
wire net_186;
wire net_46;
wire net_118;
wire n55gat;
wire net_146;
wire n96gat;
wire net_122;
wire n143gat;
wire net_7;
wire n111gat;
wire net_172;
wire net_52;
wire net_165;
wire net_13;
wire net_94;
wire net_18;
wire net_131;
wire net_114;
wire n126gat;
wire n866gat;
wire net_29;
wire net_149;
wire net_142;
wire net_31;
wire net_36;
wire net_158;
wire n189gat;
wire net_41;
wire net_3;
wire net_154;
wire n388gat;
wire net_28;
wire n153gat;
wire n391gat;
wire n448gat;
wire net_97;
wire net_182;
wire net_192;
wire net_60;
wire n101gat;
wire n59gat;
wire n149gat;
wire net_58;
wire n863gat;
wire net_82;
wire net_64;
wire net_121;
wire net_73;
wire net_177;
wire net_86;
wire net_75;
wire n447gat;
wire n106gat;
wire net_125;
wire net_107;
wire net_166;
wire net_179;
wire n152gat;
wire net_159;
wire n767gat;
wire net_61;
wire net_62;
wire n116gat;
wire net_6;
wire net_23;
wire n90gat;
wire net_117;
wire net_74;
wire n80gat;
wire net_135;
wire net_130;
wire n420gat;
wire net_147;
wire n261gat;
wire net_14;
wire net_26;
wire net_113;
wire n195gat;
wire net_32;
wire n219gat;
wire net_40;
wire n246gat;
wire n13gat;
wire n8gat;
wire net_69;
wire net_161;
wire net_141;
wire net_83;
wire net_95;
wire net_173;
wire n389gat;
wire n850gat;
wire net_78;
wire net_27;
wire n72gat;
wire net_56;
wire n874gat;
wire net_155;
wire net_191;
wire net_22;
wire net_181;
wire net_39;
wire n228gat;
wire net_2;
wire net_102;
wire net_144;
wire net_9;
wire net_59;
wire n207gat;
wire n268gat;
wire net_162;
wire net_44;
wire net_134;
wire n421gat;
wire net_45;
wire net_89;
wire n146gat;
wire n156gat;
wire net_185;
wire n75gat;
wire n450gat;
wire net_178;
wire n165gat;
wire n418gat;
wire n89gat;
wire net_152;
wire net_116;
wire n390gat;
wire net_175;
wire net_91;
wire net_55;
wire net_106;
wire net_140;
wire n449gat;
wire n210gat;
wire net_104;
wire net_148;
wire n880gat;
wire net_72;
wire net_25;
wire net_70;
wire n171gat;
wire net_194;
wire net_5;
wire net_128;
wire net_138;
wire net_184;
wire net_11;
wire n68gat;
wire n73gat;
wire n36gat;
wire net_123;
wire net_170;
wire net_68;
wire net_77;
wire net_20;
wire net_49;
wire n201gat;
wire net_15;
wire net_57;
wire n85gat;
wire net_71;
wire n267gat;
wire net_153;
wire net_156;
wire net_84;
wire net_174;
wire net_1;
wire net_92;
wire net_112;
wire net_103;
wire net_139;
wire n423gat;
wire net_43;
wire net_10;
wire net_180;
wire net_21;
wire net_169;
wire net_51;
wire net_171;
wire net_79;
wire n135gat;
wire n1gat;
wire n422gat;
wire n237gat;
wire net_143;
wire net_190;
wire n29gat;
wire net_88;
wire net_145;
wire n138gat;
wire n864gat;
wire net_81;
wire net_163;
wire n86gat;
wire net_67;
wire n121gat;
wire n42gat;
wire net_37;
wire net_188;
wire net_110;
wire net_33;
wire net_48;
wire net_8;
wire net_133;
wire n259gat;

// Start cells
NAND2_X1 inst_145 ( .ZN(net_126), .A2(net_97), .A1(n165gat) );
NAND2_X1 inst_103 ( .ZN(net_36), .A2(net_31), .A1(n42gat) );
NAND2_X1 inst_125 ( .ZN(net_73), .A2(net_72), .A1(n153gat) );
AND2_X4 inst_207 ( .ZN(net_28), .A2(n75gat), .A1(n29gat) );
NAND2_X1 inst_138 ( .ZN(net_122), .A2(net_89), .A1(n195gat) );
NAND2_X1 inst_159 ( .ZN(net_147), .A2(net_123), .A1(net_116) );
AND2_X2 inst_218 ( .A2(net_30), .ZN(n450gat), .A1(n89gat) );
XNOR2_X1 inst_15 ( .ZN(net_48), .A(net_39), .B(n207gat) );
AND4_X1 inst_197 ( .ZN(net_178), .A4(net_172), .A1(net_144), .A2(net_118), .A3(net_7) );
NAND2_X1 inst_134 ( .ZN(net_83), .A2(net_81), .A1(n177gat) );
NAND2_X1 inst_179 ( .ZN(net_191), .A2(net_188), .A1(n219gat) );
XNOR2_X1 inst_24 ( .ZN(net_182), .A(net_180), .B(net_156) );
NAND2_X1 inst_114 ( .ZN(net_85), .A2(net_55), .A1(n55gat) );
XNOR2_X1 inst_6 ( .ZN(net_25), .B(n126gat), .A(n121gat) );
AND4_X1 inst_194 ( .ZN(net_167), .A4(net_162), .A1(net_148), .A2(net_142), .A3(net_1) );
NAND2_X1 inst_131 ( .A2(net_81), .ZN(net_79), .A1(n171gat) );
NAND3_X1 inst_76 ( .A1(net_177), .A3(net_101), .A2(net_78), .ZN(n863gat) );
AND2_X4 inst_214 ( .ZN(net_151), .A2(net_123), .A1(n261gat) );
NAND2_X1 inst_180 ( .ZN(net_192), .A2(net_189), .A1(n219gat) );
NAND2_X1 inst_160 ( .A1(net_141), .ZN(net_133), .A2(net_132) );
NAND2_X1 inst_150 ( .ZN(net_103), .A2(net_102), .A1(n246gat) );
OR2_X4 inst_33 ( .A2(net_122), .A1(net_117), .ZN(net_107) );
NAND2_X1 inst_172 ( .ZN(net_176), .A2(net_175), .A1(net_138) );
NAND2_X1 inst_83 ( .ZN(net_2), .A2(n260gat), .A1(n255gat) );
OR2_X4 inst_47 ( .ZN(net_159), .A2(net_151), .A1(net_141) );
XNOR2_X1 inst_19 ( .ZN(net_158), .A(net_147), .B(n261gat) );
NAND2_X1 inst_123 ( .A2(net_72), .ZN(net_70), .A1(n149gat) );
NAND2_X1 inst_121 ( .ZN(net_68), .A2(net_67), .A1(n106gat) );
XNOR2_X1 inst_2 ( .ZN(net_20), .B(n106gat), .A(n101gat) );
XNOR2_X1 inst_8 ( .ZN(net_34), .A(net_33), .B(n42gat) );
NAND2_X1 inst_118 ( .A2(net_67), .ZN(net_64), .A1(n126gat) );
NAND2_X1 inst_86 ( .ZN(net_4), .A1(n210gat), .A2(n106gat) );
NAND2_X1 inst_153 ( .ZN(net_149), .A1(net_122), .A2(net_121) );
XNOR2_X1 inst_20 ( .ZN(net_161), .A(net_159), .B(net_149) );
OR3_X4 inst_27 ( .ZN(net_84), .A3(net_54), .A2(net_33), .A1(n268gat) );
OR2_X4 inst_38 ( .A2(net_128), .ZN(net_118), .A1(net_117) );
NAND2_X1 inst_100 ( .A2(net_27), .ZN(n421gat), .A1(n80gat) );
NOR2_X1 inst_52 ( .ZN(net_42), .A2(net_32), .A1(net_17) );
NAND2_X1 inst_90 ( .ZN(net_7), .A1(n210gat), .A2(n111gat) );
NAND2_X1 inst_140 ( .A2(net_96), .ZN(net_91), .A1(n246gat) );
AND2_X4 inst_209 ( .A2(net_18), .ZN(n447gat), .A1(n51gat) );
AND2_X4 inst_211 ( .ZN(net_52), .A2(net_45), .A1(n59gat) );
OR2_X4 inst_40 ( .ZN(net_131), .A2(net_130), .A1(net_117) );
NAND2_X1 inst_162 ( .ZN(net_142), .A2(net_141), .A1(n237gat) );
NAND2_X1 inst_167 ( .ZN(net_164), .A2(net_161), .A1(n219gat) );
NAND2_X1 inst_93 ( .ZN(net_10), .A2(n259gat), .A1(n255gat) );
NAND2_X1 inst_81 ( .ZN(net_0), .A2(n96gat), .A1(n210gat) );
NAND2_X1 inst_95 ( .ZN(net_12), .A1(n17gat), .A2(n138gat) );
XOR2_X1 inst_1 ( .Z(net_23), .B(n201gat), .A(n195gat) );
NAND3_X1 inst_72 ( .ZN(net_89), .A2(net_85), .A1(net_70), .A3(net_61) );
NAND2_X1 inst_139 ( .ZN(net_128), .A2(net_90), .A1(n189gat) );
NAND2_X1 inst_155 ( .ZN(net_153), .A1(net_126), .A2(net_105) );
NOR2_X1 inst_59 ( .ZN(net_132), .A1(net_119), .A2(net_98) );
NAND2_X1 inst_135 ( .ZN(net_111), .A2(net_86), .A1(n159gat) );
AND4_X1 inst_196 ( .ZN(net_177), .A4(net_171), .A2(net_146), .A1(net_131), .A3(net_4) );
OR2_X4 inst_44 ( .A1(net_154), .ZN(net_146), .A2(net_145) );
NOR2_X1 inst_55 ( .ZN(net_119), .A2(net_90), .A1(n189gat) );
NAND2_X1 inst_174 ( .ZN(net_181), .A2(net_180), .A1(net_124) );
NAND2_X1 inst_115 ( .A2(net_67), .ZN(net_61), .A1(n121gat) );
OR2_X4 inst_37 ( .A1(net_125), .ZN(net_115), .A2(net_114) );
AND2_X4 inst_210 ( .ZN(net_50), .A1(net_15), .A2(n447gat) );
NAND2_X1 inst_148 ( .ZN(net_101), .A2(net_100), .A1(n246gat) );
NAND2_X1 inst_164 ( .ZN(net_160), .A2(net_159), .A1(net_121) );
INV_X1 inst_191 ( .ZN(net_139), .A(net_106) );
XNOR2_X1 inst_5 ( .ZN(net_24), .B(n189gat), .A(n183gat) );
NAND2_X1 inst_157 ( .ZN(net_143), .A1(net_128), .A2(net_99) );
NAND2_X1 inst_84 ( .ZN(net_16), .A2(n8gat), .A1(n1gat) );
NOR2_X1 inst_51 ( .A2(net_32), .A1(net_16), .ZN(n418gat) );
NAND2_X1 inst_142 ( .A2(net_97), .ZN(net_93), .A1(n246gat) );
NAND3_X1 inst_80 ( .A1(net_194), .A3(net_93), .A2(net_80), .ZN(n879gat) );
NAND2_X1 inst_173 ( .ZN(net_179), .A2(net_174), .A1(n219gat) );
NAND2_X1 inst_105 ( .A2(net_42), .A1(net_36), .ZN(n419gat) );
AND2_X4 inst_213 ( .ZN(net_53), .A2(net_52), .A1(n72gat) );
NAND4_X1 inst_68 ( .A2(net_170), .A4(net_87), .A1(net_75), .A3(net_2), .ZN(n865gat) );
AND2_X2 inst_216 ( .ZN(n391gat), .A2(n86gat), .A1(n85gat) );
NAND3_X1 inst_78 ( .A1(net_190), .A3(net_91), .A2(net_79), .ZN(n880gat) );
OR2_X4 inst_42 ( .A1(net_154), .ZN(net_137), .A2(net_136) );
NAND2_X1 inst_175 ( .ZN(net_183), .A2(net_181), .A1(net_125) );
NOR2_X1 inst_53 ( .ZN(net_55), .A2(net_54), .A1(n268gat) );
AND2_X4 inst_205 ( .ZN(net_27), .A1(n59gat), .A2(n36gat) );
NAND2_X1 inst_177 ( .ZN(net_187), .A2(net_186), .A1(net_110) );
INV_X1 inst_183 ( .ZN(net_117), .A(n237gat) );
NAND2_X1 inst_133 ( .ZN(net_82), .A2(net_81), .A1(n159gat) );
XNOR2_X1 inst_26 ( .ZN(net_189), .A(net_183), .B(net_153) );
NAND2_X1 inst_151 ( .ZN(net_134), .A1(net_111), .A2(net_110) );
NAND2_X1 inst_112 ( .ZN(net_59), .A2(net_58), .A1(n153gat) );
NAND4_X1 inst_64 ( .ZN(net_95), .A2(net_84), .A4(net_68), .A1(net_59), .A3(net_6) );
NAND2_X1 inst_107 ( .ZN(net_51), .A2(net_50), .A1(n17gat) );
NAND4_X1 inst_67 ( .A2(net_167), .A4(net_103), .A1(net_77), .A3(net_9), .ZN(n850gat) );
INV_X1 inst_181 ( .ZN(net_154), .A(n228gat) );
NAND2_X1 inst_127 ( .A2(net_81), .ZN(net_75), .A1(n195gat) );
NAND4_X1 inst_70 ( .A2(net_178), .A4(net_88), .A1(net_76), .A3(net_10), .ZN(n864gat) );
INV_X1 inst_186 ( .A(net_36), .ZN(n390gat) );
NAND2_X1 inst_129 ( .A2(net_81), .ZN(net_77), .A1(n201gat) );
NAND2_X1 inst_92 ( .ZN(net_9), .A2(n267gat), .A1(n255gat) );
OR2_X4 inst_29 ( .ZN(net_110), .A2(net_86), .A1(n159gat) );
INV_X1 inst_189 ( .ZN(net_124), .A(net_104) );
XNOR2_X1 inst_17 ( .B(net_48), .A(net_47), .ZN(n768gat) );
XNOR2_X1 inst_11 ( .ZN(net_40), .B(net_26), .A(net_25) );
NAND2_X1 inst_146 ( .ZN(net_106), .A2(net_95), .A1(n177gat) );
INV_X1 inst_188 ( .A(net_119), .ZN(net_99) );
XNOR2_X1 inst_14 ( .ZN(net_47), .A(net_41), .B(n130gat) );
AND3_X4 inst_202 ( .ZN(net_45), .A3(net_37), .A1(n55gat), .A2(n13gat) );
AND2_X4 inst_206 ( .ZN(net_29), .A2(n75gat), .A1(n59gat) );
INV_X1 inst_187 ( .ZN(net_121), .A(net_98) );
NAND2_X1 inst_122 ( .ZN(net_69), .A2(net_67), .A1(n91gat) );
OR2_X4 inst_31 ( .ZN(net_129), .A2(net_100), .A1(n183gat) );
XNOR2_X1 inst_25 ( .ZN(net_188), .A(net_186), .B(net_134) );
NAND2_X1 inst_126 ( .ZN(net_74), .A2(net_72), .A1(n143gat) );
NAND2_X1 inst_158 ( .ZN(net_145), .A1(net_130), .A2(net_129) );
NAND2_X1 inst_141 ( .ZN(net_92), .A2(net_86), .A1(n246gat) );
NAND4_X1 inst_62 ( .ZN(net_96), .A2(net_84), .A4(net_65), .A1(net_56), .A3(net_12) );
AND4_X1 inst_200 ( .ZN(net_193), .A4(net_191), .A2(net_135), .A1(net_112), .A3(net_3) );
NAND2_X1 inst_110 ( .A2(net_58), .ZN(net_56), .A1(n149gat) );
NAND3_X1 inst_74 ( .ZN(net_102), .A3(net_85), .A2(net_73), .A1(net_64) );
NOR2_X1 inst_57 ( .ZN(net_114), .A2(net_97), .A1(n165gat) );
OR2_X4 inst_35 ( .A2(net_126), .A1(net_117), .ZN(net_109) );
NAND2_X1 inst_99 ( .ZN(net_15), .A1(n59gat), .A2(n156gat) );
OR2_X4 inst_48 ( .ZN(net_155), .A1(net_154), .A2(net_153) );
NAND4_X1 inst_69 ( .ZN(net_186), .A4(net_176), .A1(net_140), .A2(net_126), .A3(net_115) );
OR2_X4 inst_46 ( .A1(net_154), .ZN(net_150), .A2(net_149) );
NAND2_X1 inst_82 ( .ZN(net_1), .A1(n210gat), .A2(n121gat) );
NAND2_X1 inst_136 ( .A2(net_89), .ZN(net_87), .A1(n246gat) );
OR2_X4 inst_30 ( .ZN(net_113), .A2(net_95), .A1(n177gat) );
NAND2_X1 inst_102 ( .A2(net_27), .ZN(n422gat), .A1(n42gat) );
NAND2_X1 inst_108 ( .ZN(net_67), .A2(net_44), .A1(net_43) );
NAND2_X1 inst_165 ( .ZN(net_162), .A2(net_158), .A1(n219gat) );
OR2_X4 inst_32 ( .ZN(net_123), .A2(net_102), .A1(n201gat) );
XNOR2_X1 inst_22 ( .ZN(net_169), .A(net_163), .B(net_143) );
NAND2_X1 inst_144 ( .ZN(net_125), .A2(net_96), .A1(n171gat) );
OR2_X4 inst_34 ( .A2(net_125), .A1(net_117), .ZN(net_108) );
XNOR2_X1 inst_12 ( .ZN(net_41), .B(net_22), .A(net_21) );
AND4_X1 inst_195 ( .ZN(net_170), .A4(net_164), .A1(net_150), .A2(net_107), .A3(net_14) );
NOR2_X1 inst_56 ( .ZN(net_104), .A2(net_96), .A1(n171gat) );
NAND3_X1 inst_71 ( .ZN(net_54), .A2(net_28), .A3(n447gat), .A1(n80gat) );
XNOR2_X1 inst_21 ( .ZN(net_168), .A(net_165), .B(net_145) );
NAND2_X1 inst_104 ( .ZN(net_35), .A2(net_29), .A1(n42gat) );
NAND4_X1 inst_60 ( .ZN(net_43), .A3(net_37), .A4(net_35), .A1(n51gat), .A2(n17gat) );
AND2_X4 inst_215 ( .ZN(net_175), .A2(net_173), .A1(net_113) );
NAND2_X1 inst_169 ( .ZN(net_173), .A2(net_166), .A1(net_130) );
NAND2_X1 inst_168 ( .ZN(net_166), .A2(net_165), .A1(net_129) );
NAND2_X1 inst_97 ( .ZN(net_32), .A2(n17gat), .A1(n13gat) );
NAND2_X1 inst_161 ( .ZN(net_140), .A1(net_139), .A2(net_138) );
NAND2_X1 inst_124 ( .A2(net_72), .ZN(net_71), .A1(n146gat) );
XNOR2_X1 inst_18 ( .A(net_49), .B(net_46), .ZN(n767gat) );
XNOR2_X1 inst_16 ( .ZN(net_49), .A(net_40), .B(n135gat) );
AND2_X4 inst_208 ( .ZN(net_31), .A2(n36gat), .A1(n29gat) );
NAND2_X1 inst_88 ( .ZN(net_5), .A2(n91gat), .A1(n210gat) );
AND2_X2 inst_220 ( .A2(net_30), .ZN(n423gat), .A1(n90gat) );
XNOR2_X1 inst_3 ( .ZN(net_21), .B(n165gat), .A(n159gat) );
NAND2_X1 inst_156 ( .A2(net_139), .ZN(net_127), .A1(n237gat) );
XNOR2_X1 inst_9 ( .ZN(net_38), .B(net_20), .A(net_19) );
NAND2_X1 inst_113 ( .ZN(net_60), .A2(net_58), .A1(n143gat) );
NAND2_X1 inst_170 ( .ZN(net_171), .A2(net_168), .A1(n219gat) );
AND4_X1 inst_198 ( .ZN(net_184), .A4(net_179), .A2(net_137), .A1(net_127), .A3(net_13) );
OR2_X4 inst_50 ( .ZN(net_180), .A2(net_175), .A1(net_139) );
NAND2_X1 inst_137 ( .A2(net_90), .ZN(net_88), .A1(n246gat) );
AND4_X1 inst_199 ( .ZN(net_190), .A4(net_185), .A2(net_157), .A1(net_108), .A3(net_0) );
OR2_X4 inst_41 ( .A1(net_154), .ZN(net_135), .A2(net_134) );
NAND2_X1 inst_130 ( .A2(net_81), .ZN(net_78), .A1(n183gat) );
NAND2_X1 inst_91 ( .ZN(net_8), .A1(n8gat), .A2(n138gat) );
NAND2_X1 inst_132 ( .A2(net_81), .ZN(net_80), .A1(n165gat) );
NAND2_X1 inst_143 ( .A2(net_95), .ZN(net_94), .A1(n246gat) );
NAND2_X1 inst_176 ( .ZN(net_185), .A2(net_182), .A1(n219gat) );
NAND2_X1 inst_152 ( .ZN(net_136), .A2(net_113), .A1(net_106) );
NOR2_X1 inst_58 ( .ZN(net_138), .A1(net_114), .A2(net_104) );
OR2_X4 inst_36 ( .A1(net_117), .ZN(net_112), .A2(net_111) );
NAND2_X1 inst_147 ( .ZN(net_130), .A2(net_100), .A1(n183gat) );
NAND2_X1 inst_87 ( .ZN(net_17), .A2(n26gat), .A1(n1gat) );
NAND4_X1 inst_61 ( .ZN(net_44), .A4(net_34), .A2(n447gat), .A3(n59gat), .A1(n156gat) );
AND3_X2 inst_203 ( .A3(net_45), .ZN(n448gat), .A2(n68gat), .A1(n29gat) );
OR2_X4 inst_45 ( .A1(net_154), .ZN(net_148), .A2(net_147) );
NAND2_X1 inst_96 ( .ZN(net_13), .A1(n210gat), .A2(n101gat) );
AND2_X4 inst_212 ( .ZN(net_58), .A2(net_50), .A1(n55gat) );
NAND2_X1 inst_101 ( .A2(net_29), .ZN(n420gat), .A1(n80gat) );
XOR2_X1 inst_0 ( .Z(net_19), .B(n96gat), .A(n91gat) );
INV_X1 inst_184 ( .ZN(net_37), .A(net_16) );
XNOR2_X1 inst_10 ( .ZN(net_39), .B(net_24), .A(net_23) );
XNOR2_X1 inst_4 ( .ZN(net_22), .B(n177gat), .A(n171gat) );
NAND4_X1 inst_65 ( .ZN(net_86), .A2(net_84), .A4(net_69), .A1(net_60), .A3(net_8) );
NAND2_X1 inst_178 ( .A2(net_187), .A1(net_111), .ZN(n866gat) );
NAND2_X1 inst_89 ( .ZN(net_6), .A1(n152gat), .A2(n138gat) );
OR2_X4 inst_28 ( .ZN(net_30), .A2(n88gat), .A1(n87gat) );
NAND2_X1 inst_111 ( .A2(net_58), .ZN(net_57), .A1(n146gat) );
NAND4_X1 inst_66 ( .ZN(net_165), .A4(net_152), .A1(net_133), .A2(net_128), .A3(net_120) );
NAND2_X1 inst_117 ( .A2(net_67), .ZN(net_63), .A1(n111gat) );
NAND2_X1 inst_98 ( .ZN(net_14), .A1(n210gat), .A2(n116gat) );
INV_X1 inst_190 ( .A(net_114), .ZN(net_105) );
NAND4_X1 inst_63 ( .ZN(net_97), .A2(net_84), .A4(net_66), .A1(net_57), .A3(net_11) );
XNOR2_X1 inst_7 ( .ZN(net_26), .B(n116gat), .A(n111gat) );
AND3_X2 inst_204 ( .A3(net_52), .ZN(n449gat), .A1(n74gat), .A2(n68gat) );
INV_X1 inst_185 ( .ZN(net_18), .A(net_17) );
INV_X1 inst_182 ( .ZN(net_33), .A(n17gat) );
OR2_X4 inst_49 ( .ZN(net_157), .A2(net_156), .A1(net_154) );
NAND2_X1 inst_120 ( .A2(net_67), .ZN(net_66), .A1(n96gat) );
NAND2_X1 inst_154 ( .ZN(net_156), .A1(net_125), .A2(net_124) );
XNOR2_X1 inst_13 ( .ZN(net_46), .A(net_38), .B(n130gat) );
NAND2_X1 inst_119 ( .A2(net_67), .ZN(net_65), .A1(n101gat) );
NAND3_X1 inst_75 ( .ZN(net_100), .A3(net_85), .A2(net_74), .A1(net_63) );
INV_X1 inst_192 ( .ZN(net_141), .A(net_116) );
NAND2_X1 inst_166 ( .ZN(net_163), .A2(net_160), .A1(net_122) );
NAND2_X1 inst_116 ( .A2(net_67), .ZN(net_62), .A1(n116gat) );
NAND2_X1 inst_163 ( .ZN(net_152), .A1(net_151), .A2(net_132) );
NAND2_X1 inst_85 ( .ZN(net_3), .A2(n268gat), .A1(n210gat) );
NOR2_X1 inst_54 ( .ZN(net_98), .A2(net_89), .A1(n195gat) );
NAND3_X1 inst_79 ( .A1(net_193), .A3(net_92), .A2(net_82), .ZN(n878gat) );
NAND2_X1 inst_109 ( .ZN(net_72), .A2(net_51), .A1(n1gat) );
NAND2_X1 inst_106 ( .A2(net_42), .ZN(n446gat), .A1(n390gat) );
AND2_X2 inst_219 ( .A2(net_31), .ZN(n389gat), .A1(n80gat) );
AND4_X1 inst_201 ( .ZN(net_194), .A4(net_192), .A2(net_155), .A1(net_109), .A3(net_5) );
AND4_X1 inst_193 ( .ZN(net_81), .A4(net_53), .A1(n73gat), .A3(n68gat), .A2(n42gat) );
NAND2_X1 inst_149 ( .ZN(net_116), .A2(net_102), .A1(n201gat) );
OR2_X4 inst_43 ( .A1(net_154), .ZN(net_144), .A2(net_143) );
OR2_X4 inst_39 ( .A1(net_122), .ZN(net_120), .A2(net_119) );
NAND2_X1 inst_128 ( .A2(net_81), .ZN(net_76), .A1(n189gat) );
NAND3_X1 inst_73 ( .ZN(net_90), .A2(net_85), .A1(net_71), .A3(net_62) );
AND2_X2 inst_217 ( .A2(net_28), .ZN(n388gat), .A1(n42gat) );
XNOR2_X1 inst_23 ( .ZN(net_174), .B(net_173), .A(net_136) );
NAND2_X1 inst_171 ( .ZN(net_172), .A2(net_169), .A1(n219gat) );
NAND3_X1 inst_77 ( .A1(net_184), .A3(net_94), .A2(net_83), .ZN(n874gat) );
NAND2_X1 inst_94 ( .ZN(net_11), .A1(n51gat), .A2(n138gat) );

endmodule
