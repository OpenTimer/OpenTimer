module s349 (
B0,
A1,
B1,
A2,
A3,
blif_clk_net,
START,
B3,
A0,
blif_reset_net,
B2,
P7,
P5,
CNTVCON2,
P2,
P1,
CNTVCO2,
P0,
P6,
READY,
P3,
P4);

// Start PIs
input B0;
input A1;
input B1;
input A2;
input A3;
input blif_clk_net;
input START;
input B3;
input A0;
input blif_reset_net;
input B2;

// Start POs
output P7;
output P5;
output CNTVCON2;
output P2;
output P1;
output CNTVCO2;
output P0;
output P6;
output READY;
output P3;
output P4;

// Start wires
wire net_166;
wire net_107;
wire net_47;
wire net_179;
wire net_176;
wire net_159;
wire net_61;
wire net_137;
wire net_132;
wire net_54;
wire net_105;
wire net_62;
wire P3;
wire net_6;
wire net_129;
wire net_119;
wire net_98;
wire net_23;
wire P5;
wire net_117;
wire net_12;
wire B1;
wire net_151;
wire net_74;
wire net_53;
wire net_93;
wire net_168;
wire net_135;
wire net_130;
wire net_147;
wire net_127;
wire net_14;
wire P1;
wire net_113;
wire net_26;
wire net_76;
wire blif_clk_net;
wire net_101;
wire net_32;
wire net_111;
wire net_90;
wire net_40;
wire net_100;
wire net_85;
wire net_69;
wire net_124;
wire net_161;
wire net_141;
wire net_160;
wire net_83;
wire net_115;
wire B3;
wire net_4;
wire net_95;
wire net_17;
wire net_173;
wire net_78;
wire A1;
wire net_27;
wire net_164;
wire net_56;
wire net_87;
wire net_0;
wire net_155;
wire net_35;
wire net_16;
wire net_22;
wire net_181;
wire net_39;
wire net_157;
wire net_144;
wire net_102;
wire net_2;
wire net_59;
wire net_9;
wire net_42;
wire net_120;
wire A3;
wire net_109;
wire net_80;
wire net_65;
wire blif_reset_net;
wire net_50;
wire net_162;
wire net_96;
wire net_66;
wire net_38;
wire net_44;
wire net_167;
wire net_136;
wire net_134;
wire net_19;
wire net_89;
wire net_45;
wire net_126;
wire B0;
wire net_34;
wire net_108;
wire net_178;
wire net_150;
wire net_63;
wire P2;
wire net_152;
wire net_116;
wire net_30;
wire net_175;
wire net_91;
wire net_106;
wire net_24;
wire net_55;
wire net_99;
wire net_46;
wire net_140;
wire net_118;
wire P7;
wire net_148;
wire net_104;
wire net_146;
wire net_72;
wire net_122;
wire net_25;
wire net_7;
wire net_70;
wire P4;
wire net_172;
wire net_5;
wire net_52;
wire net_165;
wire net_128;
wire P0;
wire net_138;
wire net_13;
wire P6;
wire net_94;
wire net_11;
wire CNTVCON2;
wire net_18;
wire net_123;
wire net_131;
wire net_114;
wire CNTVCO2;
wire net_170;
wire net_29;
wire net_68;
wire net_149;
wire net_142;
wire net_77;
wire net_20;
wire net_31;
wire net_36;
wire net_49;
wire net_158;
wire net_15;
wire net_41;
wire net_57;
wire A2;
wire net_71;
wire net_153;
wire START;
wire net_156;
wire net_3;
wire net_84;
wire net_174;
wire net_154;
wire net_112;
wire net_1;
wire net_92;
wire net_103;
wire net_139;
wire net_43;
wire net_10;
wire net_180;
wire net_28;
wire net_169;
wire net_21;
wire net_51;
wire net_171;
wire net_79;
wire net_143;
wire net_97;
wire net_88;
wire net_182;
wire net_145;
wire net_60;
wire net_81;
wire net_163;
wire net_58;
wire B2;
wire net_67;
wire net_82;
wire net_64;
wire net_37;
wire net_110;
wire net_121;
wire net_73;
wire net_33;
wire net_48;
wire net_177;
wire net_8;
wire net_75;
wire net_86;
wire net_133;
wire READY;
wire A0;
wire net_125;

// Start cells
CLKBUF_X2 inst_145 ( .A(net_133), .Z(net_134) );
INV_X4 inst_103 ( .ZN(net_64), .A(net_52) );
DFFR_X2 inst_125 ( .RN(net_102), .D(net_73), .QN(net_6), .CK(net_179) );
DFFR_X1 inst_138 ( .D(net_103), .RN(net_102), .QN(net_2), .CK(net_150) );
CLKBUF_X2 inst_159 ( .A(net_147), .Z(net_148) );
NOR2_X2 inst_15 ( .ZN(net_85), .A2(net_77), .A1(START) );
DFFR_X2 inst_134 ( .RN(net_102), .D(net_87), .QN(net_13), .CK(net_146) );
CLKBUF_X2 inst_179 ( .A(blif_clk_net), .Z(net_168) );
NAND3_X2 inst_24 ( .A2(net_100), .ZN(net_99), .A3(net_95), .A1(net_61) );
INV_X2 inst_114 ( .A(net_42), .ZN(P1) );
OR2_X2 inst_6 ( .A2(net_113), .ZN(net_90), .A1(net_89) );
DFFR_X2 inst_131 ( .RN(net_102), .D(net_86), .QN(net_9), .CK(net_159) );
INV_X4 inst_76 ( .A(net_128), .ZN(net_126) );
CLKBUF_X2 inst_180 ( .A(net_168), .Z(net_169) );
CLKBUF_X2 inst_160 ( .A(net_148), .Z(net_149) );
CLKBUF_X2 inst_150 ( .A(net_138), .Z(net_139) );
NAND2_X4 inst_33 ( .ZN(net_112), .A1(net_52), .A2(net_2) );
CLKBUF_X2 inst_172 ( .A(net_137), .Z(net_161) );
INV_X4 inst_83 ( .ZN(net_56), .A(net_3) );
NAND2_X2 inst_47 ( .ZN(net_39), .A1(net_38), .A2(READY) );
NAND3_X2 inst_19 ( .ZN(net_71), .A3(net_70), .A2(net_46), .A1(P5) );
INV_X1 inst_123 ( .ZN(net_102), .A(blif_reset_net) );
INV_X2 inst_121 ( .ZN(net_111), .A(net_65) );
OR2_X4 inst_2 ( .ZN(net_40), .A2(READY), .A1(B3) );
NOR3_X2 inst_8 ( .ZN(net_80), .A1(net_78), .A3(net_51), .A2(START) );
INV_X2 inst_118 ( .ZN(net_70), .A(net_68) );
INV_X4 inst_86 ( .ZN(net_100), .A(START) );
CLKBUF_X2 inst_153 ( .A(net_141), .Z(net_142) );
NAND3_X2 inst_20 ( .A3(net_117), .ZN(net_116), .A1(net_113), .A2(P6) );
NAND3_X2 inst_27 ( .A3(net_109), .A1(net_108), .ZN(net_103), .A2(net_100) );
NAND2_X4 inst_38 ( .A1(net_105), .ZN(net_94), .A2(net_89) );
INV_X4 inst_100 ( .ZN(net_45), .A(net_32) );
NAND2_X2 inst_52 ( .ZN(net_57), .A1(net_35), .A2(net_34) );
INV_X4 inst_90 ( .ZN(net_17), .A(net_2) );
AND2_X4 inst_140 ( .A1(net_121), .ZN(net_118), .A2(net_0) );
NAND2_X4 inst_40 ( .A1(net_104), .ZN(net_97), .A2(net_66) );
CLKBUF_X2 inst_162 ( .A(net_148), .Z(net_151) );
CLKBUF_X2 inst_167 ( .A(net_146), .Z(net_156) );
INV_X4 inst_93 ( .ZN(net_18), .A(net_16) );
INV_X4 inst_81 ( .ZN(net_24), .A(net_10) );
INV_X4 inst_95 ( .ZN(net_23), .A(net_18) );
XNOR2_X2 inst_1 ( .ZN(net_79), .A(net_78), .B(net_27) );
MUX2_X2 inst_72 ( .S(net_123), .Z(net_83), .A(net_60), .B(net_38) );
CLKBUF_X3 inst_139 ( .A(net_121), .Z(P0) );
CLKBUF_X2 inst_155 ( .A(net_143), .Z(net_144) );
NAND2_X2 inst_59 ( .A2(net_128), .ZN(net_109), .A1(net_20) );
DFFR_X2 inst_135 ( .RN(net_102), .D(net_96), .QN(net_0), .CK(net_142) );
NAND2_X2 inst_44 ( .A2(net_121), .ZN(net_53), .A1(net_33) );
NAND2_X2 inst_55 ( .ZN(net_60), .A1(net_44), .A2(net_43) );
CLKBUF_X2 inst_174 ( .A(net_162), .Z(net_163) );
INV_X2 inst_115 ( .ZN(net_19), .A(P5) );
NAND2_X4 inst_37 ( .A1(net_114), .A2(net_112), .ZN(net_105) );
CLKBUF_X2 inst_148 ( .A(net_136), .Z(net_137) );
CLKBUF_X2 inst_164 ( .A(net_152), .Z(net_153) );
CLKBUF_X2 inst_191 ( .A(net_154), .Z(net_180) );
OR2_X2 inst_5 ( .ZN(net_35), .A2(READY), .A1(B0) );
CLKBUF_X2 inst_157 ( .A(net_145), .Z(net_146) );
INV_X4 inst_84 ( .ZN(net_38), .A(net_12) );
NAND2_X2 inst_51 ( .ZN(net_66), .A1(net_56), .A2(net_53) );
CLKBUF_X2 inst_142 ( .A(net_130), .Z(net_131) );
INV_X4 inst_80 ( .ZN(net_16), .A(net_8) );
CLKBUF_X2 inst_173 ( .A(net_161), .Z(net_162) );
INV_X2 inst_105 ( .A(net_128), .ZN(net_127) );
MUX2_X2 inst_68 ( .S(net_122), .Z(net_72), .B(net_33), .A(A3) );
INV_X4 inst_78 ( .ZN(net_120), .A(P0) );
NAND2_X2 inst_42 ( .ZN(net_48), .A1(net_27), .A2(net_23) );
CLKBUF_X2 inst_175 ( .A(net_139), .Z(net_164) );
NAND2_X2 inst_53 ( .ZN(net_58), .A1(net_41), .A2(net_39) );
CLKBUF_X2 inst_177 ( .A(net_165), .Z(net_166) );
CLKBUF_X2 inst_183 ( .A(net_171), .Z(net_172) );
DFFR_X2 inst_133 ( .QN(net_121), .RN(net_102), .D(net_88), .CK(net_132) );
NAND3_X2 inst_26 ( .A2(net_125), .ZN(net_108), .A3(net_107), .A1(net_106) );
CLKBUF_X2 inst_151 ( .A(net_139), .Z(net_140) );
INV_X2 inst_112 ( .A(net_38), .ZN(P2) );
NAND2_X2 inst_64 ( .ZN(net_115), .A2(net_94), .A1(net_90) );
INV_X2 inst_107 ( .A(net_114), .ZN(net_113) );
NAND2_X2 inst_67 ( .A1(net_126), .ZN(net_98), .A2(net_97) );
CLKBUF_X2 inst_181 ( .A(net_169), .Z(net_170) );
DFFR_X2 inst_127 ( .RN(net_102), .D(net_80), .QN(net_8), .CK(net_172) );
MUX2_X2 inst_70 ( .S(net_122), .Z(net_74), .B(net_21), .A(A1) );
CLKBUF_X2 inst_186 ( .A(net_174), .Z(net_175) );
DFFR_X2 inst_129 ( .RN(net_102), .D(net_85), .QN(net_10), .CK(net_163) );
INV_X4 inst_92 ( .A(net_15), .ZN(P5) );
NAND2_X4 inst_29 ( .A1(net_118), .ZN(net_68), .A2(net_30) );
CLKBUF_X2 inst_189 ( .A(net_158), .Z(net_178) );
NAND3_X4 inst_17 ( .ZN(net_49), .A2(net_24), .A3(net_16), .A1(net_9) );
NOR2_X2 inst_11 ( .ZN(net_51), .A2(net_49), .A1(net_26) );
CLKBUF_X2 inst_146 ( .A(net_134), .Z(net_135) );
CLKBUF_X2 inst_188 ( .A(net_176), .Z(net_177) );
NOR2_X2 inst_14 ( .A1(net_129), .ZN(net_81), .A2(net_70) );
CLKBUF_X2 inst_187 ( .A(net_175), .Z(net_176) );
INV_X2 inst_122 ( .A(net_94), .ZN(net_92) );
NAND2_X4 inst_31 ( .ZN(net_128), .A2(net_122), .A1(net_49) );
NAND3_X2 inst_25 ( .ZN(net_101), .A2(net_100), .A3(net_98), .A1(net_63) );
DFFR_X2 inst_126 ( .RN(net_102), .D(net_75), .QN(net_4), .CK(net_177) );
CLKBUF_X2 inst_158 ( .A(net_138), .Z(net_147) );
CLKBUF_X2 inst_141 ( .A(blif_clk_net), .Z(net_130) );
NAND2_X2 inst_62 ( .A1(net_128), .ZN(net_82), .A2(net_57) );
INV_X2 inst_110 ( .A(net_56), .ZN(P7) );
MUX2_X2 inst_74 ( .S(net_124), .Z(net_87), .B(net_69), .A(net_59) );
NAND2_X2 inst_57 ( .A2(net_128), .ZN(net_62), .A1(net_54) );
NAND2_X4 inst_35 ( .ZN(net_89), .A1(net_64), .A2(net_17) );
INV_X4 inst_99 ( .A(net_49), .ZN(READY) );
NAND2_X2 inst_48 ( .ZN(net_43), .A1(net_42), .A2(READY) );
MUX2_X2 inst_69 ( .S(net_122), .Z(net_73), .B(net_28), .A(A2) );
NAND2_X2 inst_46 ( .ZN(net_37), .A1(net_36), .A2(READY) );
INV_X4 inst_82 ( .ZN(net_21), .A(net_5) );
DFFR_X2 inst_136 ( .RN(net_102), .D(net_99), .QN(net_1), .CK(net_140) );
NAND2_X4 inst_30 ( .A1(net_121), .ZN(net_29), .A2(net_28) );
INV_X4 inst_102 ( .ZN(net_46), .A(net_45) );
INV_X2 inst_108 ( .ZN(net_33), .A(net_7) );
CLKBUF_X2 inst_165 ( .A(net_153), .Z(net_154) );
NAND2_X4 inst_32 ( .ZN(net_129), .A1(net_45), .A2(net_15) );
NAND3_X2 inst_22 ( .A2(net_127), .A3(net_116), .A1(net_115), .ZN(net_95) );
CLKBUF_X2 inst_144 ( .A(net_131), .Z(net_133) );
NAND2_X4 inst_34 ( .ZN(net_119), .A2(net_68), .A1(net_47) );
NOR2_X2 inst_12 ( .ZN(net_78), .A1(net_25), .A2(READY) );
NAND2_X2 inst_56 ( .A2(net_128), .ZN(net_61), .A1(net_19) );
MUX2_X2 inst_71 ( .S(net_122), .Z(net_75), .B(net_30), .A(A0) );
NAND3_X2 inst_21 ( .A2(net_126), .ZN(net_93), .A3(net_91), .A1(net_71) );
INV_X4 inst_104 ( .ZN(net_67), .A(net_66) );
NAND2_X2 inst_60 ( .ZN(net_69), .A2(net_68), .A1(net_55) );
CLKBUF_X2 inst_169 ( .A(net_157), .Z(net_158) );
CLKBUF_X2 inst_168 ( .A(net_156), .Z(net_157) );
INV_X4 inst_97 ( .ZN(net_25), .A(net_23) );
CLKBUF_X2 inst_161 ( .A(net_149), .Z(net_150) );
DFFR_X2 inst_124 ( .RN(net_102), .D(net_72), .QN(net_7), .CK(net_182) );
NAND3_X2 inst_18 ( .ZN(net_122), .A2(net_18), .A3(net_10), .A1(net_9) );
NOR2_X2 inst_16 ( .ZN(net_86), .A2(net_79), .A1(START) );
INV_X4 inst_88 ( .ZN(net_15), .A(net_1) );
OR2_X4 inst_3 ( .ZN(net_41), .A2(READY), .A1(B2) );
CLKBUF_X2 inst_156 ( .A(net_144), .Z(net_145) );
NOR2_X2 inst_9 ( .A2(net_48), .A1(net_14), .ZN(CNTVCO2) );
INV_X2 inst_113 ( .A(net_36), .ZN(P3) );
CLKBUF_X2 inst_170 ( .A(net_158), .Z(net_159) );
NAND2_X2 inst_50 ( .ZN(net_55), .A1(net_54), .A2(net_31) );
DFFR_X2 inst_137 ( .RN(net_102), .D(net_101), .QN(net_3), .CK(net_137) );
NAND2_X4 inst_41 ( .A2(net_110), .ZN(net_106), .A1(net_97) );
DFFR_X2 inst_130 ( .RN(net_102), .D(net_83), .QN(net_11), .CK(net_160) );
INV_X4 inst_91 ( .A(net_24), .ZN(net_14) );
DFFR_X2 inst_132 ( .RN(net_102), .D(net_84), .QN(net_12), .CK(net_155) );
CLKBUF_X2 inst_143 ( .A(net_131), .Z(net_132) );
CLKBUF_X2 inst_176 ( .A(net_164), .Z(net_165) );
CLKBUF_X2 inst_152 ( .A(net_138), .Z(net_141) );
NAND2_X2 inst_58 ( .A2(net_128), .ZN(net_63), .A1(net_56) );
NAND2_X4 inst_36 ( .A2(net_129), .A1(net_119), .ZN(net_114) );
CLKBUF_X2 inst_147 ( .A(net_135), .Z(net_136) );
INV_X4 inst_87 ( .ZN(net_42), .A(net_11) );
NAND2_X2 inst_61 ( .A2(net_125), .ZN(net_76), .A1(net_42) );
NAND2_X2 inst_45 ( .A1(net_120), .ZN(net_34), .A2(READY) );
INV_X4 inst_96 ( .ZN(net_27), .A(net_9) );
INV_X4 inst_101 ( .ZN(net_52), .A(net_29) );
XNOR2_X2 inst_0 ( .ZN(net_77), .A(net_50), .B(net_24) );
CLKBUF_X2 inst_184 ( .A(net_142), .Z(net_173) );
NOR2_X2 inst_10 ( .ZN(net_50), .A1(net_48), .A2(READY) );
OR2_X4 inst_4 ( .ZN(net_44), .A2(READY), .A1(B1) );
NAND2_X2 inst_65 ( .ZN(net_110), .A2(net_94), .A1(net_67) );
CLKBUF_X2 inst_178 ( .A(net_166), .Z(net_167) );
INV_X4 inst_89 ( .ZN(net_54), .A(net_0) );
NAND2_X4 inst_28 ( .A2(net_121), .ZN(net_22), .A1(net_21) );
INV_X2 inst_111 ( .A(net_54), .ZN(P4) );
NAND2_X2 inst_66 ( .ZN(net_107), .A2(net_92), .A1(net_65) );
INV_X2 inst_117 ( .ZN(net_26), .A(net_25) );
INV_X4 inst_98 ( .ZN(net_32), .A(net_22) );
CLKBUF_X2 inst_190 ( .A(net_178), .Z(net_179) );
NAND2_X2 inst_63 ( .ZN(net_88), .A2(net_82), .A1(net_76) );
OR2_X2 inst_7 ( .A2(net_113), .ZN(net_91), .A1(net_81) );
CLKBUF_X2 inst_185 ( .A(net_173), .Z(net_174) );
CLKBUF_X2 inst_182 ( .A(net_170), .Z(net_171) );
NAND2_X2 inst_49 ( .ZN(net_47), .A1(net_32), .A2(net_1) );
INV_X2 inst_120 ( .ZN(net_117), .A(net_64) );
CLKBUF_X2 inst_154 ( .A(net_138), .Z(net_143) );
NOR2_X2 inst_13 ( .ZN(net_65), .A1(net_56), .A2(net_53) );
INV_X2 inst_119 ( .ZN(CNTVCON2), .A(CNTVCO2) );
INV_X8 inst_75 ( .A(net_128), .ZN(net_123) );
CLKBUF_X2 inst_192 ( .A(net_180), .Z(net_181) );
CLKBUF_X2 inst_166 ( .A(net_154), .Z(net_155) );
INV_X2 inst_116 ( .ZN(net_20), .A(P6) );
CLKBUF_X2 inst_163 ( .A(net_151), .Z(net_152) );
INV_X4 inst_85 ( .ZN(net_30), .A(net_4) );
NAND2_X2 inst_54 ( .ZN(net_59), .A1(net_40), .A2(net_37) );
INV_X4 inst_79 ( .ZN(net_36), .A(net_13) );
INV_X2 inst_109 ( .ZN(net_28), .A(net_6) );
INV_X2 inst_106 ( .A(net_128), .ZN(net_125) );
CLKBUF_X2 inst_193 ( .A(net_181), .Z(net_182) );
CLKBUF_X2 inst_149 ( .A(net_130), .Z(net_138) );
NAND2_X2 inst_43 ( .A2(net_121), .ZN(net_31), .A1(net_30) );
NAND2_X4 inst_39 ( .A2(net_111), .ZN(net_104), .A1(net_94) );
DFFR_X2 inst_128 ( .RN(net_102), .D(net_74), .QN(net_5), .CK(net_167) );
MUX2_X2 inst_73 ( .S(net_123), .Z(net_84), .A(net_58), .B(net_36) );
NAND3_X2 inst_23 ( .A2(net_100), .ZN(net_96), .A3(net_93), .A1(net_62) );
CLKBUF_X2 inst_171 ( .A(net_132), .Z(net_160) );
INV_X4 inst_77 ( .A(net_128), .ZN(net_124) );
INV_X4 inst_94 ( .A(net_17), .ZN(P6) );

endmodule
