module tv80 (
x884,
x825,
x717,
x1023,
x916,
x964,
x1012,
x672,
x800,
x856,
x947,
x956,
x762,
x974,
x332,
x179,
x423,
x606,
x557,
x79,
x285,
x633,
x0,
x160,
x142,
x475,
x40,
x307,
x256,
x450,
x593,
x409,
x90,
x204,
x639,
x350,
x626,
x128,
x388,
x23,
x437,
x368,
x232,
x615,
x105,
x60);

// Start PIs
input x884;
input x825;
input x717;
input x1023;
input x916;
input x964;
input x1012;
input x672;
input x800;
input x856;
input x947;
input x956;
input x762;
input x974;

// Start POs
output x332;
output x179;
output x423;
output x606;
output x557;
output x79;
output x285;
output x633;
output x0;
output x160;
output x142;
output x475;
output x40;
output x307;
output x256;
output x450;
output x593;
output x409;
output x90;
output x204;
output x639;
output x350;
output x626;
output x128;
output x388;
output x23;
output x437;
output x368;
output x232;
output x615;
output x105;
output x60;

// Start wires
wire net_5030;
wire net_2449;
wire net_4065;
wire net_1317;
wire net_416;
wire net_215;
wire net_2394;
wire net_4854;
wire net_2418;
wire net_1382;
wire net_943;
wire net_4598;
wire net_4508;
wire net_4392;
wire net_1897;
wire net_980;
wire net_53;
wire net_3498;
wire net_2542;
wire net_1786;
wire net_1377;
wire net_4513;
wire net_3996;
wire net_4382;
wire net_1393;
wire net_2169;
wire net_1324;
wire net_4934;
wire net_2256;
wire net_4306;
wire net_264;
wire net_3904;
wire net_4122;
wire net_4315;
wire net_2207;
wire net_263;
wire net_4323;
wire net_3527;
wire net_1138;
wire net_2769;
wire net_4996;
wire net_3483;
wire net_3707;
wire net_1064;
wire net_2082;
wire net_5035;
wire net_3292;
wire net_1439;
wire x717;
wire net_4832;
wire net_4464;
wire net_4189;
wire net_1778;
wire net_508;
wire net_5098;
wire net_1090;
wire net_3685;
wire net_4285;
wire net_703;
wire net_4434;
wire net_193;
wire net_4744;
wire net_5273;
wire net_201;
wire net_5077;
wire net_2942;
wire net_3817;
wire net_3280;
wire net_4043;
wire net_3085;
wire net_2896;
wire net_3281;
wire net_4258;
wire net_4442;
wire net_3949;
wire net_3134;
wire net_1852;
wire net_1720;
wire net_1555;
wire net_3818;
wire net_3434;
wire net_2060;
wire net_2051;
wire net_2780;
wire net_4535;
wire net_4480;
wire net_789;
wire net_3756;
wire net_3244;
wire net_593;
wire net_2171;
wire net_4169;
wire net_2765;
wire net_3833;
wire net_742;
wire net_5139;
wire net_4521;
wire net_2425;
wire net_2830;
wire net_4509;
wire net_1198;
wire net_2509;
wire net_3975;
wire net_5137;
wire net_2862;
wire net_1860;
wire net_2457;
wire net_883;
wire net_2156;
wire net_1432;
wire net_4108;
wire net_1312;
wire net_2957;
wire net_4801;
wire net_446;
wire net_1516;
wire net_1712;
wire net_5290;
wire net_4314;
wire net_3063;
wire net_1083;
wire net_3546;
wire net_3343;
wire net_3423;
wire net_1499;
wire net_964;
wire net_3326;
wire net_1453;
wire net_2913;
wire net_3295;
wire net_2239;
wire net_4379;
wire net_3394;
wire net_3542;
wire net_2268;
wire net_634;
wire net_4680;
wire net_2846;
wire net_2303;
wire net_371;
wire net_3903;
wire net_4369;
wire net_1735;
wire net_2787;
wire net_2210;
wire net_4050;
wire net_2176;
wire net_1571;
wire net_4904;
wire net_2466;
wire net_4699;
wire net_997;
wire net_5090;
wire net_256;
wire net_4929;
wire net_3959;
wire net_850;
wire net_4309;
wire net_1140;
wire net_2764;
wire net_1464;
wire net_5217;
wire net_4973;
wire net_679;
wire net_1168;
wire net_2680;
wire net_3196;
wire net_308;
wire net_515;
wire net_4835;
wire net_3090;
wire net_5121;
wire net_3987;
wire net_223;
wire net_1009;
wire net_715;
wire net_2077;
wire net_890;
wire net_2219;
wire net_2745;
wire net_2546;
wire net_5084;
wire net_3965;
wire net_1876;
wire net_2471;
wire net_312;
wire net_2404;
wire net_130;
wire net_2627;
wire net_572;
wire net_5289;
wire net_5116;
wire net_147;
wire net_481;
wire net_369;
wire net_1662;
wire net_4358;
wire net_1079;
wire net_3935;
wire net_2444;
wire net_5198;
wire net_2809;
wire net_1188;
wire net_3235;
wire net_5297;
wire net_780;
wire net_4938;
wire net_3586;
wire net_3184;
wire net_1446;
wire net_541;
wire net_1251;
wire net_2391;
wire x79;
wire net_5263;
wire net_2802;
wire net_4614;
wire net_2906;
wire net_456;
wire net_155;
wire net_1697;
wire net_4222;
wire net_4163;
wire net_3850;
wire net_1753;
wire net_349;
wire net_2435;
wire net_245;
wire net_3428;
wire net_1409;
wire net_4858;
wire net_2383;
wire net_4264;
wire net_2977;
wire net_493;
wire net_3491;
wire net_1428;
wire net_987;
wire net_277;
wire net_4251;
wire net_1965;
wire net_5222;
wire net_3620;
wire net_89;
wire net_4238;
wire net_3071;
wire net_2350;
wire net_3271;
wire net_680;
wire net_338;
wire net_4494;
wire net_2998;
wire net_721;
wire net_243;
wire net_3226;
wire net_3143;
wire net_2757;
wire net_1018;
wire net_4089;
wire net_3629;
wire net_2854;
wire net_2009;
wire net_2369;
wire net_2038;
wire net_4132;
wire net_4026;
wire net_823;
wire net_4990;
wire net_106;
wire net_1380;
wire net_1676;
wire net_4788;
wire net_698;
wire net_1915;
wire net_5176;
wire net_1191;
wire net_5259;
wire net_4334;
wire net_2255;
wire net_4649;
wire net_4754;
wire net_2485;
wire net_3857;
wire net_1997;
wire net_138;
wire net_749;
wire net_1019;
wire net_1948;
wire net_1616;
wire net_1006;
wire net_2781;
wire net_4342;
wire net_2969;
wire net_1418;
wire net_3202;
wire net_4059;
wire net_2985;
wire net_537;
wire net_3056;
wire net_1713;
wire net_3614;
wire net_2668;
wire net_4684;
wire net_2677;
wire net_3252;
wire net_2775;
wire net_513;
wire x964;
wire net_3916;
wire net_163;
wire net_1576;
wire net_1421;
wire net_4496;
wire net_3407;
wire net_2736;
wire net_2127;
wire net_1280;
wire net_459;
wire net_3656;
wire net_737;
wire net_2284;
wire net_3412;
wire net_2113;
wire net_4793;
wire net_3990;
wire net_2193;
wire net_3856;
wire net_4760;
wire net_3915;
wire net_4885;
wire net_5258;
wire net_5201;
wire net_1886;
wire net_1156;
wire net_2604;
wire net_5150;
wire net_1966;
wire net_3501;
wire net_4571;
wire net_4678;
wire net_4866;
wire net_101;
wire net_1659;
wire net_1272;
wire net_326;
wire net_2381;
wire net_2109;
wire net_1770;
wire net_5059;
wire net_4001;
wire net_3505;
wire net_589;
wire net_655;
wire net_3536;
wire net_1814;
wire net_4703;
wire net_4770;
wire net_3175;
wire net_378;
wire net_2829;
wire net_724;
wire net_3309;
wire net_4815;
wire net_4099;
wire net_3142;
wire net_3036;
wire net_423;
wire net_1219;
wire net_4202;
wire net_328;
wire net_2384;
wire net_3884;
wire net_1958;
wire net_1931;
wire net_3736;
wire net_2877;
wire net_2480;
wire net_3294;
wire net_1549;
wire net_4477;
wire net_3016;
wire net_874;
wire net_2929;
wire net_1632;
wire net_3796;
wire net_1661;
wire net_1236;
wire net_4277;
wire net_818;
wire net_3749;
wire net_3674;
wire net_2746;
wire net_2700;
wire net_5024;
wire net_1211;
wire net_1183;
wire net_2594;
wire net_4248;
wire net_1488;
wire net_4966;
wire net_2812;
wire net_5244;
wire net_1684;
wire net_811;
wire net_352;
wire net_30;
wire net_3920;
wire net_1462;
wire net_436;
wire net_4674;
wire net_2837;
wire net_2017;
wire net_4993;
wire net_5154;
wire net_2824;
wire net_1777;
wire net_1926;
wire net_3115;
wire net_2735;
wire net_1641;
wire net_3518;
wire net_1621;
wire net_3680;
wire net_4919;
wire net_3984;
wire net_3615;
wire net_1702;
wire net_1103;
wire net_1035;
wire net_4403;
wire net_767;
wire net_3055;
wire net_1838;
wire x884;
wire net_4557;
wire net_131;
wire net_4656;
wire net_358;
wire net_1973;
wire net_3593;
wire net_3095;
wire net_2845;
wire net_4292;
wire net_2016;
wire net_4586;
wire net_2934;
wire net_2641;
wire net_1763;
wire net_4035;
wire net_3125;
wire net_1285;
wire net_3112;
wire net_1175;
wire net_2882;
wire net_3278;
wire net_4386;
wire net_2922;
wire net_1513;
wire net_1742;
wire net_3064;
wire net_2276;
wire net_4613;
wire net_468;
wire net_798;
wire net_5266;
wire net_3135;
wire net_73;
wire net_5165;
wire net_2059;
wire net_3370;
wire net_1899;
wire net_4746;
wire net_1336;
wire net_3947;
wire net_3441;
wire net_179;
wire net_4947;
wire net_61;
wire net_4015;
wire net_3662;
wire net_1843;
wire net_62;
wire net_3261;
wire net_534;
wire net_3793;
wire net_3336;
wire net_2289;
wire net_903;
wire net_1551;
wire net_486;
wire net_3539;
wire net_2031;
wire net_1868;
wire net_1560;
wire net_406;
wire net_4414;
wire net_4409;
wire net_4190;
wire net_2378;
wire net_3863;
wire net_3640;
wire net_3382;
wire net_4257;
wire net_1545;
wire net_748;
wire net_95;
wire net_4662;
wire net_4872;
wire net_990;
wire net_5281;
wire net_3958;
wire net_2327;
wire net_1003;
wire net_514;
wire net_2332;
wire net_3645;
wire net_3774;
wire net_1604;
wire net_2715;
wire net_1803;
wire net_1941;
wire net_524;
wire net_1134;
wire net_3899;
wire net_3742;
wire net_363;
wire net_4368;
wire net_445;
wire net_1319;
wire net_776;
wire net_4550;
wire net_3080;
wire net_2508;
wire net_44;
wire net_1650;
wire net_1582;
wire net_3748;
wire net_3149;
wire net_1675;
wire net_4016;
wire net_2247;
wire net_2333;
wire net_2213;
wire net_1368;
wire net_5067;
wire net_2575;
wire net_1248;
wire net_2291;
wire net_1097;
wire net_2238;
wire net_845;
wire net_762;
wire net_3589;
wire net_695;
wire net_4943;
wire net_2525;
wire net_1201;
wire net_3713;
wire net_556;
wire net_2671;
wire net_3330;
wire net_893;
wire net_4121;
wire net_255;
wire net_5106;
wire net_3826;
wire net_859;
wire net_620;
wire net_619;
wire net_1167;
wire net_4659;
wire net_3932;
wire net_4779;
wire net_2198;
wire net_1044;
wire net_5129;
wire net_5250;
wire net_4922;
wire net_3444;
wire net_4322;
wire net_3800;
wire net_2940;
wire net_2043;
wire net_2095;
wire net_4681;
wire net_3285;
wire net_5231;
wire net_4425;
wire net_4933;
wire net_68;
wire net_4044;
wire net_2314;
wire net_2613;
wire net_1493;
wire net_3605;
wire net_4630;
wire net_976;
wire net_4114;
wire net_2709;
wire net_865;
wire net_611;
wire net_231;
wire net_4179;
wire net_3514;
wire net_2621;
wire net_2579;
wire net_3024;
wire net_1223;
wire net_4691;
wire net_2750;
wire net_1866;
wire net_4907;
wire net_4107;
wire net_926;
wire net_4623;
wire net_3692;
wire net_3211;
wire net_2160;
wire net_3477;
wire net_4223;
wire net_391;
wire net_2297;
wire net_3325;
wire net_5040;
wire net_37;
wire net_2048;
wire net_582;
wire net_4481;
wire net_2341;
wire net_661;
wire net_4172;
wire net_3633;
wire net_3360;
wire net_2516;
wire net_2807;
wire net_4687;
wire net_1141;
wire net_3561;
wire net_4867;
wire net_3243;
wire net_1543;
wire net_1295;
wire x40;
wire net_2104;
wire net_1288;
wire net_2071;
wire net_1923;
wire x639;
wire net_4708;
wire net_1275;
wire net_210;
wire net_2766;
wire net_3771;
wire net_2417;
wire net_2300;
wire net_916;
wire net_3395;
wire net_741;
wire net_940;
wire net_4816;
wire net_4335;
wire net_851;
wire net_4411;
wire net_4857;
wire net_3719;
wire net_2426;
wire net_3789;
wire net_4937;
wire net_4199;
wire net_3310;
wire net_1043;
wire net_671;
wire x409;
wire net_2850;
wire net_770;
wire net_1005;
wire net_1059;
wire net_1630;
wire net_3891;
wire net_4918;
wire net_1454;
wire net_2956;
wire net_307;
wire net_1796;
wire net_1082;
wire net_3342;
wire net_5187;
wire net_3547;
wire net_1550;
wire net_3543;
wire net_2310;
wire net_1507;
wire net_5104;
wire net_3296;
wire net_257;
wire net_233;
wire net_474;
wire net_5138;
wire net_3459;
wire net_2656;
wire net_958;
wire net_4556;
wire net_1268;
wire net_3922;
wire net_3212;
wire net_3780;
wire net_4051;
wire net_1115;
wire net_944;
wire net_1734;
wire net_1764;
wire net_961;
wire net_3513;
wire net_4308;
wire net_4042;
wire net_2106;
wire net_3335;
wire net_3682;
wire net_5175;
wire net_4894;
wire net_3050;
wire net_1728;
wire net_63;
wire net_3327;
wire net_5091;
wire net_3956;
wire net_2667;
wire net_3456;
wire net_425;
wire net_287;
wire net_5204;
wire net_189;
wire net_4407;
wire net_1586;
wire net_2205;
wire net_3755;
wire net_480;
wire net_216;
wire net_4507;
wire net_4986;
wire net_2897;
wire x825;
wire net_433;
wire net_4443;
wire net_2881;
wire net_836;
wire net_2161;
wire net_4602;
wire net_368;
wire x105;
wire net_224;
wire net_4833;
wire net_52;
wire net_1898;
wire net_608;
wire net_1212;
wire net_3604;
wire net_370;
wire net_2000;
wire net_4383;
wire net_3706;
wire net_2984;
wire net_1120;
wire net_1020;
wire net_2848;
wire net_3282;
wire net_3122;
wire net_1169;
wire net_973;
wire net_1139;
wire net_3902;
wire net_2206;
wire net_1392;
wire net_1574;
wire net_2094;
wire net_4842;
wire net_2543;
wire net_311;
wire net_760;
wire net_2479;
wire net_2083;
wire net_3851;
wire net_873;
wire net_2488;
wire net_1811;
wire net_154;
wire net_3699;
wire net_4536;
wire net_4469;
wire net_5034;
wire net_2588;
wire net_1870;
wire net_5200;
wire net_704;
wire net_2520;
wire net_1478;
wire net_2179;
wire net_1696;
wire net_587;
wire net_1262;
wire net_2063;
wire net_3997;
wire net_4027;
wire net_192;
wire net_1739;
wire net_1356;
wire net_4505;
wire net_4213;
wire net_2912;
wire net_4393;
wire net_4140;
wire net_2197;
wire net_3816;
wire net_4131;
wire net_735;
wire net_2905;
wire net_1907;
wire net_3809;
wire net_1711;
wire net_200;
wire net_4435;
wire net_5220;
wire net_2084;
wire net_4164;
wire net_195;
wire net_5085;
wire net_1081;
wire net_1853;
wire net_2037;
wire net_2170;
wire net_1237;
wire net_1420;
wire net_4789;
wire net_2678;
wire net_4836;
wire net_4064;
wire net_4237;
wire net_4559;
wire net_3761;
wire net_3144;
wire net_699;
wire net_242;
wire net_359;
wire net_5239;
wire net_2526;
wire net_2819;
wire net_1644;
wire net_2864;
wire net_2800;
wire net_882;
wire net_1998;
wire net_1827;
wire net_4109;
wire net_3225;
wire net_1190;
wire net_3858;
wire net_2795;
wire net_1311;
wire net_4093;
wire net_4799;
wire net_2283;
wire net_1207;
wire net_1918;
wire net_2121;
wire net_2191;
wire net_3236;
wire net_3201;
wire net_3558;
wire net_2252;
wire net_555;
wire net_4755;
wire net_1613;
wire net_790;
wire net_2126;
wire net_5022;
wire net_1577;
wire net_1417;
wire net_4595;
wire net_1054;
wire x0;
wire net_2386;
wire net_2727;
wire net_2166;
wire net_3650;
wire net_2465;
wire net_5078;
wire net_2257;
wire net_3418;
wire net_3655;
wire net_2304;
wire net_898;
wire net_2968;
wire net_2643;
wire net_1593;
wire net_4416;
wire net_5015;
wire net_714;
wire net_2999;
wire net_1309;
wire net_3722;
wire net_3380;
wire net_683;
wire net_1771;
wire net_148;
wire net_1376;
wire net_5005;
wire net_4493;
wire net_1517;
wire net_5115;
wire net_4502;
wire net_1980;
wire x615;
wire net_1302;
wire net_2076;
wire net_244;
wire net_4378;
wire net_2218;
wire net_2395;
wire net_1690;
wire net_1078;
wire net_4002;
wire net_1989;
wire net_2997;
wire net_2855;
wire net_2093;
wire net_1795;
wire net_2403;
wire net_1539;
wire net_4261;
wire net_5197;
wire net_3490;
wire net_3035;
wire net_2355;
wire net_4357;
wire net_3262;
wire net_1548;
wire net_92;
wire net_394;
wire net_810;
wire net_3778;
wire net_2536;
wire net_1189;
wire net_139;
wire net_409;
wire net_2949;
wire net_3429;
wire net_1469;
wire net_3470;
wire net_4495;
wire net_4081;
wire net_88;
wire net_1708;
wire net_2436;
wire net_81;
wire net_4196;
wire net_3974;
wire net_4626;
wire net_3419;
wire net_2976;
wire net_722;
wire net_988;
wire net_1254;
wire net_3621;
wire net_5223;
wire net_621;
wire net_435;
wire net_1830;
wire net_5153;
wire net_4091;
wire net_132;
wire net_105;
wire net_5156;
wire net_2838;
wire net_1649;
wire net_1837;
wire net_5219;
wire net_1841;
wire net_1249;
wire net_4601;
wire net_2427;
wire net_3378;
wire net_1071;
wire net_3985;
wire net_3163;
wire net_5004;
wire net_4928;
wire net_4675;
wire net_327;
wire net_3877;
wire net_1701;
wire net_999;
wire net_4417;
wire net_353;
wire net_822;
wire net_1633;
wire net_5251;
wire net_4994;
wire net_3588;
wire net_1974;
wire net_1480;
wire net_319;
wire net_4963;
wire net_2670;
wire net_1743;
wire net_3046;
wire net_2597;
wire net_4952;
wire net_164;
wire net_377;
wire net_4702;
wire net_87;
wire net_1544;
wire net_288;
wire net_2649;
wire net_3096;
wire net_1629;
wire net_1459;
wire net_5265;
wire net_4400;
wire net_3277;
wire net_805;
wire net_4139;
wire net_3741;
wire net_3590;
wire net_4470;
wire net_2923;
wire net_2151;
wire net_540;
wire net_512;
wire net_2688;
wire net_2642;
wire net_1174;
wire net_1622;
wire net_891;
wire net_1109;
wire net_38;
wire net_5224;
wire net_3065;
wire net_3102;
wire net_4224;
wire net_5149;
wire net_3457;
wire net_4167;
wire net_4711;
wire net_5276;
wire net_4471;
wire net_1102;
wire net_4802;
wire net_4976;
wire net_5245;
wire net_3371;
wire net_618;
wire net_2244;
wire net_2692;
wire net_3688;
wire x368;
wire net_3777;
wire net_1875;
wire net_3420;
wire net_783;
wire net_3887;
wire net_1487;
wire net_4572;
wire net_754;
wire net_2759;
wire net_2605;
wire net_921;
wire net_3634;
wire net_550;
wire net_4957;
wire net_5238;
wire net_3308;
wire net_5178;
wire net_4543;
wire net_2835;
wire net_5086;
wire net_3991;
wire net_2192;
wire net_1533;
wire net_4871;
wire net_1240;
wire net_461;
wire net_3000;
wire net_3502;
wire net_2564;
wire net_2821;
wire net_1512;
wire net_1658;
wire net_4827;
wire net_654;
wire net_330;
wire net_858;
wire net_5025;
wire net_1330;
wire net_3506;
wire net_3007;
wire net_4275;
wire net_3015;
wire net_4487;
wire net_1785;
wire net_4766;
wire net_4771;
wire net_3174;
wire net_2876;
wire net_570;
wire net_444;
wire net_525;
wire net_844;
wire net_3829;
wire net_3646;
wire net_1496;
wire net_1210;
wire net_1067;
wire net_5058;
wire net_325;
wire net_3735;
wire net_1820;
wire net_5123;
wire net_1427;
wire net_5060;
wire net_3921;
wire net_4098;
wire net_4679;
wire net_985;
wire net_3933;
wire net_5014;
wire net_4036;
wire net_424;
wire net_1521;
wire net_4182;
wire net_1729;
wire net_3353;
wire net_1677;
wire x626;
wire net_4247;
wire net_4820;
wire net_4734;
wire net_2991;
wire net_4276;
wire net_564;
wire net_3639;
wire net_2050;
wire net_4086;
wire net_2811;
wire net_3086;
wire net_4585;
wire net_2058;
wire net_813;
wire net_3045;
wire net_1178;
wire net_4875;
wire net_2612;
wire net_1027;
wire net_2018;
wire net_3825;
wire net_5230;
wire net_2042;
wire net_340;
wire net_1408;
wire net_2510;
wire net_265;
wire net_2634;
wire net_434;
wire net_3808;
wire net_1797;
wire net_3488;
wire net_3023;
wire net_1202;
wire net_69;
wire net_1155;
wire net_4932;
wire net_4906;
wire net_4524;
wire net_925;
wire net_339;
wire net_2279;
wire net_3447;
wire net_3468;
wire net_4661;
wire net_2695;
wire net_864;
wire net_4113;
wire net_2710;
wire net_2660;
wire net_2298;
wire net_660;
wire net_3671;
wire net_102;
wire net_2313;
wire net_59;
wire net_3691;
wire net_1908;
wire net_3217;
wire net_4387;
wire net_1291;
wire net_230;
wire net_4214;
wire net_1865;
wire net_3383;
wire net_678;
wire net_5168;
wire net_3349;
wire net_4782;
wire net_1222;
wire net_3404;
wire net_928;
wire net_3810;
wire net_3914;
wire net_2578;
wire net_208;
wire net_2744;
wire net_2377;
wire net_1433;
wire net_415;
wire net_4739;
wire net_116;
wire net_4156;
wire net_3251;
wire net_2786;
wire net_347;
wire net_3794;
wire net_3440;
wire net_3358;
wire net_1776;
wire net_2145;
wire net_3368;
wire net_1335;
wire net_2574;
wire net_4014;
wire net_3311;
wire net_3531;
wire net_3747;
wire net_2212;
wire net_2132;
wire net_2292;
wire net_1880;
wire net_3862;
wire net_5103;
wire net_184;
wire net_3571;
wire net_4853;
wire net_4642;
wire net_610;
wire net_1844;
wire net_389;
wire net_3538;
wire net_902;
wire net_1867;
wire net_2344;
wire net_1323;
wire net_2650;
wire net_1949;
wire net_1506;
wire net_1583;
wire net_736;
wire net_1804;
wire net_539;
wire net_2331;
wire net_692;
wire net_4408;
wire net_1563;
wire net_5282;
wire net_4568;
wire net_4291;
wire net_3898;
wire net_4948;
wire net_4377;
wire net_3361;
wire net_1365;
wire net_1135;
wire net_5047;
wire net_1346;
wire net_43;
wire net_1942;
wire net_1801;
wire net_1400;
wire net_885;
wire net_1267;
wire net_3944;
wire net_3661;
wire net_4350;
wire net_4893;
wire net_869;
wire net_3714;
wire net_669;
wire net_937;
wire net_4077;
wire net_2441;
wire net_5131;
wire net_3517;
wire net_2349;
wire net_496;
wire net_761;
wire net_4749;
wire net_1554;
wire net_479;
wire net_1294;
wire net_2459;
wire net_2030;
wire net_3520;
wire net_1587;
wire net_5006;
wire net_1354;
wire net_4370;
wire net_4979;
wire net_2904;
wire net_796;
wire net_1308;
wire net_2249;
wire net_4332;
wire net_648;
wire net_1389;
wire net_739;
wire net_4748;
wire net_3250;
wire net_2548;
wire net_2075;
wire net_826;
wire net_1738;
wire net_3658;
wire net_548;
wire net_3359;
wire net_4985;
wire net_2402;
wire net_5082;
wire net_2624;
wire net_636;
wire net_343;
wire net_4269;
wire net_4795;
wire net_511;
wire net_3967;
wire net_4492;
wire net_1961;
wire net_5236;
wire net_4424;
wire net_1260;
wire net_4262;
wire net_4165;
wire net_2654;
wire net_2487;
wire net_4506;
wire net_2911;
wire net_1185;
wire net_1819;
wire net_5001;
wire net_239;
wire net_310;
wire net_2975;
wire net_4625;
wire net_2437;
wire net_5257;
wire net_2779;
wire net_4826;
wire net_1912;
wire net_1490;
wire net_4282;
wire net_682;
wire net_989;
wire net_1963;
wire net_1538;
wire net_108;
wire net_458;
wire net_4356;
wire net_685;
wire x388;
wire net_3560;
wire net_1007;
wire net_4052;
wire net_1579;
wire net_4772;
wire net_4616;
wire net_1292;
wire net_4786;
wire net_1999;
wire net_1014;
wire net_2796;
wire net_1444;
wire net_2679;
wire net_5016;
wire net_4024;
wire net_4686;
wire net_4082;
wire net_3410;
wire net_2111;
wire net_1946;
wire net_2733;
wire net_538;
wire net_3612;
wire net_4130;
wire net_1605;
wire net_1937;
wire net_2535;
wire net_3191;
wire net_366;
wire net_1854;
wire net_1956;
wire net_1917;
wire net_5118;
wire net_1614;
wire net_1755;
wire net_747;
wire net_1359;
wire net_2305;
wire net_1653;
wire net_2460;
wire net_2983;
wire net_3209;
wire net_4891;
wire net_2258;
wire net_198;
wire net_1647;
wire net_209;
wire net_4756;
wire net_1282;
wire net_5196;
wire net_294;
wire net_2367;
wire net_4573;
wire net_4127;
wire net_4041;
wire net_2892;
wire net_2810;
wire net_2429;
wire net_3204;
wire net_1265;
wire net_1053;
wire net_4444;
wire net_1004;
wire net_3471;
wire x232;
wire net_848;
wire net_4921;
wire net_1080;
wire net_1619;
wire net_3232;
wire net_2124;
wire net_1890;
wire net_4498;
wire net_3512;
wire net_1161;
wire net_4671;
wire x947;
wire net_82;
wire net_3228;
wire net_2282;
wire net_4501;
wire net_2430;
wire net_2357;
wire net_4461;
wire net_1395;
wire net_1546;
wire net_3481;
wire net_1589;
wire net_1046;
wire net_4363;
wire net_606;
wire net_4960;
wire net_3906;
wire net_623;
wire net_2396;
wire net_663;
wire net_1213;
wire net_1891;
wire net_2265;
wire net_5270;
wire net_5180;
wire net_3998;
wire net_579;
wire net_2445;
wire net_769;
wire net_3396;
wire net_1780;
wire net_2062;
wire net_2856;
wire net_787;
wire net_3603;
wire net_4511;
wire net_2894;
wire net_1025;
wire net_4187;
wire net_3758;
wire net_4834;
wire net_4067;
wire net_4717;
wire net_1988;
wire net_3718;
wire net_1518;
wire net_4618;
wire net_1089;
wire net_4419;
wire net_1194;
wire net_1437;
wire net_3579;
wire net_5284;
wire net_3525;
wire net_1664;
wire net_4528;
wire net_705;
wire net_2139;
wire net_1608;
wire net_4141;
wire net_506;
wire net_3769;
wire net_2948;
wire net_1910;
wire net_3775;
wire net_1036;
wire net_5146;
wire net_3544;
wire net_4537;
wire net_5229;
wire net_3034;
wire net_5096;
wire net_1196;
wire net_3973;
wire net_4394;
wire net_2493;
wire net_919;
wire net_3626;
wire net_290;
wire net_4008;
wire net_3313;
wire net_3136;
wire net_4726;
wire net_4090;
wire net_2209;
wire net_1372;
wire net_1757;
wire net_3834;
wire net_3591;
wire net_5215;
wire net_4436;
wire net_3152;
wire net_2682;
wire net_3648;
wire net_140;
wire net_740;
wire net_1722;
wire net_4072;
wire net_2329;
wire net_3790;
wire net_2150;
wire net_2008;
wire net_2065;
wire net_4267;
wire net_3183;
wire net_2927;
wire net_2808;
wire net_3908;
wire net_4856;
wire net_194;
wire net_4837;
wire net_2178;
wire net_730;
wire net_5292;
wire net_4150;
wire net_1128;
wire net_3073;
wire net_2713;
wire net_2105;
wire net_4707;
wire net_1127;
wire net_804;
wire net_1119;
wire net_3548;
wire net_1314;
wire net_957;
wire net_1287;
wire net_4312;
wire net_5299;
wire net_2726;
wire net_531;
wire net_4143;
wire net_77;
wire net_499;
wire net_3345;
wire net_2752;
wire net_49;
wire net_1340;
wire net_5140;
wire net_3123;
wire net_2955;
wire net_71;
wire net_3328;
wire net_771;
wire net_4390;
wire net_3534;
wire net_1765;
wire net_2844;
wire net_2301;
wire net_2978;
wire net_2107;
wire net_5185;
wire net_4852;
wire net_180;
wire net_3950;
wire net_4437;
wire net_51;
wire net_2774;
wire net_2420;
wire net_4028;
wire net_2860;
wire net_4367;
wire net_432;
wire net_4927;
wire net_1062;
wire net_1979;
wire net_5135;
wire net_3731;
wire net_3290;
wire net_4936;
wire net_3293;
wire x633;
wire net_1142;
wire net_1460;
wire net_1475;
wire net_1451;
wire net_4120;
wire net_3159;
wire net_67;
wire net_2240;
wire net_2416;
wire net_5065;
wire net_5008;
wire net_5188;
wire net_4803;
wire net_4590;
wire net_203;
wire net_1411;
wire net_2173;
wire net_505;
wire net_4088;
wire net_3723;
wire net_1602;
wire net_4013;
wire net_992;
wire net_237;
wire net_613;
wire net_782;
wire net_2144;
wire x593;
wire net_2236;
wire net_3744;
wire net_4635;
wire net_1095;
wire net_4729;
wire net_3443;
wire net_578;
wire net_4186;
wire net_4738;
wire net_3314;
wire net_3945;
wire net_2971;
wire net_4485;
wire net_1558;
wire net_2743;
wire net_2836;
wire net_1505;
wire net_4641;
wire net_1805;
wire net_2159;
wire net_388;
wire net_4667;
wire net_3952;
wire net_3669;
wire net_1861;
wire net_3647;
wire net_3635;
wire net_536;
wire net_4388;
wire net_455;
wire net_1332;
wire net_221;
wire net_1594;
wire net_115;
wire net_3339;
wire net_3276;
wire net_1110;
wire net_393;
wire net_442;
wire net_542;
wire x332;
wire net_408;
wire net_1832;
wire net_1026;
wire net_3246;
wire net_2215;
wire net_1845;
wire net_4562;
wire net_2573;
wire net_3087;
wire net_2376;
wire net_1520;
wire net_1821;
wire net_42;
wire net_3993;
wire net_3390;
wire net_1401;
wire net_3865;
wire net_2372;
wire net_1588;
wire net_3909;
wire net_66;
wire net_4037;
wire net_3937;
wire net_868;
wire net_1495;
wire net_2992;
wire net_3664;
wire net_5124;
wire net_3233;
wire net_443;
wire net_5029;
wire net_3522;
wire net_270;
wire net_522;
wire net_922;
wire net_2638;
wire net_668;
wire net_3079;
wire net_1584;
wire net_4992;
wire net_1990;
wire net_2330;
wire net_2264;
wire net_977;
wire net_4780;
wire net_643;
wire net_3397;
wire net_1070;
wire net_1225;
wire net_622;
wire net_812;
wire net_3587;
wire net_3762;
wire net_4391;
wire net_3687;
wire net_2857;
wire net_1107;
wire net_2767;
wire net_4920;
wire net_1338;
wire net_3874;
wire net_2045;
wire net_2053;
wire net_3384;
wire net_2180;
wire net_1203;
wire net_2869;
wire net_4242;
wire net_3332;
wire net_825;
wire net_3446;
wire net_1892;
wire net_1798;
wire net_4720;
wire net_4427;
wire net_3220;
wire net_2119;
wire net_309;
wire net_29;
wire net_1366;
wire net_837;
wire net_3469;
wire net_2615;
wire net_31;
wire net_927;
wire net_5143;
wire net_2007;
wire net_1151;
wire net_713;
wire net_5240;
wire net_693;
wire net_1519;
wire net_729;
wire net_4197;
wire net_3964;
wire net_3213;
wire net_2818;
wire net_863;
wire net_4219;
wire net_3164;
wire net_4173;
wire net_580;
wire net_2136;
wire net_904;
wire net_2339;
wire net_341;
wire net_4157;
wire net_58;
wire net_1879;
wire net_970;
wire net_488;
wire net_4909;
wire net_4941;
wire net_4221;
wire net_2319;
wire net_3044;
wire net_4845;
wire net_1532;
wire net_1160;
wire net_4475;
wire net_159;
wire net_3268;
wire net_2163;
wire net_3417;
wire net_3307;
wire net_4958;
wire net_553;
wire net_4887;
wire net_4212;
wire net_5057;
wire net_1093;
wire net_2592;
wire x128;
wire net_2875;
wire net_763;
wire net_3580;
wire net_3259;
wire net_5260;
wire net_4701;
wire net_1740;
wire net_324;
wire net_710;
wire net_462;
wire net_418;
wire net_872;
wire net_3097;
wire net_161;
wire net_5046;
wire net_3066;
wire net_3970;
wire net_3018;
wire net_2606;
wire net_173;
wire net_1486;
wire net_3880;
wire net_78;
wire net_2320;
wire net_1839;
wire net_1665;
wire net_4333;
wire net_4181;
wire net_3006;
wire net_376;
wire net_2133;
wire net_1681;
wire net_4817;
wire net_3550;
wire net_4880;
wire net_2515;
wire net_1812;
wire net_3173;
wire net_4825;
wire net_3738;
wire net_4138;
wire net_5298;
wire net_5119;
wire net_2224;
wire net_3203;
wire net_422;
wire net_4290;
wire net_4272;
wire net_1345;
wire net_1450;
wire net_561;
wire net_4899;
wire net_2659;
wire net_2589;
wire net_591;
wire net_1700;
wire net_746;
wire net_4299;
wire net_2290;
wire net_1274;
wire net_2458;
wire net_1682;
wire net_2851;
wire net_178;
wire net_3435;
wire net_2843;
wire net_3466;
wire net_2635;
wire net_5207;
wire net_3374;
wire net_3772;
wire net_4995;
wire net_3807;
wire net_4868;
wire net_2698;
wire net_809;
wire net_629;
wire net_1663;
wire net_3450;
wire net_635;
wire net_4279;
wire net_266;
wire net_1235;
wire net_2691;
wire net_1037;
wire net_3528;
wire net_4209;
wire net_2019;
wire net_4676;
wire net_350;
wire net_4270;
wire net_3019;
wire net_3460;
wire net_2351;
wire net_3117;
wire net_1350;
wire net_3482;
wire net_3198;
wire net_1626;
wire net_1648;
wire net_2822;
wire net_1258;
wire net_2982;
wire net_1623;
wire net_631;
wire net_4410;
wire net_3369;
wire net_1101;
wire net_994;
wire net_318;
wire net_3927;
wire net_4007;
wire net_1971;
wire net_4499;
wire net_4166;
wire net_2409;
wire net_4608;
wire net_3192;
wire net_1900;
wire net_1779;
wire net_2647;
wire net_5218;
wire net_670;
wire net_3340;
wire net_103;
wire net_4545;
wire net_3844;
wire net_2687;
wire net_1849;
wire net_228;
wire net_4737;
wire net_3554;
wire net_2640;
wire net_966;
wire net_4698;
wire net_3372;
wire net_4101;
wire net_1920;
wire net_2201;
wire net_3928;
wire net_1108;
wire net_2827;
wire net_2025;
wire net_2010;
wire net_3854;
wire net_2936;
wire net_1878;
wire net_4672;
wire net_755;
wire net_1723;
wire net_3890;
wire net_2900;
wire net_133;
wire net_5152;
wire net_4025;
wire net_4376;
wire net_3151;
wire net_3628;
wire net_2306;
wire net_4522;
wire net_3882;
wire net_3272;
wire net_2873;
wire net_557;
wire net_3043;
wire net_2254;
wire net_2861;
wire net_1652;
wire net_3652;
wire net_2669;
wire net_1429;
wire net_4083;
wire net_4574;
wire net_1611;
wire net_1991;
wire net_1173;
wire net_1209;
wire net_1431;
wire net_1754;
wire net_2725;
wire net_3613;
wire net_2328;
wire net_4615;
wire net_4038;
wire net_1714;
wire net_847;
wire net_727;
wire net_4787;
wire net_283;
wire net_5117;
wire net_4955;
wire net_3190;
wire net_4690;
wire net_240;
wire net_3757;
wire net_5020;
wire net_4445;
wire net_295;
wire net_344;
wire net_3951;
wire net_4757;
wire net_2269;
wire net_884;
wire net_712;
wire net_2281;
wire net_1422;
wire net_2259;
wire net_4497;
wire net_4462;
wire net_1106;
wire net_1394;
wire net_2963;
wire net_4095;
wire net_2972;
wire net_2739;
wire net_1281;
wire net_2110;
wire net_2463;
wire net_2919;
wire net_2893;
wire net_2241;
wire net_3227;
wire net_2358;
wire net_278;
wire net_3057;
wire net_1547;
wire net_4058;
wire net_4874;
wire net_571;
wire net_3509;
wire net_5122;
wire net_1162;
wire net_4935;
wire net_3934;
wire net_2443;
wire net_2472;
wire net_1307;
wire net_4514;
wire net_2790;
wire net_2742;
wire net_1877;
wire net_720;
wire net_5007;
wire net_4810;
wire net_5209;
wire net_5055;
wire net_2199;
wire net_4794;
wire net_4418;
wire net_3320;
wire net_4149;
wire net_2625;
wire net_684;
wire net_5221;
wire net_2648;
wire net_3657;
wire net_3720;
wire net_510;
wire net_1353;
wire net_1595;
wire net_114;
wire net_3581;
wire net_4049;
wire net_3776;
wire net_2653;
wire net_1300;
wire net_3432;
wire net_2974;
wire net_2960;
wire net_1252;
wire net_3895;
wire net_2734;
wire net_2782;
wire net_494;
wire net_547;
wire net_1098;
wire net_3146;
wire net_507;
wire net_1902;
wire net_238;
wire net_5237;
wire net_3074;
wire net_4283;
wire net_2438;
wire net_2600;
wire net_1911;
wire net_3022;
wire net_3563;
wire net_3461;
wire net_649;
wire net_4610;
wire net_4491;
wire net_1374;
wire net_4843;
wire net_4459;
wire net_457;
wire net_291;
wire net_1962;
wire net_2246;
wire net_772;
wire net_1964;
wire net_2494;
wire net_857;
wire net_867;
wire net_4371;
wire net_396;
wire net_3700;
wire net_107;
wire net_1277;
wire net_2661;
wire net_530;
wire net_1541;
wire net_3893;
wire net_5177;
wire net_4706;
wire net_594;
wire net_271;
wire net_3329;
wire net_673;
wire net_4268;
wire net_4075;
wire net_3611;
wire net_2064;
wire net_2797;
wire net_2852;
wire net_1721;
wire net_3846;
wire net_4633;
wire net_1925;
wire net_4402;
wire net_3549;
wire net_1445;
wire net_2074;
wire net_1909;
wire net_5256;
wire net_5274;
wire net_2577;
wire net_1410;
wire net_2954;
wire net_1073;
wire net_365;
wire net_3274;
wire net_1947;
wire net_3913;
wire net_3344;
wire net_2953;
wire net_141;
wire net_3787;
wire net_4413;
wire net_467;
wire net_879;
wire net_1810;
wire net_1118;
wire net_4313;
wire net_2910;
wire net_2415;
wire net_372;
wire net_4851;
wire net_2990;
wire net_2081;
wire net_5195;
wire x475;
wire net_4892;
wire net_803;
wire net_3165;
wire net_3595;
wire net_3197;
wire net_2788;
wire net_1348;
wire net_4965;
wire net_1476;
wire x23;
wire net_3489;
wire net_1293;
wire net_2883;
wire net_2302;
wire net_563;
wire net_1147;
wire net_3422;
wire net_199;
wire net_2789;
wire net_2681;
wire net_3835;
wire net_431;
wire net_2158;
wire net_5136;
wire net_4855;
wire net_4366;
wire net_5009;
wire net_1266;
wire net_3684;
wire net_5186;
wire net_2368;
wire net_1452;
wire net_2773;
wire net_2428;
wire net_909;
wire net_4529;
wire net_4362;
wire net_222;
wire net_4898;
wire net_152;
wire net_4520;
wire net_3105;
wire net_3999;
wire net_3966;
wire net_2895;
wire net_1788;
wire net_2138;
wire net_4301;
wire net_607;
wire net_258;
wire net_2477;
wire net_4142;
wire net_2935;
wire net_1045;
wire net_5083;
wire net_2446;
wire net_3497;
wire net_3905;
wire net_4345;
wire net_4188;
wire net_585;
wire net_4939;
wire net_3516;
wire net_3601;
wire net_4588;
wire net_4040;
wire net_1438;
wire net_4538;
wire net_4395;
wire net_3759;
wire net_3511;
wire net_374;
wire net_1143;
wire net_1987;
wire net_788;
wire x1012;
wire net_214;
wire net_3602;
wire net_249;
wire net_4527;
wire net_3578;
wire net_1088;
wire net_5283;
wire net_4716;
wire net_4144;
wire net_3885;
wire net_2079;
wire net_706;
wire net_1731;
wire net_2052;
wire net_4009;
wire net_5097;
wire net_2768;
wire net_5125;
wire net_4259;
wire net_2565;
wire net_2632;
wire net_551;
wire net_2547;
wire net_5076;
wire net_4617;
wire net_3636;
wire net_2118;
wire net_463;
wire net_4727;
wire net_2295;
wire net_5032;
wire net_1536;
wire net_1817;
wire net_197;
wire net_2560;
wire net_4168;
wire net_3478;
wire net_1498;
wire net_1381;
wire net_5017;
wire net_3709;
wire net_202;
wire net_1199;
wire net_3312;
wire net_1756;
wire net_2208;
wire net_3627;
wire net_2595;
wire net_1383;
wire net_2751;
wire net_918;
wire net_949;
wire net_4869;
wire net_450;
wire net_289;
wire net_4446;
wire net_4111;
wire net_2614;
wire net_1642;
wire net_1683;
wire net_978;
wire net_2524;
wire net_1313;
wire net_1129;
wire net_3331;
wire net_1056;
wire net_1224;
wire net_4908;
wire net_2296;
wire net_768;
wire net_3385;
wire net_4781;
wire net_357;
wire net_2044;
wire net_2181;
wire net_908;
wire net_1789;
wire net_3451;
wire net_519;
wire net_4530;
wire net_838;
wire net_3219;
wire net_2694;
wire net_3118;
wire net_2096;
wire net_4587;
wire net_2697;
wire net_4980;
wire net_2576;
wire net_3827;
wire net_2352;
wire net_1038;
wire net_1829;
wire net_4241;
wire net_1204;
wire net_2342;
wire net_3763;
wire net_3515;
wire net_5033;
wire net_662;
wire net_3214;
wire net_862;
wire net_1986;
wire net_50;
wire net_3398;
wire net_2277;
wire net_2307;
wire net_342;
wire x285;
wire net_975;
wire net_612;
wire net_4174;
wire net_4080;
wire net_738;
wire net_4325;
wire net_892;
wire net_4650;
wire net_4198;
wire net_1150;
wire net_504;
wire net_2006;
wire net_3406;
wire net_1331;
wire net_1537;
wire net_4229;
wire net_4074;
wire net_2130;
wire net_4000;
wire net_3362;
wire net_1148;
wire net_3120;
wire net_2214;
wire net_3338;
wire net_2382;
wire net_4504;
wire net_1561;
wire net_3442;
wire net_3864;
wire net_2728;
wire net_4636;
wire net_122;
wire net_417;
wire net_3269;
wire net_4421;
wire net_4092;
wire net_4389;
wire net_1940;
wire net_3337;
wire net_2662;
wire net_94;
wire net_3752;
wire net_4486;
wire net_4561;
wire net_482;
wire net_5144;
wire net_991;
wire net_3258;
wire net_3912;
wire net_149;
wire net_3088;
wire net_387;
wire net_1473;
wire net_4607;
wire net_3275;
wire net_2979;
wire net_2772;
wire net_41;
wire net_5291;
wire net_5160;
wire net_1893;
wire net_4180;
wire net_1674;
wire net_1932;
wire net_1651;
wire net_3836;
wire net_577;
wire net_3401;
wire net_2375;
wire net_5109;
wire net_1806;
wire net_3234;
wire net_2550;
wire net_797;
wire net_2347;
wire net_3545;
wire net_1957;
wire net_1363;
wire net_1799;
wire net_1869;
wire net_4053;
wire net_3806;
wire net_2684;
wire net_2572;
wire net_3972;
wire net_521;
wire net_60;
wire net_2414;
wire net_2754;
wire net_337;
wire net_267;
wire net_1585;
wire net_1846;
wire net_4476;
wire net_690;
wire net_4012;
wire net_3743;
wire net_3663;
wire net_523;
wire net_5110;
wire net_3260;
wire net_4254;
wire net_3681;
wire net_3815;
wire net_3555;
wire net_2716;
wire net_2371;
wire net_3375;
wire net_4926;
wire net_3467;
wire net_5246;
wire net_351;
wire net_4750;
wire net_4558;
wire net_4240;
wire net_4467;
wire net_3982;
wire net_1388;
wire net_2842;
wire net_5028;
wire net_4709;
wire net_3158;
wire net_2828;
wire net_1257;
wire net_939;
wire net_4721;
wire net_824;
wire net_3458;
wire net_3391;
wire net_1822;
wire net_2730;
wire net_4426;
wire net_1631;
wire net_1337;
wire net_1182;
wire net_4655;
wire net_1624;
wire net_2791;
wire net_1972;
wire net_1638;
wire net_1950;
wire net_3126;
wire net_993;
wire net_4271;
wire net_3875;
wire net_2421;
wire net_5268;
wire net_317;
wire net_856;
wire net_4901;
wire net_4804;
wire net_880;
wire net_1100;
wire net_1402;
wire net_2153;
wire net_3845;
wire net_1939;
wire net_4100;
wire net_2817;
wire net_3098;
wire net_2026;
wire net_4673;
wire net_5151;
wire net_2901;
wire net_162;
wire net_4950;
wire net_4944;
wire net_653;
wire net_1326;
wire net_3033;
wire net_5066;
wire net_134;
wire net_546;
wire net_4847;
wire net_4648;
wire net_3373;
wire net_3052;
wire net_4546;
wire net_2672;
wire net_3145;
wire net_588;
wire net_3694;
wire net_2200;
wire net_1157;
wire net_3701;
wire net_4736;
wire net_3855;
wire net_236;
wire net_487;
wire net_4974;
wire net_3883;
wire net_552;
wire net_1787;
wire net_1542;
wire net_1172;
wire net_3551;
wire net_5056;
wire net_4230;
wire net_756;
wire net_4765;
wire net_104;
wire net_1065;
wire net_5031;
wire net_4860;
wire net_2237;
wire net_3416;
wire net_72;
wire net_2566;
wire net_5166;
wire net_3953;
wire net_3795;
wire net_3100;
wire net_917;
wire net_241;
wire net_4886;
wire net_3730;
wire net_3537;
wire net_2874;
wire x142;
wire net_4597;
wire net_711;
wire net_599;
wire net_2225;
wire net_4589;
wire net_2993;
wire net_3067;
wire net_4844;
wire net_4288;
wire net_3111;
wire net_4741;
wire net_323;
wire net_963;
wire net_4700;
wire net_846;
wire net_3017;
wire net_4677;
wire net_3737;
wire net_4689;
wire net_153;
wire net_2389;
wire net_174;
wire net_2607;
wire net_562;
wire net_375;
wire net_364;
wire net_3172;
wire net_1831;
wire net_1482;
wire net_5023;
wire net_4239;
wire net_79;
wire net_3291;
wire net_2168;
wire net_3306;
wire net_2928;
wire net_2849;
wire net_1030;
wire net_1885;
wire net_4129;
wire net_1485;
wire x1023;
wire net_3245;
wire net_4873;
wire net_3171;
wire net_4298;
wire net_4773;
wire net_4201;
wire net_1247;
wire net_4273;
wire net_4137;
wire net_3673;
wire net_1969;
wire net_745;
wire net_5162;
wire net_2388;
wire net_933;
wire net_1244;
wire net_1215;
wire net_3496;
wire net_5169;
wire net_5248;
wire net_4216;
wire net_429;
wire net_129;
wire net_3377;
wire net_98;
wire net_373;
wire net_4889;
wire net_151;
wire net_356;
wire net_452;
wire net_1625;
wire net_545;
wire net_3683;
wire net_284;
wire net_1483;
wire net_2147;
wire net_560;
wire net_439;
wire net_3031;
wire net_259;
wire net_2513;
wire net_4094;
wire net_3351;
wire net_3582;
wire net_5148;
wire net_4603;
wire net_2645;
wire net_3119;
wire net_187;
wire net_1231;
wire net_3305;
wire net_4278;
wire net_2674;
wire net_160;
wire net_2872;
wire net_2432;
wire net_832;
wire net_322;
wire net_815;
wire net_1671;
wire net_4764;
wire net_420;
wire net_665;
wire net_1746;
wire net_2222;
wire net_2322;
wire net_2825;
wire net_586;
wire net_3670;
wire net_5272;
wire net_4344;
wire net_1347;
wire net_1091;
wire net_3341;
wire net_3838;
wire net_1072;
wire net_3745;
wire net_120;
wire net_4861;
wire net_292;
wire net_109;
wire net_1706;
wire net_4510;
wire net_3708;
wire net_3574;
wire net_96;
wire net_1730;
wire net_2921;
wire net_167;
wire net_3289;
wire net_5227;
wire net_4575;
wire net_651;
wire net_2931;
wire net_3114;
wire net_3415;
wire net_744;
wire net_4967;
wire net_598;
wire net_2556;
wire net_3519;
wire net_2740;
wire net_4136;
wire net_2806;
wire net_2011;
wire net_3455;
wire net_672;
wire net_4924;
wire net_777;
wire net_4806;
wire net_4818;
wire net_3157;
wire net_4483;
wire net_2820;
wire net_5212;
wire net_490;
wire net_2027;
wire net_5045;
wire net_4404;
wire net_3068;
wire net_3892;
wire net_2456;
wire net_2753;
wire net_3610;
wire net_1232;
wire net_3462;
wire net_4540;
wire net_1953;
wire net_3059;
wire net_632;
wire net_4439;
wire net_843;
wire net_3860;
wire net_3925;
wire net_464;
wire net_4473;
wire net_2841;
wire net_3847;
wire net_4582;
wire net_5089;
wire net_4200;
wire net_1977;
wire net_4547;
wire net_2100;
wire net_2938;
wire net_2122;
wire net_1171;
wire net_1540;
wire net_248;
wire net_3594;
wire net_4640;
wire net_4658;
wire net_1725;
wire net_3541;
wire net_1256;
wire net_802;
wire net_1413;
wire net_3532;
wire net_5112;
wire net_1767;
wire net_3556;
wire net_1840;
wire net_3041;
wire net_4010;
wire net_4997;
wire net_1640;
wire net_5190;
wire net_2724;
wire net_3427;
wire net_1031;
wire x606;
wire net_503;
wire net_1741;
wire net_4824;
wire net_4227;
wire net_1636;
wire net_1672;
wire net_2103;
wire net_996;
wire net_3091;
wire net_3257;
wire net_4458;
wire net_2994;
wire net_75;
wire net_959;
wire net_1334;
wire net_206;
wire net_757;
wire net_1688;
wire net_2020;
wire net_3051;
wire net_4004;
wire net_2345;
wire net_235;
wire net_2973;
wire net_3106;
wire net_2961;
wire net_5108;
wire net_4324;
wire net_4159;
wire net_2374;
wire net_2503;
wire net_4203;
wire net_2164;
wire x204;
wire net_3644;
wire net_250;
wire net_3600;
wire net_3081;
wire net_3751;
wire net_2055;
wire net_4879;
wire net_4564;
wire net_2630;
wire net_2338;
wire net_4606;
wire net_403;
wire net_1985;
wire net_3721;
wire net_2340;
wire net_3524;
wire net_32;
wire net_2616;
wire net_282;
wire net_1596;
wire net_2275;
wire net_4296;
wire net_3976;
wire net_5051;
wire net_841;
wire net_1750;
wire net_794;
wire net_2370;
wire net_2397;
wire net_2047;
wire net_3346;
wire net_2469;
wire net_2693;
wire net_528;
wire net_1012;
wire net_1404;
wire net_4878;
wire net_335;
wire net_3433;
wire net_907;
wire net_1468;
wire net_3464;
wire net_181;
wire net_4774;
wire net_3333;
wire net_39;
wire net_3076;
wire net_4694;
wire net_395;
wire net_2036;
wire net_2539;
wire net_3649;
wire net_1130;
wire net_2719;
wire net_386;
wire net_2323;
wire net_3867;
wire net_3677;
wire net_641;
wire net_4811;
wire net_1790;
wire net_4103;
wire net_2798;
wire net_5071;
wire net_4972;
wire net_3869;
wire net_1152;
wire net_1226;
wire net_2318;
wire net_3449;
wire net_4890;
wire net_1901;
wire net_3021;
wire net_1039;
wire net_3711;
wire net_1709;
wire net_3805;
wire net_4651;
wire net_400;
wire net_3942;
wire net_1935;
wire net_4580;
wire net_602;
wire net_2379;
wire net_175;
wire net_1818;
wire net_2918;
wire net_1850;
wire net_2925;
wire net_1497;
wire net_4429;
wire net_1800;
wire x450;
wire net_4634;
wire net_1855;
wire net_4882;
wire net_279;
wire net_1163;
wire net_1177;
wire net_1523;
wire net_1992;
wire net_3347;
wire net_897;
wire net_1656;
wire net_4039;
wire net_4030;
wire net_2853;
wire net_691;
wire net_2705;
wire net_5164;
wire net_615;
wire net_3273;
wire net_441;
wire net_1559;
wire net_3178;
wire net_2701;
wire net_4078;
wire net_1620;
wire net_1863;
wire net_2833;
wire net_2608;
wire net_2561;
wire net_2663;
wire net_2813;
wire net_728;
wire net_1276;
wire net_719;
wire net_170;
wire net_2519;
wire net_471;
wire net_1055;
wire net_2571;
wire net_3813;
wire net_878;
wire net_1531;
wire net_3894;
wire net_1159;
wire net_518;
wire net_861;
wire net_57;
wire net_3479;
wire net_3222;
wire net_929;
wire net_3321;
wire net_708;
wire net_2523;
wire net_3552;
wire net_4914;
wire net_696;
wire net_4210;
wire net_3954;
wire net_3216;
wire net_1565;
wire net_5262;
wire net_169;
wire net_171;
wire net_5213;
wire net_2234;
wire net_4552;
wire net_3821;
wire net_604;
wire net_967;
wire net_1527;
wire net_4503;
wire net_4420;
wire net_268;
wire net_4318;
wire net_3486;
wire net_48;
wire net_483;
wire net_3386;
wire net_4134;
wire net_4910;
wire net_1149;
wire net_1645;
wire net_2962;
wire net_4365;
wire net_176;
wire net_3638;
wire net_1298;
wire net_2570;
wire net_296;
wire net_2131;
wire net_3354;
wire net_614;
wire net_2712;
wire net_2005;
wire x350;
wire net_1123;
wire net_2771;
wire net_4897;
wire net_3194;
wire net_3572;
wire net_2228;
wire net_3020;
wire net_5141;
wire net_4740;
wire net_786;
wire net_1192;
wire net_4838;
wire net_127;
wire net_4542;
wire net_984;
wire net_1339;
wire net_3363;
wire net_3781;
wire net_4061;
wire net_1105;
wire net_906;
wire net_2172;
wire net_2422;
wire net_3156;
wire net_5205;
wire net_2482;
wire net_707;
wire net_3577;
wire x90;
wire net_652;
wire net_4457;
wire net_5039;
wire net_4361;
wire net_1815;
wire net_3840;
wire net_3782;
wire net_4850;
wire net_1856;
wire net_830;
wire net_4531;
wire net_575;
wire net_2505;
wire net_877;
wire net_1279;
wire net_1047;
wire net_2799;
wire net_4715;
wire net_3697;
wire net_3734;
wire net_4688;
wire net_2683;
wire net_2631;
wire net_4812;
wire net_4253;
wire net_2165;
wire net_3618;
wire net_4066;
wire net_3284;
wire net_4297;
wire net_1467;
wire net_1474;
wire net_1061;
wire net_2784;
wire net_3181;
wire net_765;
wire net_675;
wire net_1342;
wire net_2562;
wire net_2633;
wire net_2867;
wire net_5134;
wire net_1666;
wire net_5293;
wire net_3837;
wire net_3472;
wire net_4839;
wire net_2288;
wire net_4193;
wire net_2099;
wire net_5172;
wire net_1768;
wire net_2182;
wire net_5182;
wire net_4718;
wire net_150;
wire net_4351;
wire net_304;
wire net_4347;
wire net_2021;
wire net_1068;
wire net_1703;
wire net_186;
wire net_3983;
wire net_2495;
wire net_3693;
wire net_3814;
wire net_1050;
wire net_2072;
wire net_2760;
wire net_5100;
wire net_1316;
wire net_4751;
wire net_4319;
wire net_1872;
wire net_792;
wire net_2271;
wire net_3070;
wire net_3409;
wire net_4430;
wire net_2203;
wire net_4525;
wire net_1716;
wire net_1904;
wire net_5003;
wire net_3907;
wire net_1607;
wire net_5247;
wire net_219;
wire net_3609;
wire net_1263;
wire net_2187;
wire net_4591;
wire net_196;
wire net_2476;
wire net_3452;
wire net_913;
wire net_2067;
wire net_3130;
wire net_4518;
wire net_3387;
wire net_5183;
wire net_1479;
wire net_4330;
wire net_4019;
wire net_1639;
wire net_5267;
wire net_4152;
wire net_4126;
wire net_3094;
wire net_4289;
wire net_4549;
wire net_360;
wire net_1927;
wire net_3625;
wire net_213;
wire net_4145;
wire net_2324;
wire net_4712;
wire net_260;
wire net_4805;
wire net_947;
wire net_2947;
wire net_3137;
wire net_732;
wire net_1126;
wire net_2152;
wire net_2004;
wire net_1325;
wire net_3316;
wire net_3032;
wire net_5094;
wire net_5286;
wire net_1597;
wire net_1352;
wire net_1373;
wire net_2567;
wire net_2885;
wire net_2088;
wire net_4696;
wire net_1187;
wire net_4217;
wire net_2689;
wire net_3988;
wire net_4988;
wire net_2761;
wire net_3206;
wire net_1303;
wire net_3788;
wire net_4355;
wire net_2858;
wire net_1503;
wire net_3961;
wire net_2102;
wire net_4451;
wire net_4639;
wire net_1442;
wire net_449;
wire net_5234;
wire net_1807;
wire net_1930;
wire net_1943;
wire net_1087;
wire net_4234;
wire net_3995;
wire net_733;
wire net_887;
wire net_1894;
wire net_2431;
wire net_4054;
wire net_2308;
wire net_633;
wire net_5211;
wire net_113;
wire net_5054;
wire net_4731;
wire net_4848;
wire net_2989;
wire net_497;
wire net_1914;
wire net_4628;
wire net_40;
wire net_2770;
wire net_2408;
wire net_3889;
wire net_1424;
wire net_2636;
wire net_1414;
wire net_4375;
wire net_4153;
wire net_4412;
wire net_300;
wire net_3567;
wire net_2652;
wire net_1233;
wire net_1457;
wire net_2720;
wire net_2741;
wire net_4280;
wire net_1834;
wire net_950;
wire net_4011;
wire net_1436;
wire net_2448;
wire net_4925;
wire net_4338;
wire net_3400;
wire net_3392;
wire net_2551;
wire net_2816;
wire net_646;
wire net_2731;
wire net_1214;
wire net_2601;
wire net_3641;
wire net_866;
wire net_2891;
wire net_5194;
wire net_4220;
wire net_520;
wire net_3150;
wire net_4722;
wire net_1032;
wire net_567;
wire net_3726;
wire net_3979;
wire net_5255;
wire net_3231;
wire net_981;
wire net_272;
wire net_2401;
wire net_3939;
wire net_1024;
wire net_1566;
wire net_1590;
wire net_1305;
wire net_1612;
wire net_2354;
wire net_839;
wire net_1387;
wire net_814;
wire net_1581;
wire net_5018;
wire net_4468;
wire net_5013;
wire net_2413;
wire net_559;
wire net_4660;
wire net_345;
wire net_2792;
wire net_3042;
wire net_2128;
wire net_2965;
wire net_4785;
wire net_3930;
wire net_1717;
wire net_2586;
wire net_3299;
wire net_398;
wire net_1655;
wire net_3399;
wire net_954;
wire net_2365;
wire net_5080;
wire net_4565;
wire net_2117;
wire net_2461;
wire net_4085;
wire net_4797;
wire net_1766;
wire net_2582;
wire net_2361;
wire net_2598;
wire net_3872;
wire net_4956;
wire net_2879;
wire net_1572;
wire net_1680;
wire net_4447;
wire net_3302;
wire net_4790;
wire net_3187;
wire net_5179;
wire net_2134;
wire net_2622;
wire net_5011;
wire net_316;
wire net_4250;
wire net_84;
wire net_4961;
wire net_4184;
wire net_1759;
wire net_4900;
wire net_4647;
wire net_3764;
wire net_2262;
wire net_4022;
wire net_3011;
wire net_2087;
wire net_2541;
wire net_3689;
wire net_533;
wire net_1002;
wire net_1695;
wire net_911;
wire net_1617;
wire net_3188;
wire net_1993;
wire net_3010;
wire net_881;
wire net_2805;
wire net_1397;
wire net_2903;
wire net_4579;
wire net_568;
wire net_4474;
wire net_47;
wire net_4807;
wire net_1227;
wire x916;
wire net_1008;
wire net_4128;
wire x307;
wire net_4923;
wire net_1443;
wire net_1954;
wire net_3873;
wire net_4862;
wire net_3069;
wire net_3170;
wire net_2840;
wire net_3463;
wire net_2155;
wire net_4005;
wire net_168;
wire net_4819;
wire net_2041;
wire net_3199;
wire net_3597;
wire net_385;
wire net_5043;
wire net_269;
wire net_2609;
wire net_3193;
wire net_469;
wire net_3131;
wire net_5044;
wire net_1945;
wire net_1978;
wire net_3179;
wire net_5159;
wire net_4073;
wire net_3167;
wire net_1170;
wire net_1833;
wire net_2423;
wire net_2280;
wire net_2831;
wire net_3029;
wire net_778;
wire net_2366;
wire net_2380;
wire net_3393;
wire net_4548;
wire net_1455;
wire net_2930;
wire net_5064;
wire net_895;
wire net_5261;
wire net_4730;
wire net_1412;
wire net_4119;
wire net_1255;
wire net_1250;
wire net_3980;
wire net_1481;
wire net_995;
wire net_207;
wire net_3040;
wire net_3557;
wire net_3643;
wire net_5000;
wire net_700;
wire net_1246;
wire net_3004;
wire net_5216;
wire net_1689;
wire net_1774;
wire net_4228;
wire net_1673;
wire net_3060;
wire net_3830;
wire net_274;
wire net_2568;
wire net_3480;
wire net_321;
wire net_1075;
wire net_4135;
wire net_930;
wire net_833;
wire net_2387;
wire net_2995;
wire net_99;
wire net_3526;
wire net_2945;
wire net_4723;
wire net_2267;
wire net_934;
wire net_4758;
wire net_3103;
wire net_4249;
wire net_4769;
wire net_4896;
wire net_717;
wire net_544;
wire net_3665;
wire x956;
wire net_1399;
wire net_3630;
wire net_1824;
wire net_4888;
wire net_3350;
wire net_3402;
wire net_2223;
wire net_4763;
wire net_3553;
wire net_5074;
wire net_5161;
wire net_2673;
wire net_3500;
wire net_3166;
wire net_3304;
wire net_1245;
wire net_2549;
wire net_860;
wire net_1781;
wire net_3660;
wire net_3465;
wire net_870;
wire net_2046;
wire net_3049;
wire net_637;
wire net_2878;
wire net_2514;
wire net_2871;
wire net_2390;
wire net_3267;
wire net_2321;
wire net_4775;
wire net_2686;
wire net_3474;
wire net_2013;
wire net_817;
wire net_1509;
wire net_529;
wire net_5127;
wire net_3414;
wire net_3495;
wire net_97;
wire net_2028;
wire net_2553;
wire net_4881;
wire net_1889;
wire net_3766;
wire net_4576;
wire net_1591;
wire net_2920;
wire net_2981;
wire net_1747;
wire net_650;
wire net_1164;
wire net_2012;
wire net_121;
wire net_597;
wire net_5228;
wire net_743;
wire net_3770;
wire net_1922;
wire net_2583;
wire net_3820;
wire net_3799;
wire net_4175;
wire net_4665;
wire net_2664;
wire net_2706;
wire net_5163;
wire net_849;
wire net_603;
wire net_4913;
wire net_5294;
wire net_2451;
wire net_2602;
wire net_642;
wire net_401;
wire net_1522;
wire net_2699;
wire net_4031;
wire net_4484;
wire net_1158;
wire net_3798;
wire net_2714;
wire net_2926;
wire net_2183;
wire net_2557;
wire net_440;
wire net_758;
wire net_470;
wire net_2702;
wire net_430;
wire net_4652;
wire net_2834;
wire net_4551;
wire net_718;
wire net_83;
wire net_3943;
wire net_3129;
wire net_4998;
wire net_4438;
wire net_56;
wire net_3255;
wire net_4218;
wire net_1063;
wire net_4448;
wire net_968;
wire net_336;
wire net_1578;
wire net_2534;
wire net_4133;
wire net_2917;
wire net_3221;
wire net_1504;
wire net_697;
wire net_475;
wire net_2003;
wire net_3732;
wire net_605;
wire net_3411;
wire net_5053;
wire net_4987;
wire net_2309;
wire net_502;
wire net_2470;
wire net_1564;
wire net_3426;
wire net_1568;
wire net_3804;
wire net_5095;
wire net_924;
wire net_1526;
wire net_1884;
wire net_1333;
wire net_3919;
wire net_2348;
wire net_4112;
wire net_489;
wire net_5107;
wire net_2646;
wire net_3082;
wire net_3868;
wire net_3936;
wire net_3676;
wire net_4364;
wire net_4185;
wire net_4646;
wire net_4204;
wire net_2628;
wire net_4512;
wire net_2748;
wire net_5145;
wire net_251;
wire net_1360;
wire net_2054;
wire net_3364;
wire net_664;
wire net_128;
wire net_840;
wire net_1364;
wire net_5050;
wire net_4622;
wire net_827;
wire net_549;
wire net_4605;
wire net_2793;
wire net_4295;
wire net_411;
wire net_2137;
wire net_1836;
wire net_4563;
wire net_4310;
wire net_2337;
wire net_1369;
wire net_3430;
wire net_1862;
wire net_2317;
wire net_4695;
wire net_4244;
wire net_1013;
wire net_1530;
wire net_3075;
wire net_3583;
wire net_842;
wire net_112;
wire net_2952;
wire net_4396;
wire net_1705;
wire net_2336;
wire net_2035;
wire net_2373;
wire net_5070;
wire net_2826;
wire net_2398;
wire net_3739;
wire net_4581;
wire net_492;
wire net_3678;
wire net_4431;
wire net_2141;
wire net_2639;
wire net_3315;
wire net_2455;
wire net_1609;
wire net_402;
wire net_3453;
wire net_3695;
wire net_1327;
wire net_3448;
wire net_4047;
wire net_110;
wire net_4968;
wire net_33;
wire net_1403;
wire net_4532;
wire net_3248;
wire net_2248;
wire net_2270;
wire net_2274;
wire net_4971;
wire net_1667;
wire net_3866;
wire net_1386;
wire net_1606;
wire net_3710;
wire net_2359;
wire net_3054;
wire net_4300;
wire net_5101;
wire net_4776;
wire net_3978;
wire net_4102;
wire net_4752;
wire net_2186;
wire net_3696;
wire net_3473;
wire net_1430;
wire net_2029;
wire net_2868;
wire net_569;
wire net_2478;
wire net_3698;
wire net_2563;
wire net_4629;
wire net_2946;
wire net_2587;
wire net_4397;
wire net_1284;
wire net_3408;
wire net_4870;
wire net_630;
wire net_76;
wire net_2959;
wire net_2202;
wire net_1888;
wire net_2490;
wire net_4311;
wire net_4018;
wire net_3929;
wire net_4428;
wire net_1791;
wire net_4339;
wire net_1471;
wire net_1792;
wire net_2496;
wire net_4125;
wire net_3109;
wire net_2066;
wire net_3608;
wire net_1598;
wire net_3124;
wire net_1903;
wire net_2407;
wire net_731;
wire net_1146;
wire net_912;
wire net_4612;
wire net_4519;
wire net_1733;
wire net_4517;
wire net_2078;
wire net_779;
wire net_1928;
wire net_3841;
wire net_1328;
wire net_234;
wire net_2859;
wire net_4151;
wire net_2884;
wire net_3848;
wire net_5142;
wire net_4942;
wire net_2762;
wire net_3205;
wire net_4146;
wire net_1094;
wire net_3487;
wire net_2749;
wire net_855;
wire net_1724;
wire net_674;
wire net_3703;
wire net_4619;
wire net_303;
wire net_2089;
wire net_491;
wire net_2475;
wire net_965;
wire net_3797;
wire net_1299;
wire net_948;
wire net_2937;
wire net_3535;
wire net_1195;
wire net_2916;
wire net_421;
wire net_4743;
wire net_1396;
wire net_2502;
wire net_1104;
wire net_4069;
wire net_764;
wire net_876;
wire net_2593;
wire net_4060;
wire net_5181;
wire net_2162;
wire net_2737;
wire net_2439;
wire net_5126;
wire net_172;
wire net_5038;
wire net_4341;
wire net_2481;
wire net_4539;
wire net_1117;
wire net_1458;
wire net_4048;
wire net_4570;
wire net_3955;
wire net_905;
wire net_1060;
wire net_2617;
wire net_142;
wire net_4846;
wire net_2229;
wire net_2235;
wire net_158;
wire net_1715;
wire net_3200;
wire net_3733;
wire net_3881;
wire net_2080;
wire net_3675;
wire net_2711;
wire net_2097;
wire net_2504;
wire net_3619;
wire net_1216;
wire net_2175;
wire net_3784;
wire net_4599;
wire net_2815;
wire net_3785;
wire net_1086;
wire net_1271;
wire net_2116;
wire net_1758;
wire net_4327;
wire net_1782;
wire net_1769;
wire net_1197;
wire net_1967;
wire net_4863;
wire net_273;
wire net_1278;
wire net_5171;
wire net_1567;
wire net_4714;
wire net_576;
wire net_3182;
wire net_1654;
wire net_2098;
wire net_465;
wire net_4232;
wire net_177;
wire net_3355;
wire net_4305;
wire net_3005;
wire net_1883;
wire net_476;
wire net_2783;
wire net_2803;
wire net_382;
wire net_3058;
wire net_3301;
wire net_725;
wire net_3931;
wire net_583;
wire net_1315;
wire net_953;
wire net_894;
wire net_1074;
wire net_1058;
wire net_5208;
wire net_5019;
wire net_1423;
wire net_1871;
wire net_2902;
wire net_4719;
wire net_4977;
wire net_517;
wire net_628;
wire net_5075;
wire net_4460;
wire net_2489;
wire net_3494;
wire net_220;
wire net_1465;
wire net_293;
wire net_3666;
wire net_4982;
wire net_1938;
wire net_543;
wire net_3160;
wire net_625;
wire net_2125;
wire net_3760;
wire net_1823;
wire net_5081;
wire net_1289;
wire net_3138;
wire net_2623;
wire net_191;
wire net_261;
wire net_3576;
wire net_4331;
wire net_2909;
wire net_4953;
wire net_558;
wire net_2069;
wire net_2362;
wire net_4697;
wire net_1618;
wire net_4456;
wire net_4354;
wire net_2497;
wire net_5111;
wire net_1955;
wire net_2723;
wire net_5157;
wire net_2552;
wire net_3562;
wire net_1001;
wire net_3229;
wire net_781;
wire net_1694;
wire net_3765;
wire net_4991;
wire net_910;
wire net_5241;
wire net_3012;
wire net_3754;
wire net_2412;
wire net_185;
wire net_4023;
wire net_4265;
wire net_3989;
wire net_4450;
wire net_4158;
wire net_5285;
wire net_4631;
wire net_4321;
wire net_1984;
wire net_1994;
wire net_315;
wire net_1015;
wire net_1375;
wire net_4670;
wire net_2980;
wire net_1944;
wire net_4668;
wire net_4006;
wire net_1351;
wire net_3897;
wire net_1775;
wire net_3960;
wire net_4374;
wire net_91;
wire net_297;
wire net_346;
wire net_1535;
wire net_2400;
wire net_3992;
wire net_2287;
wire net_4211;
wire net_448;
wire net_2034;
wire net_886;
wire net_229;
wire net_3189;
wire net_4360;
wire net_4962;
wire net_1808;
wire x60;
wire net_2146;
wire net_2988;
wire net_3256;
wire net_687;
wire net_405;
wire net_3266;
wire net_4592;
wire net_4160;
wire net_1111;
wire net_4281;
wire net_2651;
wire net_5279;
wire net_3888;
wire net_3651;
wire net_3971;
wire net_3155;
wire net_3322;
wire net_2533;
wire net_1470;
wire net_3566;
wire net_4627;
wire net_4423;
wire net_1913;
wire net_4728;
wire net_831;
wire net_3596;
wire net_451;
wire net_5021;
wire net_4233;
wire net_750;
wire net_1234;
wire net_4796;
wire net_1760;
wire net_1184;
wire net_4055;
wire net_2778;
wire net_2756;
wire net_3926;
wire net_4849;
wire net_3403;
wire net_1085;
wire net_1960;
wire net_5184;
wire net_592;
wire net_3093;
wire net_647;
wire net_3247;
wire net_4759;
wire net_773;
wire net_2266;
wire net_2464;
wire net_281;
wire net_4256;
wire net_828;
wire net_3839;
wire net_4490;
wire net_1603;
wire net_2732;
wire net_5254;
wire net_5193;
wire net_5235;
wire net_3521;
wire net_1096;
wire net_795;
wire x800;
wire net_3727;
wire net_982;
wire net_5052;
wire net_1580;
wire net_1406;
wire net_54;
wire net_5287;
wire net_4205;
wire net_3896;
wire net_526;
wire net_4384;
wire net_2718;
wire net_834;
wire net_694;
wire net_1434;
wire net_2747;
wire net_3668;
wire net_4912;
wire net_5130;
wire net_1570;
wire net_974;
wire net_4946;
wire net_4645;
wire net_774;
wire net_923;
wire net_5049;
wire net_1707;
wire net_4566;
wire net_2190;
wire net_1881;
wire net_501;
wire net_111;
wire net_3679;
wire net_225;
wire net_4489;
wire net_252;
wire net_124;
wire net_3128;
wire net_3323;
wire net_4733;
wire net_2399;
wire net_4692;
wire net_901;
wire net_447;
wire net_871;
wire net_2611;
wire net_3425;
wire net_410;
wire net_1492;
wire net_390;
wire net_35;
wire net_1154;
wire net_4243;
wire net_2537;
wire net_4294;
wire net_3767;
wire net_5128;
wire net_80;
wire net_4105;
wire net_4106;
wire net_2951;
wire net_2603;
wire net_3631;
wire net_1132;
wire net_2442;
wire net_4569;
wire net_2293;
wire net_280;
wire net_3026;
wire net_495;
wire net_34;
wire net_1802;
wire net_2140;
wire net_2356;
wire net_971;
wire net_3288;
wire net_2049;
wire net_2273;
wire net_617;
wire net_2517;
wire net_2316;
wire net_2184;
wire net_554;
wire net_4176;
wire net_2755;
wire net_4653;
wire net_3740;
wire net_1678;
wire net_2703;
wire net_46;
wire net_4032;
wire net_4154;
wire net_3366;
wire net_584;
wire net_1441;
wire net_969;
wire net_1525;
wire net_2411;
wire net_3870;
wire net_165;
wire net_821;
wire net_4003;
wire net_3438;
wire net_4177;
wire net_3824;
wire net_4440;
wire net_3436;
wire net_2335;
wire net_3940;
wire net_384;
wire net_3911;
wire net_3823;
wire net_4191;
wire net_2618;
wire net_3503;
wire net_4316;
wire net_3365;
wire net_3859;
wire net_2599;
wire net_2665;
wire net_3642;
wire net_1114;
wire net_2707;
wire net_3803;
wire net_3388;
wire net_1748;
wire net_485;
wire net_4116;
wire net_3078;
wire net_3218;
wire net_4632;
wire net_2964;
wire net_3334;
wire net_3224;
wire net_64;
wire net_1719;
wire net_2232;
wire net_2343;
wire net_726;
wire net_3811;
wire net_1028;
wire net_1529;
wire net_600;
wire net_3237;
wire net_701;
wire net_125;
wire net_397;
wire net_808;
wire net_1704;
wire net_1685;
wire net_2440;
wire net_5026;
wire net_4821;
wire net_1384;
wire net_4768;
wire net_2738;
wire net_1379;
wire net_3918;
wire net_5280;
wire net_320;
wire net_4916;
wire net_1322;
wire net_2644;
wire net_2944;
wire net_1301;
wire net_986;
wire net_1242;
wire net_286;
wire net_4346;
wire net_1241;
wire net_3690;
wire net_3584;
wire net_935;
wire net_4999;
wire net_3001;
wire net_1511;
wire net_3116;
wire net_645;
wire net_426;
wire net_3121;
wire net_5203;
wire net_4841;
wire net_4621;
wire net_4340;
wire net_4071;
wire net_4954;
wire net_1634;
wire net_609;
wire net_414;
wire net_1048;
wire net_3048;
wire net_5102;
wire net_799;
wire net_3083;
wire net_3475;
wire net_4533;
wire net_1816;
wire net_2014;
wire net_1221;
wire net_4195;
wire net_1951;
wire net_4895;
wire net_331;
wire net_816;
wire net_4644;
wire net_3264;
wire net_2092;
wire net_2558;
wire net_4742;
wire net_2454;
wire net_2040;
wire net_2220;
wire net_4762;
wire net_2823;
wire net_1217;
wire net_1508;
wire net_3379;
wire net_4761;
wire net_2933;
wire net_931;
wire net_3728;
wire net_3381;
wire net_4466;
wire net_2242;
wire net_4118;
wire net_4577;
wire net_759;
wire net_4970;
wire net_1575;
wire net_4884;
wire net_3279;
wire net_657;
wire net_5042;
wire net_1727;
wire net_247;
wire net_329;
wire net_4600;
wire net_4753;
wire net_1259;
wire net_1924;
wire net_4225;
wire net_2143;
wire net_2839;
wire net_5242;
wire net_4287;
wire net_1825;
wire net_2196;
wire net_3791;
wire net_70;
wire net_3168;
wire net_3413;
wire net_5275;
wire net_1341;
wire net_962;
wire net_4541;
wire net_478;
wire net_5210;
wire net_1934;
wire x179;
wire net_3242;
wire net_1835;
wire net_596;
wire net_1848;
wire net_1261;
wire net_333;
wire net_4724;
wire net_639;
wire net_4959;
wire net_2120;
wire net_1975;
wire net_4705;
wire net_1238;
wire net_4664;
wire net_565;
wire net_2569;
wire net_2832;
wire net_4478;
wire net_1033;
wire net_2149;
wire net_3028;
wire net_3923;
wire net_2554;
wire net_1692;
wire net_4479;
wire net_5079;
wire net_2528;
wire net_2655;
wire net_5062;
wire net_3107;
wire net_4236;
wire net_1686;
wire net_1361;
wire net_367;
wire net_3303;
wire net_2450;
wire net_4813;
wire net_1842;
wire net_1208;
wire net_204;
wire net_232;
wire net_3957;
wire net_1180;
wire net_4596;
wire net_1627;
wire net_2002;
wire net_1069;
wire net_2022;
wire net_2167;
wire net_2880;
wire net_2385;
wire net_4710;
wire net_4808;
wire net_2996;
wire net_2889;
wire net_3431;
wire net_4544;
wire net_3565;
wire net_1416;
wire net_137;
wire net_3154;
wire net_4828;
wire net_2433;
wire net_4465;
wire net_532;
wire net_2501;
wire net_3530;
wire net_3622;
wire net_4029;
wire net_1601;
wire net_93;
wire net_1916;
wire net_2729;
wire net_4422;
wire net_2468;
wire net_302;
wire net_4087;
wire net_4255;
wire net_1131;
wire net_889;
wire net_1116;
wire net_348;
wire net_753;
wire net_626;
wire net_5253;
wire net_4373;
wire net_5068;
wire net_1809;
wire net_100;
wire net_686;
wire net_2195;
wire net_1615;
wire net_3421;
wire net_2814;
wire net_1691;
wire net_689;
wire net_751;
wire net_4155;
wire net_4578;
wire net_2112;
wire net_5072;
wire net_595;
wire net_2363;
wire net_1320;
wire net_1828;
wire net_1466;
wire net_3659;
wire net_5232;
wire net_5192;
wire net_157;
wire net_3724;
wire net_1710;
wire net_1228;
wire net_1205;
wire net_4593;
wire net_466;
wire net_4336;
wire net_1179;
wire net_2722;
wire net_4161;
wire net_1426;
wire net_3039;
wire net_2217;
wire net_1407;
wire net_938;
wire net_3147;
wire net_4903;
wire net_1761;
wire net_1610;
wire net_3569;
wire net_4683;
wire net_183;
wire net_3263;
wire net_4246;
wire net_1440;
wire net_4020;
wire net_1057;
wire net_2915;
wire net_4453;
wire net_1011;
wire net_1355;
wire net_800;
wire net_644;
wire net_5225;
wire net_4931;
wire net_852;
wire net_2987;
wire net_4046;
wire net_2253;
wire net_2580;
wire net_1699;
wire net_5114;
wire net_4398;
wire net_1042;
wire net_4783;
wire net_4076;
wire net_4792;
wire net_1643;
wire net_1385;
wire net_1919;
wire net_1534;
wire net_1000;
wire net_1995;
wire net_2521;
wire net_2545;
wire net_1016;
wire net_4876;
wire net_5158;
wire net_659;
wire net_3977;
wire net_4567;
wire net_1744;
wire net_899;
wire net_1010;
wire net_516;
wire net_1693;
wire net_2870;
wire net_3176;
wire net_3654;
wire net_3585;
wire net_3779;
wire net_956;
wire net_4320;
wire net_4252;
wire net_2908;
wire net_3963;
wire net_2068;
wire net_4981;
wire net_2596;
wire net_3705;
wire net_2970;
wire net_4449;
wire net_438;
wire net_2675;
wire net_2794;
wire net_2584;
wire net_1752;
wire net_314;
wire net_2250;
wire net_2527;
wire net_5278;
wire net_3013;
wire net_952;
wire net_3110;
wire net_2091;
wire net_2967;
wire net_2406;
wire net_4097;
wire net_5170;
wire net_3185;
wire net_4669;
wire net_807;
wire net_3300;
wire net_3405;
wire net_86;
wire net_3270;
wire net_2245;
wire net_4286;
wire net_3484;
wire net_2474;
wire net_945;
wire net_4380;
wire net_2530;
wire net_4231;
wire net_2101;
wire net_383;
wire net_4068;
wire net_3570;
wire net_217;
wire net_3140;
wire net_427;
wire net_135;
wire net_2785;
wire net_915;
wire net_1121;
wire net_2226;
wire net_3849;
wire net_473;
wire x423;
wire net_3599;
wire net_5099;
wire net_4329;
wire net_2777;
wire net_1049;
wire net_454;
wire net_3901;
wire net_5174;
wire x256;
wire net_1784;
wire net_1296;
wire net_709;
wire net_2484;
wire net_4326;
wire net_2863;
wire net_3507;
wire net_5199;
wire net_1165;
wire net_1066;
wire net_5167;
wire net_677;
wire net_1472;
wire net_2939;
wire net_1113;
wire net_2424;
wire net_1968;
wire net_2591;
wire net_4304;
wire net_5189;
wire net_4560;
wire net_1344;
wire net_4488;
wire net_1283;
wire net_1084;
wire net_3968;
wire net_5295;
wire net_5092;
wire net_4554;
wire net_1500;
wire net_354;
wire net_2507;
wire net_1136;
wire net_5120;
wire net_3008;
wire net_2685;
wire net_2763;
wire net_573;
wire net_2658;
wire net_2898;
wire net_1391;
wire net_2174;
wire net_5132;
wire net_784;
wire net_3356;
wire net_1772;
wire net_3529;
wire net_45;
wire net_3616;
wire net_381;
wire net_2498;
wire net_3886;
wire net_2326;
wire net_1592;
wire net_3540;
wire net_2085;
wire net_3783;
wire net_5037;
wire net_3672;
wire net_4406;
wire net_1857;
wire net_1637;
wire net_3702;
wire net_1318;
wire net_3238;
wire net_941;
wire net_55;
wire net_1557;
wire net_1514;
wire net_3852;
wire net_3092;
wire net_4555;
wire net_4349;
wire net_2070;
wire net_2311;
wire net_3575;
wire net_4611;
wire net_4124;
wire net_1599;
wire net_4984;
wire net_306;
wire net_4516;
wire net_3828;
wire net_3981;
wire net_3132;
wire net_3161;
wire net_4303;
wire net_1290;
wire net_5061;
wire net_4147;
wire net_500;
wire net_1906;
wire net_3053;
wire net_2610;
wire net_4056;
wire net_4432;
wire net_3297;
wire net_2023;
wire net_4584;
wire net_4523;
wire net_1329;
wire net_123;
wire net_5249;
wire net_1668;
wire net_527;
wire net_262;
wire net_362;
wire net_3424;
wire net_3127;
wire net_1052;
wire net_3139;
wire net_4063;
wire net_3831;
wire net_5087;
wire net_1793;
wire net_3104;
wire net_3786;
wire net_4401;
wire net_2189;
wire net_3632;
wire net_2057;
wire net_2278;
wire net_4859;
wire net_3072;
wire net_1124;
wire net_226;
wire net_1021;
wire net_5269;
wire net_1737;
wire net_143;
wire net_1859;
wire net_4964;
wire net_190;
wire net_2887;
wire net_1447;
wire net_4207;
wire net_145;
wire net_1929;
wire net_3607;
wire net_4654;
wire net_1983;
wire net_4917;
wire net_1145;
wire net_2061;
wire net_3030;
wire net_3493;
wire net_5288;
wire net_4637;
wire net_2804;
wire net_2261;
wire net_3842;
wire net_4266;
wire net_188;
wire net_1553;
wire net_3753;
wire net_1895;
wire net_3061;
wire net_509;
wire net_3319;
wire net_4975;
wire net_4353;
wire net_211;
wire net_2491;
wire net_2958;
wire net_1077;
wire net_3208;
wire net_2704;
wire net_2924;
wire net_2410;
wire net_3910;
wire net_1851;
wire net_3941;
wire net_119;
wire net_3108;
wire net_2185;
wire net_1321;
wire net_2233;
wire net_3445;
wire net_2941;
wire net_4441;
wire net_2033;
wire net_477;
wire net_3348;
wire net_4192;
wire net_2123;
wire net_4949;
wire net_1099;
wire net_2943;
wire net_3861;
wire net_2532;
wire net_90;
wire net_2315;
wire net_4583;
wire net_85;
wire net_2231;
wire net_1864;
wire net_404;
wire net_3812;
wire net_1200;
wire net_4663;
wire net_2518;
wire net_2666;
wire net_4084;
wire net_4500;
wire net_4062;
wire net_1239;
wire net_1463;
wire net_1646;
wire net_4115;
wire net_2056;
wire net_2776;
wire net_3389;
wire net_3437;
wire net_1562;
wire net_3822;
wire net_472;
wire net_2522;
wire net_4178;
wire net_1628;
wire net_1510;
wire net_65;
wire net_3476;
wire net_3077;
wire net_484;
wire net_896;
wire net_4823;
wire net_2512;
wire net_4829;
wire net_3223;
wire net_136;
wire net_1936;
wire net_1524;
wire net_4171;
wire net_3802;
wire net_1528;
wire net_126;
wire net_2708;
wire net_1749;
wire net_3367;
wire net_4915;
wire net_2211;
wire net_4784;
wire net_601;
wire net_1362;
wire net_1896;
wire net_4385;
wire net_2346;
wire net_1982;
wire net_1732;
wire net_829;
wire net_2511;
wire net_2626;
wire net_4110;
wire net_2115;
wire net_2294;
wire net_4317;
wire net_2299;
wire net_4978;
wire net_2393;
wire net_3917;
wire net_3376;
wire net_900;
wire net_1405;
wire net_3253;
wire net_1882;
wire net_413;
wire net_2001;
wire net_1491;
wire net_716;
wire net_5147;
wire net_1269;
wire net_2419;
wire net_3750;
wire net_1034;
wire net_3533;
wire net_3715;
wire net_36;
wire net_2696;
wire net_253;
wire net_276;
wire net_1449;
wire net_4293;
wire net_3439;
wire net_666;
wire net_1959;
wire net_4809;
wire net_616;
wire net_1220;
wire net_4693;
wire net_4017;
wire net_3946;
wire net_1847;
wire net_2717;
wire net_793;
wire net_1657;
wire net_460;
wire net_3084;
wire net_4945;
wire net_2353;
wire net_2272;
wire net_4206;
wire net_2334;
wire net_1367;
wire net_3994;
wire net_1133;
wire net_4104;
wire net_3287;
wire net_166;
wire net_1976;
wire net_2866;
wire net_3169;
wire net_3025;
wire net_4079;
wire net_3871;
wire net_3792;
wire net_4455;
wire net_1371;
wire net_2758;
wire net_3352;
wire net_117;
wire net_74;
wire net_5002;
wire net_1826;
wire net_3832;
wire net_205;
wire net_1286;
wire net_4609;
wire net_4704;
wire net_2142;
wire net_920;
wire net_1952;
wire net_334;
wire net_1461;
wire net_2453;
wire net_3009;
wire net_3062;
wire net_4226;
wire net_820;
wire net_3177;
wire net_4620;
wire net_380;
wire net_2847;
wire x672;
wire net_1556;
wire net_4337;
wire net_3768;
wire net_4745;
wire net_437;
wire net_1270;
wire net_3573;
wire net_4905;
wire net_2286;
wire net_566;
wire net_1552;
wire net_5063;
wire net_4940;
wire net_3878;
wire net_624;
wire net_2148;
wire net_4735;
wire net_3215;
wire net_1933;
wire net_298;
wire net_2108;
wire net_3717;
wire net_2529;
wire net_688;
wire net_4685;
wire net_3241;
wire net_998;
wire net_4732;
wire net_4657;
wire net_2157;
wire net_2555;
wire net_4864;
wire net_3504;
wire net_3027;
wire net_2405;
wire net_1687;
wire net_835;
wire net_5243;
wire net_1762;
wire net_4235;
wire net_4096;
wire net_1181;
wire net_4117;
wire x437;
wire net_1357;
wire net_638;
wire net_5214;
wire net_4822;
wire net_3986;
wire net_3637;
wire x557;
wire net_313;
wire net_932;
wire x160;
wire net_1243;
wire net_1660;
wire net_1484;
wire net_4767;
wire net_4604;
wire net_1783;
wire net_5271;
wire net_3667;
wire net_419;
wire net_1874;
wire net_1635;
wire net_972;
wire net_5027;
wire net_4840;
wire net_936;
wire net_819;
wire net_3499;
wire net_5206;
wire net_4725;
wire net_4777;
wire net_4070;
wire net_785;
wire net_3002;
wire net_1489;
wire net_854;
wire net_2619;
wire net_4343;
wire net_4215;
wire net_3141;
wire net_1670;
wire net_2221;
wire net_3746;
wire net_4274;
wire net_1349;
wire net_2801;
wire net_3265;
wire net_5264;
wire net_979;
wire net_2392;
wire net_2932;
wire net_4951;
wire net_156;
wire net_2015;
wire net_1264;
wire net_1040;
wire net_5202;
wire net_4643;
wire net_4877;
wire net_1745;
wire net_332;
wire net_4170;
wire net_1679;
wire net_3089;
wire net_3101;
wire net_4883;
wire net_3037;
wire net_3148;
wire net_4472;
wire net_1229;
wire net_656;
wire net_4800;
wire net_4463;
wire net_3876;
wire net_766;
wire net_2907;
wire net_3686;
wire net_1153;
wire net_1887;
wire net_3014;
wire net_4284;
wire net_379;
wire net_2243;
wire net_1569;
wire net_4033;
wire net_3113;
wire net_4245;
wire x856;
wire net_3454;
wire net_3133;
wire net_3047;
wire net_2559;
wire net_5113;
wire net_3969;
wire net_2657;
wire net_1358;
wire net_3729;
wire net_2629;
wire net_2486;
wire net_2251;
wire net_1698;
wire net_1017;
wire net_955;
wire net_1206;
wire net_2585;
wire net_3653;
wire net_1996;
wire net_960;
wire net_3704;
wire net_1166;
wire net_1029;
wire net_801;
wire net_412;
wire net_2620;
wire net_1718;
wire net_2581;
wire net_5093;
wire net_4798;
wire net_2986;
wire net_3162;
wire net_4791;
wire net_4348;
wire net_4034;
wire net_4526;
wire net_1873;
wire net_2129;
wire net_3801;
wire net_453;
wire net_581;
wire net_2899;
wire net_3510;
wire net_3180;
wire net_658;
wire net_3249;
wire net_2263;
wire net_734;
wire net_3624;
wire net_2544;
wire net_2090;
wire net_2325;
wire net_951;
wire net_2086;
wire net_4930;
wire net_806;
wire net_3186;
wire net_4021;
wire net_946;
wire net_1176;
wire net_5277;
wire net_2676;
wire net_2966;
wire net_4372;
wire net_1253;
wire net_4989;
wire net_2194;
wire net_2500;
wire net_1076;
wire net_3900;
wire net_1751;
wire net_5010;
wire net_3559;
wire net_4682;
wire net_4352;
wire net_681;
wire net_3153;
wire net_3508;
wire net_5155;
wire net_2434;
wire net_3564;
wire net_1448;
wire net_2032;
wire net_392;
wire net_118;
wire net_3598;
wire net_5252;
wire net_2467;
wire net_146;
wire net_2452;
wire net_3938;
wire net_3523;
wire net_4594;
wire net_4162;
wire net_3712;
wire net_1502;
wire net_4454;
wire net_4624;
wire net_428;
wire net_246;
wire net_1186;
wire net_4747;
wire net_640;
wire net_4666;
wire net_2216;
wire net_2888;
wire net_775;
wire net_1378;
wire net_752;
wire net_1773;
wire net_3773;
wire net_1600;
wire net_2531;
wire net_498;
wire net_535;
wire net_888;
wire net_3716;
wire net_676;
wire net_5191;
wire net_4263;
wire net_2721;
wire x762;
wire net_2637;
wire net_5233;
wire net_5073;
wire net_4814;
wire net_1023;
wire net_2538;
wire net_4452;
wire net_2447;
wire net_3623;
wire net_5133;
wire net_4902;
wire net_301;
wire net_2360;
wire net_3617;
wire net_299;
wire net_1343;
wire net_2285;
wire net_4260;
wire net_3492;
wire net_182;
wire net_2462;
wire net_4359;
wire net_590;
wire net_3879;
wire net_2024;
wire net_3240;
wire net_3324;
wire net_3254;
wire net_3725;
wire net_4194;
wire net_5041;
wire net_1435;
wire net_1370;
wire net_407;
wire net_3568;
wire net_1736;
wire net_3207;
wire net_4482;
wire net_4405;
wire net_2204;
wire net_5088;
wire net_2492;
wire net_2312;
wire net_4148;
wire net_1970;
wire net_5048;
wire net_1306;
wire net_4045;
wire net_1669;
wire net_3843;
wire net_1858;
wire net_1041;
wire net_2073;
wire net_3038;
wire net_2690;
wire net_2950;
wire net_3924;
wire net_5226;
wire net_4057;
wire net_791;
wire net_5105;
wire net_1419;
wire net_3239;
wire net_4778;
wire net_2188;
wire net_1051;
wire net_2364;
wire net_942;
wire net_1981;
wire net_4302;
wire net_1515;
wire net_1218;
wire net_1573;
wire net_4983;
wire net_1494;
wire x974;
wire net_4415;
wire net_361;
wire net_3286;
wire net_2890;
wire net_2154;
wire net_1726;
wire net_305;
wire net_4123;
wire net_4208;
wire net_4515;
wire net_1905;
wire net_1398;
wire net_2540;
wire net_3099;
wire net_3298;
wire net_1125;
wire net_2230;
wire net_227;
wire net_144;
wire net_4183;
wire net_4399;
wire net_1144;
wire net_1794;
wire net_3592;
wire net_4969;
wire net_4638;
wire net_1022;
wire net_1415;
wire net_3485;
wire net_2260;
wire net_2865;
wire net_3606;
wire net_2886;
wire net_3317;
wire net_1921;
wire net_702;
wire net_4328;
wire net_1477;
wire net_3195;
wire net_3210;
wire net_3853;
wire net_3318;
wire net_1230;
wire net_2135;
wire net_667;
wire net_853;
wire net_212;
wire net_914;
wire net_1193;
wire net_1425;
wire net_1122;
wire net_875;
wire net_4911;
wire net_1813;
wire net_4534;
wire net_1092;
wire net_627;
wire net_2039;
wire net_983;
wire net_355;
wire net_4713;
wire net_4307;
wire net_1456;
wire net_723;
wire net_2227;
wire net_2483;
wire net_2473;
wire net_3962;
wire net_4553;
wire net_275;
wire net_399;
wire net_5069;
wire net_4831;
wire net_2914;
wire net_1390;
wire net_218;
wire net_2590;
wire net_1112;
wire net_5173;
wire net_1273;
wire net_3283;
wire net_1137;
wire net_4433;
wire net_3948;
wire net_2114;
wire net_2506;
wire net_4830;
wire net_5012;
wire net_5036;
wire net_3230;
wire net_4865;
wire net_285;
wire net_5296;
wire net_1310;
wire net_3819;
wire net_254;
wire net_2499;
wire net_1501;
wire net_1297;
wire net_3003;
wire net_1304;
wire net_4381;
wire net_574;
wire net_2177;
wire net_3357;

// Start cells
NAND2_X2 inst_1783 ( .A1(net_1202), .A2(net_1117), .ZN(net_1062) );
CLKBUF_X2 inst_5101 ( .A(net_4473), .Z(net_5087) );
CLKBUF_X2 inst_4728 ( .A(net_4713), .Z(net_4714) );
CLKBUF_X2 inst_4385 ( .A(net_4370), .Z(net_4371) );
INV_X2 inst_2685 ( .ZN(net_1804), .A(net_1753) );
OAI21_X2 inst_481 ( .B1(net_2970), .ZN(net_2964), .B2(net_2963), .A(net_2458) );
AND2_X4 inst_4123 ( .ZN(net_4047), .A1(net_2551), .A2(net_2003) );
NAND2_X2 inst_1751 ( .ZN(net_1382), .A1(net_1228), .A2(net_321) );
CLKBUF_X2 inst_4606 ( .A(net_4591), .Z(net_4592) );
INV_X4 inst_2235 ( .ZN(net_1863), .A(net_1814) );
OAI211_X2 inst_779 ( .C1(net_3424), .A(net_3422), .ZN(net_2862), .B(net_2736), .C2(net_1351) );
CLKBUF_X2 inst_5306 ( .A(net_4455), .Z(net_5292) );
INV_X4 inst_2205 ( .ZN(net_2254), .A(net_2233) );
INV_X2 inst_2858 ( .ZN(net_330), .A(net_64) );
AND2_X4 inst_4131 ( .ZN(net_4060), .A2(net_1192), .A1(net_1188) );
OAI21_X4 inst_452 ( .B1(net_3808), .ZN(net_2790), .B2(net_2529), .A(net_2366) );
OR2_X4 inst_214 ( .ZN(net_2597), .A1(net_2212), .A2(net_742) );
INV_X2 inst_3061 ( .ZN(net_4175), .A(net_2703) );
CLKBUF_X2 inst_4228 ( .A(net_4204), .Z(net_4214) );
OAI21_X2 inst_548 ( .B2(net_2909), .B1(net_2887), .ZN(net_2883), .A(net_2466) );
AND2_X4 inst_4144 ( .ZN(net_4080), .A1(net_3627), .A2(net_246) );
CLKBUF_X2 inst_4647 ( .A(net_4632), .Z(net_4633) );
CLKBUF_X2 inst_4372 ( .A(net_4274), .Z(net_4358) );
OAI21_X2 inst_728 ( .ZN(net_713), .B2(net_587), .B1(net_584), .A(net_421) );
DFF_X2 inst_3121 ( .Q(net_3147), .D(net_2728), .CK(net_4589) );
INV_X2 inst_2780 ( .ZN(net_806), .A(net_760) );
INV_X4 inst_2485 ( .A(net_3072), .ZN(net_470) );
CLKBUF_X2 inst_4709 ( .A(net_4694), .Z(net_4695) );
AND2_X4 inst_4152 ( .A2(net_4117), .ZN(net_4100), .A1(net_1699) );
INV_X4 inst_2217 ( .ZN(net_2096), .A(net_1973) );
OAI211_X2 inst_850 ( .ZN(net_633), .B(net_632), .C1(net_449), .A(net_387), .C2(net_254) );
DFF_X1 inst_3347 ( .D(net_2756), .CK(net_4344), .Q(x79) );
DFF_X2 inst_3130 ( .D(net_3535), .QN(net_3468), .CK(net_4815) );
INV_X2 inst_2844 ( .ZN(net_388), .A(net_376) );
INV_X4 inst_2492 ( .A(net_3061), .ZN(net_735) );
AND2_X4 inst_4136 ( .ZN(net_4065), .A2(net_1586), .A1(net_1063) );
AOI22_X2 inst_3582 ( .A1(net_4063), .B1(net_4058), .B2(net_4015), .A2(net_4013), .ZN(net_1435) );
NAND4_X2 inst_1228 ( .A1(net_4111), .ZN(net_791), .A3(net_775), .A4(net_527), .A2(net_403) );
AOI22_X2 inst_3480 ( .A1(net_2675), .ZN(net_2658), .B1(net_2657), .A2(net_991), .B2(net_225) );
CLKBUF_X2 inst_4985 ( .A(net_4970), .Z(net_4971) );
CLKBUF_X2 inst_4221 ( .A(net_4206), .Z(net_4207) );
OAI21_X2 inst_521 ( .B1(net_3302), .ZN(net_2918), .B2(net_2917), .A(net_2394) );
CLKBUF_X2 inst_5164 ( .A(net_5149), .Z(net_5150) );
CLKBUF_X2 inst_4473 ( .A(net_4458), .Z(net_4459) );
NAND2_X2 inst_1685 ( .A1(net_3219), .ZN(net_1987), .A2(net_558) );
INV_X4 inst_2511 ( .A(net_3062), .ZN(net_478) );
INV_X4 inst_2438 ( .A(net_3145), .ZN(net_137) );
NAND2_X2 inst_1655 ( .A1(net_2590), .ZN(net_2185), .A2(net_2003) );
AOI22_X2 inst_3578 ( .A1(net_4060), .B1(net_4055), .ZN(net_1472), .A2(net_234), .B2(net_169) );
INV_X2 inst_2772 ( .ZN(net_861), .A(net_860) );
INV_X4 inst_2543 ( .ZN(net_3753), .A(net_3675) );
OR2_X4 inst_237 ( .ZN(net_3413), .A2(net_1126), .A1(net_1124) );
CLKBUF_X2 inst_4847 ( .A(net_4832), .Z(net_4833) );
CLKBUF_X2 inst_4818 ( .A(net_4803), .Z(net_4804) );
OAI211_X2 inst_813 ( .B(net_1628), .C1(net_1627), .ZN(net_1625), .A(net_1553), .C2(net_334) );
XNOR2_X2 inst_51 ( .A(net_3552), .ZN(net_2618), .B(net_1693) );
NAND2_X2 inst_1837 ( .ZN(net_1200), .A1(net_722), .A2(net_721) );
NOR2_X2 inst_1066 ( .A2(net_3732), .ZN(net_896), .A1(net_853) );
NOR2_X4 inst_974 ( .ZN(net_3933), .A2(net_3932), .A1(net_3722) );
DFF_X1 inst_3392 ( .D(net_1633), .CK(net_5255), .Q(x615) );
CLKBUF_X2 inst_5063 ( .A(net_4726), .Z(net_5049) );
INV_X4 inst_2342 ( .ZN(net_1717), .A(net_1381) );
CLKBUF_X2 inst_4608 ( .A(net_4564), .Z(net_4594) );
DFF_X1 inst_3291 ( .QN(net_3013), .D(net_2889), .CK(net_5224) );
INV_X4 inst_2294 ( .A(net_3723), .ZN(net_1015) );
NAND2_X2 inst_1617 ( .A1(net_2919), .ZN(net_2399), .A2(net_140) );
SDFF_X2 inst_151 ( .D(net_3611), .SE(net_2625), .SI(net_101), .Q(net_101), .CK(net_4938) );
XNOR2_X2 inst_64 ( .ZN(net_1787), .B(net_1765), .A(net_1618) );
INV_X4 inst_2256 ( .ZN(net_1211), .A(net_1156) );
NOR2_X2 inst_1001 ( .A2(net_4050), .A1(net_3504), .ZN(net_2126) );
CLKBUF_X2 inst_4821 ( .A(net_4806), .Z(net_4807) );
AND4_X4 inst_4051 ( .ZN(net_4104), .A1(net_3766), .A2(net_618), .A3(net_607), .A4(net_385) );
MUX2_X2 inst_2106 ( .S(net_2915), .A(net_2573), .Z(net_2571), .B(net_201) );
OAI21_X2 inst_743 ( .B2(net_4052), .B1(net_3694), .ZN(net_3310), .A(net_1560) );
INV_X2 inst_2723 ( .ZN(net_1504), .A(net_1503) );
AOI21_X4 inst_3931 ( .B2(net_3757), .ZN(net_3726), .A(net_3725), .B1(net_3403) );
INV_X2 inst_3033 ( .A(net_3764), .ZN(net_3565) );
CLKBUF_X2 inst_4880 ( .A(net_4865), .Z(net_4866) );
INV_X2 inst_2925 ( .A(net_3094), .ZN(net_196) );
CLKBUF_X2 inst_4265 ( .A(net_4207), .Z(net_4251) );
AOI221_X2 inst_3867 ( .B2(net_3119), .B1(net_2020), .C1(net_2019), .ZN(net_1940), .A(net_1939), .C2(x256) );
NAND2_X2 inst_1828 ( .A1(net_912), .ZN(net_828), .A2(net_526) );
NAND2_X2 inst_2072 ( .ZN(net_3990), .A2(net_3988), .A1(net_963) );
NAND2_X2 inst_1603 ( .A1(net_2969), .ZN(net_2414), .A2(net_468) );
NAND2_X2 inst_1809 ( .A2(net_1213), .ZN(net_950), .A1(net_901) );
OAI22_X2 inst_340 ( .ZN(net_3256), .A2(net_3255), .A1(net_1712), .B1(net_1711), .B2(net_1710) );
DFF_X1 inst_3388 ( .D(net_1756), .QN(net_79), .CK(net_4250) );
AOI222_X2 inst_3735 ( .B1(net_3386), .C2(net_3385), .A1(net_3384), .A2(net_1826), .ZN(net_1764), .C1(net_574), .B2(net_361) );
CLKBUF_X2 inst_5311 ( .A(net_4805), .Z(net_5297) );
INV_X2 inst_2675 ( .ZN(net_1897), .A(net_1860) );
CLKBUF_X2 inst_4280 ( .A(net_4265), .Z(net_4266) );
OR4_X2 inst_158 ( .ZN(net_2712), .A1(net_2711), .A2(net_2710), .A3(net_2709), .A4(net_50) );
SDFF_X2 inst_141 ( .SE(net_2625), .D(net_2315), .SI(net_99), .Q(net_99), .CK(net_4750) );
CLKBUF_X2 inst_4344 ( .A(net_4329), .Z(net_4330) );
INV_X4 inst_2520 ( .ZN(net_3225), .A(net_2874) );
CLKBUF_X2 inst_4244 ( .A(net_4229), .Z(net_4230) );
NAND2_X2 inst_1490 ( .A1(net_4150), .A2(net_3600), .ZN(net_2860) );
OAI21_X2 inst_507 ( .B1(net_3274), .B2(net_2969), .ZN(net_2935), .A(net_2415) );
OAI21_X2 inst_571 ( .B2(net_3428), .ZN(net_2834), .B1(net_2762), .A(net_2116) );
AOI21_X1 inst_4011 ( .ZN(net_3304), .A(net_1601), .B2(net_1600), .B1(net_64) );
CLKBUF_X2 inst_4559 ( .A(net_4544), .Z(net_4545) );
CLKBUF_X2 inst_4289 ( .A(net_4274), .Z(net_4275) );
AOI22_X2 inst_3709 ( .B2(net_4124), .A2(net_555), .ZN(net_455), .A1(net_454), .B1(net_453) );
NAND2_X2 inst_1974 ( .A1(net_3666), .ZN(net_3346), .A2(net_767) );
NAND2_X2 inst_2017 ( .A2(net_4023), .ZN(net_3649), .A1(net_3647) );
NOR3_X2 inst_884 ( .A1(net_4154), .A3(net_3175), .ZN(net_2757), .A2(net_2688) );
NOR2_X2 inst_1154 ( .ZN(net_4001), .A2(net_4000), .A1(net_3728) );
OAI21_X2 inst_711 ( .ZN(net_958), .B1(net_843), .A(net_842), .B2(net_408) );
OAI211_X2 inst_827 ( .ZN(net_1453), .A(net_1313), .B(net_1193), .C1(net_1076), .C2(net_399) );
OAI21_X2 inst_469 ( .B1(net_3509), .ZN(net_2981), .B2(net_2969), .A(net_2417) );
INV_X2 inst_3040 ( .ZN(net_3657), .A(net_3655) );
INV_X2 inst_2980 ( .A(net_3006), .ZN(net_222) );
CLKBUF_X2 inst_5197 ( .A(net_5140), .Z(net_5183) );
AND2_X4 inst_4191 ( .ZN(net_4195), .A1(net_4137), .A2(net_42) );
AOI221_X2 inst_3870 ( .B2(net_3114), .B1(net_2020), .C1(net_2019), .ZN(net_1935), .A(net_1934), .C2(x160) );
CLKBUF_X2 inst_4269 ( .A(net_4254), .Z(net_4255) );
CLKBUF_X2 inst_4640 ( .A(net_4549), .Z(net_4626) );
XOR2_X2 inst_18 ( .Z(net_3553), .B(net_3551), .A(net_1692) );
NOR3_X2 inst_915 ( .A2(net_3821), .A1(net_3674), .ZN(net_3604), .A3(net_3171) );
AND2_X4 inst_4128 ( .ZN(net_4055), .A2(net_1247), .A1(net_1192) );
CLKBUF_X2 inst_4416 ( .A(net_4401), .Z(net_4402) );
INV_X4 inst_2263 ( .ZN(net_1283), .A(net_1165) );
INV_X4 inst_2339 ( .ZN(net_963), .A(net_716) );
CLKBUF_X2 inst_4861 ( .A(net_4846), .Z(net_4847) );
CLKBUF_X2 inst_4796 ( .A(net_4781), .Z(net_4782) );
CLKBUF_X2 inst_5183 ( .A(net_4225), .Z(net_5169) );
AOI22_X2 inst_3549 ( .B1(net_4054), .A2(net_2037), .A1(net_1578), .ZN(net_1572), .B2(net_182) );
AOI22_X2 inst_3501 ( .ZN(net_2065), .A1(net_2063), .B1(net_1904), .B2(net_1401), .A2(net_1400) );
NAND4_X2 inst_1216 ( .ZN(net_1099), .A4(net_879), .A3(net_547), .A2(net_501), .A1(net_460) );
AOI21_X2 inst_3936 ( .B1(net_3882), .B2(net_3858), .A(net_2529), .ZN(net_2344) );
CLKBUF_X2 inst_4807 ( .A(net_4792), .Z(net_4793) );
NOR2_X4 inst_952 ( .ZN(net_3662), .A1(net_3106), .A2(net_283) );
AND2_X4 inst_4175 ( .ZN(net_4129), .A2(net_251), .A1(net_77) );
NAND2_X2 inst_1668 ( .A1(net_3185), .ZN(net_2090), .A2(net_212) );
CLKBUF_X2 inst_4811 ( .A(net_4796), .Z(net_4797) );
OAI21_X2 inst_721 ( .A(net_825), .ZN(net_678), .B1(net_603), .B2(net_359) );
CLKBUF_X2 inst_4741 ( .A(net_4726), .Z(net_4727) );
OAI22_X2 inst_293 ( .B2(net_3620), .A1(net_3439), .ZN(net_1809), .A2(net_1808), .B1(net_896) );
AOI222_X1 inst_3744 ( .A1(net_4189), .C1(net_3504), .B1(net_3472), .ZN(net_2317), .A2(net_396), .C2(net_387), .B2(net_282) );
INV_X2 inst_3009 ( .ZN(net_3354), .A(net_3353) );
NAND3_X2 inst_1366 ( .ZN(net_3971), .A3(net_3967), .A1(net_1058), .A2(net_877) );
CLKBUF_X2 inst_4397 ( .A(net_4382), .Z(net_4383) );
HA_X1 inst_3102 ( .S(net_274), .CO(net_273), .B(net_75), .A(net_74) );
INV_X2 inst_2695 ( .A(net_2378), .ZN(net_1689) );
AOI221_X2 inst_3860 ( .B2(net_3121), .ZN(net_2022), .B1(net_2020), .C1(net_2019), .A(net_1901), .C2(x307) );
NAND2_X2 inst_1915 ( .A2(net_3108), .ZN(net_285), .A1(net_259) );
INV_X2 inst_2794 ( .A(net_1340), .ZN(net_1324) );
NAND2_X2 inst_2063 ( .ZN(net_3925), .A2(net_3923), .A1(net_840) );
NAND4_X2 inst_1254 ( .ZN(net_3856), .A4(net_3191), .A2(net_2088), .A1(net_2087), .A3(net_1987) );
INV_X2 inst_2953 ( .A(net_3016), .ZN(net_200) );
AOI22_X2 inst_3553 ( .A1(net_4060), .B1(net_4055), .ZN(net_1497), .A2(net_197), .B2(net_175) );
CLKBUF_X2 inst_4801 ( .A(net_4786), .Z(net_4787) );
AOI22_X2 inst_3723 ( .B2(net_3972), .A1(net_3724), .ZN(net_3625), .A2(net_3621), .B1(net_1183) );
AOI22_X2 inst_3521 ( .A2(net_2203), .B1(net_2202), .B2(net_2033), .ZN(net_1925), .A1(net_1847) );
NAND2_X2 inst_1811 ( .A2(net_1105), .ZN(net_895), .A1(net_748) );
XNOR2_X2 inst_98 ( .ZN(net_664), .A(net_663), .B(net_428) );
CLKBUF_X2 inst_4544 ( .A(net_4529), .Z(net_4530) );
AOI21_X2 inst_3985 ( .A(net_3819), .B2(net_3606), .ZN(net_845), .B1(net_844) );
HA_X1 inst_3087 ( .CO(net_1875), .S(net_1743), .A(net_1570), .B(net_243) );
NAND2_X2 inst_2036 ( .A1(net_3894), .A2(net_3867), .ZN(net_3778) );
NOR2_X4 inst_959 ( .A2(net_3942), .ZN(net_3766), .A1(net_3669) );
AOI21_X2 inst_4001 ( .ZN(net_3709), .A(net_3708), .B1(net_3704), .B2(net_284) );
NAND2_X2 inst_2049 ( .ZN(net_3862), .A1(net_2084), .A2(net_1985) );
NOR4_X2 inst_868 ( .A4(net_4096), .A2(net_4001), .A1(net_1103), .ZN(net_1048), .A3(net_583) );
OR3_X4 inst_163 ( .A3(net_3443), .A2(net_2597), .ZN(net_2521), .A1(net_2303) );
OAI221_X2 inst_394 ( .C2(net_3407), .ZN(net_2358), .B1(net_2357), .C1(net_2223), .A(net_1871), .B2(net_112) );
OR2_X4 inst_201 ( .A1(net_3204), .ZN(net_2917), .A2(net_2354) );
OAI21_X2 inst_605 ( .B2(net_2815), .ZN(net_2333), .B1(net_2332), .A(net_1798) );
AOI22_X2 inst_3627 ( .A1(net_3385), .ZN(net_1101), .A2(net_721), .B2(net_641), .B1(net_261) );
NOR2_X2 inst_1084 ( .ZN(net_697), .A1(net_542), .A2(net_261) );
OAI22_X2 inst_304 ( .A2(net_3150), .A1(net_1543), .B1(net_1542), .ZN(net_1538), .B2(net_1537) );
NAND2_X2 inst_1814 ( .ZN(net_1029), .A1(net_867), .A2(net_866) );
INV_X2 inst_2799 ( .ZN(net_1026), .A(net_751) );
AND2_X4 inst_4157 ( .ZN(net_4108), .A1(net_533), .A2(net_529) );
NOR2_X2 inst_1027 ( .A2(net_4052), .ZN(net_1598), .A1(net_1438) );
CLKBUF_X2 inst_4470 ( .A(net_4455), .Z(net_4456) );
NOR2_X2 inst_1143 ( .ZN(net_3876), .A2(net_3251), .A1(net_2245) );
NAND3_X2 inst_1345 ( .ZN(net_3419), .A3(net_3418), .A2(net_3417), .A1(net_3416) );
INV_X2 inst_2947 ( .A(net_3041), .ZN(net_194) );
NAND2_X2 inst_2048 ( .ZN(net_3861), .A2(net_2104), .A1(net_2085) );
CLKBUF_X2 inst_5122 ( .A(net_5107), .Z(net_5108) );
INV_X2 inst_2948 ( .A(net_3052), .ZN(net_150) );
OAI221_X2 inst_361 ( .B1(net_4036), .C1(net_3352), .B2(net_3348), .ZN(net_2789), .A(net_2554), .C2(net_2165) );
AOI22_X2 inst_3608 ( .A1(net_4062), .B1(net_4057), .ZN(net_1409), .A2(net_462), .B2(net_461) );
DFF_X1 inst_3400 ( .Q(net_3117), .D(net_1539), .CK(net_4471) );
NOR2_X2 inst_1016 ( .A2(net_3802), .A1(net_3321), .ZN(net_1828) );
AND2_X4 inst_4147 ( .ZN(net_4084), .A1(net_963), .A2(net_414) );
NAND2_X2 inst_1538 ( .A1(net_2907), .ZN(net_2484), .A2(net_165) );
OAI211_X2 inst_848 ( .ZN(net_2717), .B(net_1998), .A(net_406), .C2(net_344), .C1(net_309) );
NAND2_X2 inst_1931 ( .ZN(net_3199), .A1(net_3198), .A2(net_205) );
CLKBUF_X2 inst_4735 ( .A(net_4720), .Z(net_4721) );
INV_X2 inst_3002 ( .ZN(net_3179), .A(net_3178) );
INV_X4 inst_2479 ( .ZN(net_290), .A(net_29) );
CLKBUF_X2 inst_4389 ( .A(net_4374), .Z(net_4375) );
INV_X4 inst_2179 ( .ZN(net_2740), .A(net_2739) );
INV_X4 inst_2578 ( .ZN(net_3600), .A(net_3599) );
OAI211_X2 inst_786 ( .C2(net_2778), .ZN(net_2761), .B(net_2674), .A(net_2651), .C1(net_2638) );
INV_X2 inst_2940 ( .A(net_3099), .ZN(net_232) );
NAND2_X2 inst_1996 ( .ZN(net_3486), .A2(net_3485), .A1(net_3484) );
NAND2_X2 inst_1554 ( .A1(net_2909), .ZN(net_2468), .A2(net_177) );
NAND2_X2 inst_1542 ( .A1(net_3207), .ZN(net_2480), .A2(net_157) );
CLKBUF_X2 inst_4511 ( .A(net_4440), .Z(net_4497) );
XOR2_X2 inst_2 ( .B(net_4180), .Z(net_1928), .A(net_1878) );
DFF_X1 inst_3340 ( .D(net_2761), .CK(net_4357), .Q(x40) );
OAI21_X2 inst_644 ( .ZN(net_2590), .B2(net_1975), .B1(net_1878), .A(net_1658) );
CLKBUF_X2 inst_4683 ( .A(net_4668), .Z(net_4669) );
CLKBUF_X2 inst_5015 ( .A(net_5000), .Z(net_5001) );
AOI22_X2 inst_3474 ( .B1(net_4039), .ZN(net_2677), .A1(net_2675), .A2(net_225), .B2(x128) );
NAND3_X1 inst_1380 ( .ZN(net_3359), .A2(net_3358), .A1(net_2550), .A3(net_1737) );
INV_X2 inst_2806 ( .A(net_1105), .ZN(net_986) );
OAI21_X2 inst_578 ( .B2(net_2912), .B1(net_2803), .ZN(net_2800), .A(net_2462) );
NOR3_X2 inst_888 ( .A2(net_4066), .ZN(net_2562), .A1(net_2524), .A3(net_2523) );
NAND2_X2 inst_1769 ( .A2(net_3789), .ZN(net_1174), .A1(net_997) );
AOI221_X2 inst_3891 ( .ZN(net_1390), .A(net_1229), .C1(net_1176), .C2(net_1124), .B1(net_656), .B2(net_432) );
AOI22_X2 inst_3625 ( .A1(net_3564), .ZN(net_964), .A2(net_963), .B1(net_957), .B2(net_408) );
AOI21_X2 inst_4008 ( .ZN(net_4159), .B1(net_2241), .A(net_2191), .B2(net_1189) );
CLKBUF_X2 inst_4834 ( .A(net_4313), .Z(net_4820) );
AOI22_X2 inst_3472 ( .B2(net_3119), .A1(net_2724), .B1(net_2722), .ZN(net_2716), .A2(net_32) );
INV_X4 inst_2581 ( .ZN(net_3620), .A(net_3619) );
CLKBUF_X2 inst_4896 ( .A(net_4881), .Z(net_4882) );
AND2_X4 inst_4110 ( .A1(net_3123), .A2(net_3103), .ZN(net_253) );
INV_X8 inst_2164 ( .ZN(net_3769), .A(net_3768) );
NAND2_X2 inst_1498 ( .ZN(net_2819), .A1(net_2774), .A2(net_2720) );
OAI221_X2 inst_432 ( .ZN(net_630), .A(net_629), .B1(net_628), .C1(net_627), .B2(net_393), .C2(net_329) );
OAI22_X2 inst_282 ( .B2(net_4041), .B1(net_2641), .A1(net_2591), .ZN(net_2527), .A2(net_2377) );
NAND3_X2 inst_1358 ( .ZN(net_3718), .A2(net_3715), .A1(net_3682), .A3(net_152) );
CLKBUF_X2 inst_4392 ( .A(net_4377), .Z(net_4378) );
CLKBUF_X2 inst_4915 ( .A(net_4900), .Z(net_4901) );
INV_X4 inst_2322 ( .ZN(net_1117), .A(net_720) );
OAI21_X2 inst_513 ( .B1(net_3274), .B2(net_3208), .ZN(net_2929), .A(net_2492) );
CLKBUF_X2 inst_4775 ( .A(net_4760), .Z(net_4761) );
DFF_X1 inst_3266 ( .QN(net_3070), .D(net_2931), .CK(net_4864) );
DFF_X2 inst_3171 ( .D(net_1949), .QN(net_124), .CK(net_5279) );
NAND2_X2 inst_1630 ( .A1(net_3581), .ZN(net_2513), .A2(net_2373) );
CLKBUF_X2 inst_4450 ( .A(net_4435), .Z(net_4436) );
NAND2_X2 inst_1586 ( .A1(net_2925), .ZN(net_2434), .A2(net_162) );
DFF_X1 inst_3385 ( .D(net_1832), .CK(net_5295), .Q(x633) );
DFF_X2 inst_3182 ( .QN(net_3125), .D(net_1804), .CK(net_4798) );
NAND2_X2 inst_1572 ( .A1(net_2912), .ZN(net_2449), .A2(net_195) );
INV_X2 inst_2866 ( .A(net_3127), .ZN(net_928) );
OAI21_X1 inst_774 ( .ZN(net_4010), .B2(net_2959), .B1(net_2893), .A(net_2504) );
INV_X4 inst_2292 ( .ZN(net_2268), .A(net_914) );
CLKBUF_X2 inst_4906 ( .A(net_4891), .Z(net_4892) );
CLKBUF_X2 inst_4256 ( .A(net_4241), .Z(net_4242) );
OAI211_X2 inst_838 ( .C1(net_1359), .ZN(net_1352), .C2(net_1351), .A(net_1233), .B(net_593) );
CLKBUF_X2 inst_5300 ( .A(net_5285), .Z(net_5286) );
INV_X2 inst_2766 ( .ZN(net_933), .A(net_870) );
CLKBUF_X2 inst_4326 ( .A(net_4308), .Z(net_4312) );
NAND2_X2 inst_1508 ( .A2(net_3600), .ZN(net_2689), .A1(net_2688) );
NAND4_X2 inst_1222 ( .ZN(net_951), .A4(net_733), .A3(net_554), .A1(net_520), .A2(net_480) );
CLKBUF_X2 inst_4978 ( .A(net_4538), .Z(net_4964) );
NAND2_X4 inst_1405 ( .A1(net_3498), .ZN(net_3238), .A2(net_2858) );
DFF_X1 inst_3407 ( .Q(net_4029), .D(net_1398), .CK(net_4500) );
AND4_X2 inst_4058 ( .ZN(net_1344), .A1(net_1343), .A4(net_1301), .A2(net_1174), .A3(net_1040) );
NOR2_X2 inst_1073 ( .ZN(net_698), .A1(net_697), .A2(net_611) );
INV_X4 inst_2323 ( .A(net_1041), .ZN(net_819) );
AOI222_X1 inst_3741 ( .A1(net_4189), .C1(net_3504), .B1(net_3472), .C2(net_3418), .ZN(net_2320), .A2(net_2033), .B2(net_179) );
INV_X2 inst_2749 ( .ZN(net_1079), .A(net_1078) );
NAND2_X4 inst_1449 ( .ZN(net_3808), .A2(net_3807), .A1(net_3537) );
XNOR2_X1 inst_127 ( .ZN(net_1732), .B(net_1608), .A(net_1597) );
CLKBUF_X2 inst_4367 ( .A(net_4307), .Z(net_4353) );
NAND2_X2 inst_2013 ( .A1(net_3913), .ZN(net_3614), .A2(net_3613) );
OR3_X2 inst_187 ( .ZN(net_3425), .A1(net_1650), .A2(net_966), .A3(net_415) );
OR2_X4 inst_206 ( .ZN(net_2965), .A2(net_2352), .A1(net_2350) );
CLKBUF_X2 inst_4506 ( .A(net_4491), .Z(net_4492) );
AOI222_X1 inst_3739 ( .B2(net_4030), .A2(net_3445), .C1(net_3242), .A1(net_3241), .B1(net_2752), .ZN(net_2635), .C2(net_2386) );
INV_X2 inst_3029 ( .ZN(net_3522), .A(net_434) );
NAND3_X4 inst_1268 ( .ZN(net_3869), .A3(net_3718), .A1(net_3683), .A2(net_3527) );
XNOR2_X2 inst_122 ( .B(net_4139), .ZN(net_4138), .A(net_818) );
INV_X2 inst_2756 ( .ZN(net_999), .A(net_998) );
OAI221_X2 inst_405 ( .C1(net_3492), .ZN(net_1947), .B2(net_1946), .A(net_1868), .B1(net_1800), .C2(net_1694) );
NAND2_X2 inst_1731 ( .A1(net_1556), .ZN(net_1554), .A2(x762) );
OAI21_X2 inst_492 ( .B1(net_3588), .B2(net_2967), .ZN(net_2950), .A(net_2405) );
CLKBUF_X2 inst_4788 ( .A(net_4773), .Z(net_4774) );
INV_X2 inst_2960 ( .A(net_3031), .ZN(net_213) );
NAND2_X2 inst_1909 ( .A2(net_3165), .ZN(net_325), .A1(net_321) );
AOI221_X2 inst_3912 ( .B2(net_4127), .A(net_4113), .ZN(net_687), .C1(net_686), .C2(net_342), .B1(net_245) );
CLKBUF_X2 inst_4318 ( .A(net_4268), .Z(net_4304) );
INV_X4 inst_2306 ( .A(net_1338), .ZN(net_837) );
CLKBUF_X2 inst_4335 ( .A(net_4320), .Z(net_4321) );
XNOR2_X2 inst_82 ( .B(net_4081), .ZN(net_1522), .A(net_1027) );
AND2_X4 inst_4187 ( .ZN(net_4183), .A1(net_2553), .A2(net_2003) );
CLKBUF_X2 inst_4239 ( .A(net_4224), .Z(net_4225) );
NAND2_X2 inst_1646 ( .ZN(net_2699), .A2(net_2169), .A1(net_2126) );
INV_X4 inst_2176 ( .ZN(net_2855), .A(net_2759) );
INV_X2 inst_2892 ( .A(net_3051), .ZN(net_146) );
NOR2_X2 inst_1121 ( .ZN(net_3414), .A2(net_3413), .A1(net_2718) );
NOR2_X2 inst_1102 ( .ZN(net_339), .A2(net_258), .A1(net_53) );
DFF_X2 inst_3161 ( .D(net_2164), .QN(net_109), .CK(net_4376) );
DFF_X2 inst_3187 ( .D(net_1742), .QN(net_266), .CK(net_4835) );
OAI22_X2 inst_307 ( .A2(net_2637), .A1(net_1543), .B1(net_1542), .ZN(net_1533), .B2(net_1532) );
INV_X2 inst_2816 ( .A(net_3733), .ZN(net_710) );
OAI21_X2 inst_702 ( .A(net_4084), .ZN(net_910), .B1(net_902), .B2(net_853) );
NAND2_X2 inst_2034 ( .ZN(net_3772), .A1(net_1809), .A2(net_360) );
NAND2_X2 inst_1505 ( .A2(net_3515), .ZN(net_2730), .A1(net_2620) );
OAI21_X2 inst_717 ( .B2(net_4000), .ZN(net_925), .B1(net_904), .A(net_702) );
OAI22_X4 inst_276 ( .A1(net_3556), .A2(net_3003), .B2(net_3000), .ZN(net_2110), .B1(net_1973) );
INV_X4 inst_2482 ( .A(net_3049), .ZN(net_495) );
INV_X2 inst_2957 ( .ZN(net_229), .A(net_112) );
DFF_X1 inst_3339 ( .D(net_2771), .CK(net_4360), .Q(x23) );
AOI222_X1 inst_3791 ( .ZN(net_985), .A2(net_984), .C1(net_983), .A1(net_638), .B1(net_599), .C2(net_333), .B2(net_225) );
INV_X2 inst_2711 ( .A(net_3437), .ZN(net_1602) );
AOI22_X2 inst_3531 ( .A1(net_3782), .B2(net_3160), .ZN(net_1883), .B1(net_1882), .A2(net_1762) );
INV_X2 inst_2753 ( .ZN(net_2189), .A(net_1044) );
AOI22_X2 inst_3672 ( .ZN(net_550), .A1(net_458), .B1(net_457), .A2(net_199), .B2(net_165) );
CLKBUF_X2 inst_5297 ( .A(net_5282), .Z(net_5283) );
XNOR2_X2 inst_91 ( .ZN(net_855), .B(net_854), .A(net_715) );
NAND2_X2 inst_1762 ( .A2(net_1394), .ZN(net_1237), .A1(net_34) );
SDFF_X2 inst_132 ( .D(net_3483), .SI(net_3024), .Q(net_3024), .SE(net_2912), .CK(net_5055) );
NAND2_X2 inst_2023 ( .ZN(net_3714), .A1(net_3712), .A2(net_976) );
INV_X2 inst_2779 ( .ZN(net_807), .A(net_761) );
AOI22_X2 inst_3686 ( .B2(net_4123), .A2(net_509), .ZN(net_494), .A1(net_493), .B1(net_492) );
AOI221_X2 inst_3842 ( .B2(net_2203), .C1(net_2202), .ZN(net_2200), .A(net_2072), .B1(net_2059), .C2(net_1791) );
CLKBUF_X2 inst_4919 ( .A(net_4904), .Z(net_4905) );
NAND2_X2 inst_1703 ( .ZN(net_1784), .A2(net_1783), .A1(net_1739) );
AOI22_X2 inst_3545 ( .B1(net_4054), .A1(net_1578), .ZN(net_1577), .A2(net_168), .B2(net_156) );
CLKBUF_X2 inst_4715 ( .A(net_4482), .Z(net_4701) );
AOI22_X2 inst_3611 ( .A1(net_4063), .B1(net_4058), .ZN(net_1406), .B2(net_176), .A2(net_163) );
INV_X2 inst_2928 ( .A(net_3126), .ZN(net_145) );
AOI221_X2 inst_3813 ( .A(net_2642), .B1(net_2641), .C1(net_2590), .ZN(net_2588), .C2(net_2581), .B2(net_280) );
OAI221_X2 inst_400 ( .B2(net_3428), .ZN(net_2284), .C1(net_2235), .B1(net_2184), .A(net_1991), .C2(net_110) );
INV_X2 inst_2991 ( .A(net_3120), .ZN(net_1541) );
OAI21_X2 inst_614 ( .A(net_3156), .ZN(net_2591), .B1(net_2293), .B2(net_2248) );
AOI22_X2 inst_3513 ( .B1(net_2625), .ZN(net_1970), .A1(net_1969), .A2(net_1837), .B2(net_152) );
NAND2_X2 inst_1896 ( .ZN(net_514), .A2(net_349), .A1(net_185) );
OR2_X2 inst_261 ( .A1(net_877), .ZN(net_863), .A2(net_745) );
NOR2_X2 inst_1031 ( .ZN(net_1578), .A1(net_1459), .A2(net_1458) );
NOR2_X4 inst_945 ( .ZN(net_3518), .A2(net_3454), .A1(net_2030) );
OR2_X2 inst_268 ( .A1(net_4137), .ZN(net_3374), .A2(net_42) );
NAND2_X2 inst_1518 ( .A1(net_3689), .ZN(net_2510), .A2(net_239) );
OAI221_X2 inst_369 ( .C1(net_3618), .ZN(net_2700), .C2(net_2699), .B2(net_2698), .B1(net_2543), .A(net_2368) );
CLKBUF_X2 inst_5161 ( .A(net_4542), .Z(net_5147) );
NAND2_X2 inst_1900 ( .A1(net_3657), .ZN(net_826), .A2(net_357) );
AOI21_X2 inst_3975 ( .B2(net_3399), .A(net_3337), .ZN(net_1159), .B1(net_995) );
OAI22_X2 inst_327 ( .A2(net_3468), .ZN(net_884), .B2(net_721), .A1(net_641), .B1(net_43) );
AOI22_X2 inst_3509 ( .B1(net_3676), .B2(net_3138), .A1(net_2012), .ZN(net_2008), .A2(net_1791) );
INV_X2 inst_2916 ( .A(net_3067), .ZN(net_244) );
NAND3_X2 inst_1286 ( .ZN(net_2261), .A1(net_2198), .A3(net_1952), .A2(net_1917) );
OR2_X2 inst_266 ( .ZN(net_3253), .A1(net_1161), .A2(net_1160) );
NAND2_X2 inst_2051 ( .ZN(net_3873), .A1(net_1982), .A2(net_177) );
AOI221_X2 inst_3853 ( .ZN(net_2061), .A(net_2060), .C1(net_2059), .C2(net_1908), .B2(net_749), .B1(net_94) );
NAND4_X2 inst_1198 ( .ZN(net_1676), .A3(net_1479), .A4(net_1478), .A1(net_1413), .A2(net_1412) );
XNOR2_X2 inst_77 ( .A(net_3379), .ZN(net_1387), .B(net_1291) );
OR3_X4 inst_171 ( .A2(net_3978), .ZN(net_882), .A3(net_881), .A1(net_707) );
HA_X1 inst_3097 ( .S(net_821), .CO(net_820), .A(net_642), .B(net_216) );
AOI22_X2 inst_3661 ( .A2(net_3027), .B2(net_3026), .A1(net_571), .B1(net_570), .ZN(net_566) );
OAI221_X2 inst_374 ( .B2(net_2733), .C1(net_2686), .ZN(net_2682), .A(net_2560), .B1(net_2332), .C2(net_2147) );
OAI21_X2 inst_502 ( .B1(net_3588), .B2(net_2959), .ZN(net_2940), .A(net_2498) );
XNOR2_X2 inst_103 ( .ZN(net_507), .A(net_372), .B(net_348) );
AOI22_X2 inst_3690 ( .B2(net_4124), .A2(net_555), .ZN(net_486), .B1(net_241), .A1(net_212) );
DFF_X1 inst_3221 ( .QN(net_3059), .D(net_2978), .CK(net_4568) );
AOI22_X2 inst_3645 ( .A1(net_4142), .B1(net_4112), .ZN(net_757), .B2(net_378), .A2(x717) );
NAND2_X2 inst_1598 ( .A1(net_2917), .ZN(net_2420), .A2(net_203) );
AOI222_X2 inst_3738 ( .C2(net_3418), .B2(net_1826), .ZN(net_977), .B1(net_677), .A1(net_626), .C1(net_578), .A2(net_225) );
OAI222_X1 inst_357 ( .C1(net_3784), .ZN(net_3362), .B2(net_3354), .A2(net_3153), .B1(net_1815), .A1(net_1814), .C2(net_117) );
INV_X2 inst_2855 ( .A(net_3657), .ZN(net_334) );
AND2_X4 inst_4092 ( .ZN(net_2849), .A1(net_2758), .A2(net_1825) );
NAND2_X2 inst_2058 ( .ZN(net_3910), .A2(net_3909), .A1(net_3908) );
OAI211_X2 inst_809 ( .A(net_3730), .ZN(net_1662), .C1(net_1617), .B(net_785), .C2(net_325) );
AOI21_X2 inst_3980 ( .A(net_4033), .ZN(net_981), .B2(net_770), .B1(net_57) );
AOI22_X2 inst_3675 ( .B2(net_555), .ZN(net_546), .A1(net_457), .A2(net_234), .B1(net_205) );
DFF_X2 inst_3152 ( .QN(net_3165), .D(net_2271), .CK(net_4805) );
AND2_X4 inst_4161 ( .ZN(net_4112), .A2(net_671), .A1(net_511) );
AOI222_X1 inst_3758 ( .A1(net_3676), .B1(net_2055), .C1(net_2054), .ZN(net_2034), .B2(net_2033), .A2(net_252), .C2(net_106) );
INV_X4 inst_2562 ( .ZN(net_3516), .A(net_3515) );
NAND4_X2 inst_1234 ( .ZN(net_869), .A3(net_557), .A1(net_524), .A2(net_490), .A4(net_465) );
NOR3_X2 inst_912 ( .ZN(net_3448), .A3(net_3447), .A2(net_3446), .A1(net_3445) );
INV_X4 inst_2398 ( .ZN(net_398), .A(net_320) );
INV_X4 inst_2595 ( .A(net_3951), .ZN(net_3727) );
NOR2_X2 inst_1022 ( .A1(net_3492), .ZN(net_1747), .A2(net_1641) );
DFF_X2 inst_3196 ( .D(net_1612), .Q(net_85), .CK(net_4797) );
INV_X4 inst_2371 ( .A(net_1126), .ZN(net_912) );
INV_X2 inst_2939 ( .A(net_3121), .ZN(net_1545) );
AOI211_X2 inst_4025 ( .ZN(net_1197), .A(net_1196), .C1(net_1135), .B(net_968), .C2(net_407) );
OAI22_X2 inst_322 ( .A1(net_2167), .A2(net_1071), .ZN(net_1021), .B2(net_433), .B1(net_135) );
NAND4_X2 inst_1223 ( .ZN(net_906), .A4(net_682), .A3(net_572), .A2(net_496), .A1(net_486) );
AOI22_X2 inst_3516 ( .B1(net_4045), .A2(net_3133), .A1(net_1955), .ZN(net_1954), .B2(net_282) );
INV_X2 inst_2785 ( .ZN(net_801), .A(net_755) );
AOI221_X2 inst_3906 ( .A(net_4090), .C2(net_1045), .ZN(net_1010), .C1(net_790), .B1(net_694), .B2(net_414) );
AND2_X2 inst_4200 ( .A1(net_3925), .ZN(net_900), .A2(net_403) );
AND2_X4 inst_4188 ( .ZN(net_4184), .A1(net_1308), .A2(net_59) );
OAI21_X2 inst_681 ( .B2(net_3974), .ZN(net_1290), .A(net_1279), .B1(net_1108) );
CLKBUF_X2 inst_4886 ( .A(net_4842), .Z(net_4872) );
AND2_X4 inst_4169 ( .ZN(net_4123), .A1(net_338), .A2(net_144) );
AOI221_X2 inst_3902 ( .ZN(net_1609), .B2(net_1011), .A(net_993), .B1(net_787), .C1(net_696), .C2(net_432) );
NAND2_X2 inst_2010 ( .A2(net_3866), .ZN(net_3582), .A1(net_3516) );
INV_X2 inst_2915 ( .A(net_3096), .ZN(net_167) );
DFF_X1 inst_3296 ( .QN(net_3008), .D(net_2884), .CK(net_5220) );
AND2_X4 inst_4181 ( .ZN(net_4142), .A1(net_1463), .A2(x1023) );
NOR4_X2 inst_871 ( .A4(net_4106), .A1(net_3429), .ZN(net_1143), .A2(net_919), .A3(net_794) );
INV_X4 inst_2315 ( .A(net_1200), .ZN(net_983) );
INV_X2 inst_2684 ( .A(net_2076), .ZN(net_1836) );
NOR2_X4 inst_962 ( .ZN(net_3787), .A2(net_3216), .A1(net_2110) );
OAI21_X2 inst_532 ( .B1(net_3195), .B2(net_2969), .ZN(net_2901), .A(net_2418) );
DFF_X2 inst_3164 ( .D(net_2162), .QN(net_61), .CK(net_4654) );
INV_X2 inst_2965 ( .A(net_3118), .ZN(net_130) );
INV_X4 inst_2382 ( .ZN(net_931), .A(net_401) );
NAND2_X2 inst_2008 ( .A1(net_3817), .ZN(net_3538), .A2(net_199) );
NOR2_X1 inst_1171 ( .ZN(net_3690), .A1(net_2307), .A2(net_70) );
OAI21_X2 inst_641 ( .ZN(net_1995), .B1(net_1993), .A(net_1895), .B2(net_1532) );
CLKBUF_X2 inst_5274 ( .A(net_4908), .Z(net_5260) );
INV_X2 inst_2969 ( .ZN(net_149), .A(net_107) );
OAI21_X2 inst_498 ( .B1(net_3588), .B2(net_2963), .ZN(net_2944), .A(net_2455) );
DFF_X1 inst_3314 ( .Q(net_3132), .D(net_2841), .CK(net_4658) );
NAND2_X2 inst_1988 ( .A1(net_3969), .A2(net_3634), .ZN(net_3432) );
CLKBUF_X2 inst_5113 ( .A(net_5098), .Z(net_5099) );
INV_X4 inst_2594 ( .ZN(net_3721), .A(net_3720) );
AND4_X4 inst_4037 ( .ZN(net_1760), .A2(net_1589), .A1(net_1055), .A3(net_1005), .A4(net_971) );
NAND2_X2 inst_1912 ( .ZN(net_293), .A1(net_290), .A2(net_250) );
AOI21_X2 inst_3976 ( .ZN(net_1156), .A(net_1155), .B1(net_1154), .B2(net_1153) );
NAND2_X2 inst_1831 ( .ZN(net_794), .A2(net_745), .A1(net_674) );
NAND3_X2 inst_1327 ( .A2(net_3713), .A3(net_3590), .ZN(net_672), .A1(net_602) );
AOI22_X2 inst_3468 ( .B2(net_3117), .A1(net_2724), .ZN(net_2723), .B1(net_2722), .A2(net_34) );
OAI222_X2 inst_350 ( .C1(net_3784), .A2(net_2165), .ZN(net_1937), .A1(net_1815), .B1(net_1814), .B2(net_327), .C2(net_116) );
INV_X4 inst_2395 ( .ZN(net_594), .A(net_358) );
OR2_X4 inst_231 ( .A1(net_3158), .ZN(net_409), .A2(net_406) );
NOR2_X2 inst_1119 ( .ZN(net_3409), .A1(net_2610), .A2(net_2385) );
DFF_X1 inst_3309 ( .QN(net_3014), .D(net_2867), .CK(net_5204) );
AOI22_X2 inst_3699 ( .B1(net_4123), .A1(net_555), .ZN(net_473), .A2(net_203), .B2(net_173) );
CLKBUF_X2 inst_5104 ( .A(net_5089), .Z(net_5090) );
CLKBUF_X2 inst_5082 ( .A(net_5067), .Z(net_5068) );
NAND4_X2 inst_1255 ( .ZN(net_3879), .A3(net_3210), .A2(net_3209), .A4(net_3205), .A1(net_2177) );
CLKBUF_X2 inst_5050 ( .A(net_4422), .Z(net_5036) );
INV_X4 inst_2317 ( .ZN(net_1652), .A(net_1637) );
NAND2_X2 inst_1791 ( .A2(net_1264), .ZN(net_993), .A1(net_882) );
NAND2_X4 inst_1452 ( .ZN(net_3831), .A2(net_3830), .A1(net_3202) );
CLKBUF_X2 inst_4925 ( .A(net_4652), .Z(net_4911) );
DFF_X1 inst_3420 ( .D(net_1358), .Q(net_32), .CK(net_4285) );
CLKBUF_X2 inst_5000 ( .A(net_4356), .Z(net_4986) );
AND3_X4 inst_4077 ( .ZN(net_4096), .A1(net_3993), .A3(net_3628), .A2(net_337) );
DFF_X2 inst_3139 ( .QN(net_2985), .D(net_2574), .CK(net_5238) );
CLKBUF_X2 inst_4457 ( .A(net_4442), .Z(net_4443) );
CLKBUF_X2 inst_5064 ( .A(net_5049), .Z(net_5050) );
OAI21_X2 inst_528 ( .B1(net_3302), .B2(net_3207), .ZN(net_2906), .A(net_2479) );
INV_X4 inst_2558 ( .ZN(net_3503), .A(net_3502) );
NOR3_X2 inst_903 ( .A2(net_1717), .ZN(net_960), .A1(net_913), .A3(net_847) );
NAND2_X2 inst_1725 ( .A1(net_2042), .ZN(net_1653), .A2(net_671) );
CLKBUF_X2 inst_4957 ( .A(net_4942), .Z(net_4943) );
NAND2_X4 inst_1396 ( .A1(net_3229), .ZN(net_1600), .A2(net_294) );
OAI222_X2 inst_352 ( .C1(net_3784), .A2(net_2272), .C2(net_1960), .ZN(net_1858), .A1(net_1815), .B1(net_1814), .B2(net_316) );
OAI211_X2 inst_846 ( .C1(net_1274), .ZN(net_892), .B(net_891), .A(net_779), .C2(net_777) );
OAI22_X2 inst_286 ( .B2(net_3164), .A2(net_2514), .ZN(net_1974), .A1(net_1843), .B1(x475) );
AOI22_X2 inst_3504 ( .B1(net_3676), .B2(net_3147), .A2(net_2033), .ZN(net_2014), .A1(net_2012) );
AOI21_X4 inst_3924 ( .B2(net_3600), .ZN(net_3482), .A(net_3481), .B1(net_3372) );
NAND2_X2 inst_1734 ( .A1(net_1556), .ZN(net_1551), .A2(x916) );
CLKBUF_X2 inst_4510 ( .A(net_4424), .Z(net_4496) );
CLKBUF_X2 inst_4646 ( .A(net_4631), .Z(net_4632) );
CLKBUF_X2 inst_4572 ( .A(net_4557), .Z(net_4558) );
CLKBUF_X2 inst_5189 ( .A(net_5174), .Z(net_5175) );
INV_X2 inst_3003 ( .A(net_3219), .ZN(net_3206) );
AOI221_X2 inst_3841 ( .B2(net_2203), .C1(net_2202), .ZN(net_2201), .A(net_2078), .B1(net_1823), .C2(net_168) );
AOI22_X2 inst_3464 ( .ZN(net_2767), .A1(net_2738), .B1(net_2711), .A2(net_1323), .B2(net_211) );
INV_X4 inst_2185 ( .ZN(net_2675), .A(net_2546) );
AND4_X4 inst_4050 ( .ZN(net_4094), .A1(net_3900), .A3(net_3395), .A4(net_513), .A2(net_386) );
NOR2_X2 inst_1044 ( .A1(net_1587), .ZN(net_1180), .A2(net_1064) );
DFF_X1 inst_3354 ( .D(net_2632), .Q(net_68), .CK(net_4262) );
INV_X4 inst_2370 ( .A(net_533), .ZN(net_430) );
CLKBUF_X2 inst_4993 ( .A(net_4978), .Z(net_4979) );
AOI221_X2 inst_3882 ( .B1(net_2020), .C1(net_2019), .ZN(net_1813), .A(net_1812), .B2(net_77), .C2(x450) );
INV_X2 inst_2811 ( .ZN(net_651), .A(net_650) );
INV_X2 inst_3014 ( .ZN(net_3401), .A(net_3011) );
CLKBUF_X2 inst_4615 ( .A(net_4600), .Z(net_4601) );
SDFF_X2 inst_137 ( .SE(net_2625), .D(net_2367), .SI(net_94), .Q(net_94), .CK(net_4961) );
OAI221_X2 inst_425 ( .C1(net_3924), .C2(net_3755), .B1(net_3566), .B2(net_3478), .ZN(net_1147), .A(net_998) );
INV_X4 inst_2567 ( .A(net_3685), .ZN(net_3533) );
DFF_X2 inst_3206 ( .QN(net_3102), .D(net_1303), .CK(net_4985) );
NAND2_X2 inst_1532 ( .A1(net_3208), .ZN(net_2490), .A2(net_596) );
OR2_X4 inst_227 ( .ZN(net_1105), .A1(net_693), .A2(net_605) );
CLKBUF_X2 inst_4303 ( .A(net_4288), .Z(net_4289) );
INV_X8 inst_2136 ( .A(net_3108), .ZN(net_337) );
AOI21_X4 inst_3927 ( .ZN(net_3583), .B1(net_3366), .A(net_3297), .B2(net_2607) );
INV_X2 inst_2891 ( .ZN(net_770), .A(x956) );
INV_X2 inst_2718 ( .A(net_3859), .ZN(net_2342) );
INV_X4 inst_2572 ( .A(net_3672), .ZN(net_3550) );
XNOR2_X2 inst_58 ( .ZN(net_2121), .B(net_1928), .A(net_1787) );
AOI22_X2 inst_3633 ( .A1(net_990), .ZN(net_876), .B1(net_874), .B2(net_721), .A2(net_371) );
AND4_X4 inst_4046 ( .A2(net_4110), .ZN(net_4075), .A4(net_3327), .A3(net_722), .A1(net_433) );
DFF_X1 inst_3365 ( .D(net_2308), .CK(net_4253), .Q(x179) );
NAND2_X4 inst_1469 ( .ZN(net_3901), .A2(net_3900), .A1(net_3899) );
DFF_X1 inst_3254 ( .QN(net_3079), .D(net_2951), .CK(net_4539) );
CLKBUF_X2 inst_5029 ( .A(net_4670), .Z(net_5015) );
NOR2_X2 inst_983 ( .ZN(net_2693), .A1(net_2624), .A2(net_2623) );
CLKBUF_X2 inst_4980 ( .A(net_4965), .Z(net_4966) );
NAND2_X2 inst_1897 ( .ZN(net_362), .A1(net_345), .A2(net_144) );
DFF_X2 inst_3159 ( .D(net_2157), .QN(net_58), .CK(net_4381) );
CLKBUF_X2 inst_5288 ( .A(net_5273), .Z(net_5274) );
INV_X4 inst_2551 ( .A(net_3686), .ZN(net_3456) );
OAI21_X2 inst_581 ( .B2(net_3207), .B1(net_2803), .ZN(net_2797), .A(net_2488) );
CLKBUF_X2 inst_4407 ( .A(net_4392), .Z(net_4393) );
XOR2_X1 inst_28 ( .Z(net_1281), .B(net_1280), .A(net_1085) );
INV_X4 inst_2424 ( .A(net_3128), .ZN(net_248) );
CLKBUF_X2 inst_4517 ( .A(net_4502), .Z(net_4503) );
CLKBUF_X2 inst_4776 ( .A(net_4761), .Z(net_4762) );
NAND2_X2 inst_1569 ( .A1(net_2912), .ZN(net_2452), .A2(net_202) );
DFF_X2 inst_3144 ( .D(net_2539), .QN(net_111), .CK(net_4395) );
INV_X2 inst_2633 ( .A(net_2670), .ZN(net_2659) );
NAND2_X2 inst_1772 ( .ZN(net_1369), .A1(net_1050), .A2(net_748) );
OAI21_X2 inst_592 ( .B1(net_2615), .ZN(net_2580), .B2(net_1529), .A(net_671) );
AOI22_X2 inst_3666 ( .B2(net_4015), .A2(net_4013), .A1(net_571), .B1(net_570), .ZN(net_561) );
NOR2_X2 inst_993 ( .A2(net_3447), .ZN(net_2299), .A1(net_2216) );
INV_X8 inst_2143 ( .ZN(net_3198), .A(net_3197) );
NAND3_X2 inst_1291 ( .ZN(net_2256), .A1(net_2199), .A3(net_1950), .A2(net_1922) );
CLKBUF_X2 inst_5177 ( .A(net_5162), .Z(net_5163) );
CLKBUF_X2 inst_5143 ( .A(net_5128), .Z(net_5129) );
INV_X8 inst_2130 ( .A(net_3613), .ZN(net_358) );
OAI221_X2 inst_359 ( .B2(net_3381), .ZN(net_2830), .B1(net_2826), .C1(net_2825), .A(net_2586), .C2(net_1516) );
CLKBUF_X2 inst_4388 ( .A(net_4373), .Z(net_4374) );
NOR2_X2 inst_1055 ( .A1(net_1132), .ZN(net_1050), .A2(net_532) );
CLKBUF_X2 inst_5096 ( .A(net_5081), .Z(net_5082) );
NAND2_X1 inst_2100 ( .ZN(net_3805), .A2(net_3803), .A1(net_3329) );
AOI21_X2 inst_3948 ( .A(net_3363), .B1(net_2238), .ZN(net_2208), .B2(net_243) );
INV_X4 inst_2284 ( .ZN(net_1656), .A(net_1120) );
NAND2_X2 inst_1962 ( .A2(net_3751), .A1(net_3694), .ZN(net_3311) );
OAI21_X2 inst_630 ( .B1(net_4044), .ZN(net_2241), .A(net_2142), .B2(net_2127) );
CLKBUF_X2 inst_5227 ( .A(net_5212), .Z(net_5213) );
CLKBUF_X2 inst_4829 ( .A(net_4814), .Z(net_4815) );
CLKBUF_X2 inst_5268 ( .A(net_5253), .Z(net_5254) );
CLKBUF_X2 inst_4757 ( .A(net_4338), .Z(net_4743) );
NAND3_X2 inst_1273 ( .ZN(net_2879), .A1(net_2864), .A2(net_2796), .A3(net_2751) );
NOR2_X4 inst_923 ( .ZN(net_2279), .A1(net_2178), .A2(net_2112) );
OAI21_X2 inst_512 ( .B1(net_3274), .B2(net_2959), .ZN(net_2930), .A(net_2500) );
CLKBUF_X2 inst_4966 ( .A(net_4381), .Z(net_4952) );
NAND3_X2 inst_1301 ( .A2(net_3406), .A3(net_1845), .ZN(net_1377), .A1(net_1376) );
CLKBUF_X2 inst_5283 ( .A(net_5268), .Z(net_5269) );
INV_X8 inst_2151 ( .A(net_3569), .ZN(net_3345) );
INV_X2 inst_2830 ( .A(net_3215), .ZN(net_440) );
OAI21_X2 inst_647 ( .ZN(net_2114), .B2(net_1852), .A(net_620), .B1(net_619) );
INV_X2 inst_3054 ( .ZN(net_3914), .A(net_3912) );
OR2_X4 inst_194 ( .ZN(net_2907), .A2(net_2354), .A1(net_2353) );
CLKBUF_X2 inst_4764 ( .A(net_4305), .Z(net_4750) );
CLKBUF_X2 inst_5137 ( .A(net_5059), .Z(net_5123) );
INV_X2 inst_2985 ( .A(net_3114), .ZN(net_1537) );
AOI222_X1 inst_3766 ( .B1(net_4048), .A1(net_1968), .ZN(net_1966), .C1(net_375), .C2(net_361), .A2(net_240), .B2(net_69) );
OAI211_X2 inst_833 ( .C1(net_1359), .ZN(net_1358), .A(net_1240), .B(net_593), .C2(net_331) );
AOI222_X1 inst_3772 ( .A2(net_2033), .ZN(net_1900), .A1(net_1863), .B1(net_1862), .C1(net_1861), .C2(net_1280), .B2(net_856) );
AND2_X2 inst_4210 ( .A1(net_4126), .ZN(net_3985), .A2(net_3979) );
INV_X4 inst_2536 ( .A(net_3867), .ZN(net_3347) );
NAND2_X2 inst_2043 ( .ZN(net_3845), .A2(net_3842), .A1(net_432) );
NOR2_X4 inst_960 ( .A2(net_3837), .ZN(net_3775), .A1(net_3574) );
CLKBUF_X2 inst_4924 ( .A(net_4909), .Z(net_4910) );
XNOR2_X2 inst_118 ( .ZN(net_3794), .B(net_3792), .A(net_1285) );
INV_X4 inst_2411 ( .ZN(net_271), .A(net_59) );
OAI221_X2 inst_442 ( .B2(net_3978), .C2(net_3634), .ZN(net_3558), .B1(net_1152), .C1(net_897), .A(net_841) );
INV_X4 inst_2507 ( .A(net_3059), .ZN(net_568) );
INV_X4 inst_2245 ( .ZN(net_1840), .A(net_1465) );
XOR2_X1 inst_38 ( .Z(net_4147), .B(net_1511), .A(net_1310) );
INV_X4 inst_2601 ( .ZN(net_3760), .A(net_3759) );
NAND2_X2 inst_2037 ( .A2(net_3959), .ZN(net_3789), .A1(net_3606) );
OAI221_X2 inst_381 ( .B2(net_2670), .C1(net_2668), .ZN(net_2639), .B1(net_2638), .C2(net_2637), .A(net_1386) );
CLKBUF_X2 inst_5237 ( .A(net_5222), .Z(net_5223) );
AOI221_X2 inst_3837 ( .B1(net_3774), .C1(net_2227), .ZN(net_2223), .C2(net_2222), .A(net_2113), .B2(net_294) );
NAND2_X2 inst_1925 ( .ZN(net_3188), .A1(net_3187), .A2(net_188) );
CLKBUF_X2 inst_4298 ( .A(net_4283), .Z(net_4284) );
NOR3_X2 inst_883 ( .ZN(net_2812), .A1(net_2770), .A2(net_2749), .A3(net_2616) );
XNOR2_X2 inst_40 ( .ZN(net_2828), .A(net_2678), .B(net_1696) );
CLKBUF_X2 inst_4437 ( .A(net_4208), .Z(net_4423) );
NAND4_X2 inst_1249 ( .A3(net_3971), .A4(net_3970), .ZN(net_3626), .A2(net_3625), .A1(net_3624) );
OAI21_X2 inst_756 ( .ZN(net_3710), .A(net_3709), .B2(net_3407), .B1(net_2229) );
AND2_X4 inst_4099 ( .A1(net_4067), .ZN(net_1365), .A2(net_996) );
CLKBUF_X2 inst_4740 ( .A(net_4725), .Z(net_4726) );
NAND2_X4 inst_1416 ( .ZN(net_3510), .A2(net_2342), .A1(net_2288) );
NAND3_X2 inst_1318 ( .ZN(net_1845), .A2(net_432), .A1(net_339), .A3(net_321) );
OAI221_X2 inst_439 ( .ZN(net_3386), .C2(net_3385), .A(net_629), .C1(net_628), .B1(net_627), .B2(net_42) );
CLKBUF_X2 inst_4597 ( .A(net_4582), .Z(net_4583) );
NAND4_X2 inst_1188 ( .A4(net_4112), .A1(net_3427), .A3(net_3406), .ZN(net_1993), .A2(net_1376) );
NOR2_X1 inst_1165 ( .A1(net_3229), .ZN(net_1373), .A2(net_69) );
CLKBUF_X2 inst_4529 ( .A(net_4514), .Z(net_4515) );
INV_X2 inst_2644 ( .ZN(net_2337), .A(net_2316) );
CLKBUF_X2 inst_4584 ( .A(net_4569), .Z(net_4570) );
NOR2_X2 inst_1070 ( .A1(net_3563), .A2(net_3549), .ZN(net_867) );
INV_X4 inst_2626 ( .ZN(net_4004), .A(net_3167) );
CLKBUF_X2 inst_4629 ( .A(net_4614), .Z(net_4615) );
INV_X4 inst_2454 ( .A(net_3090), .ZN(net_596) );
AOI22_X2 inst_3601 ( .A1(net_4062), .B1(net_4057), .ZN(net_1416), .B2(net_492), .A2(net_471) );
AOI221_X2 inst_3873 ( .B1(net_2020), .C1(net_2019), .ZN(net_1930), .A(net_1929), .B2(net_255), .C2(x423) );
CLKBUF_X2 inst_4536 ( .A(net_4521), .Z(net_4522) );
NOR2_X2 inst_992 ( .A1(net_3882), .A2(net_3516), .ZN(net_2529) );
OAI21_X2 inst_488 ( .B1(net_3588), .B2(net_2972), .ZN(net_2954), .A(net_2427) );
CLKBUF_X2 inst_5196 ( .A(net_5181), .Z(net_5182) );
OAI221_X2 inst_387 ( .B2(net_3795), .ZN(net_2602), .B1(net_2601), .C1(net_2521), .A(net_1386), .C2(net_316) );
OR2_X2 inst_254 ( .ZN(net_1334), .A1(net_1168), .A2(net_1167) );
CLKBUF_X2 inst_4601 ( .A(net_4586), .Z(net_4587) );
OAI21_X2 inst_654 ( .B2(net_2147), .ZN(net_1943), .B1(net_1815), .A(net_1803) );
NAND2_X2 inst_1673 ( .A1(net_3185), .ZN(net_2085), .A2(net_191) );
INV_X8 inst_2129 ( .A(net_3940), .ZN(net_516) );
NAND2_X4 inst_1412 ( .ZN(net_3342), .A1(net_3341), .A2(net_3288) );
NAND2_X2 inst_1708 ( .A2(net_4082), .ZN(net_1728), .A1(net_1726) );
NAND4_X2 inst_1181 ( .A1(net_3449), .ZN(net_2385), .A2(net_2384), .A3(net_1381), .A4(net_387) );
NOR2_X2 inst_1153 ( .ZN(net_3979), .A1(net_3659), .A2(net_283) );
AOI221_X2 inst_3823 ( .B2(net_3141), .A(net_2642), .B1(net_2591), .C1(net_2589), .ZN(net_2554), .C2(net_2553) );
CLKBUF_X2 inst_5045 ( .A(net_4505), .Z(net_5031) );
OAI221_X2 inst_391 ( .C2(net_3408), .ZN(net_2362), .B1(net_2361), .C1(net_2221), .A(net_1932), .B2(net_107) );
OAI21_X2 inst_661 ( .A(net_1912), .ZN(net_1723), .B2(net_1582), .B1(net_1300) );
AND2_X4 inst_4107 ( .A1(net_3108), .ZN(net_305), .A2(net_50) );
NAND2_X2 inst_1548 ( .A1(net_2961), .ZN(net_2474), .A2(net_487) );
NAND2_X2 inst_2073 ( .ZN(net_4007), .A1(net_3168), .A2(net_3167) );
INV_X2 inst_2738 ( .A(net_3229), .ZN(net_2690) );
CLKBUF_X2 inst_4682 ( .A(net_4620), .Z(net_4668) );
AOI21_X2 inst_3984 ( .B1(net_4106), .ZN(net_909), .A(net_908), .B2(net_246) );
OAI21_X2 inst_634 ( .ZN(net_2077), .B2(net_2076), .A(net_1962), .B1(net_1671) );
OAI221_X2 inst_419 ( .B2(net_3103), .C1(net_1614), .ZN(net_1249), .A(net_1119), .B1(net_1069), .C2(net_332) );
DFF_X2 inst_3122 ( .QN(net_3137), .D(net_2682), .CK(net_4585) );
NAND2_X4 inst_1477 ( .ZN(net_3942), .A2(net_3171), .A1(net_52) );
CLKBUF_X2 inst_5130 ( .A(net_5115), .Z(net_5116) );
AOI22_X2 inst_3717 ( .ZN(net_3566), .A2(net_3565), .A1(net_963), .B1(net_728), .B2(net_659) );
XOR2_X1 inst_34 ( .A(net_4136), .Z(net_3312), .B(net_1510) );
NAND2_X2 inst_1799 ( .ZN(net_941), .A1(net_830), .A2(net_601) );
XOR2_X2 inst_12 ( .Z(net_1289), .B(net_1288), .A(net_1087) );
OAI21_X2 inst_529 ( .B2(net_2965), .B1(net_2923), .ZN(net_2905), .A(net_2440) );
CLKBUF_X2 inst_4442 ( .A(net_4427), .Z(net_4428) );
NAND2_X2 inst_1528 ( .A1(net_3208), .ZN(net_2494), .A2(net_567) );
NAND2_X4 inst_1424 ( .ZN(net_3587), .A2(net_3586), .A1(net_3584) );
CLKBUF_X2 inst_5290 ( .A(net_5275), .Z(net_5276) );
CLKBUF_X2 inst_4694 ( .A(net_4441), .Z(net_4680) );
NAND3_X2 inst_1313 ( .A2(net_4080), .A3(net_3664), .ZN(net_945), .A1(net_943) );
NAND2_X4 inst_1425 ( .ZN(net_3601), .A2(net_3600), .A1(net_3597) );
OAI21_X2 inst_675 ( .ZN(net_1542), .B1(net_1340), .B2(net_1334), .A(net_671) );
AND3_X4 inst_4068 ( .A2(net_3925), .ZN(net_1057), .A3(net_1016), .A1(net_945) );
AND2_X4 inst_4116 ( .ZN(net_3996), .A1(net_3995), .A2(net_3167) );
INV_X2 inst_2886 ( .A(net_3035), .ZN(net_180) );
INV_X2 inst_2705 ( .ZN(net_1668), .A(net_1667) );
INV_X4 inst_2307 ( .A(net_2523), .ZN(net_2522) );
INV_X4 inst_2198 ( .A(net_2641), .ZN(net_2375) );
OR2_X2 inst_258 ( .A2(net_4103), .ZN(net_965), .A1(net_849) );
CLKBUF_X2 inst_5150 ( .A(net_5135), .Z(net_5136) );
INV_X4 inst_2611 ( .ZN(net_3823), .A(net_3820) );
CLKBUF_X2 inst_5004 ( .A(net_4767), .Z(net_4990) );
INV_X2 inst_2773 ( .ZN(net_846), .A(net_792) );
NAND2_X1 inst_2081 ( .A1(net_3532), .ZN(net_2853), .A2(net_2515) );
DFF_X1 inst_3261 ( .QN(net_3075), .D(net_2933), .CK(net_4871) );
INV_X4 inst_2405 ( .A(net_1173), .ZN(net_671) );
INV_X2 inst_2994 ( .A(net_3040), .ZN(net_195) );
INV_X2 inst_3023 ( .ZN(net_3451), .A(net_3171) );
NAND4_X2 inst_1243 ( .ZN(net_3353), .A1(net_739), .A2(net_560), .A3(net_494), .A4(net_472) );
INV_X1 inst_3076 ( .ZN(net_1055), .A(net_1054) );
NAND4_X2 inst_1211 ( .ZN(net_1248), .A2(net_1048), .A4(net_893), .A1(net_865), .A3(net_795) );
OAI21_X2 inst_482 ( .B1(net_2970), .ZN(net_2962), .B2(net_2961), .A(net_2473) );
AOI222_X1 inst_3751 ( .B1(net_4044), .C1(net_3114), .A1(net_2055), .C2(net_2053), .ZN(net_2052), .A2(net_2051), .B2(net_1190) );
NAND4_X2 inst_1192 ( .ZN(net_1906), .A4(net_1498), .A3(net_1496), .A1(net_1434), .A2(net_1429) );
OAI21_X2 inst_682 ( .ZN(net_1455), .A(net_1273), .B2(net_1154), .B1(net_1077) );
AOI22_X2 inst_3534 ( .A2(net_1908), .ZN(net_1771), .A1(net_1672), .B2(net_749), .B1(net_104) );
OR2_X4 inst_238 ( .ZN(net_3441), .A1(net_3196), .A2(net_262) );
DFF_X1 inst_3276 ( .QN(net_3036), .D(net_2908), .CK(net_5018) );
AOI21_X2 inst_3996 ( .B2(net_3804), .ZN(net_3369), .A(net_3330), .B1(net_3269) );
NOR2_X2 inst_1093 ( .A1(net_3755), .A2(net_530), .ZN(net_403) );
OAI21_X2 inst_539 ( .ZN(net_4008), .B2(net_2972), .B1(net_2893), .A(net_2433) );
INV_X4 inst_2222 ( .ZN(net_2043), .A(net_1869) );
CLKBUF_X2 inst_4578 ( .A(net_4563), .Z(net_4564) );
DFF_X1 inst_3333 ( .D(net_3357), .Q(net_3138), .CK(net_4642) );
NOR3_X2 inst_895 ( .A2(net_3486), .A1(net_1800), .ZN(net_1750), .A3(net_1686) );
AND4_X2 inst_4059 ( .ZN(net_3691), .A4(net_3690), .A1(net_3687), .A3(net_3309), .A2(net_3308) );
DFF_X2 inst_3109 ( .QN(net_2995), .D(net_2801), .CK(net_5104) );
DFF_X1 inst_3271 ( .QN(net_3100), .D(net_2924), .CK(net_5029) );
NAND2_X4 inst_1430 ( .ZN(net_3633), .A2(net_3632), .A1(net_3544) );
NAND2_X2 inst_1755 ( .ZN(net_1278), .A1(net_1277), .A2(net_1082) );
DFF_X1 inst_3257 ( .QN(net_3086), .D(net_2942), .CK(net_4723) );
INV_X4 inst_2240 ( .A(net_1653), .ZN(net_1603) );
NAND4_X2 inst_1210 ( .ZN(net_1260), .A2(net_1059), .A1(net_1053), .A3(net_1024), .A4(net_929) );
INV_X4 inst_2341 ( .A(net_3961), .ZN(net_1096) );
INV_X4 inst_2437 ( .A(net_3172), .ZN(net_198) );
OAI211_X2 inst_806 ( .ZN(net_1777), .C2(net_1776), .A(net_1683), .C1(net_1562), .B(net_1403) );
CLKBUF_X2 inst_4521 ( .A(net_4506), .Z(net_4507) );
AND2_X4 inst_4122 ( .ZN(net_4046), .A1(net_2594), .A2(net_2003) );
NAND2_X2 inst_1981 ( .ZN(net_3391), .A2(net_3389), .A1(net_3128) );
OAI21_X2 inst_763 ( .B1(net_3902), .ZN(net_3891), .B2(net_3890), .A(net_3889) );
INV_X4 inst_2330 ( .A(net_3524), .ZN(net_749) );
OAI21_X2 inst_491 ( .B1(net_3394), .B2(net_2967), .ZN(net_2951), .A(net_2406) );
CLKBUF_X2 inst_4943 ( .A(net_4928), .Z(net_4929) );
AOI22_X2 inst_3636 ( .A1(net_2220), .ZN(net_1160), .B1(net_1071), .A2(net_401), .B2(net_265) );
AOI222_X1 inst_3775 ( .ZN(net_1895), .C2(net_1874), .A1(net_1863), .B1(net_1862), .C1(net_1861), .A2(net_1797), .B2(net_1123) );
OAI21_X2 inst_537 ( .B1(net_3195), .B2(net_2959), .ZN(net_2896), .A(net_2503) );
CLKBUF_X2 inst_4797 ( .A(net_4782), .Z(net_4783) );
INV_X4 inst_2472 ( .A(net_3057), .ZN(net_488) );
OAI211_X2 inst_826 ( .ZN(net_2551), .A(net_1252), .C1(net_1206), .B(net_1186), .C2(net_347) );
INV_X1 inst_3086 ( .ZN(net_3998), .A(net_3996) );
AOI21_X2 inst_4002 ( .A(net_4146), .ZN(net_3730), .B2(net_788), .B1(net_675) );
INV_X2 inst_2791 ( .A(net_850), .ZN(net_789) );
CLKBUF_X2 inst_5069 ( .A(net_5054), .Z(net_5055) );
OR4_X2 inst_159 ( .A4(net_2596), .ZN(net_2270), .A1(net_2269), .A3(net_2268), .A2(net_1569) );
NOR4_X2 inst_872 ( .A3(net_1611), .ZN(net_369), .A4(net_355), .A1(net_286), .A2(net_84) );
CLKBUF_X2 inst_4419 ( .A(net_4229), .Z(net_4405) );
CLKBUF_X2 inst_5234 ( .A(net_5219), .Z(net_5220) );
NAND2_X2 inst_1667 ( .A1(net_2134), .ZN(net_2091), .A2(net_146) );
NAND3_X2 inst_1349 ( .ZN(net_3631), .A1(net_3630), .A2(net_3545), .A3(net_3542) );
AOI21_X2 inst_3950 ( .B1(net_3736), .ZN(net_1991), .A(net_1943), .B2(net_1507) );
OAI21_X4 inst_462 ( .A(net_3859), .B2(net_3791), .ZN(net_3517), .B1(net_3333) );
CLKBUF_X2 inst_4288 ( .A(net_4273), .Z(net_4274) );
NOR4_X2 inst_869 ( .A2(net_3841), .A3(net_3563), .ZN(net_970), .A1(net_809), .A4(net_700) );
INV_X2 inst_2646 ( .A(net_3875), .ZN(net_2315) );
XOR2_X2 inst_19 ( .Z(net_4036), .A(net_2517), .B(net_1709) );
AOI222_X1 inst_3745 ( .A1(net_4189), .C1(net_3504), .B1(net_3472), .C2(net_3385), .B2(net_3151), .ZN(net_2316), .A2(net_379) );
CLKBUF_X2 inst_4347 ( .A(net_4332), .Z(net_4333) );
CLKBUF_X2 inst_4268 ( .A(net_4220), .Z(net_4254) );
INV_X4 inst_2224 ( .ZN(net_2012), .A(net_1890) );
AOI221_X2 inst_3830 ( .B1(net_4189), .C1(net_2534), .ZN(net_2369), .A(net_2289), .B2(net_1797), .C2(net_267) );
CLKBUF_X2 inst_5226 ( .A(net_5211), .Z(net_5212) );
DFF_X1 inst_3267 ( .QN(net_3097), .D(net_2914), .CK(net_5039) );
DFF_X2 inst_3205 ( .D(net_1368), .QN(net_52), .CK(net_5263) );
NAND2_X2 inst_1686 ( .A1(net_3219), .ZN(net_1986), .A2(net_154) );
CLKBUF_X2 inst_4909 ( .A(x1012), .Z(net_4895) );
CLKBUF_X2 inst_5310 ( .A(net_5132), .Z(net_5296) );
NAND2_X2 inst_1914 ( .A2(net_322), .ZN(net_288), .A1(net_225) );
CLKBUF_X2 inst_4996 ( .A(net_4981), .Z(net_4982) );
NAND2_X2 inst_1975 ( .ZN(net_3348), .A1(net_2527), .A2(net_2374) );
NAND2_X2 inst_1890 ( .A1(net_4004), .ZN(net_825), .A2(net_655) );
INV_X4 inst_2308 ( .ZN(net_1719), .A(net_828) );
AND2_X4 inst_4093 ( .ZN(net_2803), .A1(net_2689), .A2(net_1907) );
OAI21_X2 inst_612 ( .B2(net_4130), .A(net_2296), .ZN(net_2295), .B1(net_1036) );
CLKBUF_X2 inst_4806 ( .A(net_4791), .Z(net_4792) );
INV_X2 inst_2879 ( .A(net_389), .ZN(net_164) );
NAND2_X2 inst_1789 ( .ZN(net_1001), .A2(net_1000), .A1(net_950) );
NAND2_X2 inst_1692 ( .A1(net_3293), .ZN(net_1978), .A2(net_242) );
AOI21_X2 inst_3986 ( .A(net_3968), .ZN(net_841), .B1(net_840), .B2(net_691) );
INV_X4 inst_2338 ( .A(net_1264), .ZN(net_740) );
AOI22_X2 inst_3475 ( .B1(net_4039), .ZN(net_2676), .A1(net_2675), .A2(net_333), .B2(x90) );
INV_X2 inst_3017 ( .ZN(net_3417), .A(net_3413) );
OAI211_X2 inst_845 ( .C2(net_3214), .ZN(net_1212), .B(net_1024), .A(net_926), .C1(net_849) );
AOI22_X2 inst_3554 ( .A1(net_4059), .B1(net_4056), .ZN(net_1496), .A2(net_227), .B2(net_181) );
INV_X4 inst_2455 ( .ZN(net_686), .A(net_245) );
NAND3_X2 inst_1367 ( .ZN(net_3980), .A2(net_3979), .A3(net_3604), .A1(net_3603) );
CLKBUF_X2 inst_5198 ( .A(net_5183), .Z(net_5184) );
CLKBUF_X2 inst_4828 ( .A(net_4813), .Z(net_4814) );
NAND2_X2 inst_2016 ( .ZN(net_3648), .A1(net_3647), .A2(net_189) );
CLKBUF_X2 inst_5218 ( .A(net_5203), .Z(net_5204) );
AOI22_X2 inst_3687 ( .B1(net_4123), .A1(net_555), .ZN(net_491), .B2(net_222), .A2(net_141) );
CLKBUF_X2 inst_4860 ( .A(net_4831), .Z(net_4846) );
INV_X4 inst_2287 ( .ZN(net_1517), .A(net_950) );
NAND2_X4 inst_1460 ( .ZN(net_3871), .A2(net_3870), .A1(net_3868) );
NAND3_X2 inst_1344 ( .ZN(net_3421), .A2(net_3420), .A1(net_3419), .A3(net_2611) );
NOR3_X2 inst_885 ( .A2(net_3151), .ZN(net_2749), .A1(net_2748), .A3(net_2746) );
INV_X2 inst_2630 ( .ZN(net_2765), .A(net_2764) );
AOI21_X1 inst_4012 ( .B2(net_4145), .ZN(net_3624), .A(net_3623), .B1(net_1212) );
INV_X2 inst_3053 ( .ZN(net_3902), .A(net_3901) );
NAND2_X4 inst_1443 ( .A2(net_3870), .ZN(net_3780), .A1(net_3779) );
NOR2_X2 inst_1028 ( .A1(net_4184), .ZN(net_1597), .A2(net_1504) );
OAI221_X2 inst_393 ( .C2(net_3407), .ZN(net_2359), .B1(net_2357), .C1(net_2234), .A(net_1813), .B2(net_106) );
AOI21_X2 inst_3935 ( .B2(net_3859), .ZN(net_2540), .A(net_2380), .B1(net_2367) );
CLKBUF_X2 inst_4810 ( .A(net_4795), .Z(net_4796) );
AOI22_X2 inst_3610 ( .A1(net_4062), .B1(net_4057), .ZN(net_1407), .A2(net_205), .B2(net_193) );
INV_X2 inst_2999 ( .ZN(net_251), .A(net_78) );
NAND2_X2 inst_1813 ( .A1(net_1107), .ZN(net_938), .A2(net_640) );
XNOR2_X2 inst_92 ( .ZN(net_1273), .B(net_987), .A(net_814) );
OAI22_X2 inst_345 ( .A2(net_3978), .B2(net_3681), .ZN(net_3561), .B1(net_408), .A1(net_403) );
NAND3_X4 inst_1271 ( .ZN(net_3994), .A2(net_3644), .A1(net_283), .A3(net_257) );
DFF_X2 inst_3103 ( .QN(net_3124), .D(net_2862), .CK(net_4691) );
INV_X4 inst_2321 ( .ZN(net_990), .A(net_777) );
DFF_X1 inst_3304 ( .QN(net_3020), .D(net_2866), .CK(net_5210) );
CLKBUF_X2 inst_5305 ( .A(net_5290), .Z(net_5291) );
AND2_X4 inst_4156 ( .ZN(net_4106), .A2(net_3664), .A1(net_583) );
OR2_X4 inst_200 ( .A1(net_3179), .ZN(net_2919), .A2(net_2354) );
CLKBUF_X2 inst_4425 ( .A(net_4410), .Z(net_4411) );
CLKBUF_X2 inst_4461 ( .A(net_4446), .Z(net_4447) );
CLKBUF_X2 inst_4373 ( .A(net_4358), .Z(net_4359) );
XNOR2_X2 inst_57 ( .ZN(net_2184), .A(net_2160), .B(net_1508) );
CLKBUF_X2 inst_4723 ( .A(net_4684), .Z(net_4709) );
AOI22_X2 inst_3655 ( .A2(net_3029), .B2(net_3028), .ZN(net_634), .A1(net_458), .B1(net_457) );
NAND2_X2 inst_1750 ( .ZN(net_1366), .A1(net_1365), .A2(net_1230) );
CLKBUF_X2 inst_5242 ( .A(net_5227), .Z(net_5228) );
INV_X4 inst_2236 ( .ZN(net_2547), .A(net_1690) );
DFF_X1 inst_3368 ( .D(net_3749), .CK(net_4441), .Q(x285) );
NAND2_X2 inst_1553 ( .A1(net_2961), .ZN(net_2469), .A2(net_196) );
INV_X2 inst_2843 ( .A(net_1274), .ZN(net_913) );
NAND2_X2 inst_1888 ( .A1(net_416), .ZN(net_397), .A2(net_357) );
AND2_X4 inst_4130 ( .ZN(net_4059), .A2(net_3339), .A1(net_1188) );
DFF_X1 inst_3379 ( .D(net_2250), .CK(net_5157), .Q(x639) );
NAND2_X2 inst_1763 ( .A2(net_1394), .ZN(net_1236), .A1(net_35) );
NAND2_X2 inst_1635 ( .A1(net_4041), .ZN(net_2247), .A2(net_220) );
NAND3_X2 inst_1307 ( .A3(net_1613), .ZN(net_1145), .A1(net_1014), .A2(net_967) );
NAND2_X2 inst_1500 ( .ZN(net_2810), .A1(net_2766), .A2(net_2721) );
INV_X2 inst_2805 ( .A(net_3922), .ZN(net_919) );
NOR2_X2 inst_1094 ( .A2(net_3128), .ZN(net_317), .A1(net_276) );
AOI22_X2 inst_3499 ( .B1(net_3219), .ZN(net_2136), .A1(net_2134), .A2(net_552), .B2(net_551) );
AND2_X4 inst_4145 ( .ZN(net_4082), .A1(net_1613), .A2(net_619) );
INV_X2 inst_2932 ( .ZN(net_255), .A(net_79) );
CLKBUF_X2 inst_4590 ( .A(net_4575), .Z(net_4576) );
NOR3_X2 inst_893 ( .A3(net_3157), .A2(net_2384), .ZN(net_2130), .A1(net_2065) );
AOI22_X2 inst_3680 ( .B1(net_4124), .A1(net_509), .ZN(net_503), .B2(net_200), .A2(net_140) );
INV_X2 inst_3048 ( .ZN(net_3744), .A(net_3743) );
CLKBUF_X2 inst_4878 ( .A(net_4863), .Z(net_4864) );
CLKBUF_X2 inst_4854 ( .A(net_4839), .Z(net_4840) );
NAND2_X2 inst_1699 ( .A1(net_3505), .ZN(net_1835), .A2(net_1834) );
OAI211_X2 inst_851 ( .A(net_4153), .ZN(net_3320), .C2(net_3319), .C1(net_3318), .B(net_3317) );
OAI211_X2 inst_831 ( .ZN(net_1361), .C1(net_1359), .A(net_1234), .B(net_593), .C2(net_318) );
XNOR2_X2 inst_50 ( .ZN(net_2621), .A(net_2531), .B(net_294) );
DFF_X1 inst_3346 ( .D(net_2755), .CK(net_4349), .Q(x60) );
OAI21_X2 inst_569 ( .B2(net_3207), .B1(net_2849), .ZN(net_2843), .A(net_2481) );
INV_X2 inst_2992 ( .A(net_3042), .ZN(net_176) );
CLKBUF_X2 inst_4264 ( .A(net_4208), .Z(net_4250) );
INV_X4 inst_2589 ( .A(net_3711), .ZN(net_3671) );
NOR2_X2 inst_1080 ( .A1(net_3958), .ZN(net_838), .A2(net_605) );
INV_X4 inst_2374 ( .A(net_3670), .ZN(net_583) );
NOR2_X2 inst_1103 ( .A1(net_3161), .ZN(net_158), .A2(net_84) );
CLKBUF_X2 inst_4430 ( .A(net_4415), .Z(net_4416) );
CLKBUF_X2 inst_4329 ( .A(net_4314), .Z(net_4315) );
NAND2_X2 inst_1650 ( .ZN(net_2154), .A1(net_2153), .A2(net_321) );
OAI21_X2 inst_549 ( .B2(net_2907), .B1(net_2887), .ZN(net_2882), .A(net_2485) );
CLKBUF_X2 inst_4708 ( .A(net_4693), .Z(net_4694) );
CLKBUF_X2 inst_4220 ( .A(net_4205), .Z(net_4206) );
NAND2_X2 inst_1497 ( .ZN(net_2820), .A1(net_2772), .A2(net_2719) );
OAI21_X2 inst_522 ( .B1(net_3302), .ZN(net_2916), .B2(net_2915), .A(net_2436) );
CLKBUF_X2 inst_5202 ( .A(net_5134), .Z(net_5188) );
CLKBUF_X2 inst_5040 ( .A(net_4273), .Z(net_5026) );
CLKBUF_X2 inst_4439 ( .A(net_4424), .Z(net_4425) );
INV_X2 inst_2872 ( .ZN(net_254), .A(net_253) );
NOR2_X2 inst_1002 ( .A1(net_3772), .ZN(net_2230), .A2(net_1746) );
INV_X2 inst_2809 ( .ZN(net_840), .A(net_680) );
OAI21_X2 inst_478 ( .ZN(net_2971), .B1(net_2970), .B2(net_2969), .A(net_2416) );
DFF_X1 inst_3380 ( .D(net_2253), .Q(net_76), .CK(net_5296) );
INV_X2 inst_2673 ( .ZN(net_1901), .A(net_1900) );
NAND2_X2 inst_1618 ( .A1(net_2919), .ZN(net_2398), .A2(net_187) );
CLKBUF_X2 inst_5062 ( .A(net_4344), .Z(net_5048) );
INV_X8 inst_2126 ( .ZN(net_509), .A(net_351) );
OAI211_X2 inst_804 ( .C1(net_2190), .ZN(net_2123), .C2(net_2122), .A(net_2013), .B(net_2000) );
DFF_X1 inst_3290 ( .QN(net_3046), .D(net_2897), .CK(net_4712) );
XOR2_X2 inst_13 ( .A(net_4074), .B(net_1148), .Z(net_1140) );
INV_X4 inst_2584 ( .ZN(net_3629), .A(net_3211) );
CLKBUF_X2 inst_4931 ( .A(net_4916), .Z(net_4917) );
AOI22_X2 inst_3600 ( .A1(net_4063), .B1(net_4058), .ZN(net_1417), .A2(net_559), .B2(net_558) );
INV_X2 inst_2765 ( .ZN(net_2165), .A(net_951) );
OAI211_X2 inst_799 ( .C1(net_2190), .ZN(net_2188), .C2(net_2187), .B(net_2056), .A(net_2009) );
AOI22_X2 inst_3481 ( .B1(net_4038), .A1(net_2675), .ZN(net_2656), .A2(net_984), .B2(net_402) );
OR2_X4 inst_219 ( .ZN(net_949), .A1(net_948), .A2(net_908) );
OAI21_X2 inst_738 ( .B2(net_3124), .ZN(net_310), .A(net_309), .B1(net_164) );
OAI21_X2 inst_719 ( .B1(net_3929), .ZN(net_724), .A(net_669), .B2(net_334) );
AND2_X4 inst_4166 ( .ZN(net_4120), .A2(net_404), .A1(net_248) );
INV_X2 inst_2755 ( .ZN(net_1003), .A(net_1002) );
CLKBUF_X2 inst_4881 ( .A(net_4866), .Z(net_4867) );
NAND2_X2 inst_1819 ( .ZN(net_871), .A1(net_817), .A2(net_766) );
AOI221_X2 inst_3868 ( .B2(net_3118), .B1(net_2020), .C1(net_2019), .ZN(net_1938), .A(net_1937), .C2(x232) );
OR2_X2 inst_255 ( .A2(net_4119), .ZN(net_1161), .A1(net_932) );
INV_X2 inst_2726 ( .A(net_2212), .ZN(net_2042) );
OAI21_X4 inst_453 ( .ZN(net_2160), .B1(net_2043), .A(net_1595), .B2(net_1505) );
NOR2_X2 inst_1134 ( .A1(net_3722), .ZN(net_3666), .A2(net_3665) );
OAI21_X2 inst_493 ( .B1(net_3394), .B2(net_2965), .ZN(net_2949), .A(net_2442) );
INV_X2 inst_2674 ( .ZN(net_1899), .A(net_1898) );
INV_X4 inst_2204 ( .A(net_3511), .ZN(net_2364) );
XOR2_X2 inst_23 ( .Z(net_4092), .A(net_681), .B(net_387) );
NOR2_X2 inst_1113 ( .A2(net_3515), .A1(net_3405), .ZN(net_3332) );
NAND2_X2 inst_1822 ( .A2(net_3900), .ZN(net_1008), .A1(net_902) );
NAND2_X2 inst_1609 ( .A1(net_2967), .ZN(net_2407), .A2(net_471) );
AND2_X4 inst_4105 ( .A1(net_4128), .A2(net_3163), .ZN(net_457) );
AOI222_X1 inst_3790 ( .B1(net_4115), .C1(net_1882), .A1(net_1385), .ZN(net_1056), .A2(net_894), .B2(net_844), .C2(net_122) );
AND2_X2 inst_4206 ( .ZN(net_3446), .A2(net_2518), .A1(net_1051) );
AOI22_X2 inst_3546 ( .B1(net_4054), .A1(net_1578), .ZN(net_1576), .A2(net_379), .B2(net_238) );
OAI221_X2 inst_408 ( .B2(net_4071), .C2(net_3123), .ZN(net_1666), .B1(net_1615), .A(net_816), .C1(net_437) );
NOR2_X2 inst_1144 ( .ZN(net_3893), .A1(net_3892), .A2(net_3867) );
CLKBUF_X2 inst_5165 ( .A(net_5132), .Z(net_5151) );
CLKBUF_X2 inst_4701 ( .A(net_4686), .Z(net_4687) );
OAI211_X2 inst_812 ( .C2(net_3755), .B(net_1628), .C1(net_1627), .ZN(net_1626), .A(net_1554) );
INV_X4 inst_2568 ( .ZN(net_3541), .A(net_3540) );
INV_X4 inst_2295 ( .A(net_1261), .ZN(net_898) );
OR3_X2 inst_179 ( .A2(net_4075), .ZN(net_2561), .A1(net_2528), .A3(net_2522) );
NAND2_X2 inst_1730 ( .A1(net_1556), .ZN(net_1555), .A2(x800) );
AOI221_X2 inst_3799 ( .ZN(net_2782), .C1(net_2781), .B1(net_2775), .A(net_2685), .C2(net_1699), .B2(net_292) );
AOI221_X2 inst_3814 ( .C1(net_3445), .A(net_2642), .ZN(net_2586), .B1(net_2584), .C2(net_2583), .B2(net_1326) );
AOI222_X2 inst_3734 ( .A2(net_1826), .ZN(net_1765), .A1(net_1387), .B2(net_991), .C2(net_920), .B1(net_624), .C1(net_580) );
AOI22_X2 inst_3532 ( .B1(net_2625), .ZN(net_1839), .A1(net_1838), .A2(net_1837), .B2(net_184) );
INV_X2 inst_3028 ( .ZN(net_3506), .A(net_3505) );
INV_X4 inst_2191 ( .ZN(net_2383), .A(net_2382) );
XNOR2_X2 inst_76 ( .A(net_3229), .ZN(net_1448), .B(net_1447) );
CLKBUF_X2 inst_5296 ( .A(net_5281), .Z(net_5282) );
AOI221_X2 inst_3854 ( .B1(net_3736), .ZN(net_2058), .C1(net_2049), .C2(net_1902), .A(net_1854), .B2(net_240) );
NOR2_X2 inst_1127 ( .A2(net_4155), .A1(net_3597), .ZN(net_3474) );
AOI22_X2 inst_3514 ( .B1(net_4045), .ZN(net_1957), .A1(net_1955), .A2(net_265), .B2(net_228) );
OR3_X4 inst_172 ( .ZN(net_2523), .A2(net_988), .A1(net_843), .A3(net_526) );
OAI221_X2 inst_362 ( .ZN(net_2783), .A(net_2726), .C1(net_2565), .B1(net_2561), .B2(net_2051), .C2(net_1537) );
CLKBUF_X2 inst_4366 ( .A(net_4351), .Z(net_4352) );
NAND2_X2 inst_1530 ( .A1(net_3208), .ZN(net_2492), .A2(net_558) );
OAI22_X4 inst_277 ( .B1(net_3871), .ZN(net_3216), .A1(net_3177), .B2(net_3002), .A2(net_3001) );
NAND2_X2 inst_1510 ( .ZN(net_2735), .A1(net_2624), .A2(net_2623) );
XNOR2_X2 inst_83 ( .ZN(net_1139), .A(net_1138), .B(net_1137) );
XNOR2_X2 inst_121 ( .ZN(net_4137), .B(net_322), .A(net_192) );
OAI22_X2 inst_306 ( .A2(net_2665), .A1(net_1543), .B1(net_1542), .ZN(net_1534), .B2(net_130) );
AND2_X4 inst_4186 ( .ZN(net_4180), .A2(net_4179), .A1(net_4178) );
NOR2_X2 inst_1065 ( .A2(net_923), .ZN(net_897), .A1(net_853) );
AND2_X4 inst_4119 ( .A2(net_4050), .ZN(net_4042), .A1(net_1959) );
CLKBUF_X2 inst_4332 ( .A(net_4317), .Z(net_4318) );
DFF_X1 inst_3386 ( .D(net_1805), .QN(net_39), .CK(net_5002) );
HA_X1 inst_3095 ( .S(net_1035), .CO(net_875), .B(net_874), .A(net_676) );
NAND2_X2 inst_1715 ( .A1(net_3492), .ZN(net_1785), .A2(net_1640) );
SDFF_X2 inst_140 ( .SE(net_2625), .D(net_2336), .SI(net_98), .Q(net_98), .CK(net_4954) );
OR2_X2 inst_267 ( .ZN(net_3355), .A2(net_3354), .A1(net_3352) );
INV_X2 inst_2824 ( .ZN(net_638), .A(net_517) );
OAI21_X2 inst_716 ( .B1(net_4125), .ZN(net_776), .A(net_775), .B2(net_644) );
CLKBUF_X2 inst_4671 ( .A(net_4656), .Z(net_4657) );
AOI22_X2 inst_3594 ( .A1(net_4059), .B1(net_4057), .ZN(net_1423), .B2(net_222), .A2(net_202) );
AND2_X4 inst_4174 ( .ZN(net_4128), .A2(net_3162), .A1(net_223) );
NAND2_X2 inst_1906 ( .ZN(net_314), .A2(net_303), .A1(net_198) );
OAI21_X2 inst_530 ( .B2(net_2963), .B1(net_2923), .ZN(net_2904), .A(net_2454) );
OAI211_X2 inst_792 ( .C2(net_2876), .ZN(net_2701), .A(net_2622), .C1(net_2621), .B(net_2139) );
NAND2_X2 inst_2024 ( .ZN(net_3719), .A2(net_3715), .A1(net_3682) );
DFF_X2 inst_3124 ( .D(net_2646), .QN(net_112), .CK(net_4396) );
INV_X2 inst_2952 ( .A(net_3101), .ZN(net_161) );
NAND3_X2 inst_1353 ( .ZN(net_3688), .A1(net_3687), .A3(net_3309), .A2(net_3308) );
INV_X4 inst_2502 ( .ZN(net_2037), .A(net_289) );
INV_X4 inst_2216 ( .ZN(net_2235), .A(net_2137) );
OAI21_X2 inst_769 ( .ZN(net_3966), .A(net_3960), .B1(net_1212), .B2(net_851) );
OR3_X4 inst_174 ( .ZN(net_627), .A3(net_389), .A2(net_344), .A1(net_309) );
NAND4_X2 inst_1200 ( .ZN(net_1767), .A3(net_1477), .A4(net_1476), .A1(net_1411), .A2(net_1410) );
INV_X2 inst_2988 ( .A(net_292), .ZN(net_142) );
CLKBUF_X2 inst_4494 ( .A(net_4479), .Z(net_4480) );
MUX2_X2 inst_2105 ( .S(net_2917), .A(net_2573), .Z(net_2572), .B(net_230) );
NAND4_X2 inst_1199 ( .ZN(net_1674), .A3(net_1495), .A4(net_1494), .A1(net_1428), .A2(net_1427) );
XOR2_X2 inst_5 ( .A(net_3492), .Z(net_1695), .B(net_1694) );
AOI21_X2 inst_3974 ( .ZN(net_1177), .A(net_1176), .B2(net_1011), .B1(net_846) );
INV_X2 inst_3021 ( .A(net_3634), .ZN(net_3440) );
OAI21_X2 inst_729 ( .A(net_629), .B1(net_628), .ZN(net_581), .B2(net_333) );
INV_X8 inst_2157 ( .A(net_3898), .ZN(net_3618) );
NAND2_X2 inst_1662 ( .ZN(net_2101), .A1(net_2099), .A2(net_241) );
CLKBUF_X2 inst_4553 ( .A(net_4538), .Z(net_4539) );
INV_X2 inst_2783 ( .ZN(net_803), .A(net_757) );
OR2_X4 inst_213 ( .A1(net_3781), .ZN(net_1815), .A2(net_711) );
OAI21_X2 inst_604 ( .B2(net_3486), .ZN(net_2334), .B1(net_2330), .A(net_1946) );
OR2_X4 inst_205 ( .ZN(net_2915), .A2(net_2354), .A1(net_2350) );
NAND2_X2 inst_1645 ( .A1(net_3190), .A2(net_3181), .ZN(net_2170) );
NAND3_X2 inst_1285 ( .ZN(net_2262), .A1(net_2204), .A3(net_1957), .A2(net_1916) );
OAI221_X2 inst_380 ( .C2(net_4088), .B2(net_2733), .C1(net_2686), .ZN(net_2652), .A(net_2588), .B1(net_2538) );
AND4_X2 inst_4057 ( .A3(net_2737), .ZN(net_1380), .A1(net_1221), .A2(net_977), .A4(net_314) );
NAND4_X2 inst_1179 ( .ZN(net_2854), .A2(net_2823), .A1(net_2812), .A3(net_2793), .A4(net_2753) );
AOI22_X2 inst_3722 ( .A2(net_4145), .ZN(net_3622), .B2(net_3621), .B1(net_845), .A1(net_743) );
OAI22_X2 inst_292 ( .A1(net_3781), .B1(net_1884), .ZN(net_1811), .A2(net_1810), .B2(net_389) );
CLKBUF_X2 inst_4311 ( .A(net_4296), .Z(net_4297) );
AOI22_X2 inst_3650 ( .ZN(net_736), .A1(net_735), .B1(net_734), .A2(net_458), .B2(net_457) );
NAND2_X2 inst_2012 ( .ZN(net_3593), .A2(net_3592), .A1(net_3591) );
AOI221_X2 inst_3911 ( .A(net_4113), .ZN(net_701), .B1(net_686), .C2(net_393), .B2(net_329), .C1(net_245) );
NAND2_X2 inst_1515 ( .ZN(net_2537), .A1(net_2367), .A2(net_2195) );
CLKBUF_X2 inst_4970 ( .A(net_4955), .Z(net_4956) );
OAI21_X2 inst_706 ( .ZN(net_873), .A(net_769), .B2(net_768), .B1(net_206) );
CLKBUF_X2 inst_5173 ( .A(net_5158), .Z(net_5159) );
NAND2_X2 inst_1782 ( .A2(net_3559), .ZN(net_2127), .A1(net_1183) );
INV_X2 inst_2951 ( .ZN(net_209), .A(net_106) );
CLKBUF_X2 inst_4472 ( .A(net_4225), .Z(net_4458) );
AOI221_X2 inst_3890 ( .B1(net_4027), .C1(net_3111), .A(net_2525), .ZN(net_1395), .B2(net_1394), .C2(net_1393) );
OAI211_X2 inst_839 ( .C1(net_1359), .ZN(net_1349), .A(net_1238), .B(net_671), .C2(net_302) );
NOR2_X2 inst_1015 ( .A1(net_1738), .ZN(net_1736), .A2(net_1632) );
CLKBUF_X2 inst_4734 ( .A(net_4719), .Z(net_4720) );
OR2_X4 inst_240 ( .A1(net_3959), .A2(net_3720), .ZN(net_3681) );
AOI21_X2 inst_3966 ( .B2(net_3968), .B1(net_1884), .ZN(net_1389), .A(net_1388) );
XNOR2_X2 inst_110 ( .ZN(net_538), .A(net_309), .B(net_47) );
AOI221_X2 inst_3899 ( .B2(net_4107), .B1(net_3561), .ZN(net_1209), .C2(net_1011), .C1(net_961), .A(net_864) );
NAND2_X2 inst_2047 ( .ZN(net_3860), .A2(net_3859), .A1(net_3857) );
DFF_X2 inst_3213 ( .D(net_807), .QN(net_327), .CK(net_4794) );
CLKBUF_X2 inst_4545 ( .A(net_4530), .Z(net_4531) );
AOI221_X2 inst_3825 ( .B1(net_3469), .B2(net_3147), .ZN(net_2536), .C1(net_2534), .A(net_2340), .C2(net_252) );
INV_X4 inst_2535 ( .A(net_3877), .ZN(net_3343) );
XNOR2_X2 inst_99 ( .A(net_729), .ZN(net_653), .B(net_387) );
CLKBUF_X2 inst_4569 ( .A(net_4554), .Z(net_4555) );
NAND2_X2 inst_1661 ( .A2(net_4019), .ZN(net_2102), .A1(net_2099) );
CLKBUF_X2 inst_4384 ( .A(net_4369), .Z(net_4370) );
NAND2_X2 inst_2059 ( .ZN(net_3908), .A1(net_3187), .A2(net_186) );
CLKBUF_X2 inst_4480 ( .A(net_4237), .Z(net_4466) );
INV_X2 inst_2949 ( .A(net_3047), .ZN(net_212) );
INV_X4 inst_2414 ( .ZN(net_276), .A(net_262) );
OAI22_X2 inst_283 ( .A1(net_3883), .A2(net_3859), .B2(net_3858), .ZN(net_2372), .B1(net_2371) );
OAI22_X2 inst_311 ( .B1(net_4077), .B2(net_3789), .ZN(net_1774), .A1(net_1050), .A2(net_877) );
DFF_X1 inst_3406 ( .Q(net_4028), .D(net_1396), .CK(net_4504) );
INV_X4 inst_2519 ( .A(net_3391), .ZN(net_3220) );
NAND2_X2 inst_1597 ( .A1(net_2925), .ZN(net_2421), .A2(net_169) );
AOI22_X2 inst_3502 ( .ZN(net_2057), .A1(net_1903), .B2(net_1719), .A2(net_1717), .B1(net_1621) );
INV_X4 inst_2203 ( .A(net_3248), .ZN(net_2543) );
AOI22_X2 inst_3473 ( .A2(net_3149), .B2(net_3113), .A1(net_2775), .B1(net_2722), .ZN(net_2713) );
OAI221_X2 inst_431 ( .B2(net_3620), .A(net_1007), .ZN(net_905), .B1(net_904), .C2(net_903), .C1(net_638) );
OAI222_X2 inst_348 ( .A2(net_2815), .ZN(net_1819), .A1(net_1818), .B1(net_1817), .C1(net_1816), .C2(net_289), .B2(net_107) );
NAND2_X2 inst_1930 ( .A2(net_4011), .ZN(net_3193), .A1(net_3186) );
NOR3_X2 inst_889 ( .ZN(net_2781), .A1(net_2528), .A2(net_1168), .A3(net_1124) );
OAI21_X2 inst_577 ( .B2(net_2915), .B1(net_2803), .ZN(net_2801), .A(net_2448) );
CLKBUF_X2 inst_5123 ( .A(net_5108), .Z(net_5109) );
INV_X2 inst_2686 ( .A(net_3407), .ZN(net_1888) );
CLKBUF_X2 inst_4975 ( .A(net_4960), .Z(net_4961) );
AOI222_X1 inst_3740 ( .C1(net_4039), .B1(net_4038), .ZN(net_2617), .A1(net_2594), .A2(net_2346), .B2(net_1523), .C2(x105) );
INV_X4 inst_2293 ( .ZN(net_2122), .A(net_906) );
CLKBUF_X2 inst_5188 ( .A(net_5173), .Z(net_5174) );
INV_X4 inst_2379 ( .A(net_3438), .ZN(net_923) );
NAND3_X2 inst_1364 ( .ZN(net_3924), .A3(net_3923), .A2(net_3627), .A1(net_963) );
AOI21_X2 inst_3938 ( .ZN(net_2330), .B1(net_2283), .B2(net_2144), .A(net_1778) );
INV_X2 inst_2865 ( .ZN(net_991), .A(net_47) );
OAI21_X2 inst_645 ( .ZN(net_1949), .B1(net_1912), .A(net_1873), .B2(net_1292) );
CLKBUF_X2 inst_4916 ( .A(net_4901), .Z(net_4902) );
CLKBUF_X2 inst_4891 ( .A(net_4224), .Z(net_4877) );
AOI22_X2 inst_3571 ( .A1(net_4059), .B1(net_4056), .ZN(net_1479), .B2(net_468), .A2(net_453) );
INV_X2 inst_3041 ( .A(net_3711), .ZN(net_3673) );
INV_X2 inst_2719 ( .ZN(net_2669), .A(net_2551) );
INV_X4 inst_2352 ( .ZN(net_618), .A(net_513) );
OR2_X2 inst_269 ( .A2(net_3447), .ZN(net_3426), .A1(net_1606) );
NAND4_X2 inst_1190 ( .ZN(net_1823), .A3(net_1493), .A4(net_1492), .A1(net_1426), .A2(net_1425) );
OAI221_X2 inst_444 ( .B1(net_4159), .ZN(net_3696), .B2(net_3407), .C1(net_2328), .A(net_1935), .C2(net_1447) );
INV_X4 inst_2544 ( .A(net_3674), .ZN(net_3667) );
OAI21_X2 inst_514 ( .B1(net_3278), .ZN(net_2928), .B2(net_2912), .A(net_2449) );
CLKBUF_X2 inst_4905 ( .A(net_4890), .Z(net_4891) );
NAND2_X2 inst_1541 ( .A1(net_3207), .ZN(net_2481), .A2(net_160) );
CLKBUF_X2 inst_4236 ( .A(net_4221), .Z(net_4222) );
OAI21_X2 inst_685 ( .B1(net_3228), .ZN(net_1310), .A(net_1259), .B2(net_260) );
XNOR2_X2 inst_63 ( .A(net_3264), .ZN(net_1902), .B(net_1526) );
XNOR2_X2 inst_119 ( .ZN(net_4074), .A(net_701), .B(net_402) );
DFF_X2 inst_3181 ( .D(net_1811), .QN(net_389), .CK(net_4837) );
NOR2_X4 inst_939 ( .ZN(net_3227), .A1(net_915), .A2(net_877) );
CLKBUF_X2 inst_4656 ( .A(net_4641), .Z(net_4642) );
NAND4_X2 inst_1233 ( .ZN(net_1637), .A4(net_550), .A3(net_545), .A1(net_503), .A2(net_473) );
INV_X2 inst_2924 ( .A(net_3002), .ZN(net_160) );
NOR2_X2 inst_1019 ( .A1(net_1815), .ZN(net_1812), .A2(net_1655) );
NAND2_X2 inst_2006 ( .A2(net_3859), .ZN(net_3534), .A1(net_3533) );
NAND2_X2 inst_1827 ( .ZN(net_779), .A1(net_778), .A2(net_777) );
OAI21_X2 inst_742 ( .B1(net_3611), .B2(net_3516), .A(net_3344), .ZN(net_3286) );
OAI221_X2 inst_427 ( .B2(net_4133), .B1(net_3733), .ZN(net_1061), .A(net_953), .C2(net_904), .C1(net_680) );
AOI221_X2 inst_3840 ( .ZN(net_2204), .B2(net_2203), .C1(net_2202), .A(net_2074), .C2(net_2037), .B1(net_1906) );
INV_X4 inst_2619 ( .A(net_3991), .ZN(net_3923) );
AOI22_X2 inst_3465 ( .B2(net_4026), .ZN(net_2753), .B1(net_2752), .A1(net_2750), .A2(net_361) );
NAND2_X2 inst_2033 ( .ZN(net_3768), .A1(net_3168), .A2(net_3108) );
INV_X8 inst_2144 ( .A(net_3871), .ZN(net_3219) );
CLKBUF_X2 inst_4481 ( .A(net_4466), .Z(net_4467) );
INV_X4 inst_2559 ( .ZN(net_3505), .A(net_3503) );
SDFF_X2 inst_138 ( .D(net_3290), .SE(net_2625), .SI(net_96), .Q(net_96), .CK(net_4957) );
CLKBUF_X2 inst_5289 ( .A(net_5274), .Z(net_5275) );
NAND2_X2 inst_1955 ( .ZN(net_3284), .A2(net_3186), .A1(net_172) );
INV_X2 inst_2810 ( .ZN(net_669), .A(net_407) );
AOI22_X2 inst_3618 ( .B1(net_3134), .ZN(net_1640), .B2(net_1071), .A1(net_1044), .A2(net_1036) );
NAND3_X4 inst_1269 ( .A3(net_4149), .ZN(net_3951), .A1(net_3950), .A2(net_3790) );
CLKBUF_X2 inst_4944 ( .A(net_4929), .Z(net_4930) );
NOR3_X2 inst_899 ( .A2(net_4072), .A3(net_3935), .ZN(net_1187), .A1(net_1054) );
OAI22_X2 inst_312 ( .A1(net_2384), .B1(net_1274), .ZN(net_1218), .A2(net_1217), .B2(net_773) );
DFF_X1 inst_3241 ( .QN(net_3045), .D(net_2957), .CK(net_5182) );
INV_X2 inst_2704 ( .ZN(net_1671), .A(net_1670) );
NAND2_X2 inst_1620 ( .A1(net_2917), .ZN(net_2396), .A2(net_166) );
CLKBUF_X2 inst_4958 ( .A(net_4487), .Z(net_4944) );
OAI22_X2 inst_309 ( .B2(net_3102), .B1(net_1884), .ZN(net_1303), .A1(net_1159), .A2(net_1090) );
DFF_X1 inst_3416 ( .D(net_1353), .Q(net_33), .CK(net_4334) );
OAI222_X2 inst_347 ( .A2(net_2815), .ZN(net_1997), .A1(net_1996), .B1(net_1817), .C1(net_1816), .C2(net_505), .B2(net_108) );
INV_X8 inst_2149 ( .ZN(net_3293), .A(net_3292) );
OAI21_X2 inst_755 ( .ZN(net_3707), .A(net_3706), .B2(net_3407), .B1(net_2228) );
CLKBUF_X2 inst_5001 ( .A(net_4590), .Z(net_4987) );
NAND2_X2 inst_1724 ( .A2(net_3490), .ZN(net_1594), .A1(net_1593) );
CLKBUF_X2 inst_4505 ( .A(net_4485), .Z(net_4491) );
INV_X4 inst_2610 ( .A(net_3823), .ZN(net_3822) );
INV_X2 inst_2694 ( .ZN(net_1716), .A(net_1680) );
NOR2_X2 inst_1043 ( .A1(net_1196), .ZN(net_1182), .A2(net_1116) );
AOI211_X2 inst_4030 ( .B(net_3916), .A(net_3656), .C1(net_889), .ZN(net_708), .C2(net_607) );
NAND2_X2 inst_1968 ( .ZN(net_3335), .A1(net_3280), .A2(net_493) );
CLKBUF_X2 inst_4817 ( .A(net_4802), .Z(net_4803) );
CLKBUF_X2 inst_4456 ( .A(net_4300), .Z(net_4442) );
CLKBUF_X2 inst_4926 ( .A(net_4911), .Z(net_4912) );
AND3_X4 inst_4078 ( .ZN(net_4098), .A3(net_3913), .A1(net_432), .A2(net_418) );
AND3_X4 inst_4067 ( .A1(net_4194), .ZN(net_1321), .A3(net_1254), .A2(net_1133) );
NAND2_X2 inst_1792 ( .ZN(net_975), .A1(net_974), .A2(net_145) );
CLKBUF_X2 inst_4426 ( .A(net_4206), .Z(net_4412) );
NAND3_X2 inst_1330 ( .A3(net_4125), .A1(net_3523), .ZN(net_711), .A2(net_407) );
CLKBUF_X2 inst_4571 ( .A(net_4556), .Z(net_4557) );
CLKBUF_X2 inst_5111 ( .A(net_5096), .Z(net_5097) );
AOI21_X4 inst_3928 ( .B2(net_3600), .ZN(net_3588), .B1(net_3587), .A(net_2186) );
DFF_X1 inst_3353 ( .D(net_2629), .QN(net_41), .CK(net_4338) );
NAND2_X2 inst_1898 ( .ZN(net_394), .A2(net_307), .A1(net_293) );
AOI22_X2 inst_3634 ( .ZN(net_932), .B1(net_931), .A1(net_869), .A2(net_401), .B2(net_252) );
AOI221_X2 inst_3883 ( .C1(net_3782), .B1(net_1882), .C2(net_1834), .ZN(net_1802), .A(net_1648), .B2(net_84) );
AOI211_X2 inst_4017 ( .ZN(net_1775), .A(net_1774), .B(net_1682), .C2(net_1383), .C1(net_1071) );
NAND2_X2 inst_1714 ( .ZN(net_2298), .A2(net_1568), .A1(net_1566) );
CLKBUF_X2 inst_4598 ( .A(net_4583), .Z(net_4584) );
CLKBUF_X2 inst_4681 ( .A(net_4548), .Z(net_4667) );
CLKBUF_X2 inst_5135 ( .A(net_5120), .Z(net_5121) );
CLKBUF_X2 inst_4777 ( .A(net_4710), .Z(net_4763) );
NAND2_X2 inst_1496 ( .ZN(net_2821), .A1(net_2776), .A2(net_2725) );
CLKBUF_X2 inst_4297 ( .A(net_4282), .Z(net_4283) );
NAND2_X2 inst_1565 ( .A1(net_2963), .ZN(net_2456), .A2(net_453) );
NOR2_X4 inst_924 ( .A2(net_3400), .A1(net_3236), .ZN(net_2280) );
CLKBUF_X2 inst_5095 ( .A(net_4483), .Z(net_5081) );
OAI22_X2 inst_287 ( .A1(net_3781), .ZN(net_1885), .B1(net_1884), .A2(net_1761), .B2(net_270) );
OAI221_X2 inst_426 ( .A(net_3731), .ZN(net_1130), .C1(net_1129), .B2(net_887), .B1(net_798), .C2(net_721) );
DFF_X2 inst_3145 ( .QN(net_3105), .D(net_2508), .CK(net_5150) );
INV_X4 inst_2577 ( .ZN(net_3595), .A(net_3592) );
CLKBUF_X2 inst_5144 ( .A(net_4572), .Z(net_5130) );
OAI21_X2 inst_648 ( .B2(net_3338), .ZN(net_1926), .A(net_1839), .B1(net_1838) );
HA_X1 inst_3094 ( .CO(net_1085), .S(net_1038), .A(net_820), .B(net_229) );
INV_X2 inst_2903 ( .A(net_3030), .ZN(net_233) );
OR2_X2 inst_270 ( .ZN(net_3737), .A1(net_3428), .A2(net_3229) );
AND4_X4 inst_4045 ( .ZN(net_4053), .A1(net_3228), .A4(net_1386), .A2(net_1115), .A3(net_1111) );
NAND2_X2 inst_1901 ( .ZN(net_353), .A1(net_350), .A2(net_144) );
CLKBUF_X2 inst_4302 ( .A(net_4287), .Z(net_4288) );
CLKBUF_X2 inst_4890 ( .A(net_4774), .Z(net_4876) );
NOR2_X2 inst_984 ( .ZN(net_2750), .A1(net_2609), .A2(net_1270) );
AOI221_X2 inst_3804 ( .C1(net_2781), .B1(net_2775), .ZN(net_2766), .A(net_2639), .B2(net_2637), .C2(net_206) );
NAND2_X2 inst_2064 ( .ZN(net_3941), .A2(net_3109), .A1(net_352) );
AND2_X4 inst_4104 ( .ZN(net_778), .A1(net_413), .A2(net_412) );
INV_X4 inst_2266 ( .ZN(net_1232), .A(net_1049) );
NAND3_X2 inst_1292 ( .A2(net_4121), .A1(net_4043), .ZN(net_2206), .A3(net_2180) );
INV_X4 inst_2552 ( .ZN(net_3471), .A(net_2126) );
CLKBUF_X2 inst_5014 ( .A(net_4999), .Z(net_5000) );
NAND2_X2 inst_1963 ( .ZN(net_3316), .A1(net_3315), .A2(net_330) );
OAI21_X2 inst_631 ( .B2(net_2525), .ZN(net_2231), .A(net_2119), .B1(net_2118) );
NOR2_X2 inst_1056 ( .A2(net_4076), .ZN(net_1108), .A1(net_661) );
CLKBUF_X2 inst_4247 ( .A(net_4232), .Z(net_4233) );
AOI22_X2 inst_3648 ( .A1(net_1011), .ZN(net_798), .B1(net_432), .A2(net_408), .B2(net_403) );
AOI22_X2 inst_3674 ( .A2(net_571), .B2(net_570), .ZN(net_547), .B1(net_235), .A1(net_232) );
INV_X4 inst_2514 ( .A(net_3886), .ZN(net_3175) );
CLKBUF_X2 inst_4988 ( .A(net_4973), .Z(net_4974) );
AOI21_X2 inst_3995 ( .ZN(net_3296), .B1(net_3295), .B2(net_2578), .A(net_2343) );
NOR2_X2 inst_1128 ( .A2(net_3568), .ZN(net_3525), .A1(net_434) );
CLKBUF_X2 inst_4211 ( .A(x1012), .Z(net_4197) );
AOI222_X1 inst_3759 ( .C1(net_4045), .ZN(net_2004), .B1(net_1968), .A1(net_1849), .A2(net_1836), .B2(net_1511), .C2(net_179) );
DFF_X1 inst_3222 ( .QN(net_3058), .D(net_2974), .CK(net_4566) );
CLKBUF_X2 inst_5074 ( .A(net_5059), .Z(net_5060) );
NAND2_X2 inst_1745 ( .ZN(net_1465), .A2(net_1386), .A1(net_1336) );
AOI221_X2 inst_3831 ( .B1(net_4189), .C1(net_2534), .ZN(net_2368), .A(net_2290), .B2(net_378), .C2(net_280) );
NAND2_X2 inst_2079 ( .ZN(net_4168), .A1(net_3736), .A2(net_73) );
XNOR2_X2 inst_102 ( .ZN(net_681), .A(net_322), .B(net_49) );
INV_X4 inst_2527 ( .ZN(net_3270), .A(net_3130) );
DFF_X1 inst_3277 ( .QN(net_3035), .D(net_2916), .CK(net_5014) );
AND3_X4 inst_4070 ( .A2(net_3819), .ZN(net_3619), .A3(net_3196), .A1(net_262) );
INV_X2 inst_2786 ( .ZN(net_2147), .A(net_800) );
NAND4_X2 inst_1224 ( .A4(net_4125), .A1(net_4097), .A3(net_3656), .ZN(net_1046), .A2(net_717) );
AOI221_X2 inst_3905 ( .A(net_4091), .B2(net_3559), .ZN(net_1019), .C2(net_1018), .B1(net_924), .C1(net_799) );
NAND2_X2 inst_1924 ( .A1(net_3817), .ZN(net_3182), .A2(net_183) );
NOR2_X1 inst_1170 ( .A2(net_4150), .ZN(net_3475), .A1(net_3271) );
INV_X4 inst_2596 ( .ZN(net_3736), .A(net_3735) );
INV_X2 inst_3022 ( .ZN(net_3442), .A(net_2303) );
OAI21_X2 inst_680 ( .B1(net_3228), .B2(net_3153), .ZN(net_1440), .A(net_1307) );
CLKBUF_X2 inst_4748 ( .A(net_4733), .Z(net_4734) );
OAI211_X2 inst_785 ( .C2(net_2778), .ZN(net_2763), .C1(net_2732), .B(net_2672), .A(net_2650) );
INV_X4 inst_2362 ( .A(net_1173), .ZN(net_593) );
DFF_X1 inst_3299 ( .D(net_3748), .Q(net_3745), .QN(net_67), .CK(net_4284) );
AND2_X4 inst_4160 ( .ZN(net_4111), .A2(net_3912), .A1(net_3900) );
DFF_X1 inst_3255 ( .QN(net_3087), .D(net_2950), .CK(net_4603) );
INV_X2 inst_2856 ( .ZN(net_2033), .A(net_260) );
NOR2_X4 inst_961 ( .ZN(net_3776), .A1(net_3346), .A2(net_3345) );
NAND2_X2 inst_1590 ( .A1(net_2972), .ZN(net_2428), .A2(net_781) );
INV_X4 inst_2318 ( .A(net_767), .ZN(net_747) );
OAI221_X2 inst_399 ( .C2(net_3407), .B1(net_2328), .ZN(net_2285), .C1(net_2208), .A(net_1936), .B2(net_70) );
CLKBUF_X2 inst_5103 ( .A(net_4830), .Z(net_5089) );
OAI21_X2 inst_527 ( .B1(net_3302), .ZN(net_2908), .B2(net_2907), .A(net_2483) );
AOI21_X2 inst_3957 ( .ZN(net_1631), .B1(net_1593), .A(net_1047), .B2(net_127) );
AOI22_X2 inst_3567 ( .A1(net_4059), .B1(net_4056), .ZN(net_1483), .B2(net_493), .A2(net_470) );
OR2_X4 inst_226 ( .ZN(net_902), .A1(net_692), .A2(net_691) );
NAND4_X2 inst_1180 ( .ZN(net_2697), .A2(net_2537), .A1(net_2341), .A3(net_2318), .A4(net_2276) );
AOI211_X2 inst_4020 ( .A(net_4091), .ZN(net_1599), .B(net_1512), .C1(net_1015), .C2(net_408) );
OAI221_X2 inst_414 ( .C1(net_4093), .ZN(net_1528), .C2(net_1381), .A(net_1231), .B1(net_1221), .B2(net_406) );
OAI21_X2 inst_531 ( .B1(net_3195), .B2(net_2972), .ZN(net_2902), .A(net_2432) );
INV_X2 inst_2737 ( .ZN(net_1309), .A(net_1308) );
INV_X4 inst_2316 ( .ZN(net_929), .A(net_763) );
OR2_X4 inst_212 ( .A1(net_3492), .A2(net_3364), .ZN(net_1740) );
INV_X2 inst_2732 ( .ZN(net_1392), .A(net_1347) );
NAND3_X2 inst_1299 ( .A1(net_3112), .ZN(net_1531), .A2(net_1337), .A3(net_671) );
OAI21_X2 inst_499 ( .B1(net_3394), .B2(net_2961), .ZN(net_2943), .A(net_2471) );
NAND2_X2 inst_1952 ( .A2(net_3578), .A1(net_3370), .ZN(net_3277) );
OAI21_X2 inst_674 ( .A(net_3793), .ZN(net_1362), .B1(net_1332), .B2(net_1041) );
CLKBUF_X2 inst_5259 ( .A(net_4436), .Z(net_5245) );
INV_X4 inst_2400 ( .ZN(net_333), .A(net_46) );
NAND2_X4 inst_1451 ( .ZN(net_3827), .A2(net_3237), .A1(net_2244) );
CLKBUF_X2 inst_4781 ( .A(net_4611), .Z(net_4767) );
AND3_X2 inst_4082 ( .A3(net_4110), .A1(net_3448), .ZN(net_2711), .A2(net_2518) );
CLKBUF_X2 inst_5023 ( .A(net_5008), .Z(net_5009) );
AOI22_X2 inst_3698 ( .B2(net_4124), .A2(net_555), .ZN(net_476), .A1(net_475), .B1(net_474) );
INV_X4 inst_2253 ( .A(net_3845), .ZN(net_1292) );
AND2_X4 inst_4155 ( .ZN(net_4105), .A1(net_3656), .A2(net_359) );
CLKBUF_X2 inst_5118 ( .A(net_5103), .Z(net_5104) );
INV_X2 inst_2966 ( .A(net_3004), .ZN(net_188) );
NAND2_X2 inst_2009 ( .A2(net_3820), .ZN(net_3545), .A1(net_3211) );
DFF_X1 inst_3246 ( .QN(net_3083), .D(net_2949), .CK(net_4555) );
INV_X2 inst_2868 ( .ZN(net_259), .A(net_50) );
OAI21_X2 inst_501 ( .B1(net_3394), .B2(net_2959), .ZN(net_2941), .A(net_2499) );
NAND2_X1 inst_2093 ( .ZN(net_415), .A2(net_281), .A1(x557) );
CLKBUF_X2 inst_4904 ( .A(net_4889), .Z(net_4890) );
NOR2_X2 inst_1081 ( .A1(net_3614), .ZN(net_613), .A2(net_436) );
DFF_X2 inst_3195 ( .QN(net_3107), .D(net_1626), .CK(net_4831) );
CLKBUF_X2 inst_4887 ( .A(net_4382), .Z(net_4873) );
INV_X4 inst_2381 ( .A(net_3789), .ZN(net_414) );
INV_X2 inst_2905 ( .A(net_3026), .ZN(net_136) );
NAND2_X2 inst_1832 ( .ZN(net_746), .A2(net_745), .A1(net_685) );
OAI21_X2 inst_570 ( .B2(net_3599), .ZN(net_2837), .B1(net_2836), .A(net_2061) );
INV_X2 inst_2819 ( .A(net_3521), .ZN(net_667) );
NAND2_X2 inst_1570 ( .A1(net_2912), .ZN(net_2451), .A2(net_200) );
CLKBUF_X2 inst_4562 ( .A(net_4254), .Z(net_4548) );
OAI21_X2 inst_640 ( .B2(net_3338), .ZN(net_2070), .A(net_1970), .B1(net_1969) );
NAND2_X2 inst_1612 ( .A1(net_2967), .ZN(net_2404), .A2(net_191) );
NAND2_X4 inst_1478 ( .A1(net_3995), .ZN(net_3943), .A2(net_3109) );
CLKBUF_X2 inst_4645 ( .A(net_4630), .Z(net_4631) );
NOR2_X2 inst_1114 ( .A2(net_3854), .ZN(net_3365), .A1(net_3286) );
OAI21_X4 inst_454 ( .B1(net_3264), .ZN(net_1869), .B2(net_1525), .A(net_1372) );
AND2_X4 inst_4163 ( .A2(net_4122), .ZN(net_4117), .A1(net_272) );
NAND2_X2 inst_1982 ( .A1(net_3881), .A2(net_3618), .ZN(net_3405) );
NAND2_X1 inst_2089 ( .A2(net_4021), .A1(net_2967), .ZN(net_2411) );
AOI22_X2 inst_3718 ( .B2(net_4099), .ZN(net_3573), .A2(net_3571), .B1(net_963), .A1(net_838) );
NAND2_X2 inst_1849 ( .ZN(net_665), .A1(net_600), .A2(net_450) );
NAND2_X2 inst_1679 ( .A1(net_3281), .ZN(net_2029), .A2(net_181) );
CLKBUF_X2 inst_4932 ( .A(net_4917), .Z(net_4918) );
NAND2_X2 inst_1976 ( .ZN(net_3352), .A1(net_2527), .A2(net_2376) );
AOI22_X2 inst_3681 ( .B1(net_4123), .A1(net_555), .ZN(net_502), .B2(net_170), .A2(net_166) );
INV_X2 inst_2744 ( .ZN(net_1195), .A(net_1144) );
INV_X4 inst_2215 ( .ZN(net_2120), .A(net_1945) );
INV_X1 inst_3077 ( .A(net_867), .ZN(net_812) );
NAND2_X2 inst_1855 ( .ZN(net_1041), .A1(net_641), .A2(net_403) );
OAI22_X2 inst_337 ( .ZN(net_429), .A2(net_347), .A1(net_344), .B2(net_263), .B1(net_47) );
CLKBUF_X2 inst_5277 ( .A(net_5262), .Z(net_5263) );
CLKBUF_X2 inst_4614 ( .A(net_4268), .Z(net_4600) );
INV_X4 inst_2384 ( .A(net_3664), .ZN(net_390) );
NAND4_X2 inst_1212 ( .ZN(net_1311), .A1(net_992), .A2(net_985), .A4(net_913), .A3(net_878) );
OAI21_X2 inst_670 ( .ZN(net_1468), .A(net_1341), .B1(net_182), .B2(net_115) );
CLKBUF_X2 inst_5224 ( .A(net_5209), .Z(net_5210) );
NAND2_X4 inst_1423 ( .ZN(net_3586), .A1(net_3585), .A2(net_2383) );
AND2_X4 inst_4180 ( .ZN(net_4140), .A2(net_3171), .A1(net_283) );
INV_X4 inst_2419 ( .ZN(net_247), .A(net_201) );
NOR2_X2 inst_1034 ( .ZN(net_1368), .A1(net_1243), .A2(net_1090) );
NAND4_X2 inst_1207 ( .A1(net_2020), .ZN(net_1628), .A4(net_321), .A3(net_258), .A2(net_53) );
AOI221_X2 inst_3901 ( .ZN(net_1204), .A(net_1203), .B1(net_1202), .C1(net_1201), .C2(net_1200), .B2(net_983) );
OAI21_X2 inst_613 ( .ZN(net_2641), .B1(net_2293), .B2(net_2246), .A(net_356) );
CLKBUF_X2 inst_4275 ( .A(net_4260), .Z(net_4261) );
CLKBUF_X2 inst_5041 ( .A(net_5026), .Z(net_5027) );
INV_X4 inst_2396 ( .ZN(net_404), .A(net_343) );
NAND2_X4 inst_1428 ( .A1(net_4002), .ZN(net_3615), .A2(net_376) );
OAI21_X2 inst_483 ( .B1(net_2970), .ZN(net_2960), .B2(net_2959), .A(net_2501) );
CLKBUF_X2 inst_5005 ( .A(net_4990), .Z(net_4991) );
INV_X2 inst_2739 ( .A(net_3931), .ZN(net_1282) );
OR2_X2 inst_259 ( .A1(net_4103), .A2(net_3670), .ZN(net_850) );
NOR2_X2 inst_1046 ( .A1(net_4156), .A2(net_3968), .ZN(net_1080) );
OR2_X4 inst_246 ( .ZN(net_4143), .A1(net_3780), .A2(net_2988) );
CLKBUF_X2 inst_4443 ( .A(net_4250), .Z(net_4429) );
CLKBUF_X2 inst_4355 ( .A(net_4340), .Z(net_4341) );
OAI21_X2 inst_635 ( .B2(net_2076), .ZN(net_2075), .A(net_1963), .B1(net_1673) );
CLKBUF_X2 inst_4707 ( .A(net_4692), .Z(net_4693) );
OAI211_X2 inst_807 ( .C2(net_3755), .ZN(net_1834), .C1(net_1513), .B(net_1197), .A(net_1187) );
CLKBUF_X2 inst_4846 ( .A(net_4494), .Z(net_4832) );
OAI21_X2 inst_705 ( .B1(net_3328), .ZN(net_890), .A(net_889), .B2(net_530) );
NOR3_X2 inst_911 ( .ZN(net_3415), .A3(net_3414), .A2(net_3412), .A1(net_3411) );
OAI21_X2 inst_519 ( .B2(net_2972), .B1(net_2923), .ZN(net_2921), .A(net_2426) );
AOI221_X2 inst_3796 ( .C2(net_3738), .B1(net_3736), .ZN(net_2856), .C1(net_2855), .A(net_1995), .B2(net_71) );
NOR3_X2 inst_909 ( .A2(net_4052), .ZN(net_3308), .A1(net_3307), .A3(net_1373) );
NOR2_X2 inst_1003 ( .ZN(net_2169), .A1(net_2129), .A2(net_2125) );
INV_X4 inst_2484 ( .A(net_3084), .ZN(net_780) );
NOR2_X2 inst_1053 ( .A2(net_4024), .ZN(net_1136), .A1(net_962) );
CLKBUF_X2 inst_5158 ( .A(net_5143), .Z(net_5144) );
INV_X2 inst_2919 ( .A(net_3137), .ZN(net_267) );
NOR3_X2 inst_894 ( .A3(net_4193), .ZN(net_1892), .A2(net_1891), .A1(net_1789) );
CLKBUF_X2 inst_5039 ( .A(net_5024), .Z(net_5025) );
INV_X4 inst_2425 ( .A(net_3123), .ZN(net_874) );
NAND2_X2 inst_1872 ( .A1(net_3713), .ZN(net_707), .A2(net_590) );
AOI22_X2 inst_3469 ( .B2(net_3116), .A1(net_2724), .B1(net_2722), .ZN(net_2721), .A2(net_35) );
NOR2_X2 inst_994 ( .A1(net_2300), .ZN(net_2296), .A2(net_1646) );
INV_X2 inst_2774 ( .ZN(net_2746), .A(net_901) );
CLKBUF_X2 inst_4577 ( .A(net_4562), .Z(net_4563) );
OR2_X4 inst_239 ( .A2(net_3640), .ZN(net_3599), .A1(net_3598) );
AOI211_X2 inst_4028 ( .A(net_4185), .C2(net_3900), .ZN(net_926), .B(net_925), .C1(net_692) );
NAND2_X2 inst_2080 ( .ZN(net_4181), .A1(net_3589), .A2(net_3184) );
NAND2_X2 inst_1879 ( .A2(net_3395), .ZN(net_637), .A1(net_407) );
NAND4_X2 inst_1193 ( .ZN(net_1667), .A3(net_1491), .A4(net_1490), .A2(net_1432), .A1(net_1424) );
NAND2_X2 inst_1625 ( .A1(net_2391), .ZN(net_2390), .A2(net_370) );
NAND2_X2 inst_1863 ( .A1(net_3156), .A2(net_1463), .ZN(net_1006) );
OAI21_X2 inst_593 ( .B1(net_2584), .ZN(net_2577), .A(net_2390), .B2(net_2114) );
INV_X4 inst_2223 ( .ZN(net_2115), .A(net_1993) );
CLKBUF_X2 inst_4522 ( .A(net_4507), .Z(net_4508) );
INV_X8 inst_2135 ( .A(net_3450), .ZN(net_513) );
OAI21_X2 inst_601 ( .B1(net_3886), .B2(net_3599), .ZN(net_2573), .A(net_1848) );
DFF_X2 inst_3119 ( .QN(net_3155), .D(net_2705), .CK(net_4489) );
CLKBUF_X2 inst_5138 ( .A(net_5123), .Z(net_5124) );
AOI222_X1 inst_3777 ( .ZN(net_1878), .A2(net_1826), .A1(net_1616), .B2(net_984), .C2(net_874), .B1(net_622), .C1(net_579) );
OAI21_X2 inst_764 ( .ZN(net_3917), .A(net_3913), .B2(net_3109), .B1(net_3106) );
NAND2_X2 inst_1773 ( .A1(net_4033), .ZN(net_1172), .A2(net_1108) );
OAI21_X2 inst_479 ( .B1(net_2970), .ZN(net_2968), .B2(net_2967), .A(net_2408) );
INV_X4 inst_2344 ( .A(net_3328), .ZN(net_788) );
NAND2_X2 inst_1547 ( .A1(net_2961), .ZN(net_2475), .A2(net_189) );
XOR2_X1 inst_29 ( .A(net_4117), .B(net_1699), .Z(net_673) );
DFF_X1 inst_3326 ( .Q(net_3110), .D(net_2829), .CK(net_4645) );
NAND2_X2 inst_1583 ( .A1(net_2915), .ZN(net_2437), .A2(net_237) );
OAI21_X1 inst_771 ( .ZN(net_4016), .B2(net_2969), .B1(net_2893), .A(net_2419) );
CLKBUF_X2 inst_4387 ( .A(net_4372), .Z(net_4373) );
INV_X4 inst_2369 ( .ZN(net_666), .A(net_397) );
INV_X8 inst_2152 ( .A(net_3531), .ZN(net_3366) );
AOI21_X2 inst_3947 ( .B1(net_4043), .A(net_2298), .ZN(net_2216), .B2(net_269) );
NAND3_X2 inst_1274 ( .ZN(net_2784), .A3(net_2715), .A2(net_2713), .A1(net_2660) );
AOI221_X2 inst_3838 ( .B1(net_3774), .C1(net_2227), .ZN(net_2221), .C2(net_2220), .A(net_2109), .B2(net_271) );
OAI21_X2 inst_538 ( .B2(net_3208), .B1(net_3195), .ZN(net_2895), .A(net_2495) );
INV_X2 inst_2831 ( .A(net_3396), .ZN(net_439) );
CLKBUF_X2 inst_4497 ( .A(net_4482), .Z(net_4483) );
CLKBUF_X2 inst_4756 ( .A(net_4741), .Z(net_4742) );
INV_X2 inst_2651 ( .ZN(net_2290), .A(net_2278) );
NAND3_X2 inst_1319 ( .A2(net_4105), .A3(net_4004), .ZN(net_785), .A1(net_784) );
NAND3_X2 inst_1300 ( .ZN(net_2815), .A2(net_1458), .A1(net_1378), .A3(net_1036) );
CLKBUF_X2 inst_5280 ( .A(net_5265), .Z(net_5266) );
CLKBUF_X2 inst_4537 ( .A(net_4522), .Z(net_4523) );
AND2_X2 inst_4201 ( .A1(net_4100), .ZN(net_772), .A2(net_82) );
XOR2_X1 inst_35 ( .A(net_4138), .Z(net_3384), .B(net_3377) );
OAI221_X2 inst_358 ( .C1(net_3352), .B2(net_3348), .ZN(net_2833), .B1(net_2816), .A(net_2564), .C2(net_2187) );
XNOR2_X2 inst_48 ( .A(net_3310), .ZN(net_2633), .B(net_2286) );
CLKBUF_X2 inst_4765 ( .A(net_4658), .Z(net_4751) );
CLKBUF_X2 inst_4462 ( .A(net_4447), .Z(net_4448) );
INV_X4 inst_2246 ( .ZN(net_1617), .A(net_1583) );
NAND2_X2 inst_1756 ( .A1(net_4064), .A2(net_4028), .ZN(net_1268) );
INV_X4 inst_2279 ( .ZN(net_1148), .A(net_922) );
OAI221_X2 inst_443 ( .B1(net_4158), .ZN(net_3695), .B2(net_3407), .C1(net_2328), .A(net_1933), .C2(net_132) );
INV_X4 inst_2600 ( .A(net_3995), .ZN(net_3755) );
NAND2_X2 inst_2038 ( .A1(net_3882), .A2(net_3880), .ZN(net_3791) );
CLKBUF_X2 inst_4259 ( .A(net_4229), .Z(net_4245) );
NAND2_X2 inst_2044 ( .A2(net_3887), .ZN(net_3849), .A1(net_3848) );
OAI21_X2 inst_655 ( .ZN(net_1931), .B1(net_1815), .A(net_1803), .B2(net_752) );
CLKBUF_X2 inst_5178 ( .A(net_5157), .Z(net_5164) );
INV_X4 inst_2274 ( .A(net_3339), .ZN(net_1192) );
NAND2_X2 inst_1700 ( .A1(net_4120), .ZN(net_1852), .A2(net_1807) );
INV_X4 inst_2571 ( .ZN(net_3543), .A(net_3542) );
CLKBUF_X2 inst_4438 ( .A(net_4274), .Z(net_4424) );
OAI21_X2 inst_695 ( .ZN(net_1458), .B1(net_1029), .B2(net_1028), .A(net_432) );
OAI21_X2 inst_730 ( .B2(net_991), .A(net_629), .B1(net_628), .ZN(net_580) );
AND4_X4 inst_4038 ( .A4(net_3973), .ZN(net_1255), .A1(net_1254), .A2(net_1253), .A3(net_748) );
OAI22_X2 inst_321 ( .A1(net_1154), .ZN(net_1027), .B1(net_1026), .B2(net_686), .A2(net_245) );
INV_X4 inst_2493 ( .A(net_2994), .ZN(net_217) );
OAI21_X2 inst_511 ( .B1(net_3274), .B2(net_2961), .ZN(net_2931), .A(net_2472) );
XNOR2_X2 inst_41 ( .ZN(net_2762), .A(net_2648), .B(net_1448) );
DFF_X2 inst_3131 ( .D(net_2619), .QN(net_114), .CK(net_4422) );
AOI22_X2 inst_3559 ( .A1(net_4059), .B1(net_4056), .ZN(net_1491), .B2(net_488), .A2(net_474) );
INV_X2 inst_2645 ( .A(net_3876), .ZN(net_2336) );
NAND2_X2 inst_1989 ( .ZN(net_3438), .A1(net_358), .A2(net_328) );
NOR2_X1 inst_1164 ( .A1(net_3554), .ZN(net_2379), .A2(net_1685) );
DFF_X2 inst_3112 ( .QN(net_2991), .D(net_2802), .CK(net_5241) );
SDFF_X2 inst_152 ( .D(net_3511), .SE(net_2514), .SI(net_103), .Q(net_103), .CK(net_4746) );
NOR2_X2 inst_1152 ( .ZN(net_3982), .A2(net_3981), .A1(net_1052) );
NAND4_X2 inst_1242 ( .ZN(net_3357), .A4(net_3356), .A3(net_3355), .A2(net_3351), .A1(net_3350) );
NAND2_X4 inst_1400 ( .A1(net_3661), .ZN(net_767), .A2(net_432) );
CLKBUF_X2 inst_5217 ( .A(net_5172), .Z(net_5203) );
CLKBUF_X2 inst_5233 ( .A(net_5218), .Z(net_5219) );
XNOR2_X2 inst_89 ( .ZN(net_936), .B(net_513), .A(net_408) );
NAND2_X2 inst_1520 ( .A1(net_2959), .ZN(net_2502), .A2(net_734) );
OAI221_X2 inst_388 ( .B2(net_2699), .C2(net_2698), .ZN(net_2542), .A(net_2369), .C1(net_2364), .B1(net_2314) );
CLKBUF_X2 inst_4600 ( .A(net_4483), .Z(net_4586) );
AOI221_X2 inst_3872 ( .B1(net_2020), .C1(net_2019), .ZN(net_1932), .A(net_1931), .B2(net_251), .C2(x437) );
NAND2_X2 inst_1535 ( .A1(net_2907), .ZN(net_2487), .A2(net_186) );
OR3_X2 inst_182 ( .ZN(net_1287), .A1(net_1168), .A3(net_1124), .A2(net_717) );
OAI211_X2 inst_788 ( .C2(net_2778), .ZN(net_2756), .C1(net_2666), .A(net_2653), .B(net_2606) );
OAI21_X2 inst_489 ( .B1(net_3394), .B2(net_2969), .ZN(net_2953), .A(net_2414) );
NOR2_X4 inst_931 ( .A1(net_3556), .A2(net_3019), .ZN(net_2027) );
DFF_X2 inst_3174 ( .D(net_1911), .Q(net_122), .CK(net_4997) );
AOI221_X2 inst_3824 ( .B2(net_3147), .A(net_2642), .B1(net_2591), .C1(net_2589), .ZN(net_2552), .C2(net_2551) );
NAND2_X2 inst_1674 ( .A1(net_2134), .ZN(net_2084), .A2(net_232) );
AOI22_X2 inst_3622 ( .B2(net_3158), .B1(net_1882), .ZN(net_1095), .A2(net_1094), .A1(net_939) );
NAND2_X2 inst_1579 ( .A1(net_2965), .ZN(net_2441), .A2(net_597) );
NAND2_X4 inst_1411 ( .A1(net_3898), .A2(net_3827), .ZN(net_3333) );
SDFF_X2 inst_149 ( .D(net_3248), .SE(net_2514), .SI(net_104), .Q(net_104), .CK(net_4747) );
OR2_X4 inst_193 ( .A1(net_3881), .A2(net_3515), .ZN(net_2366) );
XOR2_X1 inst_39 ( .Z(net_4196), .B(net_817), .A(net_766) );
AND3_X2 inst_4089 ( .A1(net_4093), .A2(net_1717), .ZN(net_859), .A3(net_40) );
NAND2_X4 inst_1415 ( .A1(net_3525), .ZN(net_3430), .A2(net_401) );
INV_X2 inst_2627 ( .A(net_3342), .ZN(net_2892) );
NAND2_X2 inst_1709 ( .A2(net_2268), .ZN(net_1727), .A1(net_1726) );
DFF_X1 inst_3301 ( .Q(net_3111), .D(net_2879), .CK(net_4523) );
INV_X4 inst_2320 ( .ZN(net_853), .A(net_683) );
DFF_X2 inst_3173 ( .D(net_1913), .QN(net_123), .CK(net_5276) );
XNOR2_X2 inst_125 ( .ZN(net_4155), .A(net_3369), .B(net_2347) );
INV_X4 inst_2534 ( .A(net_4004), .ZN(net_3319) );
INV_X4 inst_2202 ( .A(net_3857), .ZN(net_2288) );
CLKBUF_X2 inst_4770 ( .A(net_4755), .Z(net_4756) );
DFF_X2 inst_3180 ( .D(net_1819), .QN(net_107), .CK(net_4375) );
CLKBUF_X2 inst_4737 ( .A(net_4722), .Z(net_4723) );
INV_X2 inst_2987 ( .A(net_3009), .ZN(net_214) );
AOI222_X2 inst_3737 ( .B1(net_4196), .B2(net_1826), .ZN(net_1221), .A1(net_630), .C1(net_576), .C2(net_393), .A2(net_323) );
NAND2_X2 inst_1636 ( .A1(net_4041), .A2(net_3159), .ZN(net_2377) );
OAI221_X2 inst_430 ( .B1(net_3990), .C1(net_1129), .ZN(net_972), .A(net_971), .B2(net_667), .C2(net_646) );
CLKBUF_X2 inst_4599 ( .A(net_4584), .Z(net_4585) );
CLKBUF_X2 inst_4677 ( .A(net_4662), .Z(net_4663) );
OAI21_X2 inst_515 ( .B2(net_2961), .ZN(net_2927), .B1(net_2923), .A(net_2469) );
NAND2_X2 inst_1501 ( .ZN(net_2808), .A1(net_2794), .A2(net_2626) );
INV_X4 inst_2473 ( .A(net_2985), .ZN(net_147) );
DFF_X2 inst_3212 ( .D(net_801), .QN(net_289), .CK(net_4620) );
NAND2_X2 inst_1698 ( .A2(net_3506), .ZN(net_1886), .A1(net_1833) );
CLKBUF_X2 inst_5248 ( .A(net_5233), .Z(net_5234) );
INV_X4 inst_2565 ( .A(net_3631), .ZN(net_3521) );
NOR2_X4 inst_944 ( .A1(net_3983), .A2(net_3935), .ZN(net_3452) );
CLKBUF_X2 inst_4516 ( .A(net_4501), .Z(net_4502) );
INV_X2 inst_2945 ( .A(net_3053), .ZN(net_208) );
NAND2_X2 inst_1584 ( .A1(net_2915), .ZN(net_2436), .A2(net_180) );
OAI21_X2 inst_642 ( .ZN(net_1994), .B1(net_1993), .A(net_1859), .B2(net_1535) );
OAI21_X4 inst_459 ( .B1(net_4184), .ZN(net_3263), .B2(net_1608), .A(net_1503) );
INV_X2 inst_2993 ( .A(net_3020), .ZN(net_165) );
INV_X2 inst_2864 ( .A(net_3142), .ZN(net_295) );
AOI22_X2 inst_3476 ( .B1(net_4039), .A1(net_2675), .ZN(net_2674), .A2(net_1523), .B2(x40) );
NOR2_X2 inst_1018 ( .A1(net_2661), .A2(net_1905), .ZN(net_1824) );
AOI222_X1 inst_3789 ( .B1(net_4185), .C1(net_4101), .A2(net_3440), .ZN(net_1111), .C2(net_1011), .A1(net_897), .B2(net_649) );
INV_X2 inst_2933 ( .ZN(net_132), .A(net_73) );
OAI21_X2 inst_700 ( .B1(net_4088), .B2(net_3152), .ZN(net_934), .A(net_401) );
DFF_X1 inst_3393 ( .Q(net_3112), .D(net_1619), .CK(net_4473) );
OAI221_X2 inst_367 ( .B1(net_3553), .C1(net_3352), .B2(net_3348), .ZN(net_2728), .A(net_2552), .C2(net_2167) );
NOR2_X4 inst_957 ( .A1(net_4006), .A2(net_3942), .ZN(net_3713) );
NOR2_X4 inst_979 ( .ZN(net_3956), .A2(net_3954), .A1(net_3953) );
INV_X2 inst_2713 ( .A(net_3858), .ZN(net_2373) );
CLKBUF_X2 inst_4976 ( .A(net_4791), .Z(net_4962) );
NOR2_X2 inst_1008 ( .ZN(net_1782), .A2(net_1747), .A1(net_1689) );
DFF_X1 inst_3409 ( .D(net_1402), .Q(net_56), .CK(net_4819) );
CLKBUF_X2 inst_4568 ( .A(net_4553), .Z(net_4554) );
OAI21_X2 inst_559 ( .B2(net_2907), .B1(net_2871), .ZN(net_2866), .A(net_2484) );
NAND2_X2 inst_1871 ( .A2(net_3755), .ZN(net_603), .A1(net_337) );
INV_X4 inst_2296 ( .ZN(net_1586), .A(net_1064) );
AOI22_X2 inst_3591 ( .A1(net_4062), .B1(net_4057), .ZN(net_1426), .B2(net_170), .A2(net_166) );
INV_X4 inst_2300 ( .ZN(net_872), .A(net_871) );
CLKBUF_X2 inst_4964 ( .A(net_4949), .Z(net_4950) );
OAI221_X1 inst_450 ( .ZN(net_3743), .B1(net_3735), .C1(net_1993), .A(net_1898), .C2(net_1541), .B2(net_67) );
OAI21_X2 inst_520 ( .B1(net_3302), .ZN(net_2920), .B2(net_2919), .A(net_2398) );
OAI21_X2 inst_745 ( .B1(net_3430), .ZN(net_3339), .B2(net_3102), .A(net_862) );
AOI22_X2 inst_3658 ( .ZN(net_573), .A1(net_458), .B1(net_457), .B2(net_188), .A2(net_174) );
DFF_X1 inst_3405 ( .Q(net_4027), .D(net_1466), .CK(net_4508) );
AOI221_X2 inst_3888 ( .C2(net_4079), .A(net_4072), .ZN(net_1589), .C1(net_1224), .B2(net_1011), .B1(net_705) );
NAND2_X2 inst_2032 ( .A2(net_4164), .A1(net_3974), .ZN(net_3763) );
CLKBUF_X2 inst_4554 ( .A(net_4258), .Z(net_4540) );
CLKBUF_X2 inst_4258 ( .A(net_4243), .Z(net_4244) );
AND2_X4 inst_4113 ( .A2(net_3389), .ZN(net_401), .A1(net_248) );
AOI22_X2 inst_3623 ( .B1(net_3141), .ZN(net_1316), .B2(net_1071), .A2(net_1036), .A1(net_951) );
XNOR2_X2 inst_80 ( .ZN(net_1285), .B(net_1139), .A(net_1088) );
NAND2_X2 inst_2026 ( .A2(net_4162), .A1(net_4001), .ZN(net_3733) );
OAI211_X2 inst_836 ( .C2(net_3149), .C1(net_1359), .ZN(net_1354), .A(net_1239), .B(net_593) );
NAND2_X2 inst_1556 ( .A1(net_2909), .ZN(net_2466), .A2(net_222) );
AND4_X4 inst_4040 ( .A1(net_3901), .A2(net_3836), .A4(net_3547), .ZN(net_1084), .A3(net_767) );
CLKBUF_X2 inst_4334 ( .A(net_4259), .Z(net_4320) );
OR2_X4 inst_241 ( .ZN(net_3735), .A1(net_3427), .A2(net_1173) );
NOR2_X2 inst_1059 ( .ZN(net_1063), .A2(net_958), .A1(net_938) );
CLKBUF_X2 inst_5120 ( .A(net_5105), .Z(net_5106) );
CLKBUF_X2 inst_4409 ( .A(net_4394), .Z(net_4395) );
CLKBUF_X2 inst_4934 ( .A(net_4355), .Z(net_4920) );
NOR2_X2 inst_1075 ( .A2(net_3755), .ZN(net_675), .A1(net_618) );
NOR4_X2 inst_862 ( .A3(net_3777), .A2(net_3640), .ZN(net_2309), .A4(net_1325), .A1(net_1322) );
CLKBUF_X2 inst_4390 ( .A(net_4369), .Z(net_4376) );
CLKBUF_X2 inst_4358 ( .A(net_4290), .Z(net_4344) );
AOI221_X2 inst_3918 ( .B2(net_3788), .ZN(net_3570), .C2(net_3559), .A(net_1061), .C1(net_907), .B1(net_521) );
INV_X2 inst_2758 ( .A(net_1650), .ZN(net_1279) );
CLKBUF_X2 inst_4504 ( .A(net_4315), .Z(net_4490) );
NOR2_X2 inst_1116 ( .ZN(net_3389), .A1(net_3388), .A2(net_3127) );
CLKBUF_X2 inst_4328 ( .A(net_4313), .Z(net_4314) );
INV_X4 inst_2257 ( .ZN(net_1186), .A(net_1122) );
AND2_X4 inst_4173 ( .ZN(net_4127), .A1(net_3468), .A2(net_41) );
AOI222_X1 inst_3753 ( .A1(net_3676), .B1(net_2055), .C1(net_2054), .ZN(net_2040), .C2(net_821), .B2(net_378), .A2(net_280) );
NAND2_X2 inst_1764 ( .A2(net_1394), .ZN(net_1235), .A1(net_33) );
CLKBUF_X2 inst_5271 ( .A(net_4229), .Z(net_5257) );
NOR2_X2 inst_1104 ( .A2(net_4190), .A1(net_3299), .ZN(net_3184) );
NOR2_X2 inst_1159 ( .ZN(net_4097), .A1(net_526), .A2(net_380) );
INV_X4 inst_2355 ( .A(net_3997), .ZN(net_537) );
DFF_X2 inst_3136 ( .QN(net_2989), .D(net_2575), .CK(net_5153) );
OAI221_X2 inst_402 ( .C2(net_4034), .ZN(net_2300), .C1(net_2212), .B1(net_2042), .B2(net_2032), .A(net_1284) );
OAI22_X2 inst_329 ( .B1(net_3438), .ZN(net_864), .A1(net_863), .B2(net_513), .A2(net_408) );
OAI21_X2 inst_494 ( .B1(net_3588), .B2(net_2965), .ZN(net_2948), .A(net_2441) );
OAI21_X2 inst_574 ( .B2(net_2925), .ZN(net_2805), .B1(net_2803), .A(net_2434) );
NOR2_X4 inst_938 ( .A1(net_4007), .A2(net_3106), .ZN(net_376) );
INV_X4 inst_2347 ( .ZN(net_600), .A(net_541) );
AND2_X4 inst_4102 ( .A2(net_3490), .ZN(net_1837), .A1(x475) );
NAND4_X2 inst_1229 ( .A4(net_987), .A3(net_854), .ZN(net_730), .A2(net_729), .A1(net_604) );
NAND3_X2 inst_1288 ( .ZN(net_2259), .A1(net_2200), .A3(net_1953), .A2(net_1918) );
AOI221_X2 inst_3844 ( .B2(net_2203), .C1(net_2202), .ZN(net_2198), .A(net_2075), .B1(net_1767), .C2(net_378) );
CLKBUF_X2 inst_5219 ( .A(net_4457), .Z(net_5205) );
INV_X2 inst_2894 ( .A(net_3037), .ZN(net_183) );
INV_X4 inst_2358 ( .A(net_3656), .ZN(net_529) );
INV_X8 inst_2125 ( .ZN(net_641), .A(net_516) );
AOI22_X2 inst_3638 ( .ZN(net_782), .A1(net_781), .B1(net_780), .A2(net_458), .B2(net_457) );
CLKBUF_X2 inst_4365 ( .A(net_4266), .Z(net_4351) );
INV_X2 inst_2959 ( .ZN(net_258), .A(net_54) );
OAI21_X2 inst_599 ( .ZN(net_2508), .B1(net_2507), .A(net_2295), .B2(net_299) );
NOR2_X2 inst_1033 ( .A1(net_3229), .ZN(net_1443), .A2(net_294) );
NAND2_X2 inst_1683 ( .A1(net_3176), .ZN(net_2023), .A2(net_194) );
CLKBUF_X2 inst_4673 ( .A(net_4465), .Z(net_4659) );
AOI221_X2 inst_3865 ( .B1(net_2020), .C1(net_2019), .ZN(net_1944), .A(net_1943), .B2(net_206), .C2(x368) );
NAND3_X2 inst_1348 ( .A2(net_4088), .ZN(net_3485), .A3(net_3152), .A1(net_433) );
NAND2_X1 inst_2102 ( .ZN(net_4148), .A1(net_3198), .A2(net_213) );
CLKBUF_X2 inst_4908 ( .A(net_4893), .Z(net_4894) );
NAND2_X2 inst_1748 ( .A1(net_3229), .ZN(net_1437), .A2(net_68) );
OAI21_X2 inst_541 ( .ZN(net_4022), .B2(net_2961), .B1(net_2893), .A(net_2476) );
AND4_X4 inst_4047 ( .A4(net_4125), .A1(net_4097), .ZN(net_4076), .A2(net_3656), .A3(net_384) );
OAI21_X2 inst_505 ( .B1(net_3278), .ZN(net_2937), .B2(net_2917), .A(net_2393) );
NAND3_X2 inst_1365 ( .ZN(net_3970), .A3(net_3967), .A2(net_3789), .A1(net_1132) );
OR2_X4 inst_198 ( .A1(net_3179), .ZN(net_2969), .A2(net_2352) );
AND2_X4 inst_4125 ( .ZN(net_4051), .A1(net_3331), .A2(net_426) );
NAND3_X2 inst_1371 ( .ZN(net_4157), .A3(net_3999), .A1(net_3526), .A2(net_3171) );
CLKBUF_X2 inst_4321 ( .A(net_4280), .Z(net_4307) );
NAND2_X2 inst_1644 ( .A1(net_3199), .ZN(net_2171), .A2(net_2103) );
AOI22_X2 inst_3543 ( .B1(net_4054), .B2(net_3110), .ZN(net_1580), .A1(net_1578), .A2(net_396) );
OAI211_X2 inst_784 ( .C2(net_2778), .ZN(net_2771), .C1(net_2704), .B(net_2673), .A(net_2656) );
DFF_X1 inst_3237 ( .QN(net_3041), .D(net_2938), .CK(net_5194) );
NAND3_X4 inst_1264 ( .A3(net_4143), .ZN(net_3520), .A2(net_3519), .A1(net_3518) );
AOI22_X4 inst_3461 ( .A1(net_3817), .ZN(net_3209), .B1(net_3186), .A2(net_3029), .B2(net_3028) );
OAI21_X2 inst_690 ( .ZN(net_1083), .A(net_1082), .B1(net_1081), .B2(net_1026) );
CLKBUF_X2 inst_4969 ( .A(net_4928), .Z(net_4955) );
AOI22_X2 inst_3511 ( .B1(net_3676), .B2(net_3132), .A1(net_2012), .ZN(net_2006), .A2(net_396) );
CLKBUF_X2 inst_4692 ( .A(net_4660), .Z(net_4678) );
NAND2_X2 inst_2025 ( .A2(net_3947), .ZN(net_3728), .A1(net_3612) );
CLKBUF_X2 inst_4883 ( .A(net_4868), .Z(net_4869) );
INV_X4 inst_2461 ( .ZN(net_1444), .A(net_68) );
OAI21_X2 inst_732 ( .A(net_629), .B1(net_628), .ZN(net_578), .B2(net_225) );
CLKBUF_X2 inst_4717 ( .A(net_4702), .Z(net_4703) );
INV_X4 inst_2178 ( .A(net_3808), .ZN(net_2741) );
OR2_X2 inst_263 ( .A2(net_4120), .ZN(net_1776), .A1(net_586) );
OR3_X2 inst_185 ( .ZN(net_904), .A1(net_889), .A2(net_435), .A3(net_334) );
XNOR2_X2 inst_75 ( .A(net_3229), .ZN(net_1449), .B(net_70) );
OR3_X4 inst_166 ( .A2(net_4095), .ZN(net_1891), .A1(net_1012), .A3(net_56) );
AOI221_X2 inst_3815 ( .C1(net_3445), .A(net_2642), .C2(net_2594), .ZN(net_2585), .B1(net_2584), .B2(net_686) );
CLKBUF_X2 inst_4786 ( .A(net_4547), .Z(net_4772) );
XNOR2_X2 inst_79 ( .ZN(net_1329), .B(net_1221), .A(net_977) );
NAND2_X2 inst_1757 ( .A1(net_3500), .ZN(net_2125), .A2(net_1264) );
AOI221_X2 inst_3851 ( .A(net_4183), .ZN(net_2066), .C2(net_1908), .C1(net_1664), .B2(net_749), .B1(net_101) );
INV_X2 inst_2654 ( .ZN(net_2275), .A(net_2274) );
AND2_X4 inst_4118 ( .ZN(net_4039), .A1(net_2325), .A2(net_1386) );
NAND2_X2 inst_1605 ( .A1(net_2969), .ZN(net_2412), .A2(net_226) );
CLKBUF_X2 inst_4849 ( .A(net_4708), .Z(net_4835) );
CLKBUF_X2 inst_4413 ( .A(net_4398), .Z(net_4399) );
CLKBUF_X2 inst_4649 ( .A(net_4634), .Z(net_4635) );
INV_X2 inst_2975 ( .ZN(net_216), .A(net_111) );
NAND2_X2 inst_1741 ( .ZN(net_1512), .A1(net_1370), .A2(net_863) );
NOR2_X2 inst_1024 ( .A2(net_4070), .A1(net_1646), .ZN(net_1610) );
INV_X4 inst_2232 ( .ZN(net_1807), .A(net_38) );
CLKBUF_X2 inst_5308 ( .A(net_5293), .Z(net_5294) );
CLKBUF_X2 inst_4546 ( .A(net_4531), .Z(net_4532) );
NAND2_X2 inst_1658 ( .ZN(net_2105), .A1(net_1982), .A2(net_233) );
NAND2_X2 inst_1689 ( .A1(net_1982), .ZN(net_1981), .A2(net_170) );
CLKBUF_X2 inst_4475 ( .A(net_4460), .Z(net_4461) );
CLKBUF_X2 inst_4267 ( .A(net_4252), .Z(net_4253) );
AOI21_X2 inst_3965 ( .ZN(net_1452), .A(net_1318), .B1(net_1258), .B2(net_991) );
INV_X2 inst_2846 ( .ZN(net_408), .A(net_403) );
AOI22_X2 inst_3584 ( .A1(net_4063), .B1(net_4058), .B2(net_3455), .ZN(net_1433), .A2(net_201) );
CLKBUF_X2 inst_5034 ( .A(net_5019), .Z(net_5020) );
CLKBUF_X2 inst_4853 ( .A(net_4838), .Z(net_4839) );
NAND2_X4 inst_1448 ( .A1(net_3849), .ZN(net_3803), .A2(net_3517) );
OAI221_X2 inst_440 ( .B2(net_4180), .ZN(net_3465), .C2(net_3464), .C1(net_3463), .B1(net_3462), .A(net_3461) );
NAND2_X2 inst_1816 ( .A1(net_4110), .ZN(net_830), .A2(net_829) );
AOI221_X2 inst_3898 ( .B2(net_3418), .B1(net_1656), .C2(net_1288), .ZN(net_1252), .C1(net_1246), .A(net_1070) );
CLKBUF_X2 inst_5254 ( .A(net_4206), .Z(net_5240) );
CLKBUF_X2 inst_5201 ( .A(net_5150), .Z(net_5187) );
CLKBUF_X2 inst_5012 ( .A(net_4605), .Z(net_4998) );
INV_X4 inst_2373 ( .ZN(net_2642), .A(net_1386) );
CLKBUF_X2 inst_4927 ( .A(net_4912), .Z(net_4913) );
DFF_X1 inst_3381 ( .D(net_2236), .QN(net_62), .CK(net_4209) );
AOI22_X2 inst_3503 ( .B1(net_4080), .ZN(net_2032), .A2(net_1807), .A1(net_1774), .B2(net_39) );
NOR2_X2 inst_1091 ( .ZN(net_413), .A1(net_266), .A2(net_164) );
NAND2_X2 inst_1887 ( .A1(net_3929), .ZN(net_889), .A2(net_398) );
NAND3_X2 inst_1331 ( .A2(net_3395), .ZN(net_534), .A3(net_516), .A1(net_376) );
AND2_X4 inst_4138 ( .ZN(net_4067), .A1(net_3905), .A2(net_1037) );
XNOR2_X2 inst_52 ( .A(net_3311), .ZN(net_2512), .B(net_1598) );
CLKBUF_X2 inst_5059 ( .A(net_4688), .Z(net_5045) );
CLKBUF_X2 inst_4837 ( .A(net_4822), .Z(net_4823) );
OAI21_X2 inst_668 ( .A(net_4191), .ZN(net_1592), .B1(net_1389), .B2(net_786) );
DFF_X1 inst_3223 ( .QN(net_3057), .D(net_2981), .CK(net_4742) );
AOI22_X2 inst_3579 ( .A1(net_4059), .B1(net_4056), .ZN(net_1471), .B2(net_226), .A2(net_167) );
INV_X2 inst_3049 ( .A(net_3959), .ZN(net_3818) );
AND2_X4 inst_4154 ( .ZN(net_4103), .A1(net_3214), .A2(net_881) );
AOI22_X2 inst_3560 ( .A1(net_4060), .B1(net_4055), .ZN(net_1490), .B2(net_735), .A2(net_734) );
AND2_X4 inst_4159 ( .ZN(net_4110), .A2(net_3662), .A1(net_775) );
INV_X2 inst_2683 ( .ZN(net_1846), .A(net_1802) );
CLKBUF_X2 inst_4816 ( .A(net_4801), .Z(net_4802) );
NAND2_X2 inst_1672 ( .ZN(net_2086), .A1(net_2082), .A2(net_180) );
CLKBUF_X2 inst_4223 ( .A(net_4208), .Z(net_4209) );
DFF_X1 inst_3349 ( .D(net_2729), .CK(net_4343), .Q(x105) );
NAND2_X2 inst_2015 ( .A1(net_3647), .ZN(net_3646), .A2(net_492) );
DFF_X2 inst_3179 ( .D(net_1877), .Q(net_53), .CK(net_4841) );
INV_X4 inst_2545 ( .ZN(net_3445), .A(net_3444) );
INV_X2 inst_3059 ( .A(net_3994), .ZN(net_3993) );
AOI21_X2 inst_3937 ( .ZN(net_2301), .B1(net_2300), .A(net_2267), .B2(net_248) );
INV_X2 inst_2970 ( .ZN(net_224), .A(net_110) );
INV_X2 inst_2768 ( .ZN(net_918), .A(net_917) );
NAND2_X2 inst_1835 ( .A1(net_4004), .ZN(net_829), .A2(net_669) );
AND3_X2 inst_4085 ( .A1(net_1254), .ZN(net_1207), .A2(net_1037), .A3(net_899) );
NAND2_X2 inst_1910 ( .ZN(net_298), .A1(net_284), .A2(net_264) );
CLKBUF_X2 inst_4990 ( .A(net_4672), .Z(net_4976) );
CLKBUF_X2 inst_4639 ( .A(net_4624), .Z(net_4625) );
INV_X4 inst_2587 ( .ZN(net_3659), .A(net_3655) );
OAI21_X2 inst_621 ( .B1(net_2235), .ZN(net_2162), .A(net_2058), .B2(net_109) );
DFF_X2 inst_3115 ( .QN(net_2993), .D(net_2804), .CK(net_5239) );
INV_X4 inst_2560 ( .ZN(net_3508), .A(net_3507) );
DFF_X1 inst_3219 ( .QN(net_3061), .D(net_2980), .CK(net_4613) );
OAI211_X2 inst_815 ( .B(net_1628), .C1(net_1627), .ZN(net_1623), .A(net_1550), .C2(net_359) );
INV_X2 inst_3031 ( .ZN(net_3557), .A(net_3555) );
INV_X8 inst_2165 ( .A(net_3816), .ZN(net_3815) );
NOR4_X2 inst_875 ( .A3(net_4186), .ZN(net_4156), .A4(net_3788), .A1(net_969), .A2(net_706) );
NAND4_X2 inst_1257 ( .A4(net_4003), .ZN(net_3977), .A1(net_3976), .A2(net_3919), .A3(net_3811) );
DFF_X1 inst_3298 ( .QN(net_3006), .D(net_2883), .CK(net_5216) );
AOI22_X2 inst_3482 ( .A1(net_4038), .B2(net_3418), .B1(net_2657), .ZN(net_2655), .A2(net_991) );
INV_X1 inst_3081 ( .A(net_3722), .ZN(net_3547) );
NAND2_X4 inst_1387 ( .ZN(net_2839), .A2(net_2838), .A1(net_2791) );
CLKBUF_X2 inst_5187 ( .A(net_4625), .Z(net_5173) );
CLKBUF_X2 inst_5075 ( .A(net_5060), .Z(net_5061) );
NAND2_X2 inst_1991 ( .A1(net_3534), .ZN(net_3457), .A2(net_3456) );
NAND2_X2 inst_2069 ( .ZN(net_3975), .A2(net_3822), .A1(net_3721) );
INV_X4 inst_2365 ( .ZN(net_1998), .A(net_1826) );
MUX2_X2 inst_2108 ( .S(net_2909), .A(net_2573), .Z(net_2569), .B(net_148) );
AOI22_X2 inst_3572 ( .A1(net_4060), .B1(net_4055), .ZN(net_1478), .B2(net_781), .A2(net_780) );
INV_X16 inst_3066 ( .A(net_3489), .ZN(net_283) );
AND2_X4 inst_4098 ( .A2(net_1548), .ZN(net_1210), .A1(net_1023) );
INV_X4 inst_2250 ( .ZN(net_1514), .A(net_1509) );
INV_X2 inst_2978 ( .ZN(net_185), .A(net_108) );
OAI221_X2 inst_413 ( .C2(net_3720), .A(net_3570), .ZN(net_1562), .B1(net_1207), .C1(net_927), .B2(net_877) );
CLKBUF_X2 inst_5094 ( .A(net_5079), .Z(net_5080) );
INV_X4 inst_2187 ( .ZN(net_2752), .A(net_2519) );
NOR4_X2 inst_859 ( .ZN(net_1879), .A1(net_1829), .A2(net_1042), .A3(net_877), .A4(net_328) );
CLKBUF_X2 inst_4703 ( .A(net_4688), .Z(net_4689) );
INV_X2 inst_2672 ( .ZN(net_1914), .A(net_1883) );
XOR2_X2 inst_25 ( .Z(net_4139), .A(net_4137), .B(net_3385) );
DFF_X1 inst_3323 ( .D(net_4151), .Q(net_3134), .CK(net_4199) );
NAND2_X2 inst_2019 ( .ZN(net_3658), .A2(net_3655), .A1(net_279) );
CLKBUF_X2 inst_5239 ( .A(net_4356), .Z(net_5225) );
AOI22_X2 inst_3527 ( .A2(net_3134), .A1(net_1923), .B1(net_1921), .ZN(net_1917), .B2(net_207) );
CLKBUF_X2 inst_5032 ( .A(net_5017), .Z(net_5018) );
CLKBUF_X2 inst_5166 ( .A(net_5151), .Z(net_5152) );
CLKBUF_X2 inst_5186 ( .A(net_5171), .Z(net_5172) );
INV_X4 inst_2500 ( .A(net_2992), .ZN(net_227) );
XNOR2_X2 inst_69 ( .A(net_3794), .ZN(net_1621), .B(net_1289) );
CLKBUF_X2 inst_4395 ( .A(net_4380), .Z(net_4381) );
CLKBUF_X2 inst_4296 ( .A(net_4281), .Z(net_4282) );
AOI222_X1 inst_3764 ( .A2(net_3151), .C1(net_3118), .A1(net_2055), .B2(net_2054), .C2(net_2053), .ZN(net_1989), .B1(net_1571) );
INV_X2 inst_2669 ( .A(net_3504), .ZN(net_1959) );
NAND2_X2 inst_1691 ( .A1(net_1982), .ZN(net_1979), .A2(net_173) );
OAI211_X2 inst_844 ( .C2(net_4185), .ZN(net_1098), .C1(net_986), .A(net_432), .B(net_207) );
INV_X4 inst_2489 ( .A(net_3157), .ZN(net_1032) );
AOI22_X2 inst_3688 ( .B1(net_4123), .A1(net_555), .ZN(net_490), .A2(net_230), .B2(net_148) );
AOI22_X2 inst_3619 ( .ZN(net_1141), .B1(net_1131), .A1(net_1074), .A2(net_667), .B2(net_399) );
CLKBUF_X2 inst_4641 ( .A(net_4626), .Z(net_4627) );
INV_X4 inst_2340 ( .ZN(net_2376), .A(net_2374) );
OAI21_X4 inst_460 ( .ZN(net_3439), .B2(net_3438), .B1(net_3437), .A(net_3436) );
NAND2_X4 inst_1455 ( .ZN(net_3836), .A2(net_3835), .A1(net_3834) );
DFF_X2 inst_3204 ( .QN(net_3171), .D(net_1364), .CK(net_5267) );
INV_X4 inst_2497 ( .ZN(net_211), .A(net_55) );
AOI22_X2 inst_3660 ( .A1(net_571), .B1(net_570), .ZN(net_569), .A2(net_568), .B2(net_567) );
DFF_X1 inst_3421 ( .Q(net_4033), .D(net_1091), .CK(net_4852) );
CLKBUF_X2 inst_4444 ( .A(net_4429), .Z(net_4430) );
OAI21_X2 inst_560 ( .B2(net_3207), .B1(net_2871), .ZN(net_2865), .A(net_2480) );
INV_X2 inst_2679 ( .ZN(net_1876), .A(net_1822) );
XOR2_X2 inst_16 ( .A(net_4093), .B(net_3418), .Z(net_916) );
CLKBUF_X2 inst_5199 ( .A(net_5184), .Z(net_5185) );
CLKBUF_X2 inst_4230 ( .A(net_4215), .Z(net_4216) );
AOI21_X2 inst_3949 ( .B1(net_2238), .ZN(net_2194), .A(net_2168), .B2(net_1280) );
CLKBUF_X2 inst_4809 ( .A(net_4634), .Z(net_4795) );
INV_X2 inst_2808 ( .ZN(net_689), .A(net_688) );
SDFF_X2 inst_156 ( .SE(net_2625), .D(net_1834), .SI(net_87), .Q(net_87), .CK(net_4975) );
CLKBUF_X2 inst_4617 ( .A(net_4602), .Z(net_4603) );
NAND2_X2 inst_1777 ( .A1(net_4079), .ZN(net_1301), .A2(net_1089) );
NAND2_X2 inst_1802 ( .A1(net_4082), .ZN(net_1975), .A2(net_266) );
NOR2_X4 inst_950 ( .A1(net_3777), .ZN(net_3636), .A2(net_3602) );
NOR2_X2 inst_1068 ( .A1(net_1090), .ZN(net_823), .A2(x947) );
NOR3_X2 inst_886 ( .A2(net_3115), .A1(net_2748), .ZN(net_2747), .A3(net_2746) );
AOI21_X2 inst_3955 ( .ZN(net_1714), .B1(net_1604), .A(net_1547), .B2(net_717) );
INV_X2 inst_2982 ( .A(net_3110), .ZN(net_1960) );
INV_X2 inst_2693 ( .ZN(net_1729), .A(net_1661) );
DFF_X1 inst_3359 ( .D(net_2360), .CK(net_4234), .Q(x423) );
NAND4_X2 inst_1218 ( .A4(net_3984), .ZN(net_997), .A2(net_996), .A1(net_748), .A3(net_679) );
CLKBUF_X2 inst_4418 ( .A(net_4403), .Z(net_4404) );
CLKBUF_X2 inst_4468 ( .A(net_4453), .Z(net_4454) );
XNOR2_X2 inst_96 ( .ZN(net_817), .B(net_587), .A(net_585) );
INV_X2 inst_3020 ( .A(net_3763), .ZN(net_3429) );
XNOR2_X2 inst_101 ( .B(net_874), .ZN(net_617), .A(net_616) );
NAND2_X2 inst_1549 ( .A1(net_2961), .ZN(net_2473), .A2(net_478) );
CLKBUF_X2 inst_4346 ( .A(net_4331), .Z(net_4332) );
AOI22_X2 inst_3555 ( .A1(net_4059), .B1(net_4056), .ZN(net_1495), .B2(net_495), .A2(net_241) );
NAND2_X2 inst_1969 ( .ZN(net_3336), .A1(net_2099), .A2(net_470) );
INV_X2 inst_2881 ( .ZN(net_143), .A(x557) );
OAI211_X2 inst_821 ( .ZN(net_2555), .A(net_1384), .B(net_1304), .C1(net_1204), .C2(net_46) );
NOR2_X4 inst_980 ( .A1(net_3994), .ZN(net_3974), .A2(net_319) );
CLKBUF_X2 inst_4722 ( .A(net_4707), .Z(net_4708) );
OAI21_X2 inst_510 ( .B1(net_3274), .B2(net_2963), .ZN(net_2932), .A(net_2457) );
INV_X4 inst_2436 ( .ZN(net_406), .A(net_266) );
INV_X2 inst_2832 ( .A(net_616), .ZN(net_437) );
NAND2_X2 inst_1677 ( .A1(net_3185), .ZN(net_2080), .A2(net_475) );
OAI21_X2 inst_603 ( .B1(net_2597), .ZN(net_2349), .A(net_2326), .B2(net_375) );
OAI211_X2 inst_830 ( .A(net_3924), .ZN(net_1363), .C1(net_1182), .B(net_1129), .C2(net_900) );
NAND2_X2 inst_1785 ( .A2(net_1613), .A1(net_1332), .ZN(net_1203) );
OAI22_X2 inst_291 ( .A1(net_3781), .B1(net_1884), .ZN(net_1830), .A2(net_1829), .B2(net_263) );
INV_X2 inst_2878 ( .A(net_3153), .ZN(net_1791) );
CLKBUF_X2 inst_4213 ( .A(net_4198), .Z(net_4199) );
DFF_X2 inst_3150 ( .D(net_2305), .QN(net_264), .CK(net_4385) );
INV_X4 inst_2494 ( .A(net_3076), .ZN(net_737) );
OAI21_X1 inst_776 ( .A(net_3331), .ZN(net_1643), .B1(net_931), .B2(net_327) );
INV_X4 inst_2526 ( .A(net_3854), .ZN(net_3268) );
CLKBUF_X2 inst_5047 ( .A(net_5032), .Z(net_5033) );
INV_X4 inst_2286 ( .A(net_1295), .ZN(net_1052) );
NOR4_X2 inst_866 ( .A1(net_1183), .ZN(net_1133), .A3(net_1132), .A4(net_1131), .A2(net_858) );
CLKBUF_X2 inst_5313 ( .A(net_5298), .Z(net_5299) );
INV_X8 inst_2137 ( .ZN(net_322), .A(net_290) );
NAND2_X4 inst_1439 ( .A2(net_4188), .ZN(net_3715), .A1(net_3714) );
NAND2_X2 inst_1972 ( .ZN(net_3340), .A1(net_3287), .A2(net_3277) );
OAI21_X2 inst_558 ( .B2(net_2909), .B1(net_2871), .ZN(net_2867), .A(net_2465) );
AOI22_X2 inst_3640 ( .A1(net_4142), .B1(net_4112), .ZN(net_762), .B2(net_168), .A2(x856) );
OR2_X2 inst_248 ( .A1(net_3352), .ZN(net_2614), .A2(net_2272) );
NAND2_X2 inst_1613 ( .A1(net_2917), .ZN(net_2403), .A2(net_159) );
DFF_X2 inst_3107 ( .QN(net_2997), .D(net_2805), .CK(net_5247) );
CLKBUF_X2 inst_5179 ( .A(net_5164), .Z(net_5165) );
OAI221_X2 inst_389 ( .B1(net_3449), .B2(net_2661), .C1(net_2521), .ZN(net_2505), .A(net_671), .C2(net_670) );
NAND2_X2 inst_1919 ( .A1(net_3165), .ZN(net_246), .A2(net_125) );
INV_X2 inst_2712 ( .A(net_3858), .ZN(net_2838) );
NAND3_X1 inst_1382 ( .A1(net_3514), .ZN(net_3484), .A3(net_3135), .A2(net_931) );
INV_X2 inst_2795 ( .A(net_1007), .ZN(net_754) );
NOR2_X2 inst_1141 ( .A2(net_3858), .ZN(net_3852), .A1(net_3251) );
NAND2_X2 inst_1807 ( .A1(net_4082), .A2(net_1717), .ZN(net_1120) );
AOI22_X2 inst_3589 ( .A1(net_4062), .B1(net_4057), .ZN(net_1428), .A2(net_212), .B2(net_189) );
INV_X4 inst_2488 ( .ZN(net_204), .A(net_49) );
NOR2_X4 inst_932 ( .A1(net_3556), .ZN(net_2025), .A2(net_133) );
CLKBUF_X2 inst_5266 ( .A(net_5251), .Z(net_5252) );
OR3_X2 inst_180 ( .ZN(net_2217), .A1(net_2153), .A2(net_2141), .A3(net_1293) );
NOR3_X2 inst_913 ( .ZN(net_3461), .A2(net_3460), .A1(net_2747), .A3(net_2580) );
CLKBUF_X2 inst_4766 ( .A(net_4751), .Z(net_4752) );
NAND2_X2 inst_1960 ( .ZN(net_3298), .A1(net_3290), .A2(net_2874) );
CLKBUF_X2 inst_4445 ( .A(net_4430), .Z(net_4431) );
CLKBUF_X2 inst_4636 ( .A(net_4621), .Z(net_4622) );
OAI22_X2 inst_302 ( .A1(net_1543), .B1(net_1542), .ZN(net_1540), .A2(net_331), .B2(net_134) );
OAI21_X2 inst_673 ( .ZN(net_1375), .B1(net_1315), .B2(net_1314), .A(net_641) );
AOI22_X2 inst_3585 ( .A1(net_4063), .B1(net_4058), .ZN(net_1432), .A2(net_568), .B2(net_567) );
DFF_X1 inst_3287 ( .QN(net_3049), .D(net_2901), .CK(net_4968) );
OR2_X4 inst_211 ( .A1(net_3408), .A2(net_3406), .ZN(net_1803) );
INV_X4 inst_2483 ( .A(net_3093), .ZN(net_834) );
NOR2_X2 inst_1151 ( .ZN(net_3955), .A2(net_3954), .A1(net_3953) );
CLKBUF_X2 inst_4659 ( .A(net_4644), .Z(net_4645) );
DFF_X2 inst_3120 ( .Q(net_3145), .D(net_2727), .CK(net_4640) );
NAND2_X4 inst_1414 ( .A2(net_3858), .A1(net_3829), .ZN(net_3404) );
OAI21_X2 inst_561 ( .B1(net_4035), .B2(net_2876), .ZN(net_2863), .A(net_2840) );
AOI21_X2 inst_3994 ( .B2(net_3880), .A(net_3858), .ZN(net_3813), .B1(net_3290) );
OAI221_X2 inst_449 ( .ZN(net_4178), .C1(net_4177), .A(net_1826), .B1(net_1502), .C2(net_918), .B2(net_917) );
CLKBUF_X2 inst_4212 ( .A(net_4197), .Z(net_4198) );
INV_X4 inst_2505 ( .A(net_2982), .ZN(net_148) );
INV_X2 inst_2790 ( .ZN(net_795), .A(net_794) );
INV_X8 inst_2138 ( .A(net_3270), .ZN(net_3211) );
NAND2_X2 inst_1641 ( .ZN(net_3213), .A1(net_2086), .A2(net_1986) );
INV_X2 inst_2736 ( .ZN(net_1322), .A(net_1272) );
DFF_X1 inst_3249 ( .QN(net_3082), .D(net_2939), .CK(net_4542) );
OR2_X4 inst_196 ( .A1(net_3645), .ZN(net_2961), .A2(net_2352) );
CLKBUF_X2 inst_4935 ( .A(net_4920), .Z(net_4921) );
NAND2_X2 inst_1567 ( .A1(net_2963), .ZN(net_2454), .A2(net_167) );
CLKBUF_X2 inst_4489 ( .A(net_4423), .Z(net_4475) );
INV_X4 inst_2417 ( .A(net_1521), .ZN(net_1107) );
INV_X4 inst_2309 ( .A(net_1614), .ZN(net_1244) );
NAND2_X4 inst_1403 ( .A2(net_3760), .ZN(net_320), .A1(net_319) );
OAI22_X2 inst_298 ( .A1(net_3781), .A2(net_3500), .B1(net_1884), .ZN(net_1612), .B2(net_1611) );
INV_X4 inst_2180 ( .ZN(net_2649), .A(net_2602) );
NAND2_X2 inst_1856 ( .A2(net_988), .A1(net_778), .ZN(net_615) );
AOI22_X2 inst_3614 ( .ZN(net_1339), .B1(net_1338), .A1(net_1287), .B2(net_1071), .A2(net_1036) );
INV_X4 inst_2603 ( .A(net_3939), .ZN(net_3767) );
CLKBUF_X2 inst_4603 ( .A(net_4588), .Z(net_4589) );
XNOR2_X2 inst_42 ( .ZN(net_2759), .A(net_2692), .B(net_71) );
INV_X8 inst_2153 ( .ZN(net_3394), .A(net_3393) );
AND3_X2 inst_4084 ( .A1(net_4061), .ZN(net_1342), .A2(net_182), .A3(net_156) );
OAI21_X2 inst_588 ( .B2(net_3428), .ZN(net_2632), .B1(net_2512), .A(net_2117) );
NAND2_X4 inst_1479 ( .ZN(net_3949), .A1(net_3948), .A2(net_3612) );
AOI22_X2 inst_3529 ( .A1(net_1955), .B1(net_1921), .ZN(net_1915), .B2(net_371), .A2(net_252) );
NAND2_X2 inst_2040 ( .A2(net_3893), .A1(net_3869), .ZN(net_3800) );
OAI221_X2 inst_437 ( .C2(net_3123), .B2(net_874), .A(net_629), .B1(net_628), .C1(net_627), .ZN(net_622) );
CLKBUF_X2 inst_4742 ( .A(net_4603), .Z(net_4728) );
CLKBUF_X2 inst_4752 ( .A(net_4413), .Z(net_4738) );
NAND3_X2 inst_1356 ( .ZN(net_3702), .A2(net_3698), .A1(net_3389), .A3(net_317) );
NAND2_X2 inst_1706 ( .A1(net_1740), .ZN(net_1737), .A2(net_1690) );
INV_X2 inst_2628 ( .A(net_3532), .ZN(net_2852) );
CLKBUF_X2 inst_4561 ( .A(net_4546), .Z(net_4547) );
INV_X4 inst_2196 ( .ZN(net_2391), .A(net_2326) );
AOI22_X2 inst_3485 ( .A1(net_4038), .B1(net_2657), .ZN(net_2651), .A2(net_393), .B2(net_323) );
INV_X4 inst_2220 ( .ZN(net_1948), .A(net_1909) );
NOR2_X2 inst_1045 ( .ZN(net_1188), .A1(net_1068), .A2(net_1002) );
INV_X2 inst_2743 ( .ZN(net_1216), .A(net_1215) );
OR2_X2 inst_252 ( .A2(net_1507), .ZN(net_1442), .A1(net_1441) );
NOR4_X2 inst_865 ( .ZN(net_1230), .A1(net_1229), .A3(net_1228), .A2(net_1013), .A4(net_640) );
NAND2_X1 inst_2083 ( .A2(net_4011), .A1(net_2959), .ZN(net_2504) );
NOR2_X4 inst_956 ( .A1(net_3888), .ZN(net_3701), .A2(net_3615) );
NAND2_X4 inst_1470 ( .A2(net_3951), .A1(net_3921), .ZN(net_3899) );
CLKBUF_X2 inst_4684 ( .A(net_4669), .Z(net_4670) );
INV_X4 inst_2247 ( .A(net_3331), .ZN(net_1561) );
NAND4_X2 inst_1213 ( .A1(net_3174), .A4(net_3173), .ZN(net_1293), .A2(net_1108), .A3(net_955) );
INV_X1 inst_3072 ( .ZN(net_2367), .A(net_2335) );
OAI21_X2 inst_484 ( .B2(net_3208), .B1(net_2970), .ZN(net_2958), .A(net_2493) );
INV_X4 inst_2452 ( .A(net_3147), .ZN(net_135) );
CLKBUF_X2 inst_4474 ( .A(net_4459), .Z(net_4460) );
XOR2_X1 inst_32 ( .Z(net_364), .A(net_273), .B(net_76) );
OAI221_X2 inst_428 ( .B1(net_3941), .ZN(net_1288), .B2(net_987), .A(net_942), .C1(net_721), .C2(net_329) );
NAND2_X2 inst_1821 ( .A1(net_1213), .ZN(net_1000), .A2(net_371) );
DFF_X1 inst_3418 ( .D(net_1356), .Q(net_35), .CK(net_4293) );
DFF_X1 inst_3334 ( .D(net_2819), .QN(net_315), .CK(net_4319) );
OAI221_X2 inst_407 ( .B2(net_4050), .B1(net_3781), .C2(net_3159), .C1(net_1884), .ZN(net_1752), .A(net_1751) );
AOI22_X2 inst_3558 ( .A1(net_4060), .B1(net_4055), .ZN(net_1492), .A2(net_188), .B2(net_174) );
NAND4_X2 inst_1208 ( .A2(net_1719), .ZN(net_1297), .A3(net_1125), .A1(net_1102), .A4(net_982) );
XNOR2_X2 inst_97 ( .ZN(net_670), .A(net_507), .B(net_410) );
OAI21_X2 inst_616 ( .B2(net_4066), .A(net_3156), .ZN(net_2388), .B1(net_2269) );
OAI21_X1 inst_775 ( .ZN(net_2817), .B1(net_2816), .B2(net_2815), .A(net_1575) );
CLKBUF_X2 inst_4652 ( .A(net_4637), .Z(net_4638) );
OAI21_X2 inst_620 ( .B2(net_2815), .ZN(net_2164), .B1(net_2163), .A(net_1796) );
OAI21_X2 inst_652 ( .ZN(net_1832), .B2(net_1776), .A(net_1775), .B1(net_1635) );
NAND2_X2 inst_1784 ( .ZN(net_1167), .A1(net_1124), .A2(net_530) );
DFF_X2 inst_3118 ( .QN(net_3146), .D(net_2742), .CK(net_4423) );
NAND2_X2 inst_2071 ( .ZN(net_3984), .A2(net_3979), .A1(net_416) );
OAI21_X2 inst_677 ( .B2(net_2717), .ZN(net_1323), .A(net_1311), .B1(net_1025) );
SDFF_X2 inst_130 ( .D(net_3483), .SE(net_3207), .SI(net_3026), .Q(net_3026), .CK(net_5057) );
NAND2_X4 inst_1427 ( .ZN(net_3596), .A2(net_3595), .A1(net_3594) );
NAND2_X2 inst_1566 ( .A1(net_2963), .ZN(net_2455), .A2(net_497) );
NAND2_X4 inst_1409 ( .ZN(net_3299), .A2(net_3298), .A1(net_3226) );
CLKBUF_X2 inst_4662 ( .A(net_4647), .Z(net_4648) );
INV_X4 inst_2242 ( .ZN(net_2661), .A(net_2555) );
XNOR2_X2 inst_87 ( .ZN(net_1025), .A(net_855), .B(net_813) );
CLKBUF_X2 inst_5037 ( .A(net_5022), .Z(net_5023) );
INV_X2 inst_2996 ( .A(net_3038), .ZN(net_193) );
NOR2_X2 inst_1054 ( .A1(net_1132), .ZN(net_1053), .A2(net_684) );
INV_X2 inst_2918 ( .ZN(net_243), .A(net_117) );
NOR2_X4 inst_972 ( .ZN(net_3912), .A2(net_3167), .A1(net_249) );
INV_X2 inst_2721 ( .ZN(net_1634), .A(net_1562) );
NAND2_X2 inst_1671 ( .A1(net_2134), .ZN(net_2087), .A2(net_559) );
INV_X1 inst_3074 ( .A(net_3486), .ZN(net_1684) );
OAI211_X2 inst_800 ( .B(net_2302), .ZN(net_2269), .C1(net_2212), .C2(net_1517), .A(net_994) );
CLKBUF_X2 inst_5281 ( .A(net_5266), .Z(net_5267) );
NAND2_X2 inst_1843 ( .A1(net_4111), .ZN(net_679), .A2(net_590) );
CLKBUF_X2 inst_4581 ( .A(net_4532), .Z(net_4567) );
XOR2_X2 inst_10 ( .B(net_4071), .Z(net_1616), .A(net_1615) );
AOI222_X1 inst_3795 ( .B2(net_4082), .ZN(net_3793), .A1(net_3792), .A2(net_1246), .B1(net_1245), .C1(net_1244), .C2(net_396) );
XOR2_X2 inst_4 ( .B(net_3263), .Z(net_1715), .A(net_1446) );
INV_X2 inst_2884 ( .A(net_3046), .ZN(net_189) );
CLKBUF_X2 inst_4337 ( .A(net_4322), .Z(net_4323) );
OAI21_X2 inst_600 ( .B1(net_3553), .B2(net_2815), .ZN(net_2392), .A(net_1579) );
DFF_X1 inst_3272 ( .QN(net_3099), .D(net_2905), .CK(net_5025) );
CLKBUF_X2 inst_4498 ( .A(net_4483), .Z(net_4484) );
NAND4_X2 inst_1194 ( .ZN(net_1664), .A3(net_1487), .A4(net_1486), .A1(net_1421), .A2(net_1420) );
OR2_X4 inst_204 ( .A1(net_3816), .ZN(net_2972), .A2(net_2352) );
XNOR2_X2 inst_49 ( .ZN(net_2645), .A(net_2334), .B(net_1695) );
NAND2_X2 inst_1866 ( .A1(net_3702), .A2(net_3391), .ZN(net_582) );
NAND2_X2 inst_1550 ( .A1(net_2961), .ZN(net_2472), .A2(net_492) );
NAND2_X2 inst_1878 ( .A1(net_4003), .A2(net_3396), .ZN(net_541) );
CLKBUF_X2 inst_5136 ( .A(net_4820), .Z(net_5122) );
NOR3_X2 inst_910 ( .A3(net_3399), .ZN(net_3337), .A2(net_1882), .A1(net_995) );
AND2_X4 inst_4097 ( .ZN(net_1827), .A1(net_1645), .A2(net_1564) );
OAI21_X2 inst_693 ( .ZN(net_1043), .B1(net_1042), .A(net_940), .B2(net_776) );
CLKBUF_X2 inst_4731 ( .A(net_4716), .Z(net_4717) );
OAI21_X2 inst_765 ( .ZN(net_3944), .A(net_3943), .B1(net_305), .B2(net_277) );
NAND3_X2 inst_1276 ( .ZN(net_2785), .A1(net_2738), .A2(net_2737), .A3(net_1998) );
OR2_X2 inst_256 ( .A1(net_1013), .ZN(net_961), .A2(net_710) );
NAND2_X2 inst_1902 ( .A2(net_3163), .ZN(net_351), .A1(net_350) );
NOR2_X4 inst_937 ( .ZN(net_368), .A2(net_359), .A1(net_306) );
NOR3_X2 inst_908 ( .A1(net_514), .ZN(net_423), .A2(net_264), .A3(net_109) );
OAI222_X2 inst_355 ( .ZN(net_922), .B1(net_921), .C2(net_920), .A1(net_689), .C1(net_662), .A2(net_245), .B2(net_43) );
CLKBUF_X2 inst_5052 ( .A(net_5037), .Z(net_5038) );
OR2_X4 inst_218 ( .A2(net_4091), .ZN(net_1135), .A1(net_1015) );
AOI22_X2 inst_3647 ( .A1(net_4142), .B1(net_4112), .B2(net_2037), .ZN(net_755), .A2(x884) );
AOI22_X2 inst_3498 ( .A1(net_3815), .B1(net_3186), .ZN(net_2175), .A2(net_834), .B2(net_833) );
DFF_X1 inst_3422 ( .Q(net_3173), .D(net_718), .CK(net_4700) );
AOI21_X2 inst_3978 ( .ZN(net_1014), .B1(net_1013), .A(net_925), .B2(net_399) );
AOI221_X2 inst_3832 ( .ZN(net_2313), .A(net_2311), .C2(net_1908), .C1(net_1670), .B2(net_749), .B1(net_105) );
AND4_X4 inst_4039 ( .A1(net_1138), .ZN(net_1102), .A2(net_1101), .A3(net_1100), .A4(net_1092) );
AOI22_X2 inst_3693 ( .B1(net_4123), .A2(net_3023), .B2(net_3022), .A1(net_555), .ZN(net_483) );
INV_X2 inst_2967 ( .ZN(net_1699), .A(net_81) );
AOI222_X1 inst_3769 ( .B1(net_4048), .C1(net_3447), .A1(net_1968), .ZN(net_1963), .C2(net_984), .A2(net_330), .B2(net_72) );
AND4_X2 inst_4053 ( .A4(net_4180), .A1(net_3240), .ZN(net_2192), .A2(net_1878), .A3(net_1766) );
NAND2_X2 inst_2078 ( .ZN(net_4169), .A1(net_4168), .A2(net_73) );
NAND2_X2 inst_1747 ( .ZN(net_1608), .A2(net_1511), .A1(net_1310) );
CLKBUF_X2 inst_5236 ( .A(net_5221), .Z(net_5222) );
CLKBUF_X2 inst_5109 ( .A(net_5094), .Z(net_5095) );
OAI21_X2 inst_699 ( .B2(net_3153), .B1(net_1652), .ZN(net_935), .A(net_401) );
AOI221_X2 inst_3917 ( .ZN(net_3507), .C2(net_1908), .A(net_1824), .C1(net_1667), .B1(net_749), .B2(net_100) );
NAND2_X4 inst_1462 ( .ZN(net_3880), .A2(net_3810), .A1(net_3798) );
INV_X4 inst_2273 ( .A(net_3227), .ZN(net_1017) );
INV_X2 inst_2682 ( .A(net_3773), .ZN(net_1851) );
INV_X4 inst_2574 ( .A(net_3866), .ZN(net_3581) );
CLKBUF_X2 inst_4699 ( .A(net_4622), .Z(net_4685) );
INV_X4 inst_2229 ( .ZN(net_1757), .A(net_1723) );
NAND2_X2 inst_2003 ( .ZN(net_3512), .A1(net_3510), .A2(net_2364) );
CLKBUF_X2 inst_5119 ( .A(net_4666), .Z(net_5105) );
CLKBUF_X2 inst_4963 ( .A(net_4948), .Z(net_4949) );
CLKBUF_X2 inst_4749 ( .A(net_4610), .Z(net_4735) );
NOR2_X4 inst_964 ( .ZN(net_3812), .A1(net_2135), .A2(net_2111) );
INV_X2 inst_2787 ( .ZN(net_799), .A(net_798) );
DFF_X1 inst_3372 ( .D(net_2284), .QN(net_63), .CK(net_4213) );
INV_X4 inst_2599 ( .A(net_3995), .ZN(net_3754) );
INV_X4 inst_2426 ( .A(net_323), .ZN(net_250) );
NAND4_X2 inst_1245 ( .A3(net_3648), .ZN(net_3528), .A2(net_3249), .A4(net_3189), .A1(net_2090) );
INV_X4 inst_2313 ( .ZN(net_943), .A(net_774) );
AOI21_X2 inst_3971 ( .A(net_3157), .ZN(net_1276), .B1(net_1275), .B2(net_1274) );
AOI222_X1 inst_3788 ( .A2(net_1826), .ZN(net_1461), .A1(net_979), .B1(net_625), .C1(net_581), .C2(net_402), .B2(net_333) );
NAND2_X4 inst_1485 ( .ZN(net_4006), .A1(net_3397), .A2(net_3167) );
AOI22_X2 inst_3663 ( .A1(net_571), .B1(net_570), .ZN(net_564), .A2(net_180), .B2(net_154) );
INV_X2 inst_3001 ( .A(net_3131), .ZN(net_1326) );
INV_X2 inst_2818 ( .A(net_988), .ZN(net_784) );
INV_X2 inst_3008 ( .ZN(net_3305), .A(net_3304) );
DFF_X2 inst_3198 ( .QN(net_3169), .D(net_1625), .CK(net_5271) );
OAI22_X2 inst_317 ( .B2(net_3941), .A1(net_1975), .B1(net_1332), .ZN(net_1122), .A2(net_977) );
OAI21_X2 inst_750 ( .ZN(net_3427), .B2(net_3426), .A(net_3425), .B1(net_1605) );
NOR2_X2 inst_1123 ( .ZN(net_3436), .A2(net_3435), .A1(net_3433) );
INV_X2 inst_2904 ( .ZN(net_156), .A(net_115) );
CLKBUF_X2 inst_4429 ( .A(net_4414), .Z(net_4415) );
OAI22_X4 inst_278 ( .ZN(net_3774), .B2(net_3773), .B1(net_3772), .A2(net_3771), .A1(net_3770) );
INV_X4 inst_2383 ( .A(net_1071), .ZN(net_433) );
NAND2_X2 inst_1701 ( .ZN(net_2076), .A1(net_1790), .A2(net_1735) );
OAI21_X4 inst_467 ( .ZN(net_3906), .A(net_3900), .B2(net_3727), .B1(net_3562) );
AOI22_X2 inst_3677 ( .B1(net_4124), .ZN(net_524), .A1(net_509), .B2(net_242), .A2(net_147) );
AND3_X4 inst_4071 ( .ZN(net_4038), .A3(net_3559), .A1(net_2345), .A2(net_656) );
CLKBUF_X2 inst_4987 ( .A(net_4972), .Z(net_4973) );
INV_X2 inst_2963 ( .ZN(net_272), .A(net_80) );
NAND2_X2 inst_1628 ( .A2(net_3860), .A1(net_3510), .ZN(net_2515) );
NAND3_X2 inst_1329 ( .A2(net_3628), .ZN(net_1168), .A3(net_655), .A1(net_446) );
INV_X4 inst_2469 ( .ZN(net_294), .A(net_65) );
NAND4_X2 inst_1204 ( .ZN(net_1849), .A4(net_1499), .A3(net_1469), .A2(net_1435), .A1(net_1430) );
AND3_X4 inst_4066 ( .A3(net_3441), .A2(net_3156), .ZN(net_1645), .A1(net_1527) );
CLKBUF_X2 inst_4840 ( .A(net_4603), .Z(net_4826) );
OR2_X4 inst_225 ( .ZN(net_727), .A1(net_716), .A2(net_439) );
CLKBUF_X2 inst_5020 ( .A(net_4436), .Z(net_5006) );
OAI21_X2 inst_508 ( .B1(net_3274), .B2(net_2967), .ZN(net_2934), .A(net_2407) );
CLKBUF_X2 inst_4888 ( .A(net_4574), .Z(net_4874) );
CLKBUF_X2 inst_4736 ( .A(net_4286), .Z(net_4722) );
INV_X4 inst_2618 ( .ZN(net_3894), .A(net_3892) );
NOR2_X2 inst_1135 ( .ZN(net_3665), .A1(net_3615), .A2(net_530) );
CLKBUF_X2 inst_4950 ( .A(net_4935), .Z(net_4936) );
AOI22_X2 inst_3715 ( .ZN(net_3464), .A2(net_1717), .A1(net_1522), .B1(net_1137), .B2(net_912) );
OAI21_X2 inst_590 ( .B1(net_3691), .B2(net_3229), .ZN(net_2593), .A(net_72) );
INV_X4 inst_2553 ( .A(net_3644), .ZN(net_3477) );
DFF_X2 inst_3127 ( .QN(net_3144), .D(net_2681), .CK(net_4766) );
INV_X2 inst_3042 ( .A(net_3885), .ZN(net_3685) );
DFF_X1 inst_3243 ( .QN(net_3085), .D(net_2955), .CK(net_4559) );
NAND2_X2 inst_1729 ( .ZN(net_1557), .A1(net_1556), .A2(x825) );
CLKBUF_X2 inst_4531 ( .A(net_4516), .Z(net_4517) );
NOR2_X2 inst_1105 ( .A1(net_3871), .ZN(net_3218), .A2(net_3018) );
INV_X2 inst_2746 ( .A(net_3641), .ZN(net_1266) );
NOR2_X4 inst_981 ( .ZN(net_3986), .A2(net_3168), .A1(net_3106) );
NAND3_X4 inst_1266 ( .A1(net_3901), .ZN(net_3576), .A3(net_3575), .A2(net_3452) );
CLKBUF_X2 inst_4648 ( .A(net_4295), .Z(net_4634) );
NAND2_X1 inst_2094 ( .A1(net_3817), .ZN(net_3183), .A2(net_155) );
CLKBUF_X2 inst_5102 ( .A(net_5087), .Z(net_5088) );
CLKBUF_X2 inst_4872 ( .A(net_4857), .Z(net_4858) );
CLKBUF_X2 inst_4317 ( .A(net_4302), .Z(net_4303) );
OAI22_X2 inst_330 ( .A2(net_881), .ZN(net_839), .A1(net_727), .B1(net_637), .B2(net_549) );
DFF_X1 inst_3417 ( .D(net_1357), .Q(net_34), .CK(net_4465) );
AOI22_X1 inst_3733 ( .ZN(net_3865), .A1(net_3815), .B2(net_3186), .B1(net_190), .A2(net_161) );
OR3_X4 inst_165 ( .A2(net_3773), .ZN(net_2142), .A1(net_2118), .A3(net_1927) );
CLKBUF_X2 inst_4305 ( .A(net_4222), .Z(net_4291) );
AOI22_X2 inst_3491 ( .A2(net_3128), .ZN(net_2507), .B1(net_2300), .A1(net_2296), .B2(net_671) );
AOI22_X2 inst_3566 ( .A1(net_4060), .B1(net_4055), .ZN(net_1484), .B2(net_199), .A2(net_165) );
INV_X4 inst_2393 ( .A(net_1884), .ZN(net_1882) );
NAND4_X4 inst_1176 ( .A3(net_4140), .A1(net_3643), .ZN(net_3548), .A2(net_3106), .A4(net_278) );
NAND2_X2 inst_1838 ( .ZN(net_1340), .A2(net_1036), .A1(net_356) );
XNOR2_X2 inst_71 ( .A(net_1583), .ZN(net_1582), .B(net_207) );
NAND2_X4 inst_1454 ( .A2(net_4165), .ZN(net_3832), .A1(net_3753) );
AND3_X4 inst_4079 ( .ZN(net_4116), .A3(net_3662), .A2(net_528), .A1(net_337) );
NAND4_X2 inst_1232 ( .ZN(net_2220), .A3(net_556), .A2(net_510), .A4(net_459), .A1(net_443) );
DFF_X1 inst_3231 ( .QN(net_3068), .D(net_2960), .CK(net_4875) );
DFF_X2 inst_3147 ( .D(net_2392), .QN(net_113), .CK(net_4418) );
NAND2_X2 inst_1945 ( .A1(net_3815), .ZN(net_3249), .A2(net_208) );
AND2_X4 inst_4172 ( .ZN(net_4126), .A1(net_3397), .A2(net_3167) );
INV_X2 inst_2657 ( .A(net_2699), .ZN(net_2195) );
INV_X4 inst_2605 ( .ZN(net_3782), .A(net_3781) );
OAI21_X2 inst_758 ( .ZN(net_3739), .A(net_2735), .B1(net_2693), .B2(net_2690) );
OAI22_X2 inst_336 ( .B1(net_3122), .ZN(net_438), .A1(net_344), .B2(net_263), .A2(net_250) );
INV_X8 inst_2146 ( .ZN(net_3274), .A(net_3273) );
INV_X2 inst_2703 ( .ZN(net_1673), .A(net_1672) );
OAI221_X2 inst_376 ( .ZN(net_2671), .B1(net_2670), .B2(net_2669), .C1(net_2668), .A(net_1386), .C2(net_318) );
CLKBUF_X2 inst_5157 ( .A(net_4310), .Z(net_5143) );
NAND2_X2 inst_1939 ( .A2(net_3618), .ZN(net_3226), .A1(net_3225) );
DFF_X1 inst_3268 ( .QN(net_3096), .D(net_2904), .CK(net_5035) );
INV_X2 inst_2902 ( .A(net_318), .ZN(net_179) );
SDFF_X2 inst_143 ( .D(net_3882), .SE(net_2625), .SI(net_95), .Q(net_95), .CK(net_5048) );
NAND2_X2 inst_1953 ( .ZN(net_3282), .A2(net_3281), .A1(net_495) );
CLKBUF_X2 inst_5286 ( .A(net_5202), .Z(net_5272) );
CLKBUF_X2 inst_4570 ( .A(net_4234), .Z(net_4556) );
INV_X2 inst_3016 ( .ZN(net_3410), .A(net_2562) );
CLKBUF_X2 inst_4272 ( .A(net_4243), .Z(net_4258) );
NAND2_X2 inst_1958 ( .A1(net_3530), .A2(net_3513), .ZN(net_3297) );
INV_X4 inst_2337 ( .A(net_711), .ZN(net_657) );
DFF_X1 inst_3250 ( .D(net_3267), .QN(net_3090), .CK(net_4736) );
DFF_X1 inst_3240 ( .QN(net_3038), .D(net_2956), .CK(net_5186) );
NAND2_X2 inst_1778 ( .A2(net_2523), .A1(net_2518), .ZN(net_1151) );
CLKBUF_X2 inst_5174 ( .A(net_5159), .Z(net_5160) );
NAND2_X2 inst_1736 ( .A2(net_4082), .ZN(net_1530), .A1(net_1528) );
NOR2_X2 inst_1040 ( .A1(net_1458), .A2(net_1340), .ZN(net_1215) );
AOI211_X2 inst_4027 ( .C1(net_3962), .B(net_1606), .ZN(net_1034), .C2(net_928), .A(net_404) );
AOI221_X2 inst_3880 ( .A(net_4047), .C2(net_1908), .ZN(net_1848), .C1(net_1847), .B2(net_749), .B1(net_90) );
HA_X1 inst_3100 ( .S(net_643), .CO(net_642), .B(net_423), .A(net_224) );
CLKBUF_X2 inst_5042 ( .A(net_5027), .Z(net_5028) );
AND4_X4 inst_4052 ( .ZN(net_4107), .A2(net_3940), .A4(net_3395), .A3(net_594), .A1(net_376) );
CLKBUF_X2 inst_4251 ( .A(net_4236), .Z(net_4237) );
CLKBUF_X2 inst_4487 ( .A(net_4472), .Z(net_4473) );
XNOR2_X2 inst_111 ( .A(net_4132), .ZN(net_417), .B(net_402) );
NAND2_X2 inst_1596 ( .A1(net_2925), .ZN(net_2422), .A2(net_183) );
CLKBUF_X2 inst_4364 ( .A(net_4237), .Z(net_4350) );
DFF_X2 inst_3146 ( .QN(net_3127), .D(net_2509), .CK(net_5146) );
NAND2_X2 inst_1723 ( .ZN(net_1596), .A2(net_1595), .A1(net_1506) );
DFF_X1 inst_3278 ( .QN(net_3034), .D(net_2906), .CK(net_5010) );
CLKBUF_X2 inst_5145 ( .A(net_5130), .Z(net_5131) );
NAND2_X2 inst_2056 ( .ZN(net_3904), .A1(net_3901), .A2(net_3833) );
AOI222_X1 inst_3752 ( .A1(net_3676), .B1(net_2055), .C1(net_2054), .ZN(net_2041), .B2(net_1797), .C2(net_643), .A2(net_267) );
INV_X8 inst_2116 ( .ZN(net_2923), .A(net_2891) );
INV_X4 inst_2265 ( .A(net_2127), .ZN(net_2054) );
OAI22_X2 inst_284 ( .A1(net_3611), .A2(net_2838), .ZN(net_2347), .B1(net_2324), .B2(net_2323) );
CLKBUF_X2 inst_5071 ( .A(net_5056), .Z(net_5057) );
INV_X2 inst_2825 ( .ZN(net_640), .A(net_526) );
NAND2_X2 inst_1555 ( .A1(net_2909), .ZN(net_2467), .A2(net_170) );
AOI211_X2 inst_4031 ( .ZN(net_3246), .C1(net_1363), .B(net_1185), .A(net_999), .C2(net_337) );
NAND3_X2 inst_1293 ( .ZN(net_2143), .A1(net_2142), .A2(net_1890), .A3(net_1845) );
AOI221_X2 inst_3805 ( .B2(net_4031), .ZN(net_2754), .B1(net_2752), .C1(net_2710), .A(net_2505), .C2(net_145) );
INV_X4 inst_2579 ( .ZN(net_3606), .A(net_3605) );
OAI22_X2 inst_280 ( .ZN(net_2822), .A1(net_2748), .B1(net_2615), .B2(net_1214), .A2(net_901) );
OAI22_X2 inst_346 ( .A2(net_3989), .ZN(net_3964), .B2(net_3960), .B1(net_1340), .A1(net_1006) );
DFF_X2 inst_3157 ( .D(net_2179), .QN(net_44), .CK(net_4625) );
NOR2_X4 inst_978 ( .ZN(net_3957), .A1(net_3956), .A2(net_3675) );
NAND2_X2 inst_1713 ( .A1(net_3782), .ZN(net_1814), .A2(net_1271) );
INV_X2 inst_2955 ( .A(net_3050), .ZN(net_171) );
AOI21_X4 inst_3926 ( .B1(net_3957), .B2(net_3763), .ZN(net_3574), .A(net_399) );
CLKBUF_X2 inst_4527 ( .A(net_4512), .Z(net_4513) );
AOI21_X4 inst_3929 ( .B2(net_3860), .ZN(net_3591), .B1(net_3366), .A(net_2708) );
DFF_X2 inst_3137 ( .QN(net_2988), .D(net_2568), .CK(net_5095) );
CLKBUF_X2 inst_4676 ( .A(net_4661), .Z(net_4662) );
AOI221_X2 inst_3852 ( .ZN(net_2062), .A(net_2060), .C2(net_1908), .C1(net_1678), .B2(net_749), .B1(net_102) );
CLKBUF_X2 inst_4496 ( .A(net_4197), .Z(net_4482) );
INV_X4 inst_2566 ( .A(net_3568), .ZN(net_3523) );
OAI21_X2 inst_495 ( .B1(net_3278), .ZN(net_2947), .B2(net_2907), .A(net_2482) );
NOR2_X2 inst_1051 ( .ZN(net_1158), .A1(net_1035), .A2(net_751) );
NOR2_X4 inst_951 ( .ZN(net_3661), .A1(net_3660), .A2(net_346) );
NAND2_X2 inst_1864 ( .ZN(net_1381), .A2(net_588), .A1(net_406) );
AOI22_X2 inst_3603 ( .A1(net_4063), .B1(net_4058), .A2(net_3027), .B2(net_3026), .ZN(net_1414) );
DFF_X1 inst_3224 ( .QN(net_3056), .D(net_2977), .CK(net_4740) );
CLKBUF_X2 inst_4393 ( .A(net_4378), .Z(net_4379) );
INV_X2 inst_3043 ( .A(net_3889), .ZN(net_3699) );
NAND3_X2 inst_1359 ( .A3(net_3836), .ZN(net_3802), .A2(net_3801), .A1(net_1371) );
DFF_X2 inst_3188 ( .D(net_1731), .QN(net_121), .CK(net_5137) );
DFF_X2 inst_3129 ( .D(net_2697), .QN(net_43), .CK(net_4636) );
CLKBUF_X2 inst_4674 ( .A(net_4659), .Z(net_4660) );
INV_X2 inst_2893 ( .A(net_3033), .ZN(net_187) );
OAI21_X2 inst_573 ( .B2(net_2815), .ZN(net_2814), .B1(net_2813), .A(net_1573) );
AOI221_X2 inst_3797 ( .C1(net_4035), .C2(net_3738), .B1(net_3736), .ZN(net_2840), .B2(net_2623), .A(net_1992) );
XNOR2_X2 inst_100 ( .ZN(net_1291), .A(net_538), .B(net_43) );
CLKBUF_X2 inst_4352 ( .A(net_4337), .Z(net_4338) );
CLKBUF_X2 inst_4245 ( .A(net_4212), .Z(net_4231) );
NOR2_X4 inst_921 ( .A2(net_3367), .ZN(net_2890), .A1(net_2859) );
NAND2_X4 inst_1453 ( .ZN(net_3833), .A1(net_3832), .A2(net_3606) );
OAI22_X2 inst_279 ( .ZN(net_2809), .A2(net_2785), .B1(net_2764), .A1(net_2193), .B2(net_2064) );
AOI21_X2 inst_3970 ( .ZN(net_1588), .A(net_1220), .B2(net_1011), .B1(net_836) );
DFF_X1 inst_3387 ( .D(net_1777), .CK(net_5291), .Q(x626) );
INV_X2 inst_3007 ( .ZN(net_3258), .A(net_2309) );
XNOR2_X2 inst_81 ( .ZN(net_1269), .A(net_1080), .B(net_248) );
AND2_X4 inst_4185 ( .ZN(net_4149), .A1(net_3947), .A2(net_3108) );
AOI22_X2 inst_3544 ( .B1(net_4054), .A2(net_2033), .ZN(net_1579), .A1(net_1578), .B2(net_1280) );
AOI22_X2 inst_3512 ( .ZN(net_1972), .B1(net_1882), .A2(net_1879), .A1(net_1810), .B2(net_198) );
OAI211_X2 inst_790 ( .C2(net_2876), .ZN(net_2706), .A(net_2634), .C1(net_2633), .B(net_2047) );
NOR2_X2 inst_1009 ( .ZN(net_1780), .A1(net_1779), .A2(net_1778) );
NAND4_X2 inst_1206 ( .ZN(net_2067), .A3(net_1489), .A4(net_1488), .A2(net_1423), .A1(net_1422) );
INV_X2 inst_2954 ( .A(net_3012), .ZN(net_221) );
INV_X4 inst_2197 ( .A(net_3860), .ZN(net_2322) );
OAI21_X2 inst_733 ( .A(net_629), .B2(net_628), .ZN(net_577), .B1(net_204) );
AOI22_X2 inst_3466 ( .B2(net_4027), .B1(net_2752), .ZN(net_2751), .A1(net_2750), .A2(net_1523) );
NAND2_X2 inst_1959 ( .A2(net_3600), .ZN(net_3300), .A1(net_3299) );
INV_X4 inst_2582 ( .ZN(net_3627), .A(net_3620) );
SDFF_X2 inst_142 ( .SE(net_2514), .D(net_2288), .SI(net_102), .Q(net_102), .CK(net_4749) );
CLKBUF_X2 inst_4800 ( .A(net_4303), .Z(net_4786) );
CLKBUF_X2 inst_4394 ( .A(net_4379), .Z(net_4380) );
XNOR2_X2 inst_78 ( .A(net_1522), .ZN(net_1379), .B(net_1140) );
NAND2_X2 inst_1487 ( .A1(net_4155), .A2(net_3600), .ZN(net_2894) );
INV_X2 inst_2813 ( .A(net_838), .ZN(net_639) );
OR3_X4 inst_177 ( .ZN(net_3360), .A2(net_2815), .A1(net_2550), .A3(net_1737) );
OAI211_X2 inst_783 ( .ZN(net_2779), .C2(net_2778), .B(net_2676), .C1(net_2661), .A(net_2654) );
AOI22_X2 inst_3522 ( .A2(net_3141), .B2(net_3140), .ZN(net_1924), .A1(net_1923), .B1(net_1921) );
NAND2_X2 inst_1933 ( .ZN(net_3200), .A1(net_3198), .A2(net_166) );
NAND2_X2 inst_2014 ( .ZN(net_3634), .A2(net_3632), .A1(net_3543) );
CLKBUF_X2 inst_4471 ( .A(net_4355), .Z(net_4457) );
NOR2_X2 inst_1142 ( .ZN(net_3863), .A2(net_3862), .A1(net_3861) );
NAND2_X2 inst_1758 ( .A2(net_1394), .ZN(net_1241), .A1(net_31) );
CLKBUF_X2 inst_4320 ( .A(net_4305), .Z(net_4306) );
OAI21_X2 inst_615 ( .ZN(net_2325), .B1(net_2282), .B2(net_1853), .A(net_356) );
AOI221_X2 inst_3816 ( .A(net_2642), .B1(net_2641), .C2(net_2583), .ZN(net_2582), .C1(net_2581), .B2(net_287) );
INV_X2 inst_2822 ( .ZN(net_535), .A(net_534) );
INV_X4 inst_2467 ( .ZN(net_1511), .A(net_58) );
AOI221_X2 inst_3843 ( .B2(net_2203), .C1(net_2202), .ZN(net_2199), .A(net_2073), .C2(net_1797), .B1(net_1769) );
NAND3_X1 inst_1381 ( .ZN(net_3462), .A2(net_2680), .A1(net_1319), .A3(net_1217) );
NAND2_X2 inst_2031 ( .ZN(net_3762), .A1(net_3761), .A2(net_3606) );
CLKBUF_X2 inst_4386 ( .A(net_4371), .Z(net_4372) );
OAI21_X2 inst_643 ( .B1(net_1993), .ZN(net_1992), .A(net_1900), .B2(net_1545) );
CLKBUF_X2 inst_4771 ( .A(net_4756), .Z(net_4757) );
CLKBUF_X2 inst_4941 ( .A(net_4926), .Z(net_4927) );
CLKBUF_X2 inst_5133 ( .A(net_4596), .Z(net_5119) );
CLKBUF_X2 inst_4961 ( .A(net_4644), .Z(net_4947) );
CLKBUF_X2 inst_4669 ( .A(net_4536), .Z(net_4655) );
OAI22_X2 inst_338 ( .B2(net_3196), .B1(net_635), .ZN(net_420), .A2(net_381), .A1(net_210) );
INV_X4 inst_2412 ( .ZN(net_2180), .A(net_269) );
CLKBUF_X2 inst_4928 ( .A(net_4913), .Z(net_4914) );
AOI21_X2 inst_4005 ( .ZN(net_3915), .A(net_3914), .B1(net_650), .B2(net_592) );
CLKBUF_X2 inst_4323 ( .A(net_4308), .Z(net_4309) );
INV_X4 inst_2214 ( .ZN(net_2238), .A(net_2142) );
AND2_X4 inst_4146 ( .A2(net_4111), .A1(net_4102), .ZN(net_4083) );
NAND2_X2 inst_1997 ( .A2(net_3514), .ZN(net_3487), .A1(net_931) );
INV_X4 inst_2474 ( .A(net_3069), .ZN(net_732) );
NOR2_X2 inst_1017 ( .ZN(net_1731), .A1(net_1631), .A2(net_1090) );
OAI21_X2 inst_579 ( .B2(net_2909), .B1(net_2803), .ZN(net_2799), .A(net_2468) );
CLKBUF_X2 inst_5247 ( .A(net_4733), .Z(net_5233) );
AOI222_X2 inst_3736 ( .B2(net_4109), .C2(net_1791), .C1(net_1244), .ZN(net_1199), .A1(net_1198), .B1(net_1118), .A2(net_920) );
INV_X4 inst_2495 ( .A(net_3148), .ZN(net_252) );
INV_X4 inst_2297 ( .ZN(net_1103), .A(net_1046) );
AOI211_X2 inst_4019 ( .C2(net_4098), .A(net_4070), .ZN(net_1647), .B(net_1646), .C1(net_55) );
DFF_X1 inst_3341 ( .D(net_2777), .QN(net_116), .CK(net_4452) );
OAI22_X2 inst_281 ( .B1(net_3463), .A1(net_3462), .ZN(net_2770), .A2(net_1764), .B2(net_1620) );
DFF_X1 inst_3236 ( .QN(net_3042), .D(net_2946), .CK(net_5044) );
OAI21_X2 inst_698 ( .B1(net_4087), .ZN(net_2596), .A(net_1274), .B2(net_270) );
NAND2_X2 inst_1836 ( .A1(net_1107), .ZN(net_1042), .A2(net_594) );
AOI21_X2 inst_3964 ( .B2(net_3702), .A(net_3640), .ZN(net_1454), .B1(net_886) );
AOI21_X2 inst_3944 ( .B1(net_3774), .ZN(net_2226), .A(net_2149), .B2(net_330) );
DFF_X1 inst_3394 ( .Q(net_3113), .D(net_1536), .CK(net_4316) );
DFF_X1 inst_3408 ( .D(net_1399), .Q(net_36), .CK(net_4498) );
XNOR2_X2 inst_88 ( .ZN(net_979), .B(net_978), .A(net_871) );
INV_X2 inst_2863 ( .ZN(net_2181), .A(net_286) );
INV_X4 inst_2508 ( .ZN(net_239), .A(net_70) );
CLKBUF_X2 inst_4274 ( .A(net_4259), .Z(net_4260) );
CLKBUF_X2 inst_4250 ( .A(net_4235), .Z(net_4236) );
INV_X8 inst_2170 ( .ZN(net_3999), .A(net_138) );
OAI221_X2 inst_360 ( .ZN(net_2827), .B1(net_2826), .C1(net_2825), .A(net_2585), .C2(net_1519), .B2(net_645) );
AOI221_X2 inst_3897 ( .ZN(net_1304), .B1(net_1244), .C1(net_1198), .A(net_1121), .C2(net_714), .B2(net_168) );
OAI21_X1 inst_773 ( .ZN(net_4018), .B2(net_2963), .B1(net_2893), .A(net_2461) );
INV_X2 inst_2946 ( .A(net_2990), .ZN(net_177) );
AOI221_X2 inst_3908 ( .A(net_4185), .B2(net_4111), .ZN(net_1343), .C2(net_923), .C1(net_902), .B1(net_651) );
AOI22_X2 inst_3620 ( .B1(net_1244), .A1(net_1198), .ZN(net_1128), .A2(net_874), .B2(net_378) );
AOI222_X1 inst_3754 ( .A1(net_3676), .A2(net_3133), .B1(net_2055), .C1(net_2054), .ZN(net_2039), .C2(net_1038), .B2(net_396) );
OR2_X2 inst_260 ( .A2(net_3221), .A1(net_2376), .ZN(net_763) );
NOR2_X2 inst_1129 ( .ZN(net_3554), .A1(net_3551), .A2(net_3495) );
OAI211_X2 inst_837 ( .C2(net_2665), .C1(net_1359), .ZN(net_1353), .A(net_1235), .B(net_593) );
OAI21_X2 inst_744 ( .ZN(net_3325), .A(net_3324), .B2(net_3319), .B1(net_655) );
CLKBUF_X2 inst_4973 ( .A(net_4958), .Z(net_4959) );
DFF_X2 inst_3211 ( .D(net_808), .QN(net_505), .CK(net_4667) );
AOI221_X2 inst_3827 ( .B1(net_3469), .C2(net_3133), .B2(net_3132), .C1(net_2534), .ZN(net_2533), .A(net_2338) );
AND2_X4 inst_4139 ( .ZN(net_4069), .A1(net_960), .A2(net_828) );
AND2_X4 inst_4112 ( .A2(net_4131), .ZN(net_3390), .A1(net_3389) );
CLKBUF_X2 inst_4611 ( .A(net_4596), .Z(net_4597) );
CLKBUF_X2 inst_4567 ( .A(net_4552), .Z(net_4553) );
AOI221_X2 inst_3889 ( .B1(net_4026), .C1(net_3140), .A(net_2525), .ZN(net_1397), .B2(net_1394), .C2(net_1393) );
XNOR2_X2 inst_65 ( .ZN(net_1754), .A(net_1649), .B(net_1379) );
OAI21_X2 inst_536 ( .B1(net_3195), .B2(net_2961), .ZN(net_2897), .A(net_2475) );
AOI22_X2 inst_3592 ( .A1(net_4063), .B1(net_4058), .ZN(net_1425), .A2(net_219), .B2(net_160) );
INV_X4 inst_2386 ( .ZN(net_1071), .A(net_401) );
CLKBUF_X2 inst_5121 ( .A(net_4201), .Z(net_5107) );
OAI21_X2 inst_516 ( .B1(net_3302), .ZN(net_2926), .B2(net_2925), .A(net_2422) );
AOI22_X1 inst_3732 ( .ZN(net_3610), .B1(net_3219), .A1(net_2134), .A2(net_244), .B2(net_139) );
INV_X4 inst_2258 ( .ZN(net_1620), .A(net_1127) );
OR2_X4 inst_190 ( .A1(net_2615), .ZN(net_2609), .A2(net_2268) );
AND2_X4 inst_4103 ( .A1(net_920), .A2(net_449), .ZN(net_448) );
NAND3_X4 inst_1267 ( .A1(net_3928), .ZN(net_3834), .A3(net_3726), .A2(net_451) );
NAND2_X2 inst_1507 ( .A2(net_3686), .A1(net_3536), .ZN(net_2695) );
CLKBUF_X2 inst_4503 ( .A(net_4488), .Z(net_4489) );
CLKBUF_X2 inst_4907 ( .A(net_4458), .Z(net_4893) );
CLKBUF_X2 inst_4873 ( .A(net_4858), .Z(net_4859) );
NAND2_X2 inst_2027 ( .A1(net_4164), .A2(net_4162), .ZN(net_3734) );
INV_X2 inst_2926 ( .A(net_3034), .ZN(net_154) );
OAI221_X2 inst_416 ( .B1(net_4067), .ZN(net_1302), .A(net_1301), .C2(net_1228), .C1(net_1105), .B2(net_1011) );
NOR2_X2 inst_1158 ( .ZN(net_4091), .A1(net_3789), .A2(net_745) );
NAND2_X2 inst_1870 ( .A1(net_920), .ZN(net_712), .A2(net_538) );
NAND2_X2 inst_2062 ( .ZN(net_3920), .A1(net_3108), .A2(net_3107) );
AOI222_X1 inst_3786 ( .C2(net_4125), .A2(net_3755), .ZN(net_1335), .A1(net_1164), .C1(net_788), .B1(net_638), .B2(net_383) );
INV_X4 inst_2350 ( .ZN(net_1090), .A(net_671) );
NAND2_X4 inst_1406 ( .ZN(net_3273), .A1(net_3272), .A2(net_2062) );
DFF_X1 inst_3404 ( .D(net_1464), .CK(net_5248), .Q(x593) );
CLKBUF_X2 inst_5270 ( .A(net_5156), .Z(net_5256) );
OAI21_X2 inst_542 ( .ZN(net_4014), .B2(net_3208), .B1(net_2893), .A(net_2496) );
SDFF_X2 inst_128 ( .D(net_3483), .SI(net_3029), .Q(net_3029), .SE(net_2925), .CK(net_5066) );
CLKBUF_X2 inst_4319 ( .A(net_4304), .Z(net_4305) );
INV_X4 inst_2445 ( .A(net_3064), .ZN(net_518) );
CLKBUF_X2 inst_4432 ( .A(net_4417), .Z(net_4418) );
INV_X2 inst_3039 ( .ZN(net_3642), .A(net_3168) );
NOR2_X4 inst_973 ( .ZN(net_3919), .A1(net_3918), .A2(net_380) );
AOI21_X2 inst_4000 ( .ZN(net_3706), .B2(net_3705), .B1(net_3704), .A(net_3703) );
INV_X2 inst_3058 ( .ZN(net_3988), .A(net_3987) );
OAI21_X4 inst_461 ( .ZN(net_3504), .B2(net_3503), .B1(net_3500), .A(net_3156) );
DFF_X1 inst_3218 ( .D(net_3245), .QN(net_3126), .CK(net_5005) );
OAI211_X2 inst_829 ( .ZN(net_1821), .C1(net_1124), .A(net_726), .B(net_594), .C2(net_530) );
OR2_X4 inst_197 ( .A1(net_3645), .ZN(net_2909), .A2(net_2354) );
CLKBUF_X2 inst_4702 ( .A(net_4687), .Z(net_4688) );
INV_X2 inst_2958 ( .ZN(net_210), .A(net_123) );
NAND2_X2 inst_1973 ( .A1(net_3877), .A2(net_3859), .ZN(net_3344) );
HA_X1 inst_3089 ( .A(net_3492), .S(net_1709), .CO(net_1708), .B(net_1316) );
XOR2_X2 inst_24 ( .A(net_4113), .Z(net_4093), .B(net_393) );
INV_X2 inst_3051 ( .ZN(net_3840), .A(net_3835) );
INV_X2 inst_2668 ( .ZN(net_2005), .A(net_1972) );
NOR2_X2 inst_1122 ( .ZN(net_3424), .A2(net_3423), .A1(net_3412) );
DFF_X1 inst_3324 ( .D(net_2834), .Q(net_72), .CK(net_4272) );
NAND4_X2 inst_1209 ( .ZN(net_1262), .A4(net_1261), .A2(net_1060), .A3(net_1008), .A1(net_1004) );
SDFF_X2 inst_150 ( .SI(net_3174), .Q(net_3174), .SE(net_2251), .D(net_1647), .CK(net_4789) );
NAND2_X2 inst_1611 ( .A1(net_2967), .ZN(net_2405), .A2(net_462) );
CLKBUF_X2 inst_4469 ( .A(net_4454), .Z(net_4455) );
CLKBUF_X2 inst_4540 ( .A(net_4525), .Z(net_4526) );
NOR3_X2 inst_887 ( .A2(net_4066), .ZN(net_2610), .A1(net_2524), .A3(net_2522) );
CLKBUF_X2 inst_4808 ( .A(net_4793), .Z(net_4794) );
CLKBUF_X2 inst_4657 ( .A(net_4286), .Z(net_4643) );
INV_X2 inst_2981 ( .ZN(net_920), .A(net_43) );
NAND2_X2 inst_1669 ( .A1(net_3815), .ZN(net_2089), .A2(net_735) );
CLKBUF_X2 inst_4998 ( .A(net_4983), .Z(net_4984) );
CLKBUF_X2 inst_5175 ( .A(net_5160), .Z(net_5161) );
NAND2_X2 inst_1663 ( .ZN(net_2100), .A1(net_2099), .A2(net_474) );
CLKBUF_X2 inst_4406 ( .A(net_4391), .Z(net_4392) );
INV_X2 inst_2714 ( .A(net_1698), .ZN(net_1591) );
DFF_X2 inst_3162 ( .D(net_2159), .QN(net_60), .CK(net_4204) );
AOI21_X2 inst_3956 ( .B2(net_3497), .A(net_3492), .B1(net_1691), .ZN(net_1685) );
XNOR2_X2 inst_90 ( .ZN(net_917), .B(net_712), .A(net_698) );
CLKBUF_X2 inst_4316 ( .A(net_4301), .Z(net_4302) );
INV_X4 inst_2357 ( .ZN(net_854), .A(net_438) );
CLKBUF_X2 inst_4650 ( .A(net_4635), .Z(net_4636) );
NAND2_X2 inst_1801 ( .A2(net_4025), .A1(net_3430), .ZN(net_962) );
CLKBUF_X2 inst_5093 ( .A(net_5078), .Z(net_5079) );
AOI221_X2 inst_3833 ( .ZN(net_2312), .A(net_2311), .C1(net_2196), .C2(net_1908), .B2(net_749), .B1(net_97) );
OAI21_X2 inst_720 ( .ZN(net_815), .B2(net_712), .B1(net_697), .A(net_610) );
NOR2_X4 inst_958 ( .A2(net_3978), .ZN(net_3722), .A1(net_3548) );
NAND2_X2 inst_1961 ( .ZN(net_3306), .A1(net_1601), .A2(net_64) );
INV_X4 inst_2460 ( .A(net_3087), .ZN(net_462) );
NAND4_X2 inst_1217 ( .A4(net_1200), .ZN(net_1170), .A2(net_1041), .A1(net_936), .A3(net_827) );
OAI221_X2 inst_368 ( .C1(net_3352), .B2(net_3348), .ZN(net_2727), .B1(net_2618), .A(net_2595), .C2(net_2122) );
NOR2_X2 inst_1010 ( .ZN(net_2017), .A1(net_1746), .A2(net_1096) );
NAND2_X2 inst_1697 ( .ZN(net_2190), .A2(net_1927), .A1(net_1851) );
NOR4_X2 inst_867 ( .ZN(net_1076), .A1(net_1072), .A2(net_1029), .A3(net_1028), .A4(net_1018) );
INV_X2 inst_3027 ( .ZN(net_3496), .A(net_3493) );
OAI211_X2 inst_820 ( .ZN(net_1567), .A(net_1515), .B(net_1366), .C1(net_1365), .C2(net_1011) );
AOI22_X2 inst_3689 ( .B2(net_4123), .A2(net_509), .ZN(net_489), .A1(net_488), .B1(net_487) );
AOI22_X2 inst_3556 ( .A1(net_4060), .B1(net_4055), .ZN(net_1494), .B2(net_208), .A2(net_150) );
SDFF_X2 inst_157 ( .SI(net_4025), .Q(net_4025), .D(net_3320), .SE(net_2514), .CK(net_4971) );
NAND2_X4 inst_1441 ( .A1(net_3974), .A2(net_3919), .ZN(net_3764) );
INV_X2 inst_2929 ( .A(net_3005), .ZN(net_174) );
AOI22_X2 inst_3568 ( .A1(net_4060), .B1(net_4055), .ZN(net_1482), .B2(net_738), .A2(net_737) );
XNOR2_X2 inst_68 ( .A(net_1657), .ZN(net_1649), .B(net_1075) );
CLKBUF_X2 inst_4287 ( .A(net_4246), .Z(net_4273) );
NAND2_X2 inst_1966 ( .ZN(net_3328), .A2(net_3319), .A1(net_430) );
AOI221_X2 inst_3914 ( .A(net_4090), .C2(net_4004), .B2(net_3680), .ZN(net_3326), .B1(net_924), .C1(net_923) );
NAND4_X2 inst_1253 ( .ZN(net_3855), .A4(net_3646), .A3(net_3336), .A2(net_3335), .A1(net_3334) );
CLKBUF_X2 inst_4716 ( .A(net_4701), .Z(net_4702) );
INV_X4 inst_2177 ( .ZN(net_2836), .A(net_2743) );
INV_X2 inst_2793 ( .ZN(net_773), .A(net_723) );
NAND2_X2 inst_1884 ( .A1(net_590), .ZN(net_525), .A2(net_398) );
NAND2_X2 inst_2018 ( .ZN(net_3650), .A1(net_3647), .A2(net_487) );
INV_X4 inst_2435 ( .ZN(net_635), .A(net_124) );
AND2_X4 inst_4158 ( .ZN(net_4109), .A1(net_3929), .A2(net_530) );
NAND2_X2 inst_1643 ( .ZN(net_2172), .A1(net_2097), .A2(net_2023) );
CLKBUF_X2 inst_4660 ( .A(net_4568), .Z(net_4646) );
DFF_X1 inst_3410 ( .Q(net_4030), .D(net_1391), .CK(net_4496) );
NAND2_X2 inst_1690 ( .A1(net_1982), .ZN(net_1980), .A2(net_222) );
INV_X2 inst_2678 ( .ZN(net_2666), .A(net_2553) );
INV_X8 inst_2120 ( .ZN(net_721), .A(net_641) );
NAND2_X2 inst_1678 ( .ZN(net_2302), .A1(net_2114), .A2(net_369) );
CLKBUF_X2 inst_5312 ( .A(net_5297), .Z(net_5298) );
INV_X4 inst_2613 ( .ZN(net_3828), .A(net_3827) );
XOR2_X2 inst_17 ( .A(net_505), .Z(net_336), .B(net_260) );
OR2_X2 inst_249 ( .ZN(net_2565), .A1(net_2528), .A2(net_641) );
NAND3_X2 inst_1287 ( .ZN(net_2260), .A1(net_2201), .A3(net_1956), .A2(net_1919) );
INV_X4 inst_2233 ( .A(net_1866), .ZN(net_1800) );
CLKBUF_X2 inst_4231 ( .A(net_4216), .Z(net_4217) );
AOI221_X2 inst_3866 ( .B1(net_2020), .C1(net_2019), .ZN(net_1942), .A(net_1941), .B2(net_83), .C2(x350) );
INV_X4 inst_2234 ( .A(net_3784), .ZN(net_1861) );
CLKBUF_X2 inst_5253 ( .A(net_4445), .Z(net_5239) );
CLKBUF_X2 inst_5204 ( .A(net_5189), .Z(net_5190) );
CLKBUF_X2 inst_4371 ( .A(net_4356), .Z(net_4357) );
CLKBUF_X2 inst_4266 ( .A(net_4237), .Z(net_4252) );
NOR2_X1 inst_1169 ( .A2(net_3939), .A1(net_3756), .ZN(net_3396) );
NAND2_X2 inst_1649 ( .ZN(net_2156), .A2(net_2155), .A1(net_2018) );
AOI22_X2 inst_3483 ( .A1(net_4038), .B1(net_2657), .ZN(net_2654), .A2(net_984), .B2(net_402) );
NAND2_X4 inst_1480 ( .ZN(net_3948), .A2(net_3720), .A1(net_3674) );
OAI221_X2 inst_396 ( .C2(net_3407), .B1(net_2328), .ZN(net_2308), .B2(net_2307), .C1(net_2242), .A(net_2015) );
DFF_X1 inst_3382 ( .QN(net_3172), .D(net_2005), .CK(net_4856) );
DFF_X1 inst_3377 ( .D(net_2254), .Q(net_75), .CK(net_5256) );
INV_X2 inst_2877 ( .A(net_3124), .ZN(net_371) );
OAI21_X2 inst_669 ( .A(net_1884), .ZN(net_1698), .B1(net_1339), .B2(net_1173) );
CLKBUF_X2 inst_5128 ( .A(net_4216), .Z(net_5114) );
OAI21_X2 inst_664 ( .A(net_4053), .ZN(net_1682), .B2(net_1636), .B1(net_1634) );
NAND2_X2 inst_1918 ( .A2(net_3160), .ZN(net_286), .A1(net_220) );
INV_X2 inst_2845 ( .ZN(net_384), .A(net_352) );
NAND2_X4 inst_1418 ( .ZN(net_3539), .A2(net_3538), .A1(net_2106) );
NAND2_X2 inst_1740 ( .ZN(net_1615), .A1(net_1502), .A2(net_917) );
INV_X2 inst_2977 ( .ZN(net_768), .A(net_83) );
NOR2_X2 inst_1092 ( .ZN(net_340), .A1(net_339), .A2(net_297) );
AND3_X4 inst_4064 ( .A3(net_3802), .ZN(net_2203), .A1(net_1790), .A2(net_1703) );
CLKBUF_X2 inst_4427 ( .A(net_4412), .Z(net_4413) );
CLKBUF_X2 inst_4836 ( .A(net_4821), .Z(net_4822) );
NAND2_X2 inst_2001 ( .ZN(net_3500), .A1(net_1135), .A2(net_403) );
CLKBUF_X2 inst_4897 ( .A(net_4610), .Z(net_4883) );
CLKBUF_X2 inst_4635 ( .A(net_4545), .Z(net_4621) );
NAND2_X2 inst_1657 ( .A1(net_3201), .ZN(net_2111), .A2(net_1980) );
AOI221_X2 inst_3839 ( .ZN(net_2205), .B2(net_2203), .C1(net_2202), .A(net_2071), .B1(net_2067), .C2(net_379) );
NAND2_X2 inst_1844 ( .ZN(net_777), .A2(net_722), .A1(net_641) );
CLKBUF_X2 inst_5209 ( .A(net_4786), .Z(net_5195) );
NAND2_X2 inst_1913 ( .A2(net_347), .ZN(net_291), .A1(net_290) );
NAND2_X2 inst_2077 ( .ZN(net_4171), .A2(net_4170), .A1(net_2703) );
INV_X4 inst_2368 ( .A(net_3214), .ZN(net_659) );
NAND2_X2 inst_1990 ( .ZN(net_3444), .A2(net_3443), .A1(net_3442) );
INV_X2 inst_2735 ( .ZN(net_1337), .A(net_1336) );
XOR2_X1 inst_36 ( .Z(net_3546), .B(net_3545), .A(net_3196) );
INV_X2 inst_2934 ( .ZN(net_178), .A(net_120) );
INV_X2 inst_2767 ( .A(net_1029), .ZN(net_927) );
NAND3_X2 inst_1370 ( .ZN(net_3991), .A1(net_3986), .A2(net_3913), .A3(net_3912) );
CLKBUF_X2 inst_4592 ( .A(net_4449), .Z(net_4578) );
INV_X4 inst_2512 ( .A(net_3075), .ZN(net_559) );
OAI21_X4 inst_451 ( .B2(net_3599), .ZN(net_2891), .B1(net_2890), .A(net_2313) );
INV_X8 inst_2166 ( .ZN(net_3959), .A(net_3819) );
OAI211_X2 inst_797 ( .ZN(net_2250), .C1(net_2249), .A(net_1338), .B(net_593), .C2(net_445) );
NAND2_X2 inst_1495 ( .A2(net_3151), .ZN(net_2823), .A1(net_2822) );
CLKBUF_X2 inst_5051 ( .A(net_5036), .Z(net_5037) );
AND2_X4 inst_4124 ( .ZN(net_4049), .A1(net_1643), .A2(net_1642) );
INV_X16 inst_3067 ( .ZN(net_3483), .A(net_3482) );
INV_X2 inst_3032 ( .A(net_3978), .ZN(net_3559) );
CLKBUF_X2 inst_5295 ( .A(net_5280), .Z(net_5281) );
AOI22_X2 inst_3657 ( .ZN(net_595), .B1(net_555), .A1(net_457), .B2(net_213), .A2(net_172) );
NAND2_X2 inst_1998 ( .ZN(net_3493), .A2(net_3492), .A1(net_1691) );
CLKBUF_X2 inst_5307 ( .A(net_5292), .Z(net_5293) );
DFF_X1 inst_3302 ( .D(net_2875), .Q(net_71), .CK(net_4276) );
INV_X2 inst_2870 ( .A(net_3388), .ZN(net_299) );
OAI21_X2 inst_676 ( .B2(net_3964), .ZN(net_1459), .B1(net_1215), .A(net_671) );
AOI22_X2 inst_3583 ( .A1(net_4063), .B1(net_4058), .ZN(net_1434), .B2(net_217), .A2(net_153) );
DFF_X1 inst_3348 ( .D(net_2706), .Q(net_69), .CK(net_4269) );
CLKBUF_X2 inst_4933 ( .A(net_4918), .Z(net_4919) );
NOR2_X2 inst_1115 ( .ZN(net_3381), .A1(net_3380), .A2(net_588) );
CLKBUF_X2 inst_4848 ( .A(net_4833), .Z(net_4834) );
CLKBUF_X2 inst_4222 ( .A(x1012), .Z(net_4208) );
NOR4_X2 inst_874 ( .ZN(net_4152), .A3(net_3985), .A4(net_3275), .A2(net_919), .A1(net_648) );
INV_X2 inst_2976 ( .ZN(net_1797), .A(net_332) );
NOR2_X2 inst_1021 ( .ZN(net_1856), .A1(net_1815), .A2(net_1652) );
NAND2_X2 inst_1681 ( .A1(net_3281), .ZN(net_2026), .A2(net_140) );
CLKBUF_X2 inst_4859 ( .A(net_4844), .Z(net_4845) );
CLKBUF_X2 inst_4820 ( .A(net_4253), .Z(net_4806) );
NAND2_X2 inst_1684 ( .A1(net_3219), .ZN(net_1988), .A2(net_171) );
AND2_X2 inst_4204 ( .A1(net_3878), .A2(net_3858), .ZN(net_3330) );
NAND2_X4 inst_1386 ( .ZN(net_2874), .A1(net_2839), .A2(net_2824) );
CLKBUF_X2 inst_4560 ( .A(net_4545), .Z(net_4546) );
INV_X4 inst_2255 ( .ZN(net_1388), .A(net_1290) );
NAND2_X2 inst_1652 ( .ZN(net_2209), .A1(net_2029), .A2(net_1977) );
CLKBUF_X2 inst_4827 ( .A(net_4425), .Z(net_4813) );
OR2_X4 inst_217 ( .A2(net_4034), .ZN(net_1165), .A1(net_356) );
NOR2_X2 inst_1076 ( .ZN(net_702), .A2(net_614), .A1(net_613) );
OAI21_X2 inst_572 ( .ZN(net_2829), .B1(net_2828), .B2(net_2815), .A(net_1580) );
NAND2_X2 inst_1622 ( .A1(net_2917), .ZN(net_2394), .A2(net_213) );
CLKBUF_X2 inst_4852 ( .A(net_4610), .Z(net_4838) );
NAND2_X2 inst_1735 ( .A1(net_1556), .ZN(net_1550), .A2(x884) );
CLKBUF_X2 inst_5036 ( .A(net_5021), .Z(net_5022) );
OR2_X2 inst_257 ( .A2(net_3438), .ZN(net_996), .A1(net_844) );
CLKBUF_X2 inst_4616 ( .A(net_4601), .Z(net_4602) );
NAND2_X2 inst_2050 ( .ZN(net_3874), .A2(net_3873), .A1(net_3872) );
NAND2_X2 inst_2000 ( .ZN(net_3499), .A1(net_2787), .A2(net_2768) );
AOI222_X1 inst_3748 ( .C1(net_3113), .ZN(net_2237), .B1(net_2079), .A1(net_2055), .B2(net_2054), .C2(net_2053), .A2(net_282) );
CLKBUF_X2 inst_4555 ( .A(net_4540), .Z(net_4541) );
INV_X4 inst_2213 ( .ZN(net_2124), .A(net_2068) );
OAI21_X2 inst_485 ( .B1(net_3278), .ZN(net_2957), .B2(net_2925), .A(net_2421) );
NAND4_X2 inst_1195 ( .ZN(net_2059), .A3(net_1485), .A4(net_1484), .A1(net_1419), .A2(net_1418) );
OAI21_X2 inst_672 ( .ZN(net_1450), .A(net_1265), .B1(net_1152), .B2(net_1039) );
NAND2_X4 inst_1471 ( .A1(net_3992), .ZN(net_3921), .A2(net_3521) );
AOI221_X2 inst_3826 ( .B1(net_3469), .B2(net_3145), .ZN(net_2535), .C1(net_2534), .A(net_2339), .C2(net_265) );
NAND4_X2 inst_1189 ( .ZN(net_1762), .A2(net_1760), .A4(net_1609), .A1(net_1370), .A3(net_1020) );
NAND4_X2 inst_1205 ( .ZN(net_1847), .A3(net_1500), .A4(net_1497), .A1(net_1433), .A2(net_1431) );
INV_X4 inst_2360 ( .ZN(net_609), .A(net_525) );
NAND2_X2 inst_1525 ( .A1(net_2959), .ZN(net_2497), .A2(net_190) );
DFF_X1 inst_3230 ( .QN(net_3065), .D(net_2971), .CK(net_4876) );
INV_X4 inst_2248 ( .ZN(net_1383), .A(net_1382) );
CLKBUF_X2 inst_5085 ( .A(net_4926), .Z(net_5071) );
INV_X4 inst_2453 ( .A(net_3161), .ZN(net_355) );
NAND3_X2 inst_1312 ( .ZN(net_956), .A1(net_955), .A2(net_954), .A3(net_810) );
DFF_X1 inst_3281 ( .QN(net_3030), .D(net_2910), .CK(net_5176) );
OAI21_X2 inst_703 ( .A(net_1253), .ZN(net_907), .B2(net_881), .B1(net_541) );
XOR2_X1 inst_33 ( .Z(net_324), .B(net_251), .A(net_77) );
MUX2_X2 inst_2107 ( .S(net_2912), .A(net_2573), .Z(net_2570), .B(net_242) );
INV_X4 inst_2546 ( .ZN(net_3443), .A(net_2302) );
CLKBUF_X2 inst_4693 ( .A(net_4678), .Z(net_4679) );
OR2_X4 inst_232 ( .ZN(net_629), .A2(net_389), .A1(net_374) );
DFF_X1 inst_3419 ( .D(net_1360), .Q(net_31), .CK(net_4290) );
NOR2_X2 inst_1067 ( .A2(net_4103), .ZN(net_948), .A1(net_774) );
CLKBUF_X2 inst_4628 ( .A(net_4268), .Z(net_4614) );
CLKBUF_X2 inst_4787 ( .A(net_4278), .Z(net_4773) );
AOI222_X1 inst_3794 ( .B1(net_4048), .ZN(net_3750), .B2(net_3745), .C2(net_3447), .A1(net_1968), .C1(net_323), .A2(net_271) );
CLKBUF_X2 inst_4951 ( .A(net_4404), .Z(net_4937) );
NAND2_X2 inst_1824 ( .A2(net_4097), .ZN(net_901), .A1(net_690) );
AOI22_X2 inst_3716 ( .ZN(net_3479), .A2(net_1908), .A1(net_1769), .B1(net_749), .B2(net_95) );
NAND4_X2 inst_1214 ( .A2(net_4074), .A3(net_4073), .ZN(net_1149), .A1(net_1148), .A4(net_859) );
OR2_X2 inst_253 ( .ZN(net_1179), .A1(net_1178), .A2(net_605) );
NOR2_X4 inst_971 ( .ZN(net_3911), .A2(net_3910), .A1(net_3217) );
NAND2_X4 inst_1417 ( .A1(net_3804), .ZN(net_3531), .A2(net_3365) );
NAND4_X2 inst_1219 ( .ZN(net_1044), .A4(net_835), .A3(net_598), .A2(net_499), .A1(net_463) );
AOI22_X2 inst_3652 ( .B1(net_4132), .ZN(net_818), .A1(net_713), .B2(net_402), .A2(net_395) );
OAI21_X2 inst_589 ( .B2(net_2815), .ZN(net_2619), .B1(net_2618), .A(net_1572) );
CLKBUF_X2 inst_5229 ( .A(net_4690), .Z(net_5215) );
CLKBUF_X2 inst_4868 ( .A(net_4853), .Z(net_4854) );
CLKBUF_X2 inst_5043 ( .A(net_5028), .Z(net_5029) );
CLKBUF_X2 inst_4273 ( .A(net_4258), .Z(net_4259) );
CLKBUF_X2 inst_4488 ( .A(net_4206), .Z(net_4474) );
OAI21_X2 inst_602 ( .B1(net_3449), .B2(net_2669), .ZN(net_2365), .A(net_671) );
XNOR2_X2 inst_59 ( .ZN(net_2064), .A(net_2063), .B(net_1872) );
NAND2_X2 inst_1877 ( .ZN(net_447), .A1(net_401), .A2(net_396) );
INV_X4 inst_2367 ( .ZN(net_729), .A(net_429) );
SDFF_X2 inst_135 ( .D(net_3483), .SI(net_3027), .Q(net_3027), .SE(net_2915), .CK(net_5053) );
DFF_X1 inst_3335 ( .QN(net_3149), .D(net_2784), .CK(net_4486) );
DFF_X1 inst_3256 ( .QN(net_3080), .D(net_2945), .CK(net_4724) );
INV_X1 inst_3073 ( .A(net_3439), .ZN(net_1806) );
NAND2_X2 inst_1865 ( .ZN(net_903), .A2(net_775), .A1(net_723) );
XOR2_X1 inst_37 ( .Z(net_4134), .B(net_4092), .A(net_1872) );
NAND2_X2 inst_1980 ( .ZN(net_3387), .A1(net_341), .A2(net_42) );
NAND2_X2 inst_1664 ( .ZN(net_2098), .A1(net_2096), .A2(net_215) );
NAND2_X4 inst_1447 ( .ZN(net_3804), .A1(net_3803), .A2(net_3404) );
DFF_X2 inst_3117 ( .Q(net_3133), .D(net_2734), .CK(net_4593) );
INV_X2 inst_2885 ( .A(net_2999), .ZN(net_166) );
CLKBUF_X2 inst_4795 ( .A(net_4523), .Z(net_4781) );
INV_X2 inst_2632 ( .A(net_3536), .ZN(net_2620) );
INV_X4 inst_2221 ( .ZN(net_2063), .A(net_1904) );
AOI222_X1 inst_3770 ( .B1(net_4048), .C1(net_3447), .A1(net_1968), .ZN(net_1962), .A2(net_294), .C2(net_204), .B2(net_73) );
NAND2_X1 inst_2082 ( .A1(net_4154), .A2(net_3600), .ZN(net_2758) );
DFF_X1 inst_3286 ( .QN(net_3050), .D(net_2895), .CK(net_4717) );
CLKBUF_X2 inst_4225 ( .A(net_4210), .Z(net_4211) );
INV_X2 inst_2709 ( .ZN(net_2119), .A(net_2016) );
OR2_X4 inst_224 ( .A2(net_4101), .ZN(net_1131), .A1(net_656) );
CLKBUF_X2 inst_4730 ( .A(net_4715), .Z(net_4716) );
AOI22_X2 inst_3635 ( .ZN(net_1710), .B1(net_1071), .A1(net_753), .A2(net_433), .B2(net_256) );
INV_X1 inst_3075 ( .A(net_3320), .ZN(net_1564) );
CLKBUF_X2 inst_5058 ( .A(net_5043), .Z(net_5044) );
INV_X2 inst_2800 ( .ZN(net_744), .A(net_708) );
INV_X4 inst_2406 ( .ZN(net_380), .A(net_304) );
OAI21_X2 inst_766 ( .ZN(net_3961), .B1(net_3960), .A(net_3634), .B2(net_923) );
AND2_X4 inst_4141 ( .ZN(net_4077), .A1(net_702), .A2(net_606) );
DFF_X1 inst_3270 ( .QN(net_3094), .D(net_2927), .CK(net_5030) );
NAND2_X2 inst_1908 ( .A1(net_323), .A2(net_322), .ZN(net_307) );
DFF_X1 inst_3273 ( .QN(net_3098), .D(net_2922), .CK(net_5020) );
OAI211_X2 inst_801 ( .C1(net_2190), .ZN(net_2168), .C2(net_2167), .A(net_2014), .B(net_1999) );
CLKBUF_X2 inst_4591 ( .A(net_4576), .Z(net_4577) );
OAI21_X2 inst_692 ( .B1(net_3734), .A(net_1650), .ZN(net_1178), .B2(net_540) );
NAND2_X2 inst_1517 ( .A1(net_3582), .ZN(net_2578), .A2(net_2513) );
XNOR2_X2 inst_70 ( .B(net_1764), .ZN(net_1618), .A(net_1462) );
NOR4_X2 inst_870 ( .A3(net_4094), .A4(net_3549), .ZN(net_967), .A2(net_966), .A1(net_919) );
XOR2_X2 inst_11 ( .Z(net_1508), .B(net_1507), .A(net_1441) );
CLKBUF_X2 inst_4528 ( .A(net_4373), .Z(net_4514) );
OR3_X2 inst_188 ( .ZN(net_3724), .A3(net_3680), .A1(net_723), .A2(net_432) );
AOI222_X1 inst_3768 ( .B1(net_4048), .C1(net_3447), .A1(net_1968), .ZN(net_1964), .C2(net_1523), .A2(net_1507), .B2(net_71) );
NAND2_X2 inst_1619 ( .A1(net_2919), .ZN(net_2397), .A2(net_194) );
AND2_X2 inst_4207 ( .ZN(net_3460), .A1(net_3445), .A2(net_2563) );
DFF_X2 inst_3110 ( .QN(net_2994), .D(net_2797), .CK(net_5099) );
OAI221_X2 inst_441 ( .C1(net_3877), .B2(net_3685), .ZN(net_3535), .B1(net_2699), .C2(net_2698), .A(net_2370) );
INV_X2 inst_3011 ( .ZN(net_3376), .A(net_3375) );
INV_X4 inst_2276 ( .ZN(net_2213), .A(net_994) );
CLKBUF_X2 inst_5228 ( .A(net_5213), .Z(net_5214) );
INV_X2 inst_2848 ( .ZN(net_370), .A(net_369) );
INV_X4 inst_2301 ( .ZN(net_2167), .A(net_856) );
CLKBUF_X2 inst_4826 ( .A(net_4811), .Z(net_4812) );
OAI211_X2 inst_808 ( .ZN(net_1681), .B(net_1588), .C1(net_1501), .A(net_1177), .C2(net_1124) );
NAND2_X2 inst_1537 ( .A1(net_2907), .ZN(net_2485), .A2(net_221) );
OAI21_X2 inst_557 ( .B2(net_2912), .B1(net_2871), .ZN(net_2868), .A(net_2451) );
NAND2_X2 inst_2041 ( .ZN(net_3809), .A1(net_3294), .A2(net_2026) );
AOI221_X2 inst_3859 ( .C2(net_4147), .B1(net_3736), .C1(net_2049), .ZN(net_2045), .A(net_1812), .B2(net_1511) );
CLKBUF_X2 inst_5235 ( .A(net_4622), .Z(net_5221) );
AOI22_X2 inst_3593 ( .A1(net_4062), .B1(net_4057), .ZN(net_1424), .B2(net_487), .A2(net_475) );
NAND3_X1 inst_1383 ( .A3(net_3827), .ZN(net_3498), .A1(net_2787), .A2(net_2768) );
DFF_X1 inst_3279 ( .QN(net_3033), .D(net_2920), .CK(net_5085) );
OAI211_X2 inst_823 ( .A(net_3843), .ZN(net_1520), .C1(net_1369), .B(net_1195), .C2(net_1150) );
NAND2_X4 inst_1461 ( .ZN(net_3872), .A1(net_3198), .A2(net_159) );
CLKBUF_X2 inst_4589 ( .A(net_4574), .Z(net_4575) );
INV_X2 inst_2838 ( .ZN(net_605), .A(net_594) );
AOI222_X1 inst_3773 ( .A2(net_2037), .ZN(net_1898), .A1(net_1863), .B1(net_1862), .C1(net_1861), .B2(net_906), .C2(net_182) );
DFF_X1 inst_3423 ( .D(net_771), .Q(net_57), .CK(net_4695) );
DFF_X2 inst_3176 ( .D(net_1876), .Q(net_54), .CK(net_4845) );
INV_X2 inst_2833 ( .ZN(net_1351), .A(net_371) );
CLKBUF_X2 inst_4767 ( .A(net_4752), .Z(net_4753) );
NAND2_X2 inst_2042 ( .ZN(net_3830), .A2(net_1982), .A1(net_148) );
DFF_X1 inst_3325 ( .Q(net_3136), .D(net_2833), .CK(net_4649) );
AND2_X4 inst_4168 ( .A2(net_4129), .ZN(net_4122), .A1(net_255) );
OR2_X4 inst_195 ( .ZN(net_2959), .A1(net_2353), .A2(net_2352) );
CLKBUF_X2 inst_5156 ( .A(net_5141), .Z(net_5142) );
NAND2_X2 inst_1987 ( .ZN(net_3433), .A2(net_3432), .A1(net_3431) );
INV_X2 inst_2796 ( .ZN(net_2150), .A(net_753) );
NOR2_X2 inst_1150 ( .ZN(net_3947), .A1(net_3654), .A2(net_3107) );
INV_X2 inst_2729 ( .ZN(net_1399), .A(net_1355) );
NAND2_X4 inst_1413 ( .A1(net_3601), .ZN(net_3393), .A2(net_3392) );
CLKBUF_X2 inst_4914 ( .A(net_4224), .Z(net_4900) );
NAND2_X2 inst_1815 ( .A2(net_3900), .ZN(net_1261), .A1(net_853) );
AOI21_X2 inst_3993 ( .B1(net_4134), .ZN(net_3240), .A(net_3239), .B2(net_1826) );
CLKBUF_X2 inst_4780 ( .A(net_4765), .Z(net_4766) );
CLKBUF_X2 inst_5267 ( .A(net_4306), .Z(net_5253) );
CLKBUF_X2 inst_4658 ( .A(net_4643), .Z(net_4644) );
NAND2_X2 inst_1589 ( .A1(net_2972), .ZN(net_2429), .A2(net_738) );
CLKBUF_X2 inst_4535 ( .A(net_4520), .Z(net_4521) );
INV_X8 inst_2169 ( .ZN(net_3995), .A(net_3107) );
NAND3_X2 inst_1326 ( .A3(net_721), .ZN(net_683), .A1(net_609), .A2(net_435) );
CLKBUF_X2 inst_4499 ( .A(net_4484), .Z(net_4485) );
CLKBUF_X2 inst_4238 ( .A(net_4223), .Z(net_4224) );
CLKBUF_X2 inst_5275 ( .A(net_5260), .Z(net_5261) );
CLKBUF_X2 inst_4758 ( .A(net_4743), .Z(net_4744) );
OAI22_X2 inst_335 ( .ZN(net_663), .A1(net_344), .B2(net_263), .A2(net_192), .B1(net_49) );
AOI221_X2 inst_3875 ( .A(net_4046), .C2(net_1908), .ZN(net_1907), .C1(net_1906), .B2(net_749), .B1(net_91) );
INV_X2 inst_2629 ( .ZN(net_2842), .A(net_2832) );
OAI21_X2 inst_658 ( .ZN(net_1763), .B1(net_1701), .A(net_1669), .B2(net_77) );
CLKBUF_X2 inst_4520 ( .A(net_4505), .Z(net_4506) );
OAI221_X2 inst_438 ( .C2(net_987), .A(net_629), .B2(net_628), .C1(net_627), .ZN(net_621), .B1(net_387) );
NAND3_X2 inst_1341 ( .A2(net_4139), .ZN(net_3383), .A3(net_3374), .A1(net_818) );
INV_X8 inst_2154 ( .ZN(net_3492), .A(net_3491) );
OAI21_X2 inst_587 ( .B2(net_2815), .ZN(net_2646), .B1(net_2645), .A(net_1744) );
OAI21_X2 inst_666 ( .B1(net_4034), .ZN(net_2016), .A(net_1646), .B2(net_1173) );
CLKBUF_X2 inst_4602 ( .A(net_4587), .Z(net_4588) );
INV_X4 inst_2602 ( .ZN(net_3613), .A(net_3171) );
OAI22_X2 inst_324 ( .B2(net_3123), .ZN(net_1137), .B1(net_721), .A1(net_641), .A2(net_43) );
NAND2_X2 inst_1829 ( .ZN(net_1614), .A1(net_1613), .A2(net_270) );
AOI22_X2 inst_3550 ( .A1(net_4059), .B1(net_4056), .ZN(net_1500), .A2(net_242), .B2(net_147) );
XNOR2_X2 inst_109 ( .ZN(net_419), .A(net_349), .B(net_108) );
NAND4_X2 inst_1182 ( .A3(net_3193), .ZN(net_2245), .A1(net_2128), .A4(net_2102), .A2(net_2092) );
AND3_X2 inst_4083 ( .ZN(net_1590), .A1(net_1589), .A2(net_1588), .A3(net_1009) );
AOI21_X2 inst_3983 ( .B1(net_983), .ZN(net_942), .A(net_638), .B2(net_371) );
XNOR2_X2 inst_43 ( .B(net_3537), .ZN(net_2743), .A(net_2540) );
INV_X8 inst_2128 ( .ZN(net_571), .A(net_362) );
NAND2_X2 inst_1707 ( .A1(net_3321), .A2(net_3320), .ZN(net_1790) );
NAND2_X4 inst_1444 ( .ZN(net_3784), .A2(net_3783), .A1(net_3782) );
CLKBUF_X2 inst_5252 ( .A(net_5233), .Z(net_5238) );
NAND4_X2 inst_1231 ( .ZN(net_753), .A4(net_573), .A3(net_563), .A2(net_502), .A1(net_456) );
OAI221_X2 inst_375 ( .B2(net_2733), .C1(net_2686), .ZN(net_2681), .A(net_2558), .C2(net_2150), .B1(net_1996) );
AOI22_X2 inst_3490 ( .B2(net_3882), .A1(net_3881), .A2(net_3516), .ZN(net_2576), .B1(net_2381) );
NOR3_X2 inst_904 ( .ZN(net_827), .A1(net_826), .A2(net_825), .A3(net_605) );
DFF_X1 inst_3315 ( .QN(net_3150), .D(net_2842), .CK(net_4517) );
INV_X8 inst_2159 ( .ZN(net_3644), .A(net_3168) );
OAI22_X2 inst_285 ( .ZN(net_2310), .B1(net_2309), .A1(net_2274), .B2(net_975), .A2(net_974) );
NAND2_X2 inst_1830 ( .A1(net_3398), .ZN(net_969), .A2(net_810) );
AOI21_X4 inst_3923 ( .B2(net_3515), .ZN(net_2607), .B1(net_2364), .A(net_2322) );
CLKBUF_X2 inst_4831 ( .A(net_4816), .Z(net_4817) );
OAI21_X2 inst_757 ( .B2(net_4146), .B1(net_4099), .A(net_4084), .ZN(net_3731) );
OAI22_X2 inst_343 ( .ZN(net_3494), .B1(net_2122), .B2(net_1071), .A1(net_1036), .A2(net_137) );
NAND2_X2 inst_1627 ( .ZN(net_2519), .A2(net_2518), .A1(net_2389) );
CLKBUF_X2 inst_4739 ( .A(net_4211), .Z(net_4725) );
NAND2_X2 inst_1563 ( .A1(net_2963), .ZN(net_2458), .A2(net_518) );
OAI21_X2 inst_543 ( .B2(net_2925), .ZN(net_2889), .B1(net_2887), .A(net_2424) );
NOR2_X2 inst_1106 ( .A1(net_3876), .A2(net_3515), .ZN(net_3222) );
CLKBUF_X2 inst_4455 ( .A(net_4440), .Z(net_4441) );
DFF_X1 inst_3242 ( .QN(net_3044), .D(net_2947), .CK(net_5180) );
AOI221_X2 inst_3817 ( .B2(net_3136), .A(net_2642), .B1(net_2591), .C2(net_2589), .ZN(net_2564), .C1(net_2563) );
DFF_X2 inst_3138 ( .QN(net_2986), .D(net_2567), .CK(net_5152) );
NOR2_X4 inst_982 ( .ZN(net_4002), .A2(net_4000), .A1(net_3658) );
NOR2_X4 inst_929 ( .A1(net_3814), .A2(net_2989), .ZN(net_2094) );
NAND2_X2 inst_2070 ( .ZN(net_3978), .A2(net_3822), .A1(net_3721) );
NAND2_X4 inst_1397 ( .A2(net_3125), .ZN(net_1259), .A1(net_1017) );
CLKBUF_X2 inst_5065 ( .A(net_5050), .Z(net_5051) );
NAND4_X2 inst_1256 ( .ZN(net_3882), .A3(net_3210), .A2(net_3209), .A4(net_3205), .A1(net_2177) );
INV_X2 inst_2890 ( .A(net_3015), .ZN(net_203) );
OAI22_X2 inst_299 ( .B1(net_2374), .ZN(net_2293), .B2(net_1606), .A1(net_1565), .A2(net_946) );
NAND2_X2 inst_1798 ( .A2(net_3156), .ZN(net_1650), .A1(net_837) );
INV_X2 inst_2927 ( .A(net_3027), .ZN(net_133) );
DFF_X1 inst_3303 ( .QN(net_3021), .D(net_2873), .CK(net_5214) );
NAND2_X2 inst_1903 ( .A1(net_3613), .A2(net_3106), .ZN(net_346) );
CLKBUF_X2 inst_4304 ( .A(net_4289), .Z(net_4290) );
INV_X2 inst_2760 ( .A(net_1228), .ZN(net_1089) );
NAND2_X2 inst_1938 ( .A2(net_3769), .ZN(net_3215), .A1(net_590) );
INV_X4 inst_2554 ( .A(net_3976), .ZN(net_3478) );
INV_X2 inst_2745 ( .A(net_1259), .ZN(net_1193) );
NAND2_X1 inst_2095 ( .ZN(net_3368), .A2(net_3366), .A1(net_2608) );
INV_X4 inst_2604 ( .ZN(net_3779), .A(net_3778) );
CLKBUF_X2 inst_5129 ( .A(net_5114), .Z(net_5115) );
CLKBUF_X2 inst_4410 ( .A(net_4234), .Z(net_4396) );
NAND4_X2 inst_1244 ( .A2(net_3652), .ZN(net_3511), .A3(net_3194), .A4(net_2136), .A1(net_2133) );
CLKBUF_X2 inst_4995 ( .A(net_4796), .Z(net_4981) );
DFF_X1 inst_3260 ( .QN(net_3076), .D(net_2930), .CK(net_4925) );
DFF_X1 inst_3248 ( .QN(net_3084), .D(net_2941), .CK(net_4547) );
AND2_X4 inst_4190 ( .ZN(net_4189), .A1(net_4042), .A2(net_2129) );
DFF_X2 inst_3158 ( .QN(net_3129), .D(net_2156), .CK(net_5287) );
OAI21_X2 inst_582 ( .B2(net_4069), .B1(net_3230), .ZN(net_2786), .A(net_2785) );
OAI21_X2 inst_683 ( .ZN(net_1265), .B2(net_1183), .B1(net_1073), .A(net_1011) );
DFF_X1 inst_3269 ( .QN(net_3095), .D(net_2911), .CK(net_5033) );
INV_X4 inst_2186 ( .ZN(net_2657), .A(net_2545) );
NAND2_X2 inst_1944 ( .A1(net_3476), .ZN(net_3244), .A2(net_2309) );
OR2_X4 inst_210 ( .A2(net_3959), .A1(net_1891), .ZN(net_1880) );
CLKBUF_X2 inst_4515 ( .A(net_4236), .Z(net_4501) );
HA_X1 inst_3101 ( .CO(net_349), .S(net_308), .A(net_209), .B(net_149) );
MUX2_X2 inst_2110 ( .B(net_3455), .S(net_3207), .A(net_2573), .Z(net_2567) );
NAND2_X2 inst_1850 ( .A1(net_4114), .ZN(net_750), .A2(net_594) );
CLKBUF_X2 inst_4942 ( .A(net_4927), .Z(net_4928) );
AOI22_X2 inst_3477 ( .B1(net_4039), .ZN(net_2673), .A1(net_2657), .A2(net_333), .B2(x23) );
NAND2_X2 inst_1950 ( .A1(net_3600), .ZN(net_3272), .A2(net_3271) );
AOI221_X2 inst_3881 ( .C2(net_1908), .ZN(net_1825), .A(net_1824), .C1(net_1823), .B2(net_749), .B1(net_92) );
CLKBUF_X2 inst_4778 ( .A(net_4763), .Z(net_4764) );
CLKBUF_X2 inst_5287 ( .A(net_5067), .Z(net_5273) );
NAND3_X2 inst_1294 ( .A1(net_4044), .ZN(net_1961), .A3(net_1960), .A2(net_1189) );
NAND2_X2 inst_1712 ( .A1(net_1884), .ZN(net_1758), .A2(net_1585) );
CLKBUF_X2 inst_5238 ( .A(net_4359), .Z(net_5224) );
NAND2_X2 inst_2057 ( .A1(net_3915), .ZN(net_3905), .A2(net_3900) );
CLKBUF_X2 inst_4576 ( .A(net_4561), .Z(net_4562) );
DFF_X2 inst_3108 ( .QN(net_2996), .D(net_2798), .CK(net_5106) );
OAI21_X2 inst_747 ( .B2(net_4138), .ZN(net_3378), .B1(net_3377), .A(net_3376) );
OAI211_X2 inst_843 ( .B(net_3323), .ZN(net_1113), .A(net_980), .C1(net_889), .C2(net_723) );
AOI221_X2 inst_3806 ( .C2(net_4032), .ZN(net_2736), .B2(net_2612), .C1(net_2562), .A(net_2365), .B1(net_2130) );
INV_X2 inst_2853 ( .A(net_3447), .ZN(net_356) );
NAND2_X2 inst_1779 ( .A2(net_4024), .ZN(net_1191), .A1(net_1068) );
CLKBUF_X2 inst_4486 ( .A(net_4235), .Z(net_4472) );
INV_X8 inst_2115 ( .ZN(net_2970), .A(net_2903) );
CLKBUF_X2 inst_5146 ( .A(net_4368), .Z(net_5132) );
DFF_X1 inst_3251 ( .QN(net_3089), .D(net_2952), .CK(net_4734) );
XNOR2_X2 inst_112 ( .ZN(net_410), .B(net_354), .A(net_336) );
NAND2_X2 inst_1728 ( .ZN(net_1558), .A1(net_1556), .A2(x856) );
INV_X2 inst_2775 ( .A(net_996), .ZN(net_836) );
NOR3_X2 inst_916 ( .A1(net_3903), .A2(net_3890), .ZN(net_3712), .A3(net_749) );
NAND2_X2 inst_1722 ( .ZN(net_1604), .A1(net_1515), .A2(net_1344) );
OAI22_X2 inst_305 ( .A2(net_3149), .A1(net_1543), .B1(net_1542), .ZN(net_1536), .B2(net_1535) );
NAND2_X2 inst_1595 ( .A1(net_2925), .ZN(net_2423), .A2(net_199) );
AOI22_X2 inst_3665 ( .B2(net_3402), .A2(net_3401), .A1(net_571), .B1(net_570), .ZN(net_562) );
INV_X2 inst_2724 ( .ZN(net_1467), .A(net_1397) );
INV_X4 inst_2525 ( .A(net_3895), .ZN(net_3261) );
INV_X2 inst_2968 ( .ZN(net_300), .A(net_60) );
INV_X2 inst_2964 ( .ZN(net_152), .A(net_88) );
AOI22_X2 inst_3721 ( .ZN(net_3609), .A1(net_3185), .B1(net_1982), .A2(net_519), .B2(net_478) );
INV_X4 inst_2349 ( .ZN(net_2625), .A(x475) );
OAI21_X2 inst_646 ( .A(net_3256), .ZN(net_1945), .B1(net_1643), .B2(net_1642) );
CLKBUF_X2 inst_5076 ( .A(net_4207), .Z(net_5062) );
AOI211_X2 inst_4032 ( .A(net_4068), .ZN(net_3317), .B(net_1147), .C1(net_1116), .C2(net_407) );
DFF_X2 inst_3169 ( .D(net_1926), .QN(net_89), .CK(net_5093) );
NOR2_X4 inst_963 ( .ZN(net_3810), .A1(net_3809), .A2(net_3539) );
OAI221_X2 inst_382 ( .B1(net_3581), .C2(net_2699), .B2(net_2698), .ZN(net_2631), .C1(net_2630), .A(net_2533) );
INV_X4 inst_2329 ( .A(net_3661), .ZN(net_748) );
NOR3_X2 inst_907 ( .A2(net_3954), .ZN(net_656), .A3(net_641), .A1(net_637) );
NOR2_X4 inst_922 ( .ZN(net_2788), .A1(net_2741), .A2(net_2576) );
NAND2_X2 inst_1614 ( .A1(net_2919), .ZN(net_2402), .A2(net_181) );
NAND2_X2 inst_1502 ( .ZN(net_2807), .A1(net_2782), .A2(net_2723) );
INV_X2 inst_2788 ( .ZN(net_797), .A(net_796) );
AND3_X2 inst_4091 ( .A1(net_4162), .A2(net_4126), .ZN(net_3732), .A3(net_3628) );
NOR2_X2 inst_1049 ( .A1(net_4075), .A2(net_1052), .ZN(net_1051) );
AOI221_X2 inst_3907 ( .B1(net_4109), .ZN(net_992), .B2(net_991), .C1(net_990), .A(net_832), .C2(net_361) );
OR3_X4 inst_168 ( .ZN(net_1543), .A1(net_1521), .A2(net_1334), .A3(net_1071) );
CLKBUF_X2 inst_5116 ( .A(net_5101), .Z(net_5102) );
NAND2_X2 inst_1568 ( .A1(net_2912), .ZN(net_2453), .A2(net_236) );
CLKBUF_X2 inst_4575 ( .A(net_4560), .Z(net_4561) );
AOI22_X2 inst_3692 ( .B2(net_4123), .B1(net_4023), .A1(net_4017), .A2(net_509), .ZN(net_484) );
DFF_X1 inst_3366 ( .D(net_3696), .CK(net_4251), .Q(x160) );
NOR4_X2 inst_873 ( .ZN(net_3551), .A1(net_2145), .A2(net_1947), .A3(net_1801), .A4(net_1750) );
NOR2_X2 inst_991 ( .A1(net_3880), .A2(net_3859), .ZN(net_2380) );
OAI21_X2 inst_653 ( .ZN(net_1831), .A(net_1773), .B2(net_347), .B1(x475) );
AOI222_X1 inst_3767 ( .B1(net_4048), .A1(net_1968), .ZN(net_1965), .A2(net_1439), .C2(net_991), .C1(net_375), .B2(net_239) );
OAI21_X2 inst_580 ( .B2(net_2907), .B1(net_2803), .ZN(net_2798), .A(net_2487) );
OR3_X4 inst_170 ( .A3(net_4094), .A2(net_4085), .ZN(net_1072), .A1(net_1058) );
NAND2_X2 inst_1746 ( .A2(net_4005), .ZN(net_1583), .A1(net_1282) );
AOI22_X2 inst_3691 ( .B1(net_4123), .ZN(net_485), .A1(net_458), .B2(net_233), .A2(net_183) );
CLKBUF_X2 inst_4431 ( .A(net_4416), .Z(net_4417) );
DFF_X1 inst_3371 ( .D(net_2294), .CK(net_4217), .Q(x307) );
INV_X2 inst_3052 ( .ZN(net_3851), .A(net_2245) );
AOI22_X2 inst_3649 ( .ZN(net_739), .A1(net_738), .B1(net_737), .A2(net_458), .B2(net_457) );
NAND2_X2 inst_1857 ( .A2(net_3153), .ZN(net_612), .A1(net_433) );
CLKBUF_X2 inst_4609 ( .A(net_4594), .Z(net_4595) );
INV_X2 inst_2907 ( .A(net_3139), .ZN(net_287) );
AND3_X4 inst_4072 ( .A1(net_4043), .ZN(net_4040), .A2(net_2181), .A3(net_2180) );
INV_X2 inst_2656 ( .A(net_2698), .ZN(net_2240) );
INV_X2 inst_3000 ( .A(net_3024), .ZN(net_126) );
NOR2_X2 inst_1163 ( .ZN(net_4170), .A2(net_4169), .A1(net_1994) );
OAI21_X4 inst_468 ( .ZN(net_3983), .A(net_3980), .B2(net_3755), .B1(net_3615) );
NOR2_X2 inst_1099 ( .A1(net_3654), .ZN(net_278), .A2(net_138) );
CLKBUF_X2 inst_4428 ( .A(net_4218), .Z(net_4414) );
AOI22_X2 inst_3616 ( .A1(net_1518), .ZN(net_1327), .B2(net_1326), .B1(net_1146), .A2(net_1001) );
CLKBUF_X2 inst_4889 ( .A(net_4874), .Z(net_4875) );
NAND2_X2 inst_1604 ( .A1(net_2969), .ZN(net_2413), .A2(net_498) );
DFF_X1 inst_3239 ( .QN(net_3039), .D(net_2937), .CK(net_5187) );
INV_X4 inst_2314 ( .ZN(net_1385), .A(net_1042) );
INV_X4 inst_2190 ( .ZN(net_2584), .A(net_2349) );
OAI221_X2 inst_429 ( .B2(net_3789), .ZN(net_1054), .A(net_1009), .B1(net_1008), .C1(net_1007), .C2(net_526) );
INV_X2 inst_2692 ( .ZN(net_1733), .A(net_1700) );
NAND2_X2 inst_1599 ( .A1(net_2969), .ZN(net_2418), .A2(net_495) );
INV_X2 inst_2812 ( .A(net_1400), .ZN(net_645) );
CLKBUF_X2 inst_5026 ( .A(net_5011), .Z(net_5012) );
AOI22_X2 inst_3565 ( .A1(net_4059), .B1(net_4056), .ZN(net_1485), .A2(net_200), .B2(net_140) );
CLKBUF_X2 inst_4743 ( .A(net_4728), .Z(net_4729) );
DFF_X2 inst_3197 ( .QN(net_3167), .D(net_1622), .CK(net_5131) );
CLKBUF_X2 inst_4651 ( .A(net_4286), .Z(net_4637) );
XOR2_X2 inst_7 ( .B(net_3492), .Z(net_1692), .A(net_1691) );
AOI21_X2 inst_3977 ( .B2(net_3559), .A(net_1196), .ZN(net_1115), .B1(net_895) );
AOI22_X2 inst_3467 ( .B2(net_3118), .ZN(net_2725), .A1(net_2724), .B1(net_2722), .A2(net_33) );
INV_X4 inst_2593 ( .ZN(net_3717), .A(net_3715) );
INV_X16 inst_3064 ( .ZN(net_1982), .A(net_1865) );
AOI22_X2 inst_3676 ( .A1(net_571), .B1(net_570), .ZN(net_545), .A2(net_237), .B2(net_157) );
CLKBUF_X2 inst_5021 ( .A(net_5006), .Z(net_5007) );
NOR2_X2 inst_1083 ( .A1(net_3614), .ZN(net_614), .A2(net_388) );
AND3_X4 inst_4073 ( .ZN(net_4048), .A3(net_3802), .A2(net_3320), .A1(net_1645) );
OAI22_X2 inst_318 ( .A2(net_4074), .B1(net_1250), .ZN(net_1121), .A1(net_1120), .B2(net_1100) );
AOI211_X2 inst_4033 ( .C1(net_4094), .B(net_4085), .ZN(net_3839), .C2(net_3834), .A(net_969) );
NOR2_X2 inst_1136 ( .A1(net_3995), .ZN(net_3757), .A2(net_3109) );
INV_X4 inst_2466 ( .A(net_2989), .ZN(net_175) );
CLKBUF_X2 inst_5044 ( .A(net_4447), .Z(net_5030) );
INV_X2 inst_2899 ( .A(net_3018), .ZN(net_157) );
AND3_X4 inst_4065 ( .A3(net_3802), .A2(net_3321), .ZN(net_1921), .A1(net_1827) );
NAND2_X4 inst_1486 ( .ZN(net_4163), .A1(net_3713), .A2(net_3628) );
INV_X4 inst_2281 ( .ZN(net_1198), .A(net_1069) );
OAI21_X2 inst_696 ( .A(net_3907), .B1(net_3905), .B2(net_3789), .ZN(net_1022) );
NAND4_X4 inst_1175 ( .A3(net_3649), .ZN(net_3251), .A4(net_3250), .A1(net_3234), .A2(net_2093) );
DFF_X1 inst_3311 ( .D(net_2863), .QN(net_66), .CK(net_4244) );
CLKBUF_X2 inst_5256 ( .A(net_4469), .Z(net_5242) );
AND2_X4 inst_4096 ( .ZN(net_2019), .A1(net_1651), .A2(net_1650) );
CLKBUF_X2 inst_5055 ( .A(net_5040), .Z(net_5041) );
CLKBUF_X2 inst_5117 ( .A(net_5102), .Z(net_5103) );
CLKBUF_X2 inst_5081 ( .A(net_4703), .Z(net_5067) );
CLKBUF_X2 inst_4509 ( .A(net_4494), .Z(net_4495) );
CLKBUF_X2 inst_5114 ( .A(net_4537), .Z(net_5100) );
CLKBUF_X2 inst_4929 ( .A(net_4743), .Z(net_4915) );
OAI221_X2 inst_395 ( .C2(net_3408), .B1(net_2361), .ZN(net_2356), .C1(net_2226), .A(net_1942), .B2(net_111) );
OAI211_X2 inst_841 ( .C2(net_4109), .ZN(net_1258), .A(net_1257), .C1(net_1256), .B(net_1065) );
AOI21_X2 inst_3963 ( .ZN(net_1456), .B1(net_1455), .B2(net_1153), .A(net_765) );
OAI21_X2 inst_689 ( .B1(net_4004), .ZN(net_1086), .A(net_641), .B2(net_384) );
AOI21_X2 inst_3969 ( .A(net_3558), .ZN(net_1313), .B1(net_1134), .B2(net_1011) );
CLKBUF_X2 inst_4453 ( .A(net_4438), .Z(net_4439) );
INV_X4 inst_2363 ( .A(net_3954), .ZN(net_446) );
INV_X2 inst_2689 ( .A(net_3844), .ZN(net_1755) );
CLKBUF_X2 inst_4895 ( .A(net_4857), .Z(net_4881) );
AOI211_X2 inst_4029 ( .B(net_3525), .C1(net_3322), .A(net_1018), .ZN(net_865), .C2(net_594) );
NAND2_X2 inst_1629 ( .ZN(net_2341), .A1(net_2288), .A2(net_2240) );
AOI221_X2 inst_3896 ( .C1(net_4030), .A(net_2525), .C2(net_1394), .B1(net_1393), .ZN(net_1346), .B2(net_218) );
NAND2_X2 inst_1558 ( .A1(net_2909), .ZN(net_2464), .A2(net_233) );
AOI22_X2 inst_3679 ( .B1(net_4124), .ZN(net_510), .A1(net_509), .B2(net_227), .A2(net_181) );
INV_X2 inst_2906 ( .A(net_3144), .ZN(net_256) );
DFF_X1 inst_3424 ( .Q(net_4009), .D(net_4008), .CK(net_4921) );
AOI221_X2 inst_3886 ( .C2(net_1656), .ZN(net_1524), .B2(net_1523), .C1(net_1522), .B1(net_1263), .A(net_1249) );
NAND2_X2 inst_1615 ( .A1(net_2919), .ZN(net_2401), .A2(net_151) );
INV_X4 inst_2580 ( .ZN(net_3623), .A(net_3622) );
AOI22_X2 inst_3713 ( .ZN(net_3247), .A1(net_3178), .B1(net_2099), .A2(net_498), .B2(net_497) );
INV_X4 inst_2394 ( .ZN(net_379), .A(net_327) );
INV_X8 inst_2145 ( .ZN(net_3228), .A(net_3227) );
OAI21_X2 inst_709 ( .B2(net_881), .ZN(net_851), .A(net_850), .B1(net_849) );
CLKBUF_X2 inst_4574 ( .A(net_4316), .Z(net_4560) );
INV_X4 inst_2375 ( .ZN(net_1463), .A(net_511) );
NOR3_X1 inst_920 ( .A1(net_3581), .A2(net_3248), .ZN(net_2343), .A3(net_2342) );
NAND2_X2 inst_2054 ( .ZN(net_3896), .A2(net_3892), .A1(net_3867) );
CLKBUF_X2 inst_5294 ( .A(net_4341), .Z(net_5280) );
CLKBUF_X2 inst_5251 ( .A(net_5236), .Z(net_5237) );
CLKBUF_X2 inst_4422 ( .A(net_4407), .Z(net_4408) );
NAND4_X2 inst_1259 ( .ZN(net_4188), .A4(net_3699), .A2(net_3617), .A3(net_3524), .A1(net_3430) );
CLKBUF_X2 inst_5092 ( .A(net_5077), .Z(net_5078) );
CLKBUF_X2 inst_4610 ( .A(net_4595), .Z(net_4596) );
NAND2_X2 inst_1796 ( .ZN(net_998), .A1(net_839), .A2(net_432) );
CLKBUF_X2 inst_4403 ( .A(net_4388), .Z(net_4389) );
OAI21_X2 inst_535 ( .B1(net_3195), .B2(net_2963), .ZN(net_2898), .A(net_2460) );
INV_X2 inst_2889 ( .A(net_3113), .ZN(net_1535) );
NAND2_X2 inst_1670 ( .A1(net_3817), .ZN(net_2088), .A2(net_738) );
INV_X4 inst_2189 ( .A(net_2686), .ZN(net_2640) );
INV_X4 inst_2427 ( .A(net_3054), .ZN(net_487) );
AND2_X2 inst_4198 ( .ZN(net_1402), .A1(net_1296), .A2(net_671) );
OAI22_X2 inst_315 ( .A1(net_4073), .A2(net_1381), .ZN(net_1127), .B1(net_1126), .B2(net_1125) );
INV_X2 inst_2935 ( .A(net_3117), .ZN(net_131) );
OR2_X4 inst_216 ( .ZN(net_1214), .A2(net_1213), .A1(net_1151) );
DFF_X1 inst_3317 ( .QN(net_3004), .D(net_2844), .CK(net_5118) );
DFF_X1 inst_3369 ( .D(net_2285), .CK(net_4437), .Q(x204) );
CLKBUF_X2 inst_5027 ( .A(net_5012), .Z(net_5013) );
DFF_X2 inst_3113 ( .QN(net_2990), .D(net_2799), .CK(net_5199) );
NAND2_X2 inst_2060 ( .ZN(net_3909), .A1(net_3817), .A2(net_162) );
AOI22_X2 inst_3695 ( .B2(net_4124), .A1(net_4021), .B1(net_4019), .A2(net_555), .ZN(net_481) );
INV_X2 inst_2680 ( .ZN(net_1859), .A(net_1858) );
DFF_X2 inst_3168 ( .Q(net_3161), .D(net_1958), .CK(net_4762) );
INV_X4 inst_2336 ( .A(net_3734), .ZN(net_661) );
INV_X4 inst_2385 ( .ZN(net_381), .A(net_276) );
OAI221_X2 inst_415 ( .ZN(net_1318), .C1(net_1250), .A(net_1199), .B2(net_1148), .B1(net_1120), .C2(net_1101) );
AOI221_X2 inst_3855 ( .B1(net_3736), .ZN(net_2050), .C1(net_2049), .A(net_1931), .C2(net_1732), .B2(net_271) );
NAND2_X2 inst_1795 ( .ZN(net_1183), .A2(net_866), .A1(net_852) );
OAI211_X2 inst_828 ( .ZN(net_1527), .B(net_1266), .A(net_1210), .C1(net_1182), .C2(net_408) );
CLKBUF_X2 inst_4697 ( .A(net_4682), .Z(net_4683) );
DFF_X1 inst_3318 ( .QN(net_3003), .D(net_2847), .CK(net_5113) );
OR2_X4 inst_223 ( .A2(net_4107), .ZN(net_1028), .A1(net_924) );
AND2_X4 inst_4164 ( .ZN(net_4118), .A1(net_3767), .A2(net_3628) );
CLKBUF_X2 inst_5278 ( .A(net_4590), .Z(net_5264) );
INV_X4 inst_2420 ( .ZN(net_281), .A(net_246) );
NAND2_X2 inst_1561 ( .A1(net_2963), .ZN(net_2460), .A2(net_241) );
CLKBUF_X2 inst_5176 ( .A(net_4727), .Z(net_5162) );
AOI22_X2 inst_3564 ( .A1(net_4060), .B1(net_4055), .ZN(net_1486), .B2(net_732), .A2(net_731) );
MUX2_X2 inst_2104 ( .S(net_2919), .Z(net_2574), .A(net_2573), .B(net_147) );
AND2_X2 inst_4205 ( .A1(net_3480), .ZN(net_3392), .A2(net_1770) );
NAND3_X2 inst_1322 ( .A3(net_3243), .ZN(net_725), .A2(net_641), .A1(net_376) );
INV_X4 inst_2573 ( .A(net_3617), .ZN(net_3567) );
NAND2_X1 inst_2096 ( .A2(net_3870), .A1(net_3868), .ZN(net_3453) );
OAI21_X2 inst_552 ( .B2(net_2876), .ZN(net_2875), .A(net_2856), .B1(net_2855) );
INV_X2 inst_3050 ( .A(net_3820), .ZN(net_3819) );
CLKBUF_X2 inst_4793 ( .A(net_4778), .Z(net_4779) );
CLKBUF_X2 inst_4997 ( .A(net_4982), .Z(net_4983) );
AOI22_X2 inst_3493 ( .ZN(net_2233), .A1(net_2231), .B1(net_2230), .B2(net_276), .A2(net_75) );
CLKBUF_X2 inst_4622 ( .A(net_4226), .Z(net_4608) );
INV_X2 inst_3019 ( .ZN(net_3423), .A(net_2613) );
INV_X4 inst_2327 ( .ZN(net_924), .A(net_660) );
AOI221_X2 inst_3913 ( .C2(net_3196), .ZN(net_636), .C1(net_635), .A(net_420), .B2(net_381), .B1(net_210) );
NAND2_X2 inst_1564 ( .A1(net_2963), .ZN(net_2457), .A2(net_470) );
CLKBUF_X2 inst_5078 ( .A(net_5063), .Z(net_5064) );
AOI22_X2 inst_3487 ( .B1(net_4039), .A1(net_4038), .ZN(net_2606), .A2(net_204), .B2(x79) );
AOI22_X2 inst_3597 ( .A1(net_4063), .B1(net_4058), .ZN(net_1420), .A2(net_244), .B2(net_139) );
NAND2_X2 inst_1941 ( .ZN(net_3236), .A1(net_3235), .A2(net_3183) );
INV_X4 inst_2607 ( .A(net_3817), .ZN(net_3814) );
XNOR2_X2 inst_113 ( .A(net_3152), .ZN(net_372), .B(net_316) );
XOR2_X2 inst_9 ( .Z(net_1644), .A(net_1643), .B(net_1642) );
OAI222_X2 inst_356 ( .ZN(net_3969), .A2(net_3968), .B2(net_3967), .C1(net_1261), .A1(net_1141), .B1(net_896), .C2(net_414) );
DFF_X1 inst_3358 ( .D(net_2356), .CK(net_4404), .Q(x350) );
INV_X2 inst_2690 ( .ZN(net_1735), .A(net_1734) );
NAND2_X2 inst_1594 ( .A1(net_2925), .ZN(net_2424), .A2(net_155) );
NOR3_X2 inst_902 ( .A2(net_4104), .A3(net_4079), .ZN(net_989), .A1(net_740) );
AOI22_X2 inst_3489 ( .B1(net_4039), .A1(net_4038), .A2(net_3418), .ZN(net_2604), .B2(x60) );
OAI211_X4 inst_778 ( .ZN(net_3867), .C2(net_3717), .C1(net_3684), .B(net_3672), .A(net_3635) );
CLKBUF_X2 inst_4286 ( .A(net_4271), .Z(net_4272) );
NAND2_X2 inst_1544 ( .A1(net_3207), .ZN(net_2478), .A2(net_176) );
NAND2_X2 inst_1935 ( .ZN(net_3202), .A1(net_3198), .A2(net_230) );
AND3_X4 inst_4063 ( .A2(net_3770), .A1(net_3439), .ZN(net_2055), .A3(net_1808) );
INV_X4 inst_2625 ( .ZN(net_4003), .A(net_4000) );
DFF_X2 inst_3148 ( .D(net_2333), .QN(net_110), .CK(net_4390) );
INV_X8 inst_2140 ( .A(net_3281), .ZN(net_3177) );
CLKBUF_X2 inst_4761 ( .A(net_4485), .Z(net_4747) );
DFF_X1 inst_3329 ( .D(net_2814), .QN(net_119), .CK(net_4457) );
OAI211_X2 inst_781 ( .C1(net_3230), .ZN(net_2806), .A(net_2767), .B(net_2754), .C2(net_2057) );
CLKBUF_X2 inst_5180 ( .A(net_5165), .Z(net_5166) );
AND4_X4 inst_4042 ( .ZN(net_3676), .A2(net_3439), .A4(net_1845), .A1(net_1844), .A3(net_1808) );
INV_X2 inst_3026 ( .ZN(net_3490), .A(net_3104) );
AOI22_X2 inst_3696 ( .B2(net_4123), .A2(net_509), .ZN(net_480), .A1(net_479), .B1(net_478) );
NAND2_X4 inst_1442 ( .ZN(net_3777), .A2(net_3776), .A1(net_3775) );
INV_X2 inst_2847 ( .ZN(net_386), .A(net_373) );
OAI22_X2 inst_332 ( .A2(net_3214), .ZN(net_703), .B2(net_605), .A1(net_541), .B1(net_534) );
AOI22_X2 inst_3639 ( .ZN(net_764), .A2(net_621), .B1(net_577), .B2(net_387), .A1(net_204) );
NAND3_X2 inst_1289 ( .ZN(net_2258), .A1(net_2197), .A3(net_1954), .A2(net_1920) );
INV_X8 inst_2132 ( .ZN(net_359), .A(net_279) );
AOI211_X2 inst_4013 ( .ZN(net_2678), .C1(net_2599), .B(net_2598), .C2(net_1785), .A(net_1687) );
CLKBUF_X2 inst_4979 ( .A(net_4964), .Z(net_4965) );
NAND2_X2 inst_1559 ( .A1(net_2909), .ZN(net_2463), .A2(net_193) );
NAND2_X2 inst_1928 ( .ZN(net_3191), .A1(net_3186), .A2(net_737) );
NAND2_X2 inst_1967 ( .ZN(net_3334), .A2(net_3185), .A1(net_471) );
CLKBUF_X2 inst_4686 ( .A(net_4671), .Z(net_4672) );
CLKBUF_X2 inst_4485 ( .A(net_4452), .Z(net_4471) );
NOR2_X4 inst_927 ( .ZN(net_2177), .A1(net_2095), .A2(net_2031) );
CLKBUF_X2 inst_4869 ( .A(net_4854), .Z(net_4855) );
OAI21_X2 inst_752 ( .ZN(net_3502), .A(net_3501), .B1(net_1599), .B2(net_530) );
DFF_X1 inst_3245 ( .QN(net_3092), .D(net_2940), .CK(net_4737) );
XNOR2_X2 inst_73 ( .ZN(net_1510), .A(net_1509), .B(net_64) );
NAND2_X2 inst_1488 ( .ZN(net_2880), .A1(net_2860), .A2(net_1850) );
NAND2_X2 inst_1719 ( .A1(net_3492), .ZN(net_1866), .A2(net_1694) );
NAND2_X2 inst_1947 ( .ZN(net_3259), .A2(net_3258), .A1(net_3257) );
DFF_X2 inst_3202 ( .D(net_1607), .Q(net_38), .CK(net_4986) );
CLKBUF_X2 inst_4279 ( .A(net_4264), .Z(net_4265) );
OAI221_X2 inst_378 ( .B1(net_2670), .C1(net_2668), .ZN(net_2664), .B2(net_2663), .A(net_1386), .C2(net_315) );
NAND2_X2 inst_1951 ( .ZN(net_3271), .A1(net_2861), .A2(net_2853) );
NAND2_X4 inst_1384 ( .ZN(net_2903), .A1(net_2894), .A2(net_2066) );
CLKBUF_X2 inst_4690 ( .A(net_4675), .Z(net_4676) );
INV_X8 inst_2118 ( .ZN(net_2099), .A(net_1973) );
NOR3_X2 inst_890 ( .A1(net_2521), .ZN(net_2348), .A2(net_544), .A3(net_506) );
INV_X4 inst_2200 ( .ZN(net_2357), .A(net_2266) );
NAND2_X2 inst_1851 ( .A2(net_4003), .ZN(net_810), .A1(net_536) );
CLKBUF_X2 inst_4585 ( .A(net_4335), .Z(net_4571) );
CLKBUF_X2 inst_4937 ( .A(net_4922), .Z(net_4923) );
CLKBUF_X2 inst_4514 ( .A(net_4499), .Z(net_4500) );
CLKBUF_X2 inst_5048 ( .A(net_4256), .Z(net_5034) );
NOR2_X1 inst_1168 ( .A1(net_826), .A2(net_416), .ZN(net_383) );
CLKBUF_X2 inst_4356 ( .A(net_4341), .Z(net_4342) );
OR2_X2 inst_250 ( .ZN(net_1686), .A1(net_1639), .A2(net_1638) );
OAI21_X2 inst_659 ( .A(net_3491), .ZN(net_2548), .B1(net_1747), .B2(net_1317) );
CLKBUF_X2 inst_4363 ( .A(net_4348), .Z(net_4349) );
NOR2_X2 inst_1161 ( .ZN(net_4114), .A1(net_436), .A2(net_400) );
DFF_X1 inst_3362 ( .D(net_2358), .CK(net_4397), .Q(x332) );
CLKBUF_X2 inst_5273 ( .A(net_5258), .Z(net_5259) );
NAND2_X2 inst_1523 ( .A1(net_2959), .ZN(net_2499), .A2(net_780) );
INV_X4 inst_2539 ( .ZN(net_3388), .A(net_3105) );
NOR2_X2 inst_1048 ( .ZN(net_1059), .A1(net_1058), .A2(net_956) );
DFF_X2 inst_3199 ( .QN(net_3170), .D(net_1623), .CK(net_5129) );
INV_X2 inst_2797 ( .A(net_2220), .ZN(net_752) );
AOI22_X2 inst_3612 ( .A1(net_4062), .B1(net_4057), .ZN(net_1405), .B2(net_196), .A2(net_191) );
DFF_X1 inst_3431 ( .Q(net_4023), .D(net_4022), .CK(net_4894) );
NAND2_X2 inst_1581 ( .A1(net_2915), .ZN(net_2439), .A2(net_219) );
INV_X4 inst_2270 ( .ZN(net_1067), .A(net_1066) );
NAND2_X1 inst_2085 ( .A2(net_4013), .A1(net_2965), .ZN(net_2447) );
INV_X4 inst_2388 ( .A(net_3756), .ZN(net_590) );
INV_X4 inst_2401 ( .A(net_3999), .ZN(net_328) );
INV_X4 inst_2312 ( .A(net_3990), .ZN(net_908) );
CLKBUF_X2 inst_4309 ( .A(net_4294), .Z(net_4295) );
AOI22_X2 inst_3500 ( .A1(net_3178), .ZN(net_2133), .B1(net_2099), .A2(net_468), .B2(net_453) );
INV_X2 inst_2634 ( .A(net_2578), .ZN(net_2541) );
CLKBUF_X2 inst_5264 ( .A(net_5249), .Z(net_5250) );
AOI22_X2 inst_3711 ( .A1(net_3815), .ZN(net_3194), .B1(net_3186), .A2(net_781), .B2(net_780) );
INV_X4 inst_2241 ( .ZN(net_2003), .A(net_1905) );
INV_X4 inst_2182 ( .ZN(net_2680), .A(net_2609) );
OAI21_X2 inst_556 ( .B2(net_2915), .B1(net_2871), .ZN(net_2869), .A(net_2437) );
OAI21_X2 inst_650 ( .ZN(net_1877), .B2(net_1821), .A(net_1759), .B1(net_1171) );
OAI22_X2 inst_289 ( .A2(net_4092), .ZN(net_1904), .A1(net_1872), .B2(net_987), .B1(net_681) );
INV_X2 inst_2667 ( .ZN(net_2704), .A(net_2590) );
AOI22_X2 inst_3632 ( .B2(net_1523), .B1(net_1117), .ZN(net_878), .A1(net_784), .A2(net_323) );
AND2_X2 inst_4194 ( .ZN(net_2218), .A1(net_2217), .A2(net_1226) );
NOR2_X2 inst_987 ( .ZN(net_2724), .A1(net_2528), .A2(net_2523) );
OAI221_X2 inst_420 ( .A(net_1257), .C1(net_1256), .ZN(net_1205), .B1(net_959), .B2(net_646), .C2(net_638) );
OAI21_X2 inst_679 ( .B1(net_3228), .ZN(net_1441), .A(net_1307), .B2(net_332) );
CLKBUF_X2 inst_5147 ( .A(net_4736), .Z(net_5133) );
INV_X2 inst_3006 ( .ZN(net_3242), .A(net_3240) );
AOI21_X2 inst_3992 ( .B2(net_3853), .B1(net_3806), .ZN(net_3223), .A(net_3222) );
DFF_X1 inst_3265 ( .QN(net_3071), .D(net_2934), .CK(net_4923) );
DFF_X1 inst_3364 ( .D(net_2331), .QN(net_64), .CK(net_4226) );
NAND3_X2 inst_1351 ( .A1(net_3836), .ZN(net_3641), .A3(net_3639), .A2(net_3547) );
XNOR2_X2 inst_44 ( .ZN(net_2816), .A(net_2636), .B(net_1707) );
CLKBUF_X2 inst_4433 ( .A(net_4415), .Z(net_4419) );
DFF_X1 inst_3300 ( .D(net_2877), .Q(net_73), .CK(net_4280) );
OAI221_X2 inst_371 ( .C2(net_4089), .B2(net_2733), .ZN(net_2687), .C1(net_2686), .A(net_2557), .B1(net_2163) );
NAND3_X2 inst_1305 ( .A3(net_4076), .A1(net_1178), .ZN(net_1175), .A2(net_1046) );
OAI22_X2 inst_314 ( .B2(net_3627), .ZN(net_1144), .A1(net_1143), .B1(net_1142), .A2(net_668) );
OAI221_X2 inst_435 ( .B1(net_920), .A(net_629), .B2(net_628), .C1(net_627), .ZN(net_624), .C2(net_43) );
DFF_X1 inst_3225 ( .QN(net_3055), .D(net_2979), .CK(net_4607) );
CLKBUF_X2 inst_4962 ( .A(net_4947), .Z(net_4948) );
AOI221_X2 inst_3822 ( .B2(net_3143), .A(net_2642), .B1(net_2591), .C1(net_2589), .ZN(net_2556), .C2(net_2555) );
OAI21_X2 inst_597 ( .B2(net_3978), .ZN(net_2546), .A(net_2345), .B1(net_1253) );
CLKBUF_X2 inst_4593 ( .A(net_4578), .Z(net_4579) );
DFF_X1 inst_3307 ( .QN(net_3016), .D(net_2868), .CK(net_5205) );
CLKBUF_X2 inst_4619 ( .A(net_4604), .Z(net_4605) );
NAND2_X2 inst_1587 ( .A1(net_2972), .ZN(net_2432), .A2(net_208) );
NAND4_X2 inst_1185 ( .A1(net_3772), .ZN(net_2153), .A2(net_2042), .A3(net_1891), .A4(net_1097) );
AOI222_X1 inst_3787 ( .A2(net_4105), .C2(net_3656), .ZN(net_1286), .A1(net_1086), .B1(net_890), .C1(net_678), .B2(net_359) );
CLKBUF_X2 inst_4982 ( .A(net_4967), .Z(net_4968) );
OAI21_X2 inst_628 ( .B1(net_2190), .ZN(net_2148), .B2(net_2147), .A(net_2041) );
AOI22_X2 inst_3684 ( .B2(net_4124), .A2(net_509), .ZN(net_499), .A1(net_498), .B1(net_497) );
NAND2_X2 inst_1923 ( .A1(net_3817), .ZN(net_3181), .A2(net_169) );
INV_X2 inst_2748 ( .ZN(net_1110), .A(net_1109) );
INV_X2 inst_3013 ( .A(net_3429), .ZN(net_3398) );
CLKBUF_X2 inst_4744 ( .A(net_4729), .Z(net_4730) );
OAI21_X2 inst_472 ( .B1(net_3509), .ZN(net_2978), .B2(net_2965), .A(net_2445) );
CLKBUF_X2 inst_4533 ( .A(net_4518), .Z(net_4519) );
OAI221_X2 inst_447 ( .ZN(net_3792), .C1(net_988), .B2(net_987), .A(net_876), .B1(net_720), .C2(net_40) );
AOI22_X2 inst_3642 ( .A1(net_4142), .B1(net_4112), .B2(net_1791), .ZN(net_760), .A2(x800) );
OAI21_X4 inst_457 ( .ZN(net_3229), .B1(net_3228), .A(net_1307), .B2(net_316) );
CLKBUF_X2 inst_5087 ( .A(net_5072), .Z(net_5073) );
NAND2_X2 inst_1738 ( .A1(net_2212), .ZN(net_1646), .A2(x1023) );
INV_X4 inst_2623 ( .ZN(net_3958), .A(net_3441) );
INV_X2 inst_2802 ( .ZN(net_728), .A(net_727) );
AND2_X4 inst_4171 ( .ZN(net_4125), .A1(net_3450), .A2(net_359) );
NAND2_X4 inst_1391 ( .ZN(net_2173), .A1(net_2083), .A2(net_1984) );
HA_X1 inst_3092 ( .S(net_1526), .CO(net_1525), .A(net_1306), .B(net_61) );
OAI21_X2 inst_665 ( .B2(net_3149), .ZN(net_1619), .A(net_1531), .B1(net_1465) );
CLKBUF_X2 inst_4843 ( .A(net_4369), .Z(net_4829) );
INV_X2 inst_2734 ( .ZN(net_1384), .A(net_1333) );
CLKBUF_X2 inst_4920 ( .A(net_4905), .Z(net_4906) );
DFF_X1 inst_3395 ( .Q(net_3119), .D(net_1540), .CK(net_4311) );
NOR2_X2 inst_1130 ( .A2(net_3764), .ZN(net_3563), .A1(net_526) );
AOI22_X2 inst_3538 ( .A1(net_1794), .B1(net_1793), .ZN(net_1744), .B2(net_396), .A2(net_229) );
OAI211_X2 inst_855 ( .ZN(net_3748), .C2(net_3747), .B(net_3744), .A(net_3742), .C1(net_3739) );
NAND2_X2 inst_2039 ( .ZN(net_3797), .A1(net_3203), .A2(net_1979) );
AOI222_X1 inst_3755 ( .A1(net_3676), .B1(net_2055), .C1(net_2054), .ZN(net_2038), .B2(net_2037), .C2(net_308), .A2(net_265) );
SDFF_X2 inst_146 ( .D(net_3883), .SE(net_2514), .SI(net_91), .Q(net_91), .CK(net_4945) );
DFF_X1 inst_3233 ( .QN(net_3063), .D(net_2968), .CK(net_4931) );
AOI21_X2 inst_3999 ( .B2(net_3777), .B1(net_3711), .ZN(net_3635), .A(net_749) );
NAND4_X2 inst_1196 ( .ZN(net_1678), .A3(net_1483), .A4(net_1482), .A1(net_1417), .A2(net_1416) );
OAI22_X2 inst_326 ( .B1(net_3619), .ZN(net_930), .A1(net_929), .A2(net_928), .B2(net_299) );
OAI211_X2 inst_817 ( .C1(net_1764), .ZN(net_1726), .A(net_1620), .B(net_1112), .C2(net_406) );
CLKBUF_X2 inst_4295 ( .A(net_4245), .Z(net_4281) );
INV_X4 inst_2194 ( .ZN(net_2531), .A(net_2306) );
DFF_X1 inst_3428 ( .Q(net_4017), .D(net_4016), .CK(net_4906) );
OAI21_X2 inst_518 ( .B2(net_3208), .B1(net_2923), .ZN(net_2922), .A(net_2489) );
NAND3_X2 inst_1363 ( .ZN(net_3888), .A1(net_3698), .A2(net_3390), .A3(net_317) );
CLKBUF_X2 inst_4851 ( .A(net_4836), .Z(net_4837) );
DFF_X1 inst_3336 ( .D(net_3361), .QN(net_117), .CK(net_4456) );
AOI221_X2 inst_3863 ( .B2(net_3116), .B1(net_2020), .C1(net_2019), .ZN(net_2015), .A(net_1896), .C2(x179) );
DFF_X1 inst_3293 ( .QN(net_3011), .D(net_2885), .CK(net_5122) );
INV_X4 inst_2345 ( .A(net_3789), .ZN(net_1011) );
INV_X2 inst_2837 ( .A(net_627), .ZN(net_588) );
AOI222_X1 inst_3793 ( .ZN(net_3677), .A1(net_3676), .B1(net_2055), .C1(net_2054), .B2(net_1791), .C2(net_515), .A2(net_287) );
XNOR2_X2 inst_108 ( .A(net_3818), .ZN(net_427), .B(net_122) );
NAND2_X2 inst_1845 ( .ZN(net_720), .A1(net_641), .A2(net_407) );
CLKBUF_X2 inst_4799 ( .A(net_4441), .Z(net_4785) );
AOI222_X1 inst_3778 ( .ZN(net_1798), .C2(net_1797), .B1(net_1795), .A1(net_1794), .C1(net_1793), .B2(net_1045), .A2(net_224) );
AOI22_X2 inst_3602 ( .A1(net_4059), .B1(net_4057), .A2(net_3024), .B2(net_3022), .ZN(net_1415) );
CLKBUF_X2 inst_5260 ( .A(net_5245), .Z(net_5246) );
AOI21_X2 inst_3940 ( .A(net_2525), .ZN(net_2255), .B1(net_2217), .B2(net_2154) );
CLKBUF_X2 inst_5190 ( .A(net_5175), .Z(net_5176) );
NAND3_X2 inst_1354 ( .ZN(net_3687), .A1(net_3305), .A2(net_2161), .A3(net_1436) );
NAND2_X4 inst_1429 ( .A2(net_3823), .ZN(net_3630), .A1(net_3629) );
NOR2_X4 inst_970 ( .ZN(net_3881), .A2(net_3880), .A1(net_3879) );
NAND3_X2 inst_1278 ( .ZN(net_2825), .A2(net_2597), .A1(net_2577), .A3(net_914) );
AOI222_X1 inst_3763 ( .C1(net_3121), .A1(net_2055), .B1(net_2054), .C2(net_2053), .ZN(net_1999), .B2(net_1281), .A2(net_179) );
OAI21_X2 inst_638 ( .B2(net_2076), .ZN(net_2072), .A(net_1965), .B1(net_1679) );
OAI21_X2 inst_586 ( .ZN(net_2792), .B1(net_2609), .A(net_2391), .B2(net_1275) );
OAI21_X2 inst_749 ( .ZN(net_3403), .B2(net_3124), .B1(net_3108), .A(net_296) );
CLKBUF_X2 inst_5220 ( .A(net_4940), .Z(net_5206) );
NOR2_X2 inst_1030 ( .ZN(net_1795), .A1(net_1459), .A2(net_1036) );
INV_X8 inst_2127 ( .ZN(net_555), .A(net_353) );
INV_X4 inst_2591 ( .A(net_3720), .ZN(net_3680) );
INV_X2 inst_2649 ( .A(net_3883), .ZN(net_2371) );
CLKBUF_X2 inst_5008 ( .A(net_4993), .Z(net_4994) );
DFF_X1 inst_3275 ( .QN(net_3037), .D(net_2926), .CK(net_5179) );
NAND2_X4 inst_1466 ( .A1(net_3933), .ZN(net_3890), .A2(net_767) );
NAND2_X2 inst_1726 ( .A1(net_3599), .ZN(net_1905), .A2(net_1568) );
INV_X2 inst_2841 ( .ZN(net_521), .A(net_399) );
CLKBUF_X2 inst_5221 ( .A(net_5206), .Z(net_5207) );
NAND3_X2 inst_1373 ( .ZN(net_4173), .A1(net_4172), .A3(net_4168), .A2(net_3737) );
INV_X4 inst_2268 ( .ZN(net_1548), .A(net_1022) );
INV_X2 inst_2652 ( .ZN(net_2289), .A(net_2277) );
NAND4_X2 inst_1203 ( .ZN(net_1670), .A3(net_1471), .A4(net_1470), .A1(net_1405), .A2(net_1404) );
INV_X4 inst_2458 ( .A(net_3115), .ZN(net_2637) );
AOI221_X2 inst_3828 ( .B1(net_3469), .B2(net_3141), .C1(net_2534), .ZN(net_2532), .A(net_2337), .C2(net_295) );
OAI22_X2 inst_296 ( .B2(net_3163), .A2(net_2514), .A1(net_1808), .ZN(net_1697), .B1(x475) );
OAI211_X2 inst_802 ( .C1(net_2190), .ZN(net_2166), .C2(net_2165), .A(net_2010), .B(net_1989) );
NOR3_X2 inst_905 ( .A1(net_4113), .A3(net_3387), .A2(net_920), .ZN(net_688) );
DFF_X2 inst_3155 ( .D(net_2255), .QN(net_125), .CK(net_4800) );
DFF_X2 inst_3134 ( .D(net_2627), .QN(net_42), .CK(net_4807) );
CLKBUF_X2 inst_4370 ( .A(net_4355), .Z(net_4356) );
NOR2_X2 inst_1006 ( .A1(net_1807), .ZN(net_1805), .A2(net_1090) );
NAND2_X2 inst_1985 ( .A2(net_4141), .ZN(net_3420), .A1(net_3416) );
CLKBUF_X2 inst_4214 ( .A(net_4197), .Z(net_4200) );
AOI221_X2 inst_3834 ( .ZN(net_2251), .C1(net_2249), .B2(net_1636), .C2(net_1294), .A(net_1227), .B1(net_861) );
AND4_X4 inst_4043 ( .ZN(net_4041), .A3(net_3160), .A1(net_2114), .A4(net_158), .A2(net_85) );
AOI21_X2 inst_3943 ( .B1(net_3774), .ZN(net_2229), .A(net_2146), .B2(net_240) );
AOI22_X2 inst_3651 ( .ZN(net_733), .A1(net_732), .B1(net_731), .A2(net_458), .B2(net_457) );
NAND2_X2 inst_1759 ( .A2(net_1394), .ZN(net_1240), .A1(net_32) );
INV_X4 inst_2615 ( .ZN(net_3859), .A(net_3858) );
INV_X4 inst_2532 ( .ZN(net_3307), .A(net_3306) );
CLKBUF_X2 inst_5134 ( .A(net_5119), .Z(net_5120) );
INV_X4 inst_2463 ( .A(net_3073), .ZN(net_493) );
AOI22_X2 inst_3463 ( .B2(net_4078), .A2(net_3140), .ZN(net_2793), .A1(net_2792), .B1(net_2707) );
CLKBUF_X2 inst_4753 ( .A(net_4738), .Z(net_4739) );
AND4_X2 inst_4055 ( .ZN(net_1761), .A1(net_1760), .A2(net_1548), .A4(net_1264), .A3(net_1225) );
NAND4_X2 inst_1247 ( .ZN(net_3572), .A4(net_3571), .A3(net_1385), .A1(net_1011), .A2(net_618) );
NAND2_X4 inst_1464 ( .ZN(net_3884), .A2(net_3812), .A1(net_2280) );
CLKBUF_X2 inst_5284 ( .A(net_5269), .Z(net_5270) );
CLKBUF_X2 inst_4947 ( .A(net_4932), .Z(net_4933) );
CLKBUF_X2 inst_5031 ( .A(net_5016), .Z(net_5017) );
NAND2_X2 inst_1493 ( .A2(net_3884), .ZN(net_2831), .A1(net_2795) );
NAND3_X2 inst_1308 ( .A3(net_1261), .ZN(net_1134), .A1(net_1053), .A2(net_915) );
CLKBUF_X2 inst_4733 ( .A(net_4718), .Z(net_4719) );
XNOR2_X2 inst_85 ( .B(net_4119), .ZN(net_1748), .A(net_932) );
INV_X1 inst_3070 ( .A(net_3463), .ZN(net_2707) );
CLKBUF_X2 inst_4588 ( .A(net_4524), .Z(net_4574) );
INV_X2 inst_2998 ( .A(net_3066), .ZN(net_139) );
INV_X4 inst_2612 ( .ZN(net_3824), .A(net_3769) );
AND2_X4 inst_4184 ( .A2(net_4162), .ZN(net_4146), .A1(net_3729) );
AND4_X4 inst_4049 ( .ZN(net_4089), .A3(net_562), .A4(net_548), .A2(net_491), .A1(net_477) );
CLKBUF_X2 inst_5067 ( .A(net_5052), .Z(net_5053) );
INV_X2 inst_2702 ( .ZN(net_1675), .A(net_1674) );
INV_X2 inst_2910 ( .ZN(net_1447), .A(net_72) );
CLKBUF_X2 inst_4670 ( .A(net_4655), .Z(net_4656) );
AOI211_X2 inst_4022 ( .C1(net_4084), .C2(net_3915), .ZN(net_1299), .B(net_1110), .A(net_944) );
NAND3_X2 inst_1362 ( .ZN(net_3878), .A3(net_3877), .A2(net_3876), .A1(net_3875) );
DFF_X1 inst_3238 ( .QN(net_3040), .D(net_2928), .CK(net_5191) );
OAI22_X2 inst_290 ( .A1(net_3781), .B1(net_1884), .ZN(net_1864), .A2(net_1714), .B2(net_322) );
SDFF_X2 inst_145 ( .D(net_3866), .SE(net_2625), .SI(net_105), .Q(net_105), .CK(net_4946) );
NAND2_X2 inst_1978 ( .ZN(net_3377), .A1(net_978), .A2(net_872) );
OR2_X2 inst_272 ( .ZN(net_3801), .A1(net_3318), .A2(net_513) );
CLKBUF_X2 inst_4718 ( .A(net_4208), .Z(net_4704) );
INV_X2 inst_2854 ( .A(net_3669), .ZN(net_543) );
INV_X2 inst_3030 ( .ZN(net_3542), .A(net_3540) );
MUX2_X2 inst_2112 ( .A(net_3999), .B(net_3734), .Z(net_1243), .S(net_1178) );
CLKBUF_X2 inst_4594 ( .A(net_4579), .Z(net_4580) );
OAI211_X2 inst_814 ( .B(net_1628), .C1(net_1627), .ZN(net_1624), .A(net_1551), .C2(net_513) );
INV_X2 inst_3036 ( .ZN(net_3589), .A(net_3587) );
INV_X4 inst_2230 ( .ZN(net_1829), .A(net_1681) );
CLKBUF_X2 inst_5203 ( .A(net_5188), .Z(net_5189) );
AND2_X4 inst_4133 ( .ZN(net_4062), .A2(net_3339), .A1(net_1136) );
NAND2_X4 inst_1458 ( .ZN(net_3853), .A2(net_3852), .A1(net_3851) );
AOI22_X2 inst_3471 ( .B2(net_3121), .A1(net_2724), .B1(net_2722), .ZN(net_2719), .A2(net_30) );
OAI211_X2 inst_789 ( .C2(net_2778), .ZN(net_2755), .C1(net_2684), .A(net_2658), .B(net_2604) );
NAND2_X2 inst_1806 ( .A1(net_4082), .ZN(net_1250), .A2(net_912) );
NAND2_X2 inst_1810 ( .ZN(net_1132), .A2(net_899), .A1(net_695) );
NAND2_X2 inst_1860 ( .A2(net_4125), .ZN(net_650), .A1(net_609) );
INV_X4 inst_2275 ( .ZN(net_1196), .A(net_1005) );
NAND2_X2 inst_1885 ( .ZN(net_517), .A2(net_516), .A1(net_403) );
NAND2_X4 inst_1437 ( .ZN(net_3684), .A1(net_3682), .A2(net_86) );
OAI211_X2 inst_822 ( .ZN(net_1657), .A(net_1331), .C2(net_1330), .B(net_1277), .C1(net_1079) );
CLKBUF_X2 inst_4341 ( .A(net_4326), .Z(net_4327) );
NOR2_X2 inst_1125 ( .ZN(net_3454), .A1(net_3453), .A2(net_2986) );
CLKBUF_X2 inst_4885 ( .A(net_4710), .Z(net_4871) );
OAI21_X2 inst_609 ( .B2(net_2815), .ZN(net_2305), .B1(net_2304), .A(net_1792) );
CLKBUF_X2 inst_4477 ( .A(net_4462), .Z(net_4463) );
INV_X4 inst_2533 ( .ZN(net_3313), .A(net_1436) );
INV_X4 inst_2391 ( .ZN(net_412), .A(net_363) );
OAI211_X2 inst_795 ( .C2(net_4069), .ZN(net_2603), .C1(net_2601), .A(net_2387), .B(net_218) );
INV_X4 inst_2496 ( .A(net_2996), .ZN(net_186) );
INV_X4 inst_2239 ( .A(net_1817), .ZN(net_1794) );
XOR2_X1 inst_27 ( .Z(net_1446), .A(net_1445), .B(net_300) );
INV_X4 inst_2491 ( .A(net_3091), .ZN(net_597) );
NAND2_X2 inst_1639 ( .ZN(net_2183), .A2(net_2155), .A1(net_2069) );
CLKBUF_X2 inst_4381 ( .A(net_4236), .Z(net_4367) );
CLKBUF_X2 inst_4446 ( .A(net_4431), .Z(net_4432) );
OAI21_X2 inst_619 ( .ZN(net_2283), .B1(net_2152), .A(net_1799), .B2(net_1738) );
INV_X2 inst_2671 ( .A(net_3772), .ZN(net_2118) );
CLKBUF_X2 inst_5155 ( .A(net_4725), .Z(net_5141) );
NAND2_X2 inst_1654 ( .A2(net_4017), .A1(net_3280), .ZN(net_2128) );
CLKBUF_X2 inst_4547 ( .A(net_4532), .Z(net_4533) );
CLKBUF_X2 inst_5230 ( .A(net_5215), .Z(net_5216) );
OAI21_X2 inst_639 ( .B2(net_2076), .ZN(net_2071), .A(net_1966), .B1(net_1665) );
NAND3_X2 inst_1355 ( .ZN(net_3694), .A1(net_3687), .A2(net_3309), .A3(net_3306) );
NOR3_X4 inst_877 ( .A3(net_3969), .A1(net_3626), .ZN(net_3437), .A2(net_1321) );
SDFF_X2 inst_155 ( .SI(net_4024), .Q(net_4024), .SE(net_2514), .D(net_1784), .CK(net_4936) );
CLKBUF_X2 inst_4858 ( .A(net_4843), .Z(net_4844) );
AOI21_X2 inst_3939 ( .A(net_2300), .ZN(net_2267), .B1(net_2212), .B2(net_248) );
CLKBUF_X2 inst_5309 ( .A(net_5294), .Z(net_5295) );
XNOR2_X2 inst_55 ( .ZN(net_2332), .A(net_2283), .B(net_1780) );
INV_X8 inst_2167 ( .ZN(net_3870), .A(net_3869) );
INV_X4 inst_2280 ( .A(net_1256), .ZN(net_1201) );
NAND2_X2 inst_2076 ( .A2(net_4175), .ZN(net_4167), .A1(net_4166) );
CLKBUF_X2 inst_4248 ( .A(net_4233), .Z(net_4234) );
NAND2_X2 inst_1651 ( .A1(net_2597), .A2(net_2302), .ZN(net_2214) );
AND2_X4 inst_4127 ( .ZN(net_4054), .A2(net_1328), .A1(net_1216) );
INV_X4 inst_2481 ( .A(net_3151), .ZN(net_2665) );
CLKBUF_X2 inst_4285 ( .A(net_4270), .Z(net_4271) );
NOR2_X2 inst_1137 ( .A2(net_3954), .A1(net_3953), .ZN(net_3761) );
OAI22_X2 inst_323 ( .B1(net_2717), .A2(net_1274), .ZN(net_1245), .B2(net_987), .A1(net_831) );
NOR2_X2 inst_1162 ( .ZN(net_4166), .A1(net_1994), .A2(net_73) );
NAND2_X4 inst_1389 ( .A1(net_3537), .ZN(net_2739), .A2(net_2530) );
INV_X2 inst_2973 ( .A(net_3025), .ZN(net_129) );
INV_X16 inst_3065 ( .ZN(net_530), .A(net_337) );
OAI21_X2 inst_715 ( .A(net_1264), .ZN(net_1229), .B1(net_658), .B2(net_652) );
OAI211_X2 inst_793 ( .ZN(net_2692), .B(net_2691), .C2(net_2690), .C1(net_2511), .A(net_2510) );
NAND2_X4 inst_1433 ( .ZN(net_3669), .A1(net_3654), .A2(net_3107) );
NAND2_X2 inst_1494 ( .ZN(net_2824), .A1(net_2790), .A2(net_2323) );
CLKBUF_X2 inst_5206 ( .A(net_4306), .Z(net_5192) );
CLKBUF_X2 inst_5213 ( .A(net_4917), .Z(net_5199) );
NAND2_X2 inst_1894 ( .A2(net_513), .ZN(net_436), .A1(net_377) );
CLKBUF_X2 inst_4815 ( .A(net_4276), .Z(net_4801) );
AOI22_X2 inst_3525 ( .A2(net_3143), .A1(net_1923), .B1(net_1921), .ZN(net_1919), .B2(net_301) );
CLKBUF_X2 inst_4643 ( .A(net_4628), .Z(net_4629) );
NAND2_X2 inst_1999 ( .ZN(net_3491), .A2(net_3331), .A1(net_447) );
NAND2_X2 inst_1682 ( .A1(net_3176), .ZN(net_2024), .A2(net_187) );
CLKBUF_X2 inst_5077 ( .A(net_5062), .Z(net_5063) );
INV_X2 inst_2733 ( .ZN(net_1391), .A(net_1346) );
NAND3_X2 inst_1340 ( .ZN(net_3373), .A1(net_3371), .A3(net_2836), .A2(net_2757) );
NAND2_X4 inst_1481 ( .ZN(net_3967), .A2(net_3959), .A1(net_3958) );
OAI21_X2 inst_475 ( .B1(net_3509), .ZN(net_2975), .B2(net_2959), .A(net_2502) );
CLKBUF_X2 inst_4738 ( .A(net_4308), .Z(net_4724) );
CLKBUF_X2 inst_4412 ( .A(net_4242), .Z(net_4398) );
XOR2_X1 inst_31 ( .A(net_4129), .Z(net_382), .B(net_255) );
INV_X2 inst_2701 ( .ZN(net_1677), .A(net_1676) );
AOI22_X2 inst_3505 ( .B1(net_3676), .B2(net_3145), .A2(net_2037), .ZN(net_2013), .A1(net_2012) );
DFF_X2 inst_3165 ( .D(net_2070), .QN(net_88), .CK(net_5142) );
DFF_X2 inst_3217 ( .D(net_805), .QN(net_332), .CK(net_4616) );
OAI21_X2 inst_575 ( .B2(net_2919), .ZN(net_2804), .B1(net_2803), .A(net_2402) );
CLKBUF_X2 inst_4331 ( .A(net_4197), .Z(net_4317) );
CLKBUF_X2 inst_4376 ( .A(net_4361), .Z(net_4362) );
AOI22_X2 inst_3537 ( .A1(net_1794), .B1(net_1793), .ZN(net_1745), .B2(net_378), .A2(net_216) );
CLKBUF_X2 inst_4705 ( .A(net_4690), .Z(net_4691) );
CLKBUF_X2 inst_4556 ( .A(net_4541), .Z(net_4542) );
OAI21_X2 inst_627 ( .B2(net_4088), .B1(net_2190), .ZN(net_2149), .A(net_2040) );
CLKBUF_X2 inst_4725 ( .A(net_4710), .Z(net_4711) );
DFF_X1 inst_3352 ( .QN(net_3123), .D(net_2700), .CK(net_4820) );
OAI22_X2 inst_344 ( .ZN(net_3552), .A1(net_3551), .A2(net_3496), .B2(net_3492), .B1(net_1691) );
NAND2_X2 inst_1833 ( .A2(net_3627), .ZN(net_1129), .A1(net_614) );
CLKBUF_X2 inst_5301 ( .A(net_5286), .Z(net_5287) );
INV_X8 inst_2122 ( .ZN(net_723), .A(net_435) );
INV_X2 inst_3044 ( .ZN(net_3703), .A(net_1857) );
AOI22_X2 inst_3520 ( .B1(net_4045), .B2(net_3115), .A1(net_1955), .ZN(net_1950), .A2(net_267) );
AOI22_X2 inst_3573 ( .A1(net_4059), .B1(net_4056), .ZN(net_1477), .A2(net_215), .B2(net_187) );
OAI21_X2 inst_623 ( .B1(net_2235), .ZN(net_2158), .A(net_2050), .B2(net_107) );
NOR2_X2 inst_1072 ( .A1(net_2525), .ZN(net_718), .A2(x964) );
AOI22_X2 inst_3580 ( .A1(net_4060), .B1(net_4055), .ZN(net_1470), .A2(net_190), .B2(net_161) );
AOI221_X2 inst_3818 ( .A(net_2642), .B1(net_2641), .C2(net_2581), .C1(net_2563), .ZN(net_2560), .B2(net_267) );
NAND2_X2 inst_1621 ( .A1(net_2917), .ZN(net_2395), .A2(net_141) );
NAND2_X2 inst_1993 ( .ZN(net_3463), .A2(net_2680), .A1(net_2596) );
NAND3_X2 inst_1338 ( .A3(net_3343), .ZN(net_3288), .A1(net_3287), .A2(net_3277) );
INV_X4 inst_2430 ( .A(net_3079), .ZN(net_454) );
INV_X1 inst_3080 ( .A(net_3135), .ZN(net_280) );
CLKBUF_X2 inst_4952 ( .A(net_4937), .Z(net_4938) );
INV_X4 inst_2434 ( .A(net_3055), .ZN(net_475) );
DFF_X1 inst_3226 ( .QN(net_3054), .D(net_2976), .CK(net_4564) );
AOI22_X1 inst_3731 ( .B1(net_4054), .B2(net_1874), .A2(net_1797), .A1(net_1578), .ZN(net_1575) );
NOR2_X2 inst_1107 ( .A1(net_3871), .ZN(net_3233), .A2(net_136) );
AOI22_X2 inst_3617 ( .B1(net_3156), .B2(net_1636), .ZN(net_1325), .A1(net_1324), .A2(net_1228) );
CLKBUF_X2 inst_4839 ( .A(net_4819), .Z(net_4825) );
NAND3_X1 inst_1377 ( .A2(net_3321), .A1(net_1827), .ZN(net_1773), .A3(net_1772) );
NAND2_X2 inst_2028 ( .ZN(net_3742), .A2(net_3741), .A1(net_3739) );
DFF_X2 inst_3125 ( .QN(net_3139), .D(net_2696), .CK(net_4577) );
INV_X4 inst_2201 ( .ZN(net_2361), .A(net_2265) );
CLKBUF_X2 inst_4253 ( .A(net_4238), .Z(net_4239) );
OAI21_X2 inst_722 ( .B2(net_3387), .ZN(net_921), .A(net_662), .B1(net_311) );
INV_X2 inst_2776 ( .ZN(net_832), .A(net_831) );
OAI21_X2 inst_760 ( .ZN(net_3751), .B2(net_3745), .A(net_3229), .B1(net_2623) );
OAI21_X2 inst_746 ( .B1(net_4187), .ZN(net_3367), .B2(net_3366), .A(net_2579) );
NAND2_X2 inst_1696 ( .A2(net_3229), .ZN(net_2876), .A1(net_2049) );
CLKBUF_X2 inst_4232 ( .A(net_4202), .Z(net_4218) );
CLKBUF_X2 inst_4270 ( .A(net_4255), .Z(net_4256) );
INV_X4 inst_2267 ( .ZN(net_2272), .A(net_1099) );
INV_X2 inst_3010 ( .ZN(net_3372), .A(net_3371) );
CLKBUF_X2 inst_4911 ( .A(net_4896), .Z(net_4897) );
CLKBUF_X2 inst_4525 ( .A(net_4510), .Z(net_4511) );
AND2_X4 inst_4115 ( .A2(net_4131), .ZN(net_3616), .A1(net_3220) );
DFF_X2 inst_3133 ( .D(net_2628), .QN(net_40), .CK(net_4808) );
AOI22_X2 inst_3727 ( .ZN(net_3747), .B1(net_3746), .A2(net_3745), .A1(net_3738), .B2(net_67) );
NAND2_X2 inst_1577 ( .A1(net_2965), .ZN(net_2443), .A2(net_559) );
NAND2_X2 inst_1687 ( .A1(net_3219), .ZN(net_1985), .A2(net_235) );
NOR2_X2 inst_1110 ( .A1(net_3752), .ZN(net_3309), .A2(net_1443) );
NAND2_X2 inst_1970 ( .A2(net_3399), .ZN(net_3338), .A1(x475) );
INV_X4 inst_2588 ( .ZN(net_3668), .A(net_3521) );
AOI21_X2 inst_3989 ( .ZN(net_1058), .A(net_881), .B1(net_707), .B2(net_541) );
INV_X2 inst_2873 ( .A(net_3109), .ZN(net_249) );
CLKBUF_X2 inst_4665 ( .A(net_4650), .Z(net_4651) );
INV_X4 inst_2442 ( .A(net_3071), .ZN(net_471) );
AOI22_X2 inst_3569 ( .B1(net_4062), .A1(net_4056), .A2(net_3025), .B2(net_3023), .ZN(net_1481) );
NAND2_X2 inst_2066 ( .ZN(net_3960), .A2(net_3959), .A1(net_3958) );
DFF_X1 inst_3411 ( .D(net_1392), .Q(net_51), .CK(net_4495) );
INV_X4 inst_2524 ( .ZN(net_3262), .A(net_3261) );
NAND2_X4 inst_1446 ( .A2(net_3893), .A1(net_3870), .ZN(net_3799) );
OAI221_X2 inst_390 ( .C2(net_3408), .ZN(net_2363), .B1(net_2361), .C1(net_2225), .A(net_1944), .B2(net_110) );
INV_X4 inst_2421 ( .A(net_3103), .ZN(net_261) );
CLKBUF_X2 inst_4842 ( .A(net_4827), .Z(net_4828) );
NAND2_X2 inst_1742 ( .ZN(net_1595), .A1(net_1440), .A2(net_1439) );
CLKBUF_X2 inst_4466 ( .A(net_4451), .Z(net_4452) );
NOR2_X2 inst_1062 ( .A1(net_3661), .ZN(net_1037), .A2(net_705) );
INV_X2 inst_2663 ( .A(net_3186), .ZN(net_2353) );
INV_X2 inst_2875 ( .ZN(net_303), .A(net_207) );
DFF_X1 inst_3289 ( .QN(net_3048), .D(net_2898), .CK(net_4714) );
CLKBUF_X2 inst_4779 ( .A(net_4764), .Z(net_4765) );
OAI221_X2 inst_401 ( .C2(net_3428), .ZN(net_2236), .B1(net_2235), .C1(net_2044), .A(net_1990), .B2(net_264) );
INV_X4 inst_2302 ( .A(net_3430), .ZN(net_1908) );
DFF_X2 inst_3175 ( .D(net_1864), .QN(net_29), .CK(net_4679) );
DFF_X1 inst_3389 ( .D(net_1729), .QN(net_80), .CK(net_4249) );
DFF_X2 inst_3210 ( .D(net_804), .QN(net_316), .CK(net_4672) );
INV_X4 inst_2447 ( .A(net_2995), .ZN(net_153) );
OAI211_X2 inst_782 ( .ZN(net_2780), .C2(net_2778), .B(net_2677), .C1(net_2669), .A(net_2655) );
CLKBUF_X2 inst_5200 ( .A(net_5185), .Z(net_5186) );
INV_X2 inst_2642 ( .ZN(net_2339), .A(net_2319) );
INV_X2 inst_2869 ( .ZN(net_301), .A(net_50) );
CLKBUF_X2 inst_4653 ( .A(net_4638), .Z(net_4639) );
XOR2_X2 inst_6 ( .A(net_3497), .B(net_3492), .Z(net_1693) );
INV_X4 inst_2486 ( .A(net_3080), .ZN(net_453) );
INV_X4 inst_2410 ( .A(net_3106), .ZN(net_306) );
CLKBUF_X2 inst_4465 ( .A(net_4450), .Z(net_4451) );
CLKBUF_X2 inst_4865 ( .A(net_4850), .Z(net_4851) );
CLKBUF_X2 inst_5250 ( .A(net_5235), .Z(net_5236) );
XNOR2_X2 inst_123 ( .ZN(net_4150), .A(net_3805), .B(net_2811) );
NOR2_X4 inst_930 ( .A1(net_3557), .ZN(net_2030), .A2(net_247) );
CLKBUF_X2 inst_4803 ( .A(net_4788), .Z(net_4789) );
INV_X8 inst_2160 ( .ZN(net_3645), .A(net_1982) );
NOR2_X4 inst_935 ( .A1(net_3324), .ZN(net_435), .A2(net_359) );
CLKBUF_X2 inst_5181 ( .A(net_5166), .Z(net_5167) );
CLKBUF_X2 inst_4772 ( .A(net_4205), .Z(net_4758) );
CLKBUF_X2 inst_4634 ( .A(net_4497), .Z(net_4620) );
INV_X4 inst_2298 ( .ZN(net_1092), .A(net_824) );
OR3_X4 inst_167 ( .ZN(net_1912), .A1(net_1587), .A3(net_1586), .A2(net_1583) );
INV_X2 inst_2944 ( .A(net_3045), .ZN(net_169) );
NOR2_X2 inst_1026 ( .A1(net_1646), .ZN(net_1607), .A2(net_1367) );
NAND3_X2 inst_1320 ( .A1(net_4100), .ZN(net_769), .A3(net_768), .A2(net_206) );
CLKBUF_X2 inst_5011 ( .A(net_4896), .Z(net_4997) );
CLKBUF_X2 inst_4913 ( .A(net_4898), .Z(net_4899) );
AOI221_X2 inst_3874 ( .A(net_4046), .ZN(net_1909), .C2(net_1908), .C1(net_1674), .B2(net_749), .B1(net_99) );
NAND4_X2 inst_1251 ( .A2(net_3911), .ZN(net_3846), .A4(net_3812), .A3(net_3787), .A1(net_3786) );
CLKBUF_X2 inst_5246 ( .A(net_5231), .Z(net_5232) );
XNOR2_X2 inst_95 ( .ZN(net_978), .A(net_713), .B(net_417) );
DFF_X1 inst_3376 ( .D(net_2258), .QN(net_49), .CK(net_4476) );
CLKBUF_X2 inst_4874 ( .A(net_4859), .Z(net_4860) );
INV_X4 inst_2475 ( .ZN(net_323), .A(net_45) );
INV_X2 inst_2921 ( .A(net_3125), .ZN(net_231) );
INV_X2 inst_2862 ( .ZN(net_361), .A(net_192) );
OAI22_X2 inst_331 ( .B2(net_3468), .ZN(net_824), .B1(net_721), .A1(net_641), .A2(net_40) );
AOI21_X2 inst_4009 ( .ZN(net_4160), .B1(net_2243), .A(net_2132), .B2(net_156) );
CLKBUF_X2 inst_4900 ( .A(net_4885), .Z(net_4886) );
INV_X4 inst_2172 ( .ZN(net_2893), .A(net_2880) );
INV_X4 inst_2353 ( .ZN(net_549), .A(net_418) );
OAI21_X2 inst_667 ( .ZN(net_1817), .B1(net_1451), .B2(net_1340), .A(net_1328) );
INV_X2 inst_2762 ( .A(net_3326), .ZN(net_968) );
INV_X2 inst_2896 ( .A(net_3032), .ZN(net_215) );
CLKBUF_X2 inst_4454 ( .A(net_4439), .Z(net_4440) );
NOR2_X2 inst_997 ( .A2(net_3874), .A1(net_3831), .ZN(net_2182) );
NOR4_X2 inst_857 ( .A4(net_4075), .A2(net_4040), .ZN(net_2281), .A3(net_2213), .A1(net_1569) );
CLKBUF_X2 inst_4901 ( .A(net_4886), .Z(net_4887) );
CLKBUF_X2 inst_4824 ( .A(net_4809), .Z(net_4810) );
INV_X2 inst_2691 ( .A(net_3770), .ZN(net_1844) );
AOI22_X2 inst_3590 ( .A1(net_4063), .B1(net_4058), .ZN(net_1427), .B2(net_171), .A2(net_146) );
NAND2_X2 inst_1511 ( .A2(net_3738), .ZN(net_2622), .A1(net_2621) );
CLKBUF_X2 inst_4315 ( .A(net_4300), .Z(net_4301) );
AND2_X4 inst_4179 ( .ZN(net_4136), .A1(net_2161), .A2(net_1436) );
OAI221_X2 inst_365 ( .ZN(net_2734), .B2(net_2733), .C1(net_2732), .C2(net_2731), .B1(net_2645), .A(net_2643) );
AOI21_X2 inst_4006 ( .ZN(net_3931), .B2(net_3930), .B1(net_1167), .A(net_843) );
XNOR2_X2 inst_67 ( .A(net_1718), .ZN(net_1660), .B(net_1456) );
CLKBUF_X2 inst_4243 ( .A(net_4228), .Z(net_4229) );
NOR2_X4 inst_954 ( .ZN(net_3686), .A1(net_3533), .A2(net_3515) );
DFF_X2 inst_3203 ( .Q(net_3157), .D(net_1549), .CK(net_4825) );
CLKBUF_X2 inst_4974 ( .A(net_4959), .Z(net_4960) );
CLKBUF_X2 inst_5073 ( .A(net_5058), .Z(net_5059) );
NAND2_X2 inst_1504 ( .A2(net_3332), .ZN(net_2768), .A1(net_2739) );
INV_X4 inst_2476 ( .A(net_2997), .ZN(net_162) );
DFF_X1 inst_3403 ( .Q(net_4026), .D(net_1467), .CK(net_4509) );
CLKBUF_X2 inst_5084 ( .A(net_5069), .Z(net_5070) );
NAND2_X2 inst_1823 ( .A1(net_4102), .A2(net_4097), .ZN(net_954) );
OR2_X4 inst_202 ( .ZN(net_2963), .A2(net_2352), .A1(net_2351) );
NAND3_X2 inst_1310 ( .A1(net_1279), .ZN(net_1104), .A2(net_1103), .A3(net_1045) );
INV_X4 inst_2212 ( .ZN(net_2263), .A(net_2143) );
DFF_X1 inst_3280 ( .QN(net_3032), .D(net_2913), .CK(net_5083) );
NAND2_X4 inst_1401 ( .ZN(net_451), .A1(net_391), .A2(net_303) );
CLKBUF_X2 inst_4491 ( .A(net_4399), .Z(net_4477) );
CLKBUF_X2 inst_4502 ( .A(net_4443), .Z(net_4488) );
INV_X2 inst_2823 ( .ZN(net_532), .A(net_531) );
CLKBUF_X2 inst_4830 ( .A(net_4206), .Z(net_4816) );
NAND2_X2 inst_2030 ( .A1(net_3995), .ZN(net_3756), .A2(net_3655) );
AOI221_X2 inst_3807 ( .ZN(net_2726), .B1(net_2714), .C2(net_2659), .C1(net_2590), .B2(net_2051), .A(net_1173) );
NOR2_X2 inst_1069 ( .A1(net_2525), .ZN(net_771), .A2(net_770) );
XOR2_X1 inst_30 ( .A(net_4122), .Z(net_512), .B(net_272) );
SDFF_X2 inst_136 ( .D(net_3533), .SE(net_2514), .SI(net_92), .Q(net_92), .CK(net_4963) );
OAI21_X2 inst_610 ( .B2(net_4121), .ZN(net_2352), .A(net_2299), .B1(net_2298) );
AOI22_X2 inst_3541 ( .A1(net_2042), .ZN(net_1605), .B2(net_1463), .B1(net_1453), .A2(net_1377) );
NOR2_X2 inst_1036 ( .A1(net_1340), .ZN(net_1336), .A2(net_1287) );
OR2_X4 inst_233 ( .A1(net_3156), .ZN(net_1884), .A2(net_1173) );
NAND2_X2 inst_1526 ( .A2(net_4015), .A1(net_3208), .ZN(net_2496) );
INV_X4 inst_2547 ( .ZN(net_3447), .A(net_3156) );
CLKBUF_X2 inst_4637 ( .A(net_4622), .Z(net_4623) );
NOR2_X2 inst_1047 ( .ZN(net_1254), .A1(net_1074), .A2(net_898) );
CLKBUF_X2 inst_5167 ( .A(net_4238), .Z(net_5153) );
XNOR2_X2 inst_60 ( .ZN(net_2044), .A(net_2043), .B(net_1596) );
AOI221_X2 inst_3850 ( .A(net_4183), .ZN(net_2068), .C1(net_2067), .C2(net_1908), .B2(net_749), .B1(net_93) );
AOI22_X2 inst_3700 ( .B2(net_4124), .A2(net_555), .ZN(net_472), .A1(net_471), .B1(net_470) );
CLKBUF_X2 inst_4613 ( .A(net_4598), .Z(net_4599) );
NAND2_X2 inst_1858 ( .ZN(net_1264), .A2(net_666), .A1(net_522) );
NAND2_X2 inst_1786 ( .A1(net_2596), .ZN(net_2384), .A2(net_266) );
INV_X4 inst_2376 ( .ZN(net_591), .A(net_411) );
AOI221_X2 inst_3846 ( .B1(net_3736), .ZN(net_2139), .C1(net_2137), .A(net_1870), .B2(net_294), .C2(net_229) );
NAND3_X2 inst_1334 ( .A3(net_3395), .A1(net_528), .ZN(net_442), .A2(net_416) );
CLKBUF_X2 inst_4360 ( .A(net_4345), .Z(net_4346) );
OAI21_X2 inst_496 ( .B1(net_3278), .B2(net_3207), .ZN(net_2946), .A(net_2478) );
NOR4_X2 inst_860 ( .A3(net_3486), .ZN(net_1801), .A1(net_1800), .A4(net_1799), .A2(net_1779) );
OAI21_X2 inst_563 ( .B2(net_2919), .ZN(net_2850), .B1(net_2849), .A(net_2401) );
AOI21_X2 inst_3962 ( .ZN(net_1460), .B1(net_1278), .A(net_1223), .B2(net_1222) );
NOR2_X4 inst_943 ( .ZN(net_3371), .A2(net_3291), .A1(net_2788) );
AOI22_X2 inst_3478 ( .B1(net_4039), .A1(net_2675), .ZN(net_2672), .A2(net_204), .B2(x0) );
AOI222_X1 inst_3749 ( .ZN(net_2069), .B1(net_2017), .C1(net_2016), .A1(net_1893), .A2(net_1881), .C2(net_276), .B2(net_274) );
INV_X4 inst_2620 ( .ZN(net_3927), .A(net_3926) );
CLKBUF_X2 inst_4711 ( .A(net_4696), .Z(net_4697) );
INV_X2 inst_2782 ( .ZN(net_804), .A(net_758) );
NAND2_X2 inst_1964 ( .ZN(net_3315), .A2(net_3314), .A1(net_2161) );
NAND2_X2 inst_1633 ( .A2(net_3516), .A1(net_3248), .ZN(net_2679) );
NAND2_X2 inst_1765 ( .A2(net_1394), .ZN(net_1234), .A1(net_30) );
NAND3_X4 inst_1262 ( .A1(net_3554), .ZN(net_2549), .A3(net_2378), .A2(net_1788) );
CLKBUF_X2 inst_5303 ( .A(net_5288), .Z(net_5289) );
OR2_X2 inst_265 ( .A2(net_3166), .ZN(net_363), .A1(net_322) );
AOI22_X2 inst_3720 ( .ZN(net_3608), .A1(net_3178), .B1(net_2099), .B2(net_518), .A2(net_479) );
NAND2_X2 inst_2005 ( .ZN(net_3532), .A2(net_3531), .A1(net_3530) );
NAND2_X2 inst_2055 ( .ZN(net_3903), .A2(net_3901), .A1(net_3430) );
AOI221_X2 inst_3856 ( .B1(net_3736), .C1(net_2049), .ZN(net_2048), .A(net_1929), .C2(net_1715), .B2(net_300) );
OAI21_X2 inst_544 ( .B2(net_2919), .ZN(net_2888), .B1(net_2887), .A(net_2400) );
OAI21_X2 inst_736 ( .A(net_629), .B1(net_628), .ZN(net_574), .B2(net_361) );
CLKBUF_X2 inst_5091 ( .A(net_5076), .Z(net_5077) );
DFF_X1 inst_3262 ( .QN(net_3074), .D(net_2929), .CK(net_4870) );
OR3_X2 inst_178 ( .ZN(net_2857), .A1(net_2835), .A2(net_2809), .A3(net_2806) );
CLKBUF_X2 inst_4566 ( .A(net_4551), .Z(net_4552) );
CLKBUF_X2 inst_4402 ( .A(net_4387), .Z(net_4388) );
OAI21_X2 inst_734 ( .A(net_629), .B1(net_628), .ZN(net_576), .B2(net_323) );
NAND3_X2 inst_1282 ( .ZN(net_2686), .A2(net_2377), .A3(net_2376), .A1(net_2375) );
NOR2_X2 inst_1077 ( .A1(net_3733), .A2(net_3681), .ZN(net_648) );
NOR2_X2 inst_1148 ( .A1(net_3926), .A2(net_3106), .ZN(net_418) );
AOI221_X2 inst_3919 ( .ZN(net_3843), .B2(net_3842), .B1(net_3841), .C2(net_3789), .C1(net_1369), .A(net_933) );
AOI21_X2 inst_3954 ( .ZN(net_1730), .B1(net_1594), .B2(net_1104), .A(net_1090) );
INV_X2 inst_2757 ( .ZN(net_2187), .A(net_1123) );
OR2_X4 inst_222 ( .A2(net_3997), .ZN(net_1295), .A1(net_877) );
NAND2_X2 inst_1932 ( .A2(net_3869), .A1(net_3261), .ZN(net_3197) );
AOI22_X2 inst_3704 ( .B1(net_4124), .A1(net_509), .ZN(net_464), .B2(net_215), .A2(net_187) );
CLKBUF_X2 inst_4350 ( .A(net_4335), .Z(net_4336) );
AOI22_X2 inst_3587 ( .A1(net_4062), .B1(net_4057), .B2(net_4023), .A2(net_4021), .ZN(net_1430) );
NOR2_X2 inst_1052 ( .A1(net_1154), .ZN(net_1078), .A2(net_1033) );
NAND3_X2 inst_1280 ( .A2(net_3449), .ZN(net_2709), .A3(net_2521), .A1(net_2519) );
NAND3_X2 inst_1302 ( .A1(net_4061), .ZN(net_1341), .A2(net_182), .A3(net_115) );
NAND2_X2 inst_1648 ( .ZN(net_2161), .A1(net_2160), .A2(net_1442) );
OAI211_X2 inst_842 ( .ZN(net_1208), .A(net_1109), .B(net_1010), .C1(net_909), .C2(net_667) );
NOR2_X2 inst_1079 ( .A1(net_3984), .ZN(net_692), .A2(net_385) );
NAND2_X2 inst_2068 ( .ZN(net_3973), .A2(net_3967), .A1(net_923) );
AOI21_X4 inst_3925 ( .B2(net_3600), .ZN(net_3509), .A(net_3508), .B1(net_3342) );
OAI21_X2 inst_551 ( .B1(net_4176), .A(net_4174), .ZN(net_2877), .B2(net_2876) );
INV_X4 inst_2606 ( .ZN(net_3785), .A(net_3662) );
CLKBUF_X2 inst_4314 ( .A(net_4282), .Z(net_4300) );
NAND2_X1 inst_2101 ( .ZN(net_3806), .A1(net_3803), .A2(net_3404) );
INV_X4 inst_2523 ( .ZN(net_3257), .A(net_2310) );
OAI21_X2 inst_506 ( .B1(net_3274), .B2(net_2972), .ZN(net_2936), .A(net_2429) );
OAI222_X2 inst_353 ( .A1(net_2815), .B1(net_1817), .C1(net_1816), .ZN(net_1749), .A2(net_1748), .C2(net_260), .B2(net_106) );
AOI221_X2 inst_3808 ( .C1(net_2724), .ZN(net_2715), .B1(net_2714), .A(net_2525), .B2(net_282), .C2(net_37) );
NAND2_X2 inst_1940 ( .A1(net_3280), .ZN(net_3231), .A2(net_488) );
SDFF_X2 inst_134 ( .D(net_3483), .SI(net_3022), .Q(net_3022), .SE(net_2909), .CK(net_5198) );
INV_X4 inst_2409 ( .ZN(net_1401), .A(net_312) );
DFF_X1 inst_3322 ( .QN(net_2998), .D(net_2845), .CK(net_5200) );
NOR2_X2 inst_1085 ( .ZN(net_444), .A1(net_340), .A2(net_281) );
NAND3_X2 inst_1323 ( .ZN(net_1007), .A1(net_723), .A2(net_528), .A3(net_334) );
DFF_X1 inst_3425 ( .Q(net_4011), .D(net_4010), .CK(net_4919) );
CLKBUF_X2 inst_4632 ( .A(net_4617), .Z(net_4618) );
INV_X4 inst_2328 ( .ZN(net_1018), .A(net_685) );
INV_X2 inst_2655 ( .A(net_3611), .ZN(net_2324) );
OR4_X2 inst_160 ( .A3(net_3771), .A4(net_2054), .ZN(net_1890), .A2(net_1844), .A1(net_1806) );
NAND2_X2 inst_1720 ( .A2(net_1884), .ZN(net_1651), .A1(net_1646) );
AND4_X4 inst_4041 ( .A3(net_3934), .ZN(net_3640), .A4(net_3639), .A2(net_3575), .A1(net_1084) );
AOI22_X2 inst_3701 ( .B2(net_4123), .A2(net_509), .ZN(net_469), .A1(net_468), .B1(net_467) );
DFF_X1 inst_3357 ( .D(net_3710), .CK(net_4408), .Q(x409) );
XOR2_X2 inst_8 ( .B(net_4051), .Z(net_1818), .A(net_1163) );
INV_X2 inst_2912 ( .A(net_3014), .ZN(net_173) );
OAI21_X2 inst_762 ( .ZN(net_3841), .A(net_3840), .B2(net_3620), .B1(net_810) );
OAI221_X2 inst_370 ( .B2(net_2733), .ZN(net_2696), .C1(net_2686), .A(net_2582), .B1(net_2304), .C2(net_1652) );
INV_X2 inst_3025 ( .ZN(net_3466), .A(net_331) );
NAND3_X4 inst_1265 ( .A3(net_4144), .ZN(net_3524), .A2(net_3523), .A1(net_3522) );
NAND2_X1 inst_2090 ( .A2(net_3777), .ZN(net_1565), .A1(net_1322) );
NOR2_X4 inst_965 ( .ZN(net_3825), .A1(net_3824), .A2(net_281) );
DFF_X1 inst_3370 ( .D(net_2287), .CK(net_4222), .Q(x232) );
CLKBUF_X2 inst_4530 ( .A(net_4515), .Z(net_4516) );
NAND3_X2 inst_1321 ( .A2(net_3767), .A1(net_963), .ZN(net_774), .A3(net_543) );
NOR2_X2 inst_1012 ( .A2(net_3961), .ZN(net_1893), .A1(net_1746) );
CLKBUF_X2 inst_5255 ( .A(net_5240), .Z(net_5241) );
NOR3_X2 inst_901 ( .A1(net_1650), .ZN(net_1047), .A2(net_1046), .A3(net_1045) );
NAND2_X2 inst_1956 ( .ZN(net_3294), .A1(net_3293), .A2(net_200) );
AOI22_X2 inst_3492 ( .B1(net_3469), .B2(net_3138), .A1(net_2534), .ZN(net_2276), .A2(net_287) );
OAI21_X2 inst_751 ( .ZN(net_3495), .B1(net_3494), .A(net_3493), .B2(net_3491) );
DFF_X2 inst_3149 ( .QN(net_3128), .D(net_2355), .CK(net_5145) );
CLKBUF_X2 inst_4283 ( .A(net_4268), .Z(net_4269) );
INV_X4 inst_2403 ( .ZN(net_326), .A(net_325) );
INV_X4 inst_2471 ( .ZN(net_138), .A(net_52) );
AOI211_X2 inst_4034 ( .ZN(net_4153), .B(net_1208), .C1(net_1196), .A(net_1066), .C2(net_407) );
OAI221_X2 inst_377 ( .B1(net_2670), .C1(net_2668), .ZN(net_2667), .B2(net_2666), .C2(net_2665), .A(net_593) );
CLKBUF_X2 inst_4948 ( .A(net_4933), .Z(net_4934) );
CLKBUF_X2 inst_4760 ( .A(net_4745), .Z(net_4746) );
NAND2_X2 inst_1934 ( .ZN(net_3201), .A1(net_3198), .A2(net_141) );
AOI21_X2 inst_3946 ( .B1(net_3774), .ZN(net_2219), .A(net_2151), .B2(net_300) );
HA_X1 inst_3098 ( .CO(net_766), .S(net_677), .B(net_504), .A(net_452) );
DFF_X1 inst_3244 ( .QN(net_3093), .D(net_2954), .CK(net_4784) );
AOI221_X2 inst_3916 ( .B1(net_3504), .ZN(net_3470), .C1(net_3469), .A(net_3467), .C2(net_3143), .B2(net_402) );
AOI221_X1 inst_3920 ( .C1(net_3241), .B2(net_3132), .B1(net_2591), .C2(net_2589), .ZN(net_2566), .A(net_1090) );
AOI221_X2 inst_3821 ( .A(net_2642), .B1(net_2641), .C1(net_2581), .ZN(net_2557), .C2(net_2553), .B2(net_295) );
INV_X2 inst_3018 ( .ZN(net_3418), .A(net_40) );
INV_X1 inst_3078 ( .A(net_3478), .ZN(net_649) );
CLKBUF_X2 inst_5013 ( .A(net_4825), .Z(net_4999) );
CLKBUF_X2 inst_4623 ( .A(net_4532), .Z(net_4609) );
CLKBUF_X2 inst_5054 ( .A(net_4480), .Z(net_5040) );
AOI221_X2 inst_3835 ( .B1(net_3774), .ZN(net_2234), .C1(net_2227), .A(net_2107), .B2(net_1511), .C2(net_869) );
CLKBUF_X2 inst_4627 ( .A(net_4612), .Z(net_4613) );
NAND2_X1 inst_2097 ( .A2(net_3876), .A1(net_3875), .ZN(net_3577) );
CLKBUF_X2 inst_4484 ( .A(net_4469), .Z(net_4470) );
NOR2_X4 inst_928 ( .A1(net_3283), .ZN(net_2095), .A2(net_129) );
XNOR2_X2 inst_107 ( .A(net_3123), .B(net_3103), .ZN(net_428) );
INV_X8 inst_2117 ( .A(net_3520), .ZN(net_2292) );
NOR2_X2 inst_990 ( .A1(net_2641), .ZN(net_2581), .A2(net_2377) );
DFF_X2 inst_3140 ( .QN(net_2984), .D(net_2570), .CK(net_5237) );
CLKBUF_X2 inst_4710 ( .A(net_4620), .Z(net_4696) );
NAND2_X2 inst_1539 ( .A1(net_2907), .ZN(net_2483), .A2(net_172) );
INV_X2 inst_2662 ( .ZN(net_2107), .A(net_2034) );
AOI22_X2 inst_3628 ( .ZN(net_1138), .A2(net_721), .B2(net_641), .B1(net_387), .A1(net_261) );
NAND2_X2 inst_1718 ( .ZN(net_2144), .A1(net_1639), .A2(net_1638) );
NOR2_X2 inst_1050 ( .A2(net_3559), .A1(net_1228), .ZN(net_1039) );
INV_X4 inst_2366 ( .ZN(net_911), .A(net_891) );
CLKBUF_X2 inst_4642 ( .A(net_4627), .Z(net_4628) );
CLKBUF_X2 inst_5049 ( .A(net_5034), .Z(net_5035) );
DFF_X1 inst_3316 ( .QN(net_3005), .D(net_2851), .CK(net_5201) );
NAND3_X2 inst_1296 ( .ZN(net_1663), .A1(net_1584), .A2(net_1335), .A3(net_1286) );
CLKBUF_X2 inst_4661 ( .A(net_4646), .Z(net_4647) );
CLKBUF_X2 inst_4411 ( .A(net_4274), .Z(net_4397) );
NAND2_X2 inst_1852 ( .A1(net_4164), .A2(net_4116), .ZN(net_695) );
AOI22_X2 inst_3671 ( .A2(net_571), .B2(net_570), .ZN(net_553), .A1(net_552), .B1(net_551) );
DFF_X1 inst_3282 ( .QN(net_3031), .D(net_2918), .CK(net_5172) );
AOI211_X2 inst_4014 ( .ZN(net_2526), .A(net_2525), .B(net_2348), .C1(net_2303), .C2(net_207) );
CLKBUF_X2 inst_4605 ( .A(net_4590), .Z(net_4591) );
AOI22_X2 inst_3694 ( .B1(net_4124), .A2(net_509), .ZN(net_482), .B2(net_195), .A1(net_194) );
AND3_X4 inst_4074 ( .A3(net_4116), .ZN(net_4070), .A2(net_4001), .A1(net_1036) );
CLKBUF_X2 inst_4513 ( .A(net_4256), .Z(net_4499) );
AOI222_X1 inst_3783 ( .B2(net_2020), .C1(net_1840), .ZN(net_1700), .A1(net_1699), .A2(net_1698), .B1(net_673), .C2(net_142) );
NAND2_X2 inst_1557 ( .A1(net_2909), .ZN(net_2465), .A2(net_173) );
CLKBUF_X2 inst_4882 ( .A(net_4530), .Z(net_4868) );
INV_X4 inst_2399 ( .A(net_528), .ZN(net_385) );
INV_X2 inst_2698 ( .ZN(net_1683), .A(net_1682) );
NAND4_X2 inst_1237 ( .A2(net_3993), .A1(net_3713), .A4(net_3657), .ZN(net_2374), .A3(net_403) );
DFF_X1 inst_3412 ( .D(net_1354), .Q(net_37), .CK(net_4468) );
CLKBUF_X2 inst_4698 ( .A(net_4683), .Z(net_4684) );
CLKBUF_X2 inst_4452 ( .A(net_4324), .Z(net_4438) );
INV_X4 inst_2518 ( .ZN(net_3204), .A(net_3198) );
CLKBUF_X2 inst_5152 ( .A(net_4874), .Z(net_5138) );
NAND2_X2 inst_1616 ( .A1(net_2919), .ZN(net_2400), .A2(net_214) );
NAND2_X2 inst_2075 ( .ZN(net_4165), .A1(net_4164), .A2(net_3974) );
INV_X2 inst_3062 ( .ZN(net_4177), .A(net_1502) );
DFF_X1 inst_3310 ( .QN(net_3017), .D(net_2872), .CK(net_5163) );
NAND2_X2 inst_1911 ( .A2(net_3108), .ZN(net_296), .A1(net_207) );
AND2_X4 inst_4151 ( .A1(net_4118), .A2(net_4116), .ZN(net_4099) );
NAND2_X2 inst_1825 ( .A1(net_4099), .A2(net_3900), .ZN(net_899) );
OAI21_X2 inst_585 ( .B2(net_3428), .ZN(net_2702), .B1(net_2587), .A(net_2046) );
NAND2_X2 inst_1606 ( .A1(net_2967), .ZN(net_2410), .A2(net_212) );
INV_X2 inst_2851 ( .ZN(net_342), .A(net_341) );
CLKBUF_X2 inst_5100 ( .A(net_4501), .Z(net_5086) );
CLKBUF_X2 inst_5126 ( .A(net_4453), .Z(net_5112) );
OAI221_X2 inst_410 ( .A(net_3572), .C1(net_1884), .ZN(net_1549), .B1(net_1548), .B2(net_1521), .C2(net_1032) );
OAI22_X2 inst_316 ( .B1(net_3136), .ZN(net_1705), .A1(net_1123), .A2(net_1071), .B2(net_1036) );
CLKBUF_X2 inst_5107 ( .A(net_4309), .Z(net_5093) );
NOR2_X1 inst_1174 ( .ZN(net_4194), .A1(net_1212), .A2(net_743) );
NOR2_X2 inst_1023 ( .A1(net_3492), .ZN(net_1687), .A2(net_1640) );
OAI221_X2 inst_383 ( .C1(net_3875), .B2(net_2699), .C2(net_2698), .ZN(net_2629), .A(net_2535), .B1(net_2371) );
INV_X4 inst_2428 ( .A(net_3083), .ZN(net_552) );
CLKBUF_X2 inst_5115 ( .A(net_5100), .Z(net_5101) );
AND2_X4 inst_4132 ( .ZN(net_4061), .A2(net_1280), .A1(net_1085) );
DFF_X2 inst_3186 ( .QN(net_3104), .D(net_1730), .CK(net_5140) );
OAI21_X2 inst_678 ( .B1(net_3228), .B2(net_3152), .ZN(net_1509), .A(net_1307) );
NOR2_X2 inst_1124 ( .A2(net_3958), .ZN(net_3435), .A1(net_3434) );
AND3_X2 inst_4086 ( .A1(net_1517), .ZN(net_1060), .A3(net_965), .A2(net_797) );
AOI222_X1 inst_3762 ( .C1(net_3120), .A1(net_2055), .B1(net_2054), .C2(net_2053), .ZN(net_2000), .B2(net_1345), .A2(net_228) );
OAI211_X2 inst_854 ( .ZN(net_3363), .C2(net_3354), .C1(net_2190), .A(net_2008), .B(net_2001) );
DFF_X1 inst_3259 ( .QN(net_3077), .D(net_2936), .CK(net_4930) );
CLKBUF_X2 inst_4359 ( .A(net_4259), .Z(net_4345) );
INV_X4 inst_2555 ( .A(net_3653), .ZN(net_3488) );
DFF_X1 inst_3375 ( .D(net_2261), .QN(net_48), .CK(net_4513) );
OR2_X4 inst_234 ( .A1(net_3468), .ZN(net_341), .A2(net_329) );
CLKBUF_X2 inst_5293 ( .A(net_5278), .Z(net_5279) );
AOI22_X2 inst_3678 ( .B2(net_4124), .A2(net_555), .ZN(net_520), .A1(net_519), .B1(net_518) );
CLKBUF_X2 inst_5240 ( .A(net_5225), .Z(net_5226) );
AOI21_X2 inst_3979 ( .B1(net_4079), .ZN(net_1040), .A(net_986), .B2(net_528) );
NAND2_X2 inst_1946 ( .A2(net_4015), .ZN(net_3250), .A1(net_3219) );
AOI22_X2 inst_3714 ( .A2(net_3966), .B1(net_3661), .ZN(net_3434), .A1(net_1255), .B2(net_667) );
CLKBUF_X2 inst_5285 ( .A(net_5270), .Z(net_5271) );
NAND3_X2 inst_1304 ( .A3(net_1613), .A1(net_1548), .ZN(net_1315), .A2(net_857) );
DFF_X1 inst_3429 ( .Q(net_4019), .D(net_4018), .CK(net_4903) );
NAND3_X2 inst_1328 ( .A3(net_3395), .ZN(net_1024), .A2(net_666), .A1(net_539) );
OAI21_X2 inst_688 ( .A(net_1257), .B1(net_1256), .ZN(net_1184), .B2(net_819) );
NAND2_X2 inst_1749 ( .ZN(net_1372), .A1(net_1305), .A2(net_240) );
INV_X4 inst_2549 ( .ZN(net_3450), .A(net_3106) );
DFF_X1 inst_3292 ( .QN(net_3012), .D(net_2882), .CK(net_5126) );
NAND2_X2 inst_1776 ( .ZN(net_1106), .A2(net_1105), .A1(net_989) );
AOI22_X2 inst_3641 ( .A1(net_4142), .B1(net_4112), .ZN(net_761), .B2(net_379), .A2(x825) );
CLKBUF_X2 inst_4894 ( .A(net_4879), .Z(net_4880) );
CLKBUF_X2 inst_5024 ( .A(net_5009), .Z(net_5010) );
INV_X4 inst_2335 ( .ZN(net_668), .A(net_667) );
INV_X4 inst_2387 ( .ZN(net_1386), .A(net_1173) );
NOR3_X1 inst_919 ( .A1(net_3463), .A3(net_3103), .ZN(net_2745), .A2(net_2717) );
CLKBUF_X2 inst_4391 ( .A(net_4229), .Z(net_4377) );
OAI21_X2 inst_598 ( .B2(net_3127), .ZN(net_2509), .B1(net_2507), .A(net_2297) );
NAND2_X2 inst_1916 ( .ZN(net_632), .A1(net_253), .A2(net_43) );
DFF_X2 inst_3156 ( .QN(net_3130), .D(net_2183), .CK(net_5289) );
INV_X2 inst_2747 ( .A(net_1275), .ZN(net_1146) );
OAI211_X2 inst_840 ( .ZN(net_1263), .A(net_1257), .C1(net_1256), .C2(net_1117), .B(net_1062) );
NAND2_X2 inst_1624 ( .ZN(net_2615), .A1(net_2391), .A2(net_2302) );
NAND4_X2 inst_1220 ( .ZN(net_1123), .A4(net_782), .A3(net_553), .A2(net_469), .A1(net_455) );
NAND2_X4 inst_1456 ( .A1(net_3906), .ZN(net_3837), .A2(net_3836) );
INV_X4 inst_2181 ( .A(net_3230), .ZN(net_2738) );
NAND2_X2 inst_1797 ( .A1(net_2522), .ZN(net_994), .A2(net_947) );
DFF_X2 inst_3167 ( .QN(net_3164), .D(net_1974), .CK(net_4966) );
CLKBUF_X2 inst_4408 ( .A(net_4393), .Z(net_4394) );
INV_X2 inst_2708 ( .ZN(net_1751), .A(net_1648) );
CLKBUF_X2 inst_5154 ( .A(net_5139), .Z(net_5140) );
CLKBUF_X2 inst_4294 ( .A(net_4279), .Z(net_4280) );
AND2_X2 inst_4195 ( .A2(net_1946), .ZN(net_1781), .A1(net_1684) );
AOI22_X2 inst_3530 ( .B1(net_2017), .ZN(net_1894), .A1(net_1893), .A2(net_1880), .B2(net_128) );
CLKBUF_X2 inst_5009 ( .A(net_4994), .Z(net_4995) );
CLKBUF_X2 inst_4785 ( .A(net_4770), .Z(net_4771) );
CLKBUF_X2 inst_4440 ( .A(net_4425), .Z(net_4426) );
INV_X4 inst_2592 ( .ZN(net_3682), .A(net_3636) );
OAI22_X2 inst_325 ( .A1(net_4089), .B2(net_3142), .ZN(net_1642), .A2(net_931), .B1(net_433) );
CLKBUF_X2 inst_4769 ( .A(net_4402), .Z(net_4755) );
NAND4_X2 inst_1197 ( .ZN(net_1769), .A3(net_1481), .A4(net_1480), .A2(net_1415), .A1(net_1414) );
DFF_X2 inst_3116 ( .QN(net_3154), .D(net_2760), .CK(net_4684) );
CLKBUF_X2 inst_4378 ( .A(net_4363), .Z(net_4364) );
NOR2_X4 inst_955 ( .A1(net_3821), .ZN(net_3698), .A2(net_3543) );
AND2_X2 inst_4199 ( .A1(net_4061), .ZN(net_1345), .A2(net_114) );
XNOR2_X2 inst_114 ( .A(net_3153), .ZN(net_354), .B(net_332) );
INV_X4 inst_2278 ( .A(net_2596), .ZN(net_2518) );
CLKBUF_X2 inst_4866 ( .A(net_4851), .Z(net_4852) );
OAI21_X2 inst_617 ( .B2(net_3407), .ZN(net_2266), .A(net_2264), .B1(net_2263) );
AND2_X4 inst_4150 ( .ZN(net_4095), .A1(net_636), .A2(net_427) );
OAI21_X2 inst_534 ( .B1(net_3195), .B2(net_2965), .ZN(net_2899), .A(net_2446) );
CLKBUF_X2 inst_4420 ( .A(net_4405), .Z(net_4406) );
NOR2_X2 inst_1057 ( .A1(net_3838), .A2(net_3567), .ZN(net_976) );
CLKBUF_X2 inst_5191 ( .A(net_4908), .Z(net_5177) );
INV_X2 inst_2842 ( .A(net_3941), .ZN(net_391) );
CLKBUF_X2 inst_5193 ( .A(net_5178), .Z(net_5179) );
NAND2_X1 inst_2084 ( .A2(net_4019), .A1(net_2963), .ZN(net_2461) );
INV_X2 inst_2836 ( .A(net_825), .ZN(net_607) );
AOI222_X1 inst_3792 ( .ZN(net_3323), .A2(net_3319), .B2(net_826), .C2(net_825), .A1(net_724), .B1(net_618), .C1(net_528) );
CLKBUF_X2 inst_4336 ( .A(net_4321), .Z(net_4322) );
OAI21_X2 inst_748 ( .B2(net_4195), .ZN(net_3375), .A(net_3374), .B1(net_818) );
INV_X2 inst_2839 ( .A(net_3468), .ZN(net_402) );
CLKBUF_X2 inst_4582 ( .A(net_4567), .Z(net_4568) );
INV_X2 inst_2770 ( .ZN(net_886), .A(net_885) );
CLKBUF_X2 inst_4573 ( .A(net_4558), .Z(net_4559) );
CLKBUF_X2 inst_4526 ( .A(net_4511), .Z(net_4512) );
OAI211_X2 inst_803 ( .C1(net_2190), .ZN(net_2132), .C2(net_2131), .A(net_2011), .B(net_2002) );
CLKBUF_X2 inst_4587 ( .A(net_4572), .Z(net_4573) );
NAND2_X2 inst_1986 ( .A2(net_4142), .ZN(net_3428), .A1(net_3427) );
INV_X2 inst_2909 ( .ZN(net_206), .A(net_82) );
CLKBUF_X2 inst_4732 ( .A(net_4465), .Z(net_4718) );
NAND2_X2 inst_1949 ( .A2(net_3281), .ZN(net_3265), .A1(net_147) );
INV_X4 inst_2348 ( .A(net_707), .ZN(net_589) );
DFF_X2 inst_3135 ( .QN(net_2987), .D(net_2571), .CK(net_5156) );
AOI211_X2 inst_4021 ( .ZN(net_1371), .C2(net_1228), .B(net_1194), .A(net_1130), .C1(net_949) );
OAI21_X2 inst_701 ( .A(net_3925), .B2(net_3478), .ZN(net_1116), .B1(net_699) );
OAI21_X2 inst_662 ( .B1(net_4100), .ZN(net_1841), .B2(net_1701), .A(net_1591) );
INV_X2 inst_2911 ( .ZN(net_2286), .A(net_69) );
NAND2_X2 inst_1533 ( .A1(net_3208), .ZN(net_2489), .A2(net_235) );
INV_X4 inst_2380 ( .A(net_3633), .ZN(net_432) );
AOI22_X2 inst_3495 ( .B2(net_3818), .A1(net_2231), .B1(net_2230), .ZN(net_2224), .A2(net_74) );
CLKBUF_X2 inst_5261 ( .A(net_5246), .Z(net_5247) );
NAND2_X2 inst_1859 ( .A2(net_3440), .A1(net_923), .ZN(net_608) );
CLKBUF_X2 inst_5080 ( .A(net_5065), .Z(net_5066) );
CLKBUF_X2 inst_4666 ( .A(net_4651), .Z(net_4652) );
NAND2_X4 inst_1465 ( .ZN(net_3886), .A1(net_2292), .A2(net_2210) );
CLKBUF_X2 inst_5030 ( .A(net_5015), .Z(net_5016) );
XNOR2_X2 inst_53 ( .A(net_3876), .B(net_3515), .ZN(net_2811) );
CLKBUF_X2 inst_5265 ( .A(net_5250), .Z(net_5251) );
NOR2_X2 inst_1007 ( .ZN(net_2202), .A1(net_1790), .A2(net_1734) );
INV_X2 inst_2815 ( .A(net_3755), .ZN(net_1045) );
AND2_X2 inst_4208 ( .ZN(net_3501), .A1(net_1187), .A2(net_741) );
AOI22_X2 inst_3605 ( .A1(net_4063), .B1(net_4058), .ZN(net_1412), .A2(net_552), .B2(net_551) );
INV_X4 inst_2614 ( .ZN(net_3842), .A(net_3834) );
DFF_X1 inst_3337 ( .Q(net_3141), .D(net_2789), .CK(net_4771) );
CLKBUF_X2 inst_5066 ( .A(net_5051), .Z(net_5052) );
CLKBUF_X2 inst_4215 ( .A(net_4200), .Z(net_4201) );
OAI21_X2 inst_651 ( .B2(net_3492), .ZN(net_2598), .A(net_2548), .B1(net_1741) );
AND3_X2 inst_4090 ( .ZN(net_3467), .A3(net_3466), .A1(net_2129), .A2(net_2126) );
NOR2_X2 inst_999 ( .A2(net_4049), .ZN(net_2152), .A1(net_2120) );
MUX2_X2 inst_2111 ( .A(net_1774), .Z(net_1403), .S(net_1228), .B(net_321) );
INV_X2 inst_2883 ( .A(net_987), .ZN(net_387) );
NOR2_X2 inst_1157 ( .ZN(net_4081), .A1(net_765), .A2(net_371) );
NAND2_X2 inst_1846 ( .ZN(net_742), .A1(net_613), .A2(net_414) );
INV_X8 inst_2139 ( .A(net_3177), .ZN(net_3176) );
CLKBUF_X2 inst_4278 ( .A(net_4263), .Z(net_4264) );
NAND2_X4 inst_1463 ( .A1(net_3911), .ZN(net_3883), .A2(net_3303) );
OR3_X2 inst_186 ( .ZN(net_3351), .A2(net_3348), .A1(net_2550), .A3(net_1737) );
CLKBUF_X2 inst_4271 ( .A(net_4256), .Z(net_4257) );
AOI22_X2 inst_3528 ( .A2(net_3145), .A1(net_1923), .B1(net_1921), .ZN(net_1916), .B2(net_686) );
OAI21_X2 inst_759 ( .ZN(net_3741), .A(net_3740), .B1(net_2876), .B2(net_67) );
INV_X1 inst_3071 ( .A(net_3691), .ZN(net_2506) );
NAND2_X2 inst_2061 ( .ZN(net_3918), .A1(net_3653), .A2(net_3107) );
AOI22_X2 inst_3685 ( .B2(net_4123), .A2(net_509), .ZN(net_496), .A1(net_495), .B1(net_189) );
CLKBUF_X2 inst_4255 ( .A(net_4240), .Z(net_4241) );
NOR4_X2 inst_863 ( .ZN(net_1515), .A2(net_1262), .A1(net_1260), .A4(net_1248), .A3(net_1145) );
NAND2_X4 inst_1472 ( .A2(net_4003), .A1(net_3992), .ZN(net_3922) );
CLKBUF_X2 inst_4261 ( .A(net_4203), .Z(net_4247) );
NAND2_X4 inst_1385 ( .ZN(net_2878), .A1(net_2831), .A2(net_2808) );
NAND2_X2 inst_1573 ( .A1(net_2915), .ZN(net_2448), .A2(net_153) );
NAND4_X2 inst_1183 ( .A4(net_3650), .A3(net_3192), .ZN(net_2207), .A2(net_2089), .A1(net_2080) );
AOI222_X1 inst_3784 ( .B1(net_2020), .C1(net_1840), .A1(net_1698), .ZN(net_1680), .B2(net_324), .A2(net_251), .C2(net_228) );
NAND2_X4 inst_1390 ( .A1(net_3188), .A2(net_3180), .ZN(net_2178) );
AOI22_X2 inst_3586 ( .A1(net_4062), .B1(net_4057), .ZN(net_1431), .A2(net_230), .B2(net_148) );
OR2_X4 inst_229 ( .ZN(net_988), .A2(net_516), .A1(net_384) );
INV_X4 inst_2282 ( .ZN(net_1202), .A(net_959) );
NAND2_X2 inst_1489 ( .ZN(net_2861), .A1(net_2852), .A2(net_2516) );
CLKBUF_X2 inst_5272 ( .A(net_5257), .Z(net_5258) );
CLKBUF_X2 inst_4992 ( .A(net_4977), .Z(net_4978) );
INV_X4 inst_2415 ( .A(net_3122), .ZN(net_1523) );
CLKBUF_X2 inst_4689 ( .A(net_4674), .Z(net_4675) );
INV_X4 inst_2262 ( .ZN(net_1166), .A(net_1095) );
DFF_X1 inst_3288 ( .QN(net_3047), .D(net_2900), .CK(net_4772) );
CLKBUF_X2 inst_4981 ( .A(net_4242), .Z(net_4967) );
NOR2_X2 inst_1160 ( .ZN(net_4113), .A1(net_1326), .A2(net_449) );
NAND2_X4 inst_1394 ( .A1(net_3219), .ZN(net_1984), .A2(net_176) );
INV_X8 inst_2131 ( .A(net_3642), .ZN(net_357) );
NAND2_X2 inst_1808 ( .A1(net_4082), .ZN(net_1332), .A2(net_911) );
NOR2_X2 inst_988 ( .ZN(net_2355), .A1(net_2301), .A2(net_1090) );
NAND2_X2 inst_1876 ( .ZN(net_450), .A1(net_411), .A2(net_390) );
OR3_X4 inst_169 ( .ZN(net_1701), .A1(net_1232), .A3(net_1173), .A2(net_947) );
OAI221_X2 inst_421 ( .C1(net_3560), .ZN(net_1194), .A(net_1057), .B1(net_964), .B2(net_877), .C2(net_408) );
CLKBUF_X2 inst_4954 ( .A(net_4939), .Z(net_4940) );
NAND3_X2 inst_1315 ( .A1(net_4087), .ZN(net_974), .A3(net_619), .A2(x475) );
CLKBUF_X2 inst_5035 ( .A(net_4325), .Z(net_5021) );
OAI21_X2 inst_555 ( .B2(net_2917), .B1(net_2871), .ZN(net_2870), .A(net_2420) );
CLKBUF_X2 inst_4759 ( .A(net_4744), .Z(net_4745) );
OAI211_X2 inst_816 ( .C2(net_3319), .B(net_1628), .C1(net_1627), .ZN(net_1622), .A(net_1558) );
INV_X4 inst_2392 ( .A(net_3324), .ZN(net_416) );
CLKBUF_X2 inst_4308 ( .A(net_4235), .Z(net_4294) );
CLKBUF_X2 inst_4678 ( .A(net_4581), .Z(net_4664) );
INV_X2 inst_2798 ( .ZN(net_1655), .A(net_869) );
AOI22_X2 inst_3667 ( .A1(net_571), .B1(net_570), .ZN(net_560), .A2(net_559), .B2(net_558) );
NAND4_X2 inst_1184 ( .ZN(net_2179), .A1(net_2004), .A4(net_1971), .A2(net_1925), .A3(net_1915) );
CLKBUF_X2 inst_4434 ( .A(net_4419), .Z(net_4420) );
CLKBUF_X2 inst_4685 ( .A(net_4670), .Z(net_4671) );
CLKBUF_X2 inst_4967 ( .A(net_4952), .Z(net_4953) );
OAI21_X2 inst_656 ( .B2(net_2150), .ZN(net_1929), .B1(net_1815), .A(net_1803) );
XNOR2_X2 inst_45 ( .ZN(net_2813), .A(net_2600), .B(net_1786) );
NOR2_X2 inst_1108 ( .A1(net_3808), .ZN(net_3291), .A2(net_2344) );
CLKBUF_X2 inst_5148 ( .A(net_5133), .Z(net_5134) );
CLKBUF_X2 inst_5140 ( .A(net_5125), .Z(net_5126) );
OAI21_X4 inst_458 ( .B2(net_4051), .ZN(net_3254), .A(net_3253), .B1(net_1162) );
HA_X1 inst_3093 ( .S(net_1163), .CO(net_1162), .A(net_1161), .B(net_1160) );
NAND2_X2 inst_1562 ( .A1(net_2963), .ZN(net_2459), .A2(net_474) );
AND2_X4 inst_4148 ( .ZN(net_4086), .A2(net_2374), .A1(net_711) );
CLKBUF_X2 inst_4618 ( .A(net_4282), .Z(net_4604) );
CLKBUF_X2 inst_4534 ( .A(net_4495), .Z(net_4520) );
NAND2_X2 inst_1922 ( .A1(net_3817), .ZN(net_3180), .A2(net_174) );
DFF_X1 inst_3361 ( .D(net_2359), .CK(net_4400), .Q(x450) );
OAI21_X2 inst_741 ( .ZN(net_3279), .B1(net_3278), .B2(net_2915), .A(net_2435) );
DFF_X2 inst_3170 ( .Q(net_3160), .D(net_1914), .CK(net_4998) );
DFF_X1 inst_3232 ( .QN(net_3064), .D(net_2964), .CK(net_4873) );
AOI21_X2 inst_3991 ( .B1(net_4190), .B2(net_3600), .ZN(net_3195), .A(net_1948) );
DFF_X1 inst_3343 ( .D(net_2780), .CK(net_4352), .Q(x128) );
NAND3_X2 inst_1350 ( .A3(net_3762), .ZN(net_3638), .A1(net_3637), .A2(net_3452) );
AND2_X4 inst_4140 ( .ZN(net_4072), .A1(net_1131), .A2(net_432) );
INV_X2 inst_3012 ( .ZN(net_3385), .A(net_42) );
INV_X2 inst_2635 ( .A(net_2601), .ZN(net_2520) );
NAND2_X2 inst_1543 ( .A1(net_3207), .ZN(net_2479), .A2(net_154) );
INV_X2 inst_2828 ( .A(net_3702), .ZN(net_441) );
CLKBUF_X2 inst_4219 ( .A(net_4202), .Z(net_4205) );
INV_X2 inst_2801 ( .ZN(net_1314), .A(net_742) );
NOR2_X2 inst_1118 ( .ZN(net_3422), .A2(net_3421), .A1(net_3415) );
INV_X4 inst_2303 ( .A(net_1028), .ZN(net_852) );
CLKBUF_X2 inst_4745 ( .A(net_4730), .Z(net_4731) );
DFF_X1 inst_3363 ( .D(net_2363), .CK(net_4227), .Q(x368) );
AOI221_X2 inst_3877 ( .B1(net_2020), .C1(net_2019), .ZN(net_1857), .A(net_1856), .B2(net_1699), .C2(x388) );
INV_X2 inst_2666 ( .A(net_2230), .ZN(net_2155) );
OAI21_X2 inst_473 ( .B1(net_3509), .ZN(net_2977), .B2(net_2963), .A(net_2459) );
NOR2_X2 inst_1131 ( .ZN(net_3578), .A1(net_3577), .A2(net_2373) );
NAND3_X2 inst_1357 ( .ZN(net_3716), .A2(net_3715), .A1(net_3682), .A3(net_87) );
OAI21_X2 inst_691 ( .A(net_1650), .ZN(net_1049), .B1(net_1006), .B2(net_608) );
INV_X4 inst_2211 ( .A(net_3241), .ZN(net_2732) );
AOI222_X1 inst_3771 ( .A1(net_4065), .C1(net_1882), .ZN(net_1873), .A2(net_1662), .B1(net_1385), .B2(net_941), .C2(net_635) );
INV_X1 inst_3083 ( .A(net_3938), .ZN(net_3639) );
NAND2_X2 inst_1695 ( .A1(net_2264), .ZN(net_2137), .A2(net_1993) );
OAI21_X2 inst_770 ( .ZN(net_4182), .B2(net_4181), .B1(net_3260), .A(net_3259) );
OAI21_X2 inst_565 ( .B2(net_2915), .B1(net_2849), .ZN(net_2847), .A(net_2439) );
CLKBUF_X2 inst_5302 ( .A(net_4594), .Z(net_5288) );
OAI21_X2 inst_622 ( .B1(net_2235), .ZN(net_2159), .A(net_2048), .B2(net_108) );
NAND2_X2 inst_1971 ( .A2(net_3877), .ZN(net_3341), .A1(net_3340) );
NAND2_X4 inst_1404 ( .A2(net_4021), .ZN(net_3234), .A1(net_3185) );
CLKBUF_X2 inst_4476 ( .A(net_4301), .Z(net_4462) );
INV_X2 inst_2989 ( .A(net_3100), .ZN(net_190) );
AOI22_X2 inst_3479 ( .A1(net_3241), .B2(net_3112), .B1(net_2781), .ZN(net_2660), .A2(net_2659) );
OAI221_X2 inst_409 ( .ZN(net_2594), .B1(net_1614), .C1(net_1613), .A(net_1530), .B2(net_289), .C2(net_250) );
INV_X4 inst_2288 ( .ZN(net_1125), .A(net_884) );
NAND3_X2 inst_1339 ( .ZN(net_3361), .A2(net_3360), .A1(net_3359), .A3(net_1574) );
CLKBUF_X2 inst_4284 ( .A(net_4216), .Z(net_4270) );
CLKBUF_X2 inst_4971 ( .A(net_4956), .Z(net_4957) );
CLKBUF_X2 inst_4704 ( .A(net_4613), .Z(net_4690) );
CLKBUF_X2 inst_4724 ( .A(net_4709), .Z(net_4710) );
CLKBUF_X2 inst_4841 ( .A(net_4826), .Z(net_4827) );
NAND2_X2 inst_1834 ( .A1(net_4105), .ZN(net_842), .A2(net_513) );
CLKBUF_X2 inst_4467 ( .A(net_4391), .Z(net_4453) );
AOI22_X2 inst_3575 ( .A1(net_4059), .B1(net_4056), .ZN(net_1475), .B2(net_498), .A2(net_497) );
CLKBUF_X2 inst_4493 ( .A(net_4474), .Z(net_4479) );
AOI22_X2 inst_3506 ( .B1(net_3676), .B2(net_3143), .A1(net_2012), .ZN(net_2011), .A2(net_168) );
AOI22_X2 inst_3654 ( .B2(net_4011), .A2(net_4009), .ZN(net_654), .A1(net_458), .B1(net_457) );
NOR2_X4 inst_977 ( .A1(net_3939), .ZN(net_3936), .A2(net_281) );
INV_X4 inst_2228 ( .A(net_1893), .ZN(net_1789) );
AOI22_X2 inst_3574 ( .A1(net_4060), .B1(net_4055), .ZN(net_1476), .B2(net_183), .A2(net_172) );
OAI21_X2 inst_768 ( .B2(net_4131), .B1(net_4086), .ZN(net_3963), .A(net_3960) );
OAI21_X2 inst_663 ( .A(net_3229), .ZN(net_2691), .B1(net_1559), .B2(net_69) );
INV_X8 inst_2121 ( .ZN(net_877), .A(net_432) );
CLKBUF_X2 inst_4802 ( .A(net_4787), .Z(net_4788) );
CLKBUF_X2 inst_4850 ( .A(net_4583), .Z(net_4836) );
OAI22_X2 inst_297 ( .A1(net_3487), .ZN(net_1738), .B1(net_1637), .B2(net_612), .A2(net_287) );
DFF_X1 inst_3227 ( .QN(net_3067), .D(net_2966), .CK(net_4887) );
NAND2_X4 inst_1395 ( .A2(net_3869), .A1(net_3868), .ZN(net_1865) );
INV_X4 inst_2477 ( .A(net_3063), .ZN(net_519) );
CLKBUF_X2 inst_4838 ( .A(net_4516), .Z(net_4824) );
INV_X4 inst_2188 ( .ZN(net_2612), .A(net_2524) );
AOI22_X2 inst_3494 ( .B2(net_3543), .ZN(net_2232), .A1(net_2231), .B1(net_2230), .A2(net_76) );
CLKBUF_X2 inst_4224 ( .A(net_4205), .Z(net_4210) );
NAND2_X2 inst_1875 ( .A1(net_3619), .ZN(net_947), .A2(net_299) );
DFF_X1 inst_3351 ( .D(net_2701), .QN(net_65), .CK(net_4239) );
NAND2_X2 inst_1867 ( .A1(net_3713), .ZN(net_849), .A2(net_543) );
DFF_X2 inst_3190 ( .QN(net_3156), .D(net_1704), .CK(net_4989) );
OR3_X4 inst_162 ( .ZN(net_2778), .A1(net_2325), .A2(net_2206), .A3(net_1173) );
DFF_X1 inst_3308 ( .QN(net_3015), .D(net_2870), .CK(net_5168) );
INV_X4 inst_2290 ( .A(net_938), .ZN(net_937) );
DFF_X1 inst_3397 ( .D(net_1563), .CK(net_5252), .Q(x606) );
CLKBUF_X2 inst_4421 ( .A(net_4406), .Z(net_4407) );
INV_X2 inst_2829 ( .ZN(net_601), .A(net_424) );
AOI221_X2 inst_3819 ( .A(net_2642), .B1(net_2641), .C1(net_2581), .ZN(net_2559), .C2(net_2551), .B2(net_252) );
CLKBUF_X2 inst_4233 ( .A(net_4218), .Z(net_4219) );
AOI22_X2 inst_3668 ( .B2(net_3455), .A1(net_571), .B1(net_570), .ZN(net_557), .A2(net_201) );
CLKBUF_X2 inst_5070 ( .A(net_4474), .Z(net_5056) );
CLKBUF_X2 inst_4912 ( .A(net_4897), .Z(net_4898) );
AOI21_X2 inst_3968 ( .ZN(net_1370), .A(net_1315), .B1(net_1314), .B2(net_517) );
DFF_X1 inst_3342 ( .Q(net_3143), .D(net_2769), .CK(net_4599) );
CLKBUF_X2 inst_4825 ( .A(net_4810), .Z(net_4811) );
CLKBUF_X2 inst_4633 ( .A(net_4618), .Z(net_4619) );
NOR2_X2 inst_1098 ( .A2(net_3162), .ZN(net_350), .A1(net_223) );
INV_X4 inst_2621 ( .ZN(net_3940), .A(net_3109) );
AND2_X4 inst_4149 ( .A1(net_4186), .ZN(net_4087), .A2(net_3521) );
AOI221_X2 inst_3895 ( .C2(net_1394), .B1(net_1393), .ZN(net_1347), .A(net_1173), .B2(net_207), .C1(net_51) );
INV_X4 inst_2443 ( .A(net_3088), .ZN(net_497) );
OAI21_X2 inst_723 ( .B2(net_3619), .ZN(net_647), .B1(net_641), .A(net_537) );
OAI22_X2 inst_303 ( .A1(net_1543), .B1(net_1542), .ZN(net_1539), .A2(net_292), .B2(net_131) );
OAI21_X2 inst_618 ( .B2(net_3408), .ZN(net_2265), .A(net_2264), .B1(net_2263) );
INV_X4 inst_2444 ( .A(net_3086), .ZN(net_461) );
AOI221_X2 inst_3893 ( .C2(net_4029), .C1(net_1394), .B1(net_1393), .ZN(net_1350), .A(net_1173), .B2(net_686) );
NAND2_X2 inst_1647 ( .A1(net_3774), .ZN(net_2328), .A2(net_1888) );
DFF_X1 inst_3263 ( .QN(net_3073), .D(net_2935), .CK(net_4867) );
INV_X2 inst_3057 ( .ZN(net_3952), .A(net_3948) );
NAND3_X2 inst_1275 ( .ZN(net_2764), .A1(net_2738), .A2(net_2737), .A3(net_1826) );
INV_X4 inst_2462 ( .A(net_3085), .ZN(net_781) );
OAI21_X2 inst_474 ( .B1(net_3509), .ZN(net_2976), .B2(net_2961), .A(net_2474) );
XOR2_X1 inst_26 ( .Z(net_1910), .A(net_1875), .B(net_1874) );
NAND2_X2 inst_2067 ( .ZN(net_3965), .A2(net_3960), .A1(net_930) );
OAI21_X2 inst_626 ( .B1(net_2190), .ZN(net_2151), .B2(net_2150), .A(net_2036) );
NAND3_X1 inst_1376 ( .A3(net_2691), .ZN(net_2648), .A1(net_2647), .A2(net_2506) );
INV_X2 inst_2882 ( .ZN(net_240), .A(net_61) );
INV_X2 inst_2777 ( .A(net_3907), .ZN(net_811) );
CLKBUF_X2 inst_4864 ( .A(net_4831), .Z(net_4850) );
INV_X4 inst_2446 ( .A(net_3065), .ZN(net_479) );
CLKBUF_X2 inst_5046 ( .A(net_5031), .Z(net_5032) );
AOI222_X1 inst_3765 ( .B1(net_4048), .C1(net_3447), .A1(net_1968), .ZN(net_1967), .C2(net_333), .A2(net_300), .B2(net_68) );
NAND2_X2 inst_1659 ( .ZN(net_2104), .A1(net_1982), .A2(net_196) );
CLKBUF_X2 inst_4218 ( .A(net_4203), .Z(net_4204) );
OAI211_X2 inst_798 ( .ZN(net_2191), .C1(net_2190), .C2(net_2189), .B(net_2052), .A(net_2007) );
CLKBUF_X2 inst_5210 ( .A(net_5195), .Z(net_5196) );
OAI221_X2 inst_398 ( .C2(net_3407), .B1(net_2328), .ZN(net_2287), .B2(net_2286), .C1(net_2239), .A(net_1938) );
CLKBUF_X2 inst_4340 ( .A(net_4325), .Z(net_4326) );
OAI221_X2 inst_436 ( .C2(net_3103), .A(net_629), .B1(net_628), .C1(net_627), .ZN(net_623), .B2(net_261) );
NAND2_X4 inst_1434 ( .ZN(net_3672), .A1(net_3671), .A2(net_3636) );
NAND2_X2 inst_1886 ( .A2(net_3418), .ZN(net_587), .A1(net_365) );
AOI22_X2 inst_3705 ( .B2(net_4123), .A2(net_555), .ZN(net_463), .A1(net_462), .B1(net_461) );
CLKBUF_X2 inst_5053 ( .A(net_5038), .Z(net_5039) );
INV_X4 inst_2231 ( .ZN(net_1872), .A(net_1666) );
CLKBUF_X2 inst_4349 ( .A(net_4239), .Z(net_4335) );
SDFF_X2 inst_144 ( .D(net_3886), .SE(net_2625), .SI(net_90), .Q(net_90), .CK(net_4951) );
NAND2_X4 inst_1457 ( .ZN(net_3838), .A2(net_3836), .A1(net_3637) );
NAND2_X4 inst_1438 ( .A1(net_3891), .ZN(net_3711), .A2(net_3700) );
NAND2_X2 inst_1818 ( .A2(net_3627), .A1(net_1463), .ZN(net_1338) );
AOI22_X2 inst_3662 ( .A1(net_571), .B1(net_570), .ZN(net_565), .B2(net_176), .A2(net_163) );
NAND2_X2 inst_1766 ( .A2(net_4032), .A1(net_1394), .ZN(net_1233) );
INV_X2 inst_2670 ( .ZN(net_2638), .A(net_2563) );
NOR3_X4 inst_880 ( .A3(net_3822), .ZN(net_3790), .A1(net_3785), .A2(net_357) );
CLKBUF_X2 inst_4857 ( .A(net_4842), .Z(net_4843) );
INV_X2 inst_2974 ( .ZN(net_1189), .A(net_119) );
NAND2_X2 inst_1895 ( .A1(net_4128), .ZN(net_367), .A2(net_144) );
INV_X2 inst_2681 ( .ZN(net_1853), .A(net_1852) );
INV_X2 inst_2730 ( .ZN(net_1398), .A(net_1350) );
CLKBUF_X2 inst_4548 ( .A(net_4281), .Z(net_4534) );
OAI21_X2 inst_737 ( .ZN(net_445), .B2(net_343), .B1(net_248), .A(x639) );
CLKBUF_X2 inst_4447 ( .A(net_4432), .Z(net_4433) );
NOR3_X4 inst_876 ( .ZN(net_2599), .A1(net_2549), .A2(net_2547), .A3(net_1706) );
INV_X2 inst_2979 ( .A(net_3021), .ZN(net_199) );
CLKBUF_X2 inst_4727 ( .A(net_4343), .Z(net_4713) );
OAI21_X2 inst_545 ( .B2(net_2917), .B1(net_2887), .ZN(net_2886), .A(net_2395) );
AOI21_X2 inst_3972 ( .ZN(net_1231), .A(net_1093), .B1(net_704), .B2(net_323) );
NAND2_X4 inst_1388 ( .ZN(net_2787), .A1(net_2740), .A2(net_2373) );
INV_X4 inst_2433 ( .ZN(net_396), .A(net_316) );
INV_X2 inst_2699 ( .A(net_3321), .ZN(net_1783) );
AOI22_X2 inst_3517 ( .B1(net_4045), .A1(net_1955), .ZN(net_1953), .A2(net_287), .B2(net_142) );
OAI21_X2 inst_562 ( .B2(net_2925), .ZN(net_2851), .B1(net_2849), .A(net_2425) );
INV_X4 inst_2480 ( .ZN(net_393), .A(net_41) );
NAND3_X2 inst_1372 ( .ZN(net_4174), .A3(net_4173), .A2(net_4171), .A1(net_4167) );
DFF_X1 inst_3396 ( .Q(net_3116), .D(net_1533), .CK(net_4309) );
NAND3_X2 inst_1360 ( .A3(net_3881), .ZN(net_3829), .A2(net_3828), .A1(net_3618) );
OAI21_X4 inst_466 ( .A(net_3858), .ZN(net_3848), .B2(net_3847), .B1(net_3846) );
INV_X2 inst_2761 ( .ZN(net_1153), .A(net_1033) );
AOI21_X2 inst_3981 ( .A(net_3916), .ZN(net_980), .B1(net_646), .B2(net_523) );
CLKBUF_X2 inst_4953 ( .A(net_4301), .Z(net_4939) );
NOR2_X2 inst_989 ( .A1(net_2591), .ZN(net_2589), .A2(net_2247) );
CLKBUF_X2 inst_5205 ( .A(net_5190), .Z(net_5191) );
INV_X4 inst_2283 ( .A(net_1250), .ZN(net_1246) );
INV_X2 inst_3038 ( .ZN(net_3632), .A(net_3630) );
NOR4_X2 inst_858 ( .A4(net_3796), .ZN(net_2274), .A1(net_2192), .A2(net_1659), .A3(net_1312) );
AOI22_X2 inst_3659 ( .ZN(net_572), .A1(net_571), .B1(net_570), .B2(net_171), .A2(net_146) );
AOI22_X2 inst_3604 ( .A1(net_4062), .B1(net_4057), .ZN(net_1413), .B2(net_467), .A2(net_454) );
NOR2_X2 inst_1109 ( .A2(net_3874), .ZN(net_3303), .A1(net_2209) );
AOI221_X2 inst_3864 ( .B1(net_4048), .C2(net_3147), .B2(net_2623), .ZN(net_1971), .C1(net_1923), .A(net_1831) );
CLKBUF_X2 inst_4415 ( .A(net_4333), .Z(net_4401) );
AND2_X2 inst_4209 ( .ZN(net_3972), .A1(net_3967), .A2(net_3478) );
INV_X2 inst_3037 ( .A(net_3973), .ZN(net_3621) );
XNOR2_X2 inst_54 ( .A(net_2543), .ZN(net_2382), .B(net_2342) );
INV_X4 inst_2468 ( .A(net_3077), .ZN(net_738) );
INV_X2 inst_2936 ( .A(net_3166), .ZN(net_344) );
NAND3_X2 inst_1314 ( .A2(net_4108), .ZN(net_894), .A3(net_829), .A1(net_783) );
NAND2_X4 inst_1420 ( .A1(net_3788), .ZN(net_3569), .A2(net_3521) );
NAND2_X4 inst_1482 ( .ZN(net_3976), .A2(net_3975), .A1(net_3679) );
CLKBUF_X2 inst_4260 ( .A(net_4245), .Z(net_4246) );
NOR2_X2 inst_1156 ( .ZN(net_4058), .A2(net_3339), .A1(net_1191) );
DFF_X1 inst_3378 ( .D(net_2252), .Q(net_74), .CK(net_5299) );
CLKBUF_X2 inst_5214 ( .A(net_5007), .Z(net_5200) );
AOI22_X2 inst_3484 ( .B2(net_3385), .A1(net_2675), .B1(net_2657), .ZN(net_2653), .A2(net_361) );
AND3_X4 inst_4062 ( .A3(net_3802), .ZN(net_1923), .A1(net_1827), .A2(net_1783) );
NOR2_X4 inst_942 ( .ZN(net_3289), .A2(net_3285), .A1(net_2174) );
CLKBUF_X2 inst_4626 ( .A(net_4611), .Z(net_4612) );
AND2_X4 inst_4108 ( .ZN(net_3590), .A2(net_3106), .A1(net_283) );
NAND3_X2 inst_1295 ( .A2(net_2054), .ZN(net_1889), .A1(net_1888), .A3(net_514) );
NAND2_X2 inst_1880 ( .ZN(net_881), .A1(net_398), .A2(net_368) );
CLKBUF_X2 inst_4794 ( .A(net_4779), .Z(net_4780) );
OR2_X2 inst_262 ( .A1(net_663), .A2(net_632), .ZN(net_631) );
AOI221_X2 inst_3829 ( .B1(net_4189), .C1(net_2534), .ZN(net_2370), .A(net_2291), .C2(net_256), .B2(net_168) );
AOI22_X2 inst_3630 ( .B1(net_4114), .A2(net_1094), .A1(net_963), .ZN(net_887), .B2(net_838) );
CLKBUF_X2 inst_4675 ( .A(net_4660), .Z(net_4661) );
OAI21_X2 inst_497 ( .B1(net_3394), .B2(net_2963), .ZN(net_2945), .A(net_2456) );
CLKBUF_X2 inst_4501 ( .A(net_4238), .Z(net_4487) );
INV_X4 inst_2195 ( .ZN(net_2389), .A(net_2327) );
CLKBUF_X2 inst_4252 ( .A(net_4237), .Z(net_4238) );
NOR2_X2 inst_1035 ( .A2(net_4080), .A1(net_1774), .ZN(net_1367) );
INV_X8 inst_2168 ( .ZN(net_3950), .A(net_3949) );
NAND3_X2 inst_1335 ( .A3(net_1401), .ZN(net_405), .A2(net_371), .A1(net_344) );
AOI221_X2 inst_3845 ( .B2(net_2203), .C1(net_2202), .ZN(net_2197), .B1(net_2196), .A(net_2077), .C2(net_396) );
AOI22_X2 inst_3637 ( .ZN(net_835), .A1(net_834), .B1(net_833), .A2(net_458), .B2(net_457) );
CLKBUF_X2 inst_5168 ( .A(net_4492), .Z(net_5154) );
DFF_X2 inst_3128 ( .QN(net_3148), .D(net_2683), .CK(net_4570) );
NAND2_X2 inst_1883 ( .ZN(net_1217), .A2(net_412), .A1(net_164) );
CLKBUF_X2 inst_4322 ( .A(net_4307), .Z(net_4308) );
NOR2_X2 inst_1078 ( .A2(net_4004), .ZN(net_644), .A1(net_618) );
INV_X4 inst_2517 ( .A(net_3543), .ZN(net_3196) );
AOI22_X2 inst_3621 ( .A1(net_1246), .A2(net_1137), .ZN(net_1119), .B1(net_1118), .B2(net_1117) );
NOR4_X2 inst_864 ( .A1(net_4064), .A2(net_1518), .ZN(net_1320), .A3(net_1319), .A4(net_793) );
OAI221_X2 inst_418 ( .C1(net_1332), .ZN(net_1251), .B1(net_1250), .B2(net_1138), .A(net_1128), .C2(net_646) );
XNOR2_X2 inst_86 ( .B(net_4073), .ZN(net_1075), .A(net_916) );
AND2_X4 inst_4183 ( .ZN(net_4145), .A1(net_3967), .A2(net_3620) );
NOR2_X4 inst_949 ( .A1(net_3701), .ZN(net_3617), .A2(net_3616) );
DFF_X1 inst_3283 ( .QN(net_3053), .D(net_2902), .CK(net_4780) );
AOI22_X2 inst_3557 ( .A1(net_4059), .B1(net_4056), .ZN(net_1493), .A2(net_236), .B2(net_151) );
NOR2_X2 inst_1039 ( .A1(net_1521), .A2(net_1170), .ZN(net_1169) );
NAND2_X2 inst_1992 ( .ZN(net_3458), .A2(net_2329), .A1(net_2321) );
AOI21_X2 inst_3961 ( .B1(net_4067), .ZN(net_1501), .A(net_1302), .B2(net_1298) );
OAI21_X2 inst_714 ( .B2(net_3789), .A(net_3733), .B1(net_810), .ZN(net_809) );
AOI22_X2 inst_3730 ( .ZN(net_4179), .B2(net_1523), .B1(net_623), .A1(net_575), .A2(net_261) );
INV_X2 inst_2895 ( .A(net_3098), .ZN(net_235) );
INV_X2 inst_3005 ( .ZN(net_3239), .A(net_764) );
AOI22_X2 inst_3598 ( .A1(net_4062), .B1(net_4057), .ZN(net_1419), .A2(net_203), .B2(net_173) );
AND4_X4 inst_4048 ( .ZN(net_4088), .A1(net_595), .A4(net_564), .A2(net_485), .A3(net_464) );
NAND2_X2 inst_1826 ( .A1(net_947), .ZN(net_786), .A2(net_671) );
MUX2_X2 inst_2109 ( .S(net_2907), .A(net_2573), .Z(net_2568), .B(net_197) );
AOI21_X2 inst_4003 ( .ZN(net_3752), .B2(net_3745), .A(net_3229), .B1(net_2623) );
NAND2_X2 inst_2020 ( .A2(net_3767), .A1(net_3766), .ZN(net_3670) );
CLKBUF_X2 inst_5033 ( .A(net_4249), .Z(net_5019) );
NOR2_X2 inst_1061 ( .ZN(net_939), .A1(net_938), .A2(net_399) );
CLKBUF_X2 inst_4361 ( .A(net_4346), .Z(net_4347) );
NAND4_X4 inst_1177 ( .ZN(net_3887), .A4(net_3886), .A3(net_3885), .A2(net_3884), .A1(net_3883) );
INV_X4 inst_2326 ( .ZN(net_957), .A(net_699) );
INV_X2 inst_2820 ( .ZN(net_717), .A(net_530) );
INV_X4 inst_2548 ( .ZN(net_3449), .A(net_3445) );
XNOR2_X2 inst_72 ( .B(net_3124), .A(net_1583), .ZN(net_1581) );
INV_X4 inst_2404 ( .A(net_3920), .ZN(net_352) );
CLKBUF_X2 inst_5127 ( .A(net_5112), .Z(net_5113) );
NAND2_X2 inst_1578 ( .A1(net_2965), .ZN(net_2442), .A2(net_552) );
NAND2_X2 inst_1634 ( .A2(net_3156), .ZN(net_2303), .A1(net_2215) );
NAND2_X2 inst_1666 ( .A2(net_4009), .A1(net_3817), .ZN(net_2092) );
AOI22_X2 inst_3542 ( .ZN(net_1584), .A1(net_1583), .B1(net_744), .B2(net_513), .A2(net_297) );
OAI21_X2 inst_735 ( .B2(net_1523), .A(net_629), .B1(net_628), .ZN(net_575) );
NAND2_X2 inst_1529 ( .A1(net_3208), .ZN(net_2493), .A2(net_139) );
XNOR2_X2 inst_115 ( .ZN(net_348), .A(net_327), .B(net_289) );
CLKBUF_X2 inst_4612 ( .A(net_4323), .Z(net_4598) );
NAND2_X2 inst_1653 ( .ZN(net_2135), .A1(net_2028), .A2(net_1976) );
CLKBUF_X2 inst_4691 ( .A(net_4676), .Z(net_4677) );
AOI22_X2 inst_3726 ( .A1(net_4107), .ZN(net_3723), .A2(net_3680), .B1(net_1018), .B2(net_521) );
CLKBUF_X2 inst_4638 ( .A(net_4623), .Z(net_4624) );
INV_X2 inst_3045 ( .ZN(net_3705), .A(net_264) );
NAND2_X2 inst_1582 ( .A2(net_3401), .A1(net_2915), .ZN(net_2438) );
INV_X2 inst_2984 ( .A(net_3007), .ZN(net_141) );
OR3_X4 inst_175 ( .ZN(net_628), .A2(net_389), .A1(net_309), .A3(net_263) );
DFF_X1 inst_3258 ( .QN(net_3078), .D(net_2943), .CK(net_4537) );
CLKBUF_X2 inst_5010 ( .A(net_4995), .Z(net_4996) );
NAND2_X2 inst_1737 ( .A2(net_2268), .ZN(net_1529), .A1(net_1528) );
NAND2_X2 inst_1805 ( .A1(net_4082), .ZN(net_959), .A2(net_913) );
NAND2_X2 inst_1840 ( .A2(net_4111), .ZN(net_1213), .A1(net_690) );
INV_X2 inst_2995 ( .ZN(net_127), .A(net_121) );
AOI22_X2 inst_3563 ( .A1(net_4059), .B1(net_4056), .ZN(net_1487), .A2(net_518), .B2(net_479) );
SDFF_X2 inst_133 ( .D(net_3483), .SI(net_3023), .Q(net_3023), .SE(net_2917), .CK(net_5161) );
NAND3_X4 inst_1263 ( .A3(net_3965), .ZN(net_2212), .A1(net_1269), .A2(net_1034) );
CLKBUF_X2 inst_4541 ( .A(net_4526), .Z(net_4527) );
INV_X2 inst_2752 ( .ZN(net_1124), .A(net_641) );
DFF_X1 inst_3330 ( .D(net_2820), .QN(net_318), .CK(net_4325) );
NOR2_X2 inst_1149 ( .ZN(net_3934), .A2(net_3932), .A1(net_3221) );
NAND2_X2 inst_1721 ( .A1(net_3320), .ZN(net_1739), .A2(net_360) );
NAND2_X4 inst_1445 ( .A1(net_3922), .A2(net_3826), .ZN(net_3788) );
NAND3_X2 inst_1281 ( .A2(net_4101), .A3(net_3559), .ZN(net_2545), .A1(net_2345) );
NAND2_X2 inst_1509 ( .A2(net_3738), .ZN(net_2634), .A1(net_2633) );
HA_X1 inst_3088 ( .S(net_1713), .CO(net_1712), .A(net_1711), .B(net_1710) );
AOI21_X2 inst_3990 ( .B1(net_3984), .A(net_3438), .ZN(net_705), .B2(net_442) );
XNOR2_X2 inst_126 ( .ZN(net_4190), .B(net_3224), .A(net_3223) );
AOI222_X1 inst_3782 ( .C2(net_3466), .B1(net_2020), .C1(net_1840), .ZN(net_1722), .A1(net_1698), .B2(net_382), .A2(net_255) );
CLKBUF_X2 inst_4719 ( .A(net_4704), .Z(net_4705) );
NAND2_X2 inst_1512 ( .ZN(net_2611), .A1(net_2610), .A2(net_1000) );
AOI221_X2 inst_3887 ( .C1(net_4064), .C2(net_4029), .ZN(net_1519), .B1(net_1518), .B2(net_1517), .A(net_1320) );
CLKBUF_X2 inst_5160 ( .A(net_4498), .Z(net_5146) );
NAND2_X2 inst_1631 ( .A1(net_3883), .A2(net_3858), .ZN(net_2321) );
CLKBUF_X2 inst_4353 ( .A(net_4279), .Z(net_4339) );
AOI21_X2 inst_3934 ( .ZN(net_2613), .B1(net_2612), .A(net_2388), .B2(net_1276) );
NOR2_X4 inst_948 ( .A2(net_3764), .ZN(net_3562), .A1(net_3478) );
NOR2_X2 inst_1140 ( .A1(net_3994), .ZN(net_3811), .A2(net_319) );
NOR2_X2 inst_1086 ( .A1(net_641), .ZN(net_431), .A2(net_334) );
INV_X2 inst_2643 ( .ZN(net_2338), .A(net_2317) );
NAND2_X2 inst_1688 ( .A1(net_3219), .ZN(net_1983), .A2(net_567) );
INV_X4 inst_2299 ( .A(net_3620), .ZN(net_1228) );
NAND2_X2 inst_1800 ( .A1(net_4081), .ZN(net_1082), .A2(net_245) );
CLKBUF_X2 inst_4773 ( .A(net_4758), .Z(net_4759) );
OAI221_X2 inst_448 ( .ZN(net_4151), .B1(net_3352), .C2(net_3348), .C1(net_2813), .A(net_2592), .B2(net_2189) );
CLKBUF_X2 inst_5292 ( .A(net_5277), .Z(net_5278) );
NOR3_X2 inst_914 ( .ZN(net_3473), .A2(net_3373), .A1(net_3238), .A3(net_2878) );
CLKBUF_X2 inst_4921 ( .A(net_4203), .Z(net_4907) );
CLKBUF_X2 inst_5170 ( .A(net_5155), .Z(net_5156) );
CLKBUF_X2 inst_5182 ( .A(net_5167), .Z(net_5168) );
CLKBUF_X2 inst_4380 ( .A(net_4365), .Z(net_4366) );
NAND2_X2 inst_2002 ( .A2(net_3858), .ZN(net_3513), .A1(net_3512) );
OAI221_X2 inst_384 ( .C1(net_3876), .B1(net_3175), .B2(net_2699), .C2(net_2698), .ZN(net_2628), .A(net_2536) );
NAND2_X2 inst_1642 ( .ZN(net_2174), .A1(net_2098), .A2(net_2024) );
NAND4_X2 inst_1252 ( .ZN(net_3847), .A2(net_2292), .A1(net_2280), .A4(net_2279), .A3(net_2182) );
OAI21_X2 inst_608 ( .B1(net_4136), .A(net_3316), .ZN(net_2306), .B2(net_1514) );
NAND3_X2 inst_1343 ( .ZN(net_3411), .A3(net_3410), .A1(net_3409), .A2(net_2613) );
AOI221_X2 inst_3800 ( .C1(net_2781), .ZN(net_2776), .B1(net_2775), .A(net_2667), .B2(net_2665), .C2(net_272) );
OAI211_X2 inst_834 ( .C1(net_1359), .ZN(net_1357), .A(net_1237), .B(net_671), .C2(net_292) );
INV_X2 inst_2920 ( .A(net_2984), .ZN(net_242) );
AND4_X2 inst_4054 ( .ZN(net_1766), .A1(net_1765), .A2(net_1764), .A4(net_1461), .A3(net_1380) );
NOR2_X4 inst_966 ( .ZN(net_3835), .A2(net_3633), .A1(net_3548) );
OR2_X4 inst_199 ( .A1(net_3204), .ZN(net_2967), .A2(net_2352) );
NAND4_X2 inst_1246 ( .ZN(net_3529), .A4(net_3282), .A1(net_2101), .A2(net_2091), .A3(net_1988) );
INV_X2 inst_2961 ( .A(net_3150), .ZN(net_2051) );
DFF_X2 inst_3185 ( .D(net_1763), .Q(net_77), .CK(net_4461) );
CLKBUF_X2 inst_4679 ( .A(net_4664), .Z(net_4665) );
INV_X4 inst_2209 ( .A(net_2377), .ZN(net_2246) );
INV_X4 inst_2506 ( .A(net_2987), .ZN(net_201) );
INV_X2 inst_2722 ( .ZN(net_1506), .A(net_1505) );
NAND4_X2 inst_1238 ( .A4(net_3153), .A3(net_3152), .ZN(net_544), .A1(net_332), .A2(net_316) );
INV_X8 inst_2171 ( .ZN(net_4164), .A(net_4163) );
CLKBUF_X2 inst_5245 ( .A(net_5230), .Z(net_5231) );
CLKBUF_X2 inst_4875 ( .A(net_4532), .Z(net_4861) );
CLKBUF_X2 inst_4557 ( .A(net_4385), .Z(net_4543) );
AOI22_X2 inst_3607 ( .A1(net_4062), .B1(net_4057), .ZN(net_1410), .B2(net_233), .A2(net_213) );
NAND2_X2 inst_2029 ( .ZN(net_3740), .A1(net_3738), .A2(net_67) );
DFF_X1 inst_3402 ( .Q(net_3120), .D(net_1544), .CK(net_4299) );
NOR2_X2 inst_1011 ( .ZN(net_2264), .A1(net_1863), .A2(net_1861) );
AND2_X4 inst_4114 ( .ZN(net_3469), .A1(net_2126), .A2(net_2125) );
OAI21_X2 inst_540 ( .ZN(net_4020), .B2(net_2967), .B1(net_2893), .A(net_2411) );
CLKBUF_X2 inst_4936 ( .A(net_4555), .Z(net_4922) );
OAI221_X2 inst_404 ( .B1(net_3781), .B2(net_3506), .ZN(net_1958), .C1(net_1884), .A(net_1751), .C2(net_355) );
INV_X4 inst_2356 ( .A(net_4005), .ZN(net_536) );
NOR2_X2 inst_998 ( .A2(net_3233), .ZN(net_3210), .A1(net_2025) );
DFF_X2 inst_3209 ( .QN(net_4034), .D(net_823), .CK(net_4823) );
DFF_X2 inst_3160 ( .D(net_2158), .QN(net_59), .CK(net_4207) );
INV_X2 inst_2861 ( .ZN(net_321), .A(net_125) );
XNOR2_X2 inst_66 ( .B(net_3492), .ZN(net_1696), .A(net_1242) );
AOI22_X2 inst_3615 ( .ZN(net_1331), .A2(net_1330), .A1(net_1211), .B1(net_1083), .B2(net_1035) );
CLKBUF_X2 inst_4814 ( .A(net_4799), .Z(net_4800) );
DFF_X2 inst_3216 ( .D(net_802), .QN(net_260), .CK(net_4619) );
OAI33_X1 inst_273 ( .ZN(net_1654), .A1(net_1653), .A2(net_1283), .B3(net_1173), .A3(net_791), .B2(net_246), .B1(x557) );
CLKBUF_X2 inst_5090 ( .A(net_4337), .Z(net_5076) );
OR2_X4 inst_192 ( .A1(net_3445), .ZN(net_2524), .A2(net_2388) );
NAND2_X2 inst_1965 ( .A2(net_4004), .ZN(net_3324), .A1(net_3106) );
AOI221_X2 inst_3915 ( .ZN(net_3356), .B2(net_3138), .A(net_2642), .B1(net_2591), .C2(net_2589), .C1(net_2583) );
OAI221_X2 inst_366 ( .ZN(net_2729), .A(net_2617), .B1(net_2546), .C1(net_2545), .C2(net_329), .B2(net_250) );
INV_X4 inst_2418 ( .A(net_3108), .ZN(net_319) );
INV_X2 inst_2715 ( .ZN(net_1560), .A(net_1559) );
CLKBUF_X2 inst_4242 ( .A(net_4204), .Z(net_4228) );
AOI22_X2 inst_3540 ( .ZN(net_1635), .A1(net_1634), .B2(net_1228), .A2(net_1089), .B1(net_1071) );
AND2_X4 inst_4126 ( .ZN(net_4052), .A1(net_2690), .A2(net_1444) );
AND2_X4 inst_4178 ( .ZN(net_4135), .A1(net_2185), .A2(net_1768) );
AOI22_X2 inst_3547 ( .B1(net_4054), .A2(net_1791), .A1(net_1578), .ZN(net_1574), .B2(net_243) );
NAND2_X2 inst_1574 ( .A1(net_2965), .ZN(net_2446), .A2(net_146) );
INV_X4 inst_2413 ( .A(net_322), .ZN(net_309) );
DFF_X1 inst_3285 ( .QN(net_3051), .D(net_2899), .CK(net_4860) );
CLKBUF_X2 inst_4746 ( .A(net_4731), .Z(net_4732) );
OR2_X4 inst_228 ( .ZN(net_1613), .A2(net_903), .A1(net_658) );
OAI21_X2 inst_486 ( .B1(net_3278), .ZN(net_2956), .B2(net_2909), .A(net_2463) );
NAND4_X2 inst_1240 ( .ZN(net_3232), .A3(net_3231), .A2(net_2100), .A1(net_2081), .A4(net_1983) );
NOR2_X2 inst_1025 ( .A1(net_3781), .ZN(net_1648), .A2(net_1609) );
OAI21_X2 inst_707 ( .ZN(net_857), .B1(net_709), .B2(net_684), .A(net_414) );
CLKBUF_X2 inst_4655 ( .A(net_4430), .Z(net_4641) );
AOI22_X2 inst_3670 ( .A2(net_571), .B2(net_570), .ZN(net_554), .A1(net_244), .B1(net_139) );
CLKBUF_X2 inst_4460 ( .A(net_4258), .Z(net_4446) );
OR2_X4 inst_244 ( .ZN(net_3945), .A2(net_3109), .A1(net_3107) );
CLKBUF_X2 inst_5262 ( .A(net_5239), .Z(net_5248) );
INV_X2 inst_2804 ( .ZN(net_1094), .A(net_725) );
CLKBUF_X2 inst_5131 ( .A(net_5116), .Z(net_5117) );
NAND2_X2 inst_1521 ( .A1(net_2959), .ZN(net_2501), .A2(net_731) );
INV_X4 inst_2576 ( .ZN(net_3594), .A(net_3591) );
INV_X1 inst_3079 ( .ZN(net_3358), .A(net_2815) );
INV_X2 inst_2631 ( .ZN(net_2694), .A(net_2693) );
CLKBUF_X2 inst_4845 ( .A(net_4830), .Z(net_4831) );
NAND3_X2 inst_1306 ( .ZN(net_1150), .A2(net_1143), .A1(net_1142), .A3(net_970) );
OAI21_X1 inst_772 ( .ZN(net_4012), .B2(net_2965), .B1(net_2893), .A(net_2447) );
INV_X4 inst_2563 ( .A(net_3858), .ZN(net_3515) );
AOI221_X2 inst_3810 ( .B2(net_3133), .ZN(net_2643), .A(net_2642), .B1(net_2641), .C1(net_2640), .C2(net_2222) );
NAND2_X4 inst_1407 ( .ZN(net_3287), .A1(net_3252), .A2(net_2838) );
AOI22_X2 inst_3682 ( .B2(net_4123), .A2(net_555), .ZN(net_501), .B1(net_196), .A1(net_191) );
CLKBUF_X2 inst_4940 ( .A(net_4413), .Z(net_4926) );
CLKBUF_X2 inst_4523 ( .A(net_4482), .Z(net_4509) );
CLKBUF_X2 inst_4583 ( .A(net_4557), .Z(net_4569) );
INV_X2 inst_2636 ( .ZN(net_2516), .A(net_2515) );
CLKBUF_X2 inst_4870 ( .A(net_4855), .Z(net_4856) );
OAI221_X2 inst_445 ( .B1(net_4160), .ZN(net_3697), .B2(net_3407), .C1(net_2328), .A(net_1940), .C2(net_1444) );
CLKBUF_X2 inst_5192 ( .A(net_5177), .Z(net_5178) );
XNOR2_X2 inst_93 ( .ZN(net_813), .A(net_664), .B(net_653) );
AOI22_X2 inst_3606 ( .A1(net_4063), .B1(net_4058), .ZN(net_1411), .A2(net_180), .B2(net_154) );
CLKBUF_X2 inst_4832 ( .A(net_4817), .Z(net_4818) );
OAI21_X2 inst_606 ( .B2(net_3428), .B1(net_3312), .ZN(net_2331), .A(net_2138) );
INV_X2 inst_2942 ( .A(net_3019), .ZN(net_237) );
CLKBUF_X2 inst_5089 ( .A(net_5074), .Z(net_5075) );
AOI222_X1 inst_3761 ( .C1(net_3117), .A1(net_2055), .B2(net_2054), .C2(net_2053), .ZN(net_2001), .B1(net_1743), .A2(net_142) );
CLKBUF_X2 inst_5099 ( .A(net_5084), .Z(net_5085) );
CLKBUF_X2 inst_4595 ( .A(net_4580), .Z(net_4581) );
OAI211_X2 inst_853 ( .A(net_4108), .C1(net_3913), .B(net_3669), .ZN(net_3322), .C2(net_3319) );
SDFF_X2 inst_139 ( .D(net_3343), .SE(net_2514), .SI(net_100), .Q(net_100), .CK(net_4754) );
OAI21_X2 inst_657 ( .B2(net_4088), .ZN(net_1941), .B1(net_1815), .A(net_1803) );
NAND2_X2 inst_1675 ( .ZN(net_2083), .A1(net_2082), .A2(net_163) );
OAI21_X2 inst_584 ( .B1(net_4037), .B2(net_2815), .ZN(net_2744), .A(net_1577) );
CLKBUF_X2 inst_4550 ( .A(net_4535), .Z(net_4536) );
NAND3_X2 inst_1316 ( .A1(net_4096), .A2(net_3713), .ZN(net_995), .A3(net_947) );
NAND2_X1 inst_2098 ( .ZN(net_3605), .A1(net_3541), .A2(net_3270) );
OAI21_X2 inst_470 ( .B1(net_3509), .ZN(net_2980), .B2(net_2972), .A(net_2431) );
AOI22_X2 inst_3551 ( .A1(net_4060), .B1(net_4055), .A2(net_4011), .B2(net_4009), .ZN(net_1499) );
NAND2_X2 inst_1921 ( .A1(net_3156), .ZN(net_1521), .A2(x1023) );
CLKBUF_X2 inst_5149 ( .A(net_5134), .Z(net_5135) );
CLKBUF_X2 inst_4237 ( .A(net_4211), .Z(net_4223) );
CLKBUF_X2 inst_4490 ( .A(net_4475), .Z(net_4476) );
SDFF_X2 inst_148 ( .D(net_3827), .SE(net_2514), .SI(net_97), .Q(net_97), .CK(net_4943) );
NAND2_X2 inst_1752 ( .ZN(net_1312), .A2(net_1311), .A1(net_1114) );
OAI21_X2 inst_554 ( .B2(net_2919), .ZN(net_2872), .B1(net_2871), .A(net_2399) );
CLKBUF_X2 inst_4293 ( .A(net_4278), .Z(net_4279) );
NAND4_X2 inst_1187 ( .A3(net_4049), .A4(net_2144), .ZN(net_1868), .A1(net_1867), .A2(net_1866) );
OR2_X4 inst_191 ( .A2(net_4040), .A1(net_2714), .ZN(net_2528) );
CLKBUF_X2 inst_4333 ( .A(net_4318), .Z(net_4319) );
NOR2_X2 inst_1063 ( .A2(net_4104), .A1(net_4083), .ZN(net_1009) );
INV_X2 inst_2700 ( .ZN(net_1679), .A(net_1678) );
NAND2_X2 inst_1917 ( .A2(net_389), .A1(net_322), .ZN(net_312) );
INV_X2 inst_2638 ( .ZN(net_2387), .A(net_2386) );
DFF_X1 inst_3252 ( .QN(net_3081), .D(net_2953), .CK(net_4732) );
CLKBUF_X2 inst_4565 ( .A(net_4319), .Z(net_4551) );
CLKBUF_X2 inst_4538 ( .A(net_4512), .Z(net_4524) );
CLKBUF_X2 inst_5212 ( .A(net_5197), .Z(net_5198) );
CLKBUF_X2 inst_4955 ( .A(net_4940), .Z(net_4941) );
CLKBUF_X2 inst_4755 ( .A(net_4691), .Z(net_4741) );
DFF_X1 inst_3235 ( .D(net_3279), .QN(net_3043), .CK(net_5047) );
CLKBUF_X2 inst_5276 ( .A(net_5261), .Z(net_5262) );
NOR2_X1 inst_1167 ( .A2(net_514), .ZN(net_425), .A1(net_284) );
AOI221_X2 inst_3879 ( .A(net_4047), .C2(net_1908), .ZN(net_1850), .C1(net_1849), .B2(net_749), .B1(net_98) );
CLKBUF_X2 inst_5269 ( .A(net_5254), .Z(net_5255) );
NAND2_X1 inst_2087 ( .A1(net_2972), .ZN(net_2430), .A2(net_732) );
INV_X4 inst_2184 ( .ZN(net_2775), .A(net_2561) );
NAND3_X2 inst_1303 ( .A3(net_3497), .A1(net_1691), .ZN(net_1317), .A2(net_1316) );
NOR3_X2 inst_892 ( .ZN(net_2345), .A1(net_2325), .A2(net_2282), .A3(net_1173) );
NAND2_X2 inst_1623 ( .A1(net_2917), .ZN(net_2393), .A2(net_205) );
INV_X2 inst_2665 ( .ZN(net_2350), .A(net_2134) );
AND3_X2 inst_4088 ( .A3(net_3627), .ZN(net_944), .A1(net_943), .A2(net_591) );
NOR2_X2 inst_1132 ( .ZN(net_3643), .A2(net_3168), .A1(net_3167) );
CLKBUF_X2 inst_4922 ( .A(net_4907), .Z(net_4908) );
CLKBUF_X2 inst_4464 ( .A(net_4449), .Z(net_4450) );
AND2_X4 inst_4100 ( .A2(net_4034), .ZN(net_1097), .A1(net_1096) );
NOR2_X4 inst_968 ( .ZN(net_3875), .A2(net_3529), .A1(net_3528) );
OAI211_X2 inst_819 ( .A(net_3487), .ZN(net_1946), .B(net_934), .C2(net_433), .C1(net_280) );
CLKBUF_X2 inst_4700 ( .A(net_4685), .Z(net_4686) );
DFF_X1 inst_3320 ( .QN(net_3001), .D(net_2850), .CK(net_5070) );
CLKBUF_X2 inst_4441 ( .A(net_4426), .Z(net_4427) );
NAND2_X4 inst_1468 ( .ZN(net_3898), .A1(net_3897), .A2(net_3289) );
NAND2_X2 inst_1803 ( .A1(net_4082), .ZN(net_1256), .A2(net_778) );
NAND2_X2 inst_1516 ( .A2(net_4040), .ZN(net_2670), .A1(net_2668) );
AOI222_X1 inst_3776 ( .C1(net_3115), .B2(net_2020), .ZN(net_1842), .A1(net_1841), .C2(net_1840), .B1(net_772), .A2(net_206) );
DFF_X2 inst_3153 ( .D(net_2262), .QN(net_45), .CK(net_4413) );
OAI221_X2 inst_386 ( .B1(net_3449), .B2(net_2666), .ZN(net_2616), .C1(net_2615), .C2(net_1727), .A(net_1386) );
INV_X2 inst_2814 ( .ZN(net_646), .A(net_638) );
INV_X4 inst_2617 ( .ZN(net_3889), .A(net_3888) );
NOR2_X4 inst_936 ( .A2(net_3755), .ZN(net_407), .A1(net_337) );
AOI221_X2 inst_3809 ( .ZN(net_2644), .A(net_2642), .B1(net_2641), .C1(net_2640), .C2(net_2220), .B2(net_265) );
AOI21_X2 inst_4004 ( .ZN(net_3844), .B2(net_3842), .A(net_1721), .B1(net_1228) );
AOI21_X2 inst_3942 ( .ZN(net_2239), .B1(net_2238), .A(net_2166), .B2(net_238) );
INV_X16 inst_3068 ( .ZN(net_3817), .A(net_3799) );
CLKBUF_X2 inst_5225 ( .A(net_4471), .Z(net_5211) );
INV_X4 inst_2277 ( .A(net_1081), .ZN(net_973) );
INV_X2 inst_2778 ( .ZN(net_808), .A(net_762) );
CLKBUF_X2 inst_5223 ( .A(net_5208), .Z(net_5209) );
AOI221_X2 inst_3798 ( .ZN(net_2832), .A(net_2783), .C1(net_2781), .B1(net_2724), .C2(net_83), .B2(net_36) );
CLKBUF_X2 inst_5232 ( .A(net_5217), .Z(net_5218) );
AND2_X4 inst_4109 ( .A1(net_3164), .A2(net_3162), .ZN(net_345) );
AND2_X2 inst_4192 ( .ZN(net_2608), .A2(net_2607), .A1(net_2544) );
INV_X2 inst_2962 ( .A(net_2998), .ZN(net_170) );
INV_X2 inst_3004 ( .A(net_3615), .ZN(net_3221) );
AOI222_X1 inst_3780 ( .A2(net_3705), .B1(net_1795), .A1(net_1794), .C1(net_1793), .ZN(net_1792), .C2(net_1791), .B2(net_717) );
INV_X2 inst_2647 ( .A(net_3880), .ZN(net_2335) );
CLKBUF_X2 inst_4672 ( .A(net_4657), .Z(net_4658) );
OAI211_X2 inst_811 ( .ZN(net_1629), .B(net_1628), .C1(net_1627), .A(net_1555), .C2(net_530) );
OR2_X4 inst_208 ( .A2(net_3447), .ZN(net_2714), .A1(net_2281) );
AND2_X2 inst_4202 ( .A2(net_3662), .ZN(net_690), .A1(net_609) );
INV_X4 inst_2456 ( .A(net_3089), .ZN(net_498) );
AOI222_X1 inst_3774 ( .C2(net_2051), .B2(net_2020), .ZN(net_1860), .A1(net_1841), .C1(net_1840), .B1(net_873), .A2(net_83) );
INV_X2 inst_2710 ( .A(net_1799), .ZN(net_1632) );
NOR2_X2 inst_1058 ( .A2(net_4024), .A1(net_1908), .ZN(net_1002) );
INV_X2 inst_2887 ( .A(net_505), .ZN(net_168) );
CLKBUF_X2 inst_5282 ( .A(net_4869), .Z(net_5268) );
AOI221_X2 inst_3909 ( .B1(net_4106), .C1(net_3563), .A(net_3546), .C2(net_3478), .ZN(net_870), .B2(net_281) );
NAND2_X2 inst_1869 ( .ZN(net_610), .A1(net_542), .A2(net_261) );
NOR3_X2 inst_897 ( .A2(net_3783), .ZN(net_1376), .A1(net_1271), .A3(net_657) );
DFF_X1 inst_3360 ( .D(net_2362), .CK(net_4230), .Q(x437) );
AOI21_X2 inst_3945 ( .B1(net_3774), .ZN(net_2225), .A(net_2148), .B2(net_1507) );
CLKBUF_X2 inst_4984 ( .A(net_4969), .Z(net_4970) );
NAND4_X2 inst_1201 ( .ZN(net_1672), .A3(net_1475), .A4(net_1474), .A1(net_1409), .A2(net_1408) );
NAND2_X4 inst_1473 ( .ZN(net_3926), .A1(net_3168), .A2(net_268) );
NAND2_X2 inst_1788 ( .ZN(net_1066), .A2(net_1016), .A1(net_910) );
NAND3_X4 inst_1272 ( .ZN(net_3997), .A2(net_3996), .A3(net_3765), .A1(net_3243) );
AND2_X4 inst_4182 ( .ZN(net_4144), .A2(net_4130), .A1(net_3128) );
OAI21_X2 inst_636 ( .A(net_3750), .B2(net_2076), .ZN(net_2074), .B1(net_1675) );
OAI21_X2 inst_632 ( .ZN(net_2079), .A(net_1961), .B2(net_1960), .B1(net_1189) );
XOR2_X2 inst_0 ( .Z(net_2538), .A(net_2330), .B(net_1781) );
INV_X2 inst_2852 ( .A(net_374), .ZN(net_335) );
NAND2_X2 inst_1927 ( .ZN(net_3190), .A1(net_3186), .A2(net_234) );
OR3_X2 inst_184 ( .ZN(net_606), .A3(net_605), .A1(net_601), .A2(net_523) );
NAND2_X2 inst_1847 ( .ZN(net_680), .A2(net_640), .A1(net_414) );
AOI21_X2 inst_3973 ( .B2(net_1330), .ZN(net_1219), .A(net_1155), .B1(net_1078) );
NAND2_X2 inst_1907 ( .A2(net_1326), .A1(net_686), .ZN(net_311) );
OAI221_X2 inst_433 ( .B2(net_3418), .A(net_629), .B1(net_628), .C1(net_627), .ZN(net_626), .C2(net_40) );
NAND2_X2 inst_1983 ( .A1(net_4095), .ZN(net_3406), .A2(net_297) );
CLKBUF_X2 inst_4939 ( .A(net_4924), .Z(net_4925) );
AOI221_X2 inst_3836 ( .B1(net_3774), .ZN(net_2228), .C1(net_2227), .A(net_2108), .C2(net_1637), .B2(net_1439) );
INV_X4 inst_2192 ( .A(net_2714), .ZN(net_2668) );
NAND2_X2 inst_1948 ( .ZN(net_3266), .A2(net_3265), .A1(net_1978) );
MUX2_X2 inst_2114 ( .Z(net_3380), .S(net_3379), .A(net_1401), .B(net_1400) );
INV_X2 inst_2784 ( .ZN(net_802), .A(net_756) );
CLKBUF_X2 inst_4216 ( .A(net_4201), .Z(net_4202) );
XNOR2_X2 inst_106 ( .B(net_3122), .ZN(net_542), .A(net_309) );
OAI221_X2 inst_422 ( .ZN(net_1185), .A(net_1067), .B2(net_719), .B1(net_716), .C2(net_693), .C1(net_667) );
INV_X4 inst_2583 ( .A(net_3918), .ZN(net_3628) );
INV_X4 inst_2243 ( .ZN(net_1808), .A(net_1520) );
NAND2_X4 inst_1475 ( .A1(net_3977), .ZN(net_3938), .A2(net_3937) );
NAND2_X4 inst_1426 ( .ZN(net_3597), .A2(net_3596), .A1(net_3593) );
CLKBUF_X2 inst_4812 ( .A(net_4487), .Z(net_4798) );
HA_X1 inst_3090 ( .A(net_3492), .S(net_1707), .CO(net_1706), .B(net_1705) );
NAND2_X2 inst_1637 ( .A1(net_4042), .ZN(net_2698), .A2(net_2169) );
AOI21_X2 inst_3997 ( .ZN(net_3560), .B2(net_3559), .B1(net_957), .A(net_848) );
NAND3_X2 inst_1352 ( .A1(net_3719), .ZN(net_3683), .A2(net_3672), .A3(net_3399) );
CLKBUF_X2 inst_5241 ( .A(net_5226), .Z(net_5227) );
CLKBUF_X2 inst_4377 ( .A(net_4213), .Z(net_4363) );
INV_X4 inst_2261 ( .ZN(net_1393), .A(net_1359) );
CLKBUF_X2 inst_4879 ( .A(net_4296), .Z(net_4865) );
CLKBUF_X2 inst_4383 ( .A(net_4368), .Z(net_4369) );
CLKBUF_X2 inst_4301 ( .A(net_4286), .Z(net_4287) );
CLKBUF_X2 inst_4695 ( .A(net_4680), .Z(net_4681) );
AND2_X4 inst_4142 ( .ZN(net_4078), .A2(net_847), .A1(net_663) );
DFF_X1 inst_3390 ( .D(net_1733), .QN(net_81), .CK(net_4428) );
INV_X2 inst_2930 ( .ZN(net_1280), .A(net_113) );
CLKBUF_X2 inst_5106 ( .A(net_5091), .Z(net_5092) );
NAND2_X4 inst_1410 ( .A1(net_3858), .ZN(net_3331), .A2(net_931) );
CLKBUF_X2 inst_4790 ( .A(net_4775), .Z(net_4776) );
CLKBUF_X2 inst_4307 ( .A(net_4292), .Z(net_4293) );
INV_X2 inst_2859 ( .ZN(net_302), .A(net_301) );
CLKBUF_X2 inst_4991 ( .A(net_4976), .Z(net_4977) );
OAI221_X2 inst_397 ( .C2(net_3407), .B1(net_2328), .ZN(net_2294), .C1(net_2194), .A(net_2022), .B2(net_66) );
AOI222_X1 inst_3756 ( .A1(net_3676), .B1(net_2055), .C1(net_2054), .ZN(net_2036), .C2(net_419), .A2(net_256), .B2(net_168) );
OAI21_X2 inst_504 ( .B1(net_3278), .ZN(net_2938), .B2(net_2919), .A(net_2397) );
CLKBUF_X2 inst_4424 ( .A(net_4409), .Z(net_4410) );
DFF_X2 inst_3192 ( .QN(net_3109), .D(net_1630), .CK(net_4834) );
CLKBUF_X2 inst_5006 ( .A(net_4822), .Z(net_4992) );
NAND2_X2 inst_1733 ( .A1(net_1556), .ZN(net_1552), .A2(x672) );
NAND3_X2 inst_1297 ( .A2(net_1821), .ZN(net_1585), .A3(net_1386), .A1(net_1170) );
AOI221_X2 inst_3900 ( .C2(net_3941), .ZN(net_1206), .A(net_1203), .B1(net_1202), .C1(net_1201), .B2(net_599) );
DFF_X2 inst_3194 ( .QN(net_3106), .D(net_1624), .CK(net_5132) );
NOR3_X2 inst_918 ( .ZN(net_4101), .A2(net_3954), .A1(net_637), .A3(net_516) );
INV_X4 inst_2199 ( .A(net_3882), .ZN(net_2314) );
CLKBUF_X2 inst_4751 ( .A(net_4501), .Z(net_4737) );
AOI221_X2 inst_3884 ( .ZN(net_1720), .C1(net_1718), .C2(net_1656), .A(net_1362), .B1(net_1184), .B2(net_204) );
CLKBUF_X2 inst_4246 ( .A(net_4231), .Z(net_4232) );
NOR2_X1 inst_1173 ( .ZN(net_4193), .A2(net_3543), .A1(net_432) );
AOI221_X2 inst_3904 ( .A(net_4090), .B2(net_3680), .B1(net_1028), .ZN(net_1020), .C1(net_746), .C2(net_521) );
INV_X2 inst_2908 ( .A(net_3095), .ZN(net_191) );
CLKBUF_X2 inst_5019 ( .A(net_5004), .Z(net_5005) );
NAND2_X4 inst_1393 ( .A2(net_4013), .A1(net_2134), .ZN(net_2093) );
NAND2_X2 inst_2074 ( .ZN(net_4068), .A1(net_3836), .A2(net_3547) );
AOI211_X1 inst_4035 ( .A(net_3958), .B(net_3621), .ZN(net_3318), .C2(net_963), .C1(net_905) );
NAND2_X2 inst_1862 ( .ZN(net_592), .A1(net_591), .A2(net_590) );
AOI22_X2 inst_3519 ( .B1(net_4045), .B2(net_3151), .A1(net_1955), .ZN(net_1951), .A2(net_295) );
CLKBUF_X2 inst_4823 ( .A(net_4806), .Z(net_4809) );
NAND4_X2 inst_1236 ( .A3(net_4125), .A2(net_3900), .ZN(net_745), .A4(net_431), .A1(net_386) );
OR2_X4 inst_221 ( .A1(net_4081), .ZN(net_1033), .A2(net_245) );
AND3_X4 inst_4075 ( .A3(net_4162), .A2(net_4118), .ZN(net_4085), .A1(net_3900) );
CLKBUF_X2 inst_5112 ( .A(net_5097), .Z(net_5098) );
DFF_X1 inst_3313 ( .QN(net_2999), .D(net_2848), .CK(net_5202) );
AOI22_X2 inst_3562 ( .A1(net_4060), .B1(net_4055), .ZN(net_1488), .A2(net_221), .B2(net_155) );
CLKBUF_X2 inst_4893 ( .A(net_4878), .Z(net_4879) );
CLKBUF_X2 inst_5153 ( .A(net_5138), .Z(net_5139) );
INV_X4 inst_2334 ( .ZN(net_765), .A(net_633) );
INV_X4 inst_2429 ( .A(net_2991), .ZN(net_159) );
INV_X4 inst_2210 ( .ZN(net_2282), .A(net_2206) );
OAI21_X2 inst_754 ( .B1(net_4103), .A(net_3764), .ZN(net_3564), .B2(net_439) );
CLKBUF_X2 inst_4791 ( .A(net_4776), .Z(net_4777) );
INV_X2 inst_2937 ( .A(net_3048), .ZN(net_241) );
CLKBUF_X2 inst_5028 ( .A(net_5013), .Z(net_5014) );
INV_X4 inst_2590 ( .ZN(net_3678), .A(net_3270) );
INV_X2 inst_2913 ( .A(net_3119), .ZN(net_134) );
OAI21_X2 inst_687 ( .B1(net_3228), .A(net_1307), .ZN(net_1305), .B2(net_327) );
NAND2_X2 inst_1774 ( .A1(net_2213), .A2(net_1884), .ZN(net_1394) );
INV_X4 inst_2319 ( .ZN(net_866), .A(net_703) );
CLKBUF_X2 inst_5025 ( .A(net_4513), .Z(net_5011) );
DFF_X1 inst_3295 ( .QN(net_3009), .D(net_2888), .CK(net_5223) );
NOR2_X2 inst_985 ( .ZN(net_2600), .A1(net_2599), .A2(net_2598) );
CLKBUF_X2 inst_5057 ( .A(net_5042), .Z(net_5043) );
INV_X4 inst_2225 ( .ZN(net_2129), .A(net_1835) );
INV_X4 inst_2513 ( .ZN(net_1611), .A(net_85) );
AND3_X4 inst_4061 ( .A3(net_3320), .ZN(net_1968), .A1(net_1828), .A2(net_1645) );
INV_X4 inst_2254 ( .ZN(net_2020), .A(net_1701) );
CLKBUF_X2 inst_4459 ( .A(net_4444), .Z(net_4445) );
INV_X2 inst_2923 ( .A(net_3001), .ZN(net_151) );
INV_X2 inst_2707 ( .ZN(net_2663), .A(net_2594) );
NOR2_X2 inst_1117 ( .A1(net_3654), .ZN(net_3395), .A2(net_283) );
AOI211_X2 inst_4015 ( .C1(net_3554), .ZN(net_2517), .C2(net_2378), .A(net_1747), .B(net_1685) );
AOI21_X2 inst_3958 ( .B2(net_3441), .ZN(net_1703), .B1(net_1527), .A(net_375) );
NAND2_X2 inst_2007 ( .A2(net_3887), .A1(net_3848), .ZN(net_3537) );
INV_X2 inst_2725 ( .ZN(net_1466), .A(net_1395) );
CLKBUF_X2 inst_5141 ( .A(net_4252), .Z(net_5127) );
AOI22_X2 inst_3644 ( .A1(net_4142), .B1(net_4112), .ZN(net_758), .B2(net_396), .A2(x672) );
NAND2_X2 inst_1610 ( .A1(net_2967), .ZN(net_2406), .A2(net_454) );
OAI22_X2 inst_334 ( .ZN(net_515), .A1(net_514), .A2(net_298), .B1(net_284), .B2(net_264) );
CLKBUF_X2 inst_4620 ( .A(net_4605), .Z(net_4606) );
OAI211_X2 inst_805 ( .C2(net_3845), .ZN(net_1913), .C1(net_1912), .A(net_1820), .B(net_1755) );
AOI22_X2 inst_3707 ( .ZN(net_459), .A1(net_458), .B1(net_457), .B2(net_186), .A2(net_162) );
OAI222_X2 inst_354 ( .B1(net_2717), .A1(net_1126), .ZN(net_1093), .A2(net_1092), .C2(net_988), .C1(net_891), .B2(net_854) );
NOR2_X2 inst_1145 ( .ZN(net_3897), .A1(net_3213), .A2(net_3212) );
NOR2_X2 inst_1042 ( .A2(net_4025), .ZN(net_1247), .A1(net_1003) );
CLKBUF_X2 inst_4492 ( .A(net_4477), .Z(net_4478) );
OAI221_X2 inst_373 ( .B1(net_2733), .C1(net_2686), .ZN(net_2683), .A(net_2559), .B2(net_1748), .C2(net_1655) );
INV_X2 inst_3056 ( .ZN(net_3930), .A(net_3929) );
NAND2_X2 inst_1868 ( .ZN(net_662), .A2(net_449), .A1(net_245) );
OAI21_X2 inst_595 ( .B2(net_2815), .ZN(net_2539), .B1(net_2538), .A(net_1745) );
INV_X4 inst_2609 ( .A(net_3823), .ZN(net_3821) );
XOR2_X2 inst_22 ( .Z(net_4073), .A(net_687), .B(net_42) );
CLKBUF_X2 inst_5002 ( .A(net_4987), .Z(net_4988) );
NAND2_X2 inst_1717 ( .A1(net_3492), .ZN(net_2378), .A2(net_1641) );
INV_X4 inst_2556 ( .ZN(net_3489), .A(net_3170) );
HA_X1 inst_3099 ( .S(net_751), .CO(net_676), .A(net_448), .B(net_261) );
NAND2_X2 inst_1704 ( .A1(net_1834), .ZN(net_1833), .A2(net_360) );
CLKBUF_X2 inst_4604 ( .A(net_4519), .Z(net_4590) );
INV_X2 inst_2901 ( .A(net_3146), .ZN(net_265) );
OAI21_X2 inst_767 ( .ZN(net_3962), .A(net_3960), .B2(net_3620), .B1(net_763) );
CLKBUF_X2 inst_4688 ( .A(net_4673), .Z(net_4674) );
OR4_X2 inst_161 ( .A4(net_3955), .ZN(net_1073), .A1(net_1072), .A2(net_969), .A3(net_812) );
DFF_X1 inst_3356 ( .D(net_3707), .CK(net_4411), .Q(x388) );
CLKBUF_X2 inst_4798 ( .A(net_4783), .Z(net_4784) );
AOI221_X2 inst_3849 ( .B1(net_3736), .C2(net_3114), .ZN(net_2116), .C1(net_2115), .A(net_1934), .B2(net_72) );
OAI21_X2 inst_718 ( .B1(net_3670), .B2(net_3214), .A(net_748), .ZN(net_743) );
NOR2_X2 inst_1029 ( .A1(net_2212), .ZN(net_1569), .A2(net_954) );
AOI211_X2 inst_4024 ( .A(net_3438), .ZN(net_1220), .B(net_1089), .C1(net_1007), .C2(net_903) );
INV_X4 inst_2408 ( .ZN(net_313), .A(net_285) );
NAND3_X2 inst_1324 ( .A3(net_3619), .A1(net_1168), .ZN(net_706), .A2(net_531) );
CLKBUF_X2 inst_4310 ( .A(net_4225), .Z(net_4296) );
OAI22_X2 inst_342 ( .B1(net_3871), .A1(net_3556), .ZN(net_3400), .A2(net_3011), .B2(net_3010) );
OAI21_X2 inst_526 ( .B1(net_3302), .ZN(net_2910), .B2(net_2909), .A(net_2464) );
INV_X8 inst_2147 ( .A(net_3580), .ZN(net_3278) );
NAND4_X4 inst_1178 ( .ZN(net_3937), .A4(net_3936), .A3(net_3766), .A2(net_3664), .A1(net_3521) );
OAI21_X4 inst_463 ( .B1(net_3878), .A(net_3858), .B2(net_3611), .ZN(net_3530) );
NAND2_X1 inst_2091 ( .A1(net_3430), .ZN(net_862), .A2(net_184) );
NAND2_X2 inst_1534 ( .A1(net_3207), .ZN(net_2488), .A2(net_217) );
DFF_X2 inst_3104 ( .D(net_2857), .QN(net_50), .CK(net_4689) );
CLKBUF_X2 inst_4667 ( .A(net_4652), .Z(net_4653) );
AOI221_X2 inst_3820 ( .A(net_2642), .B1(net_2641), .C1(net_2581), .ZN(net_2558), .C2(net_2555), .B2(net_256) );
OAI22_X2 inst_319 ( .B1(net_3143), .ZN(net_1641), .A2(net_1071), .B2(net_1036), .A1(net_952) );
NAND2_X4 inst_1450 ( .A2(net_3859), .ZN(net_3807), .A1(net_2335) );
INV_X4 inst_2422 ( .ZN(net_984), .A(net_48) );
DFF_X2 inst_3123 ( .QN(net_3135), .D(net_2652), .CK(net_4581) );
OAI21_X2 inst_649 ( .B1(net_4180), .ZN(net_2563), .B2(net_1975), .A(net_1524) );
INV_X8 inst_2158 ( .A(net_3938), .ZN(net_3637) );
AOI22_X2 inst_3725 ( .ZN(net_3652), .B1(net_3647), .A1(net_3185), .B2(net_467), .A2(net_454) );
NAND2_X2 inst_1711 ( .A2(net_4034), .ZN(net_1746), .A1(net_1603) );
INV_X4 inst_2597 ( .ZN(net_3738), .A(net_3737) );
DFF_X1 inst_3426 ( .Q(net_4013), .D(net_4012), .CK(net_4914) );
OAI21_X2 inst_500 ( .B1(net_3588), .B2(net_2961), .ZN(net_2942), .A(net_2470) );
NAND2_X2 inst_1592 ( .A1(net_2972), .ZN(net_2426), .A2(net_161) );
NAND2_X2 inst_1770 ( .ZN(net_1171), .A2(net_1170), .A1(net_1107) );
CLKBUF_X2 inst_5185 ( .A(net_5170), .Z(net_5171) );
NAND2_X2 inst_1575 ( .A1(net_2965), .ZN(net_2445), .A2(net_568) );
NOR2_X2 inst_995 ( .ZN(net_2271), .A1(net_2211), .A2(net_1090) );
OAI21_X2 inst_550 ( .B2(net_3207), .B1(net_2887), .ZN(net_2881), .A(net_2477) );
NAND2_X2 inst_2052 ( .ZN(net_3885), .A1(net_3787), .A2(net_2279) );
DFF_X1 inst_3413 ( .Q(net_4031), .D(net_1349), .CK(net_4708) );
CLKBUF_X2 inst_4483 ( .A(net_4353), .Z(net_4469) );
INV_X4 inst_2470 ( .A(net_2983), .ZN(net_230) );
NAND4_X2 inst_1258 ( .ZN(net_4005), .A1(net_3656), .A4(net_3167), .A3(net_513), .A2(net_359) );
DFF_X2 inst_3141 ( .QN(net_2982), .D(net_2569), .CK(net_5232) );
AOI221_X1 inst_3921 ( .ZN(net_3795), .B1(net_3792), .B2(net_1719), .C1(net_1718), .C2(net_1717), .A(net_1245) );
NAND2_X2 inst_1957 ( .A2(net_3869), .A1(net_3779), .ZN(net_3292) );
CLKBUF_X2 inst_5151 ( .A(net_5136), .Z(net_5137) );
AOI221_X2 inst_3857 ( .B1(net_3736), .C2(net_3118), .C1(net_2115), .ZN(net_2047), .A(net_1937), .B2(net_69) );
NOR2_X2 inst_1060 ( .A1(net_1908), .ZN(net_1568), .A2(net_749) );
NAND2_X4 inst_1419 ( .A1(net_3713), .A2(net_3656), .ZN(net_3568) );
NOR3_X2 inst_900 ( .ZN(net_1091), .A3(net_1090), .A1(net_981), .A2(net_297) );
INV_X2 inst_2661 ( .A(net_3677), .ZN(net_2108) );
CLKBUF_X2 inst_4949 ( .A(net_4934), .Z(net_4935) );
CLKBUF_X2 inst_4624 ( .A(net_4609), .Z(net_4610) );
INV_X4 inst_2501 ( .A(net_3068), .ZN(net_731) );
AOI22_X2 inst_3548 ( .B1(net_4054), .A1(net_1578), .ZN(net_1573), .B2(net_1189), .A2(net_378) );
INV_X2 inst_2807 ( .ZN(net_696), .A(net_695) );
OAI21_X2 inst_594 ( .A(net_3582), .ZN(net_2544), .B2(net_2543), .B1(net_2513) );
CLKBUF_X2 inst_4435 ( .A(net_4420), .Z(net_4421) );
INV_X2 inst_2983 ( .A(net_315), .ZN(net_228) );
NAND2_X2 inst_1632 ( .ZN(net_2326), .A1(net_2270), .A2(net_356) );
INV_X4 inst_2175 ( .ZN(net_2791), .A(net_2790) );
CLKBUF_X2 inst_4241 ( .A(net_4218), .Z(net_4227) );
NOR2_X4 inst_925 ( .ZN(net_2244), .A2(net_2171), .A1(net_2170) );
INV_X4 inst_2193 ( .A(net_2778), .ZN(net_2346) );
INV_X4 inst_2378 ( .ZN(net_523), .A(net_368) );
NOR2_X2 inst_1120 ( .ZN(net_3412), .A1(net_2718), .A2(net_2717) );
NAND2_X2 inst_1536 ( .A1(net_2907), .ZN(net_2486), .A2(net_188) );
NOR3_X4 inst_881 ( .ZN(net_3798), .A1(net_3797), .A3(net_3218), .A2(net_2027) );
AOI221_X2 inst_3876 ( .B2(net_3112), .B1(net_2020), .C1(net_2019), .ZN(net_1871), .A(net_1870), .C2(x332) );
DFF_X2 inst_3184 ( .QN(net_3159), .D(net_1752), .CK(net_4757) );
AOI221_X2 inst_3848 ( .B1(net_3736), .C2(net_3119), .ZN(net_2117), .C1(net_2115), .A(net_1939), .B2(net_68) );
NAND4_X2 inst_1225 ( .ZN(net_856), .A4(net_654), .A3(net_561), .A1(net_484), .A2(net_481) );
NOR2_X4 inst_947 ( .A2(net_3869), .ZN(net_3555), .A1(net_3262) );
OAI21_X2 inst_731 ( .B1(net_984), .A(net_629), .B2(net_628), .ZN(net_579) );
AOI22_X2 inst_3706 ( .B2(net_4124), .A2(net_509), .ZN(net_460), .A1(net_226), .B1(net_167) );
INV_X4 inst_2459 ( .A(net_3056), .ZN(net_474) );
OAI22_X2 inst_301 ( .ZN(net_1544), .A1(net_1543), .B1(net_1542), .B2(net_1541), .A2(net_315) );
OAI221_X2 inst_363 ( .B1(net_4037), .C1(net_3352), .B2(net_3348), .ZN(net_2769), .A(net_2556), .C2(net_2131) );
INV_X8 inst_2141 ( .A(net_3204), .ZN(net_3185) );
OR2_X2 inst_247 ( .ZN(net_2826), .A1(net_2825), .A2(net_2384) );
CLKBUF_X2 inst_4551 ( .A(net_4536), .Z(net_4537) );
CLKBUF_X2 inst_4313 ( .A(net_4298), .Z(net_4299) );
OAI221_X2 inst_403 ( .C2(net_3959), .ZN(net_2140), .C1(net_2119), .B2(net_2118), .B1(net_1894), .A(net_593) );
CLKBUF_X2 inst_4714 ( .A(net_4699), .Z(net_4700) );
CLKBUF_X2 inst_4706 ( .A(net_4590), .Z(net_4692) );
CLKBUF_X2 inst_4348 ( .A(net_4333), .Z(net_4334) );
INV_X2 inst_2728 ( .ZN(net_1438), .A(net_1437) );
NAND2_X2 inst_1588 ( .A1(net_2972), .ZN(net_2431), .A2(net_735) );
AOI221_X2 inst_3801 ( .C1(net_2781), .B1(net_2775), .ZN(net_2774), .A(net_2664), .B2(net_315), .C2(net_251) );
AND2_X4 inst_4177 ( .ZN(net_4131), .A1(net_3104), .A2(net_121) );
INV_X2 inst_2956 ( .A(net_3097), .ZN(net_226) );
CLKBUF_X2 inst_4713 ( .A(net_4698), .Z(net_4699) );
AOI22_X2 inst_3729 ( .ZN(net_4176), .A1(net_4175), .B1(net_2703), .A2(net_132), .B2(net_73) );
OAI221_X2 inst_412 ( .ZN(net_1718), .A(net_1460), .C1(net_1455), .B2(net_1273), .B1(net_1219), .C2(net_1033) );
INV_X4 inst_2516 ( .A(net_3780), .ZN(net_3187) );
INV_X2 inst_2650 ( .A(net_3470), .ZN(net_2291) );
CLKBUF_X2 inst_4508 ( .A(net_4493), .Z(net_4494) );
INV_X8 inst_2155 ( .ZN(net_3556), .A(net_3555) );
NAND2_X2 inst_1506 ( .A1(net_3530), .A2(net_3510), .ZN(net_2708) );
OAI21_X4 inst_464 ( .B1(net_3904), .B2(net_3638), .ZN(net_3602), .A(net_582) );
OAI22_X2 inst_341 ( .ZN(net_3364), .A1(net_3353), .B2(net_3138), .A2(net_1071), .B1(net_1036) );
AOI222_X1 inst_3785 ( .C1(net_3151), .B1(net_2020), .C2(net_1840), .A2(net_1698), .ZN(net_1661), .B2(net_512), .A1(net_272) );
DFF_X2 inst_3189 ( .D(net_1654), .CK(net_4991), .QN(x557) );
DFF_X2 inst_3163 ( .QN(net_3820), .D(net_2140), .CK(net_5283) );
INV_X4 inst_2504 ( .ZN(net_184), .A(net_89) );
INV_X4 inst_2359 ( .ZN(net_527), .A(net_523) );
AOI22_X2 inst_3702 ( .B1(net_4124), .A2(net_3025), .B2(net_3024), .A1(net_509), .ZN(net_466) );
OAI21_X2 inst_684 ( .B1(net_3228), .ZN(net_1445), .A(net_1307), .B2(net_505) );
CLKBUF_X2 inst_4354 ( .A(net_4339), .Z(net_4340) );
DFF_X1 inst_3374 ( .D(net_2259), .QN(net_47), .CK(net_4478) );
CLKBUF_X2 inst_4400 ( .A(net_4361), .Z(net_4386) );
DFF_X2 inst_3177 ( .D(net_1846), .Q(net_84), .CK(net_4996) );
NAND3_X2 inst_1361 ( .ZN(net_3866), .A3(net_3865), .A2(net_3864), .A1(net_3863) );
CLKBUF_X2 inst_4930 ( .A(net_4915), .Z(net_4916) );
DFF_X1 inst_3401 ( .Q(net_3114), .D(net_1538), .CK(net_4470) );
AOI221_X2 inst_3811 ( .B2(net_3145), .A(net_2642), .ZN(net_2595), .C2(net_2594), .B1(net_2591), .C1(net_2589) );
AOI22_X2 inst_3653 ( .ZN(net_682), .A1(net_458), .B1(net_457), .A2(net_208), .B2(net_150) );
CLKBUF_X2 inst_4968 ( .A(net_4953), .Z(net_4954) );
CLKBUF_X2 inst_4463 ( .A(net_4202), .Z(net_4449) );
INV_X4 inst_2208 ( .ZN(net_2248), .A(net_2247) );
NOR2_X2 inst_1138 ( .ZN(net_3765), .A2(net_3477), .A1(net_358) );
AND2_X4 inst_4162 ( .ZN(net_4115), .A1(net_1107), .A2(net_923) );
NAND4_X2 inst_1241 ( .A2(net_3651), .ZN(net_3248), .A1(net_3247), .A4(net_2176), .A3(net_2175) );
NOR2_X2 inst_1038 ( .ZN(net_1224), .A1(net_1089), .A2(net_775) );
CLKBUF_X2 inst_5171 ( .A(net_4390), .Z(net_5157) );
INV_X4 inst_2174 ( .ZN(net_2795), .A(net_2794) );
NOR2_X4 inst_940 ( .ZN(net_3237), .A2(net_2173), .A1(net_2172) );
NOR2_X2 inst_1004 ( .A1(net_2684), .ZN(net_2060), .A2(net_1905) );
DFF_X2 inst_3201 ( .D(net_1592), .QN(net_120), .CK(net_4988) );
AOI22_X2 inst_3595 ( .A1(net_4063), .B1(net_4058), .B2(net_3402), .A2(net_3401), .ZN(net_1422) );
OR2_X4 inst_189 ( .A2(net_2607), .ZN(net_2579), .A1(net_2578) );
CLKBUF_X2 inst_4876 ( .A(net_4861), .Z(net_4862) );
XOR2_X2 inst_14 ( .A(net_1125), .B(net_1101), .Z(net_1088) );
INV_X4 inst_2450 ( .A(net_3060), .ZN(net_734) );
CLKBUF_X2 inst_4362 ( .A(net_4347), .Z(net_4348) );
XNOR2_X2 inst_62 ( .ZN(net_1903), .A(net_1754), .B(net_1660) );
INV_X4 inst_2325 ( .A(net_3547), .ZN(net_700) );
CLKBUF_X2 inst_4696 ( .A(net_4681), .Z(net_4682) );
CLKBUF_X2 inst_4369 ( .A(net_4354), .Z(net_4355) );
AOI222_X1 inst_3743 ( .A1(net_4189), .C1(net_3504), .B1(net_3472), .ZN(net_2318), .A2(net_1791), .C2(net_920), .B2(net_142) );
OR2_X2 inst_251 ( .A2(net_4131), .ZN(net_1927), .A1(net_1808) );
INV_X2 inst_2860 ( .A(net_3165), .ZN(net_297) );
CLKBUF_X2 inst_5194 ( .A(net_4524), .Z(net_5180) );
NOR2_X2 inst_1074 ( .ZN(net_694), .A1(net_693), .A2(net_639) );
NOR3_X4 inst_879 ( .A2(net_3946), .A3(net_3940), .ZN(net_3725), .A1(net_3108) );
AOI21_X2 inst_4007 ( .ZN(net_4158), .B2(net_3110), .A(net_2273), .B1(net_2241) );
NAND2_X2 inst_1552 ( .A1(net_2961), .ZN(net_2470), .A2(net_461) );
NAND2_X2 inst_1524 ( .A1(net_2959), .ZN(net_2498), .A2(net_833) );
CLKBUF_X2 inst_4789 ( .A(net_4774), .Z(net_4775) );
CLKBUF_X2 inst_4977 ( .A(net_4962), .Z(net_4963) );
CLKBUF_X2 inst_4482 ( .A(net_4467), .Z(net_4468) );
CLKBUF_X2 inst_4291 ( .A(net_4198), .Z(net_4277) );
NAND2_X2 inst_1602 ( .A1(net_2969), .ZN(net_2415), .A2(net_493) );
NOR2_X4 inst_969 ( .ZN(net_3877), .A1(net_3232), .A2(net_2207) );
CLKBUF_X2 inst_4903 ( .A(net_4888), .Z(net_4889) );
OAI21_X2 inst_629 ( .B2(net_4089), .B1(net_2190), .ZN(net_2146), .A(net_2035) );
NOR2_X2 inst_1100 ( .A2(net_3108), .ZN(net_277), .A1(net_218) );
INV_X4 inst_2528 ( .ZN(net_3275), .A(net_647) );
OAI211_X2 inst_791 ( .C1(net_3449), .ZN(net_2705), .C2(net_2704), .A(net_2605), .B(net_2526) );
NAND2_X2 inst_2021 ( .ZN(net_3693), .A1(net_3688), .A2(net_70) );
CLKBUF_X2 inst_4917 ( .A(net_4902), .Z(net_4903) );
CLKBUF_X2 inst_4379 ( .A(net_4364), .Z(net_4365) );
NOR3_X2 inst_898 ( .ZN(net_1223), .A1(net_1222), .A2(net_1158), .A3(net_1081) );
DFF_X1 inst_3383 ( .D(net_1887), .QN(net_82), .CK(net_4433) );
NAND2_X2 inst_1977 ( .A1(net_3804), .ZN(net_3370), .A2(net_3268) );
NAND2_X2 inst_1793 ( .A1(net_3905), .A2(net_1105), .ZN(net_1074) );
NAND4_X2 inst_1191 ( .A2(net_4053), .A3(net_1776), .A1(net_1634), .ZN(net_1633), .A4(net_1382) );
CLKBUF_X2 inst_4227 ( .A(net_4212), .Z(net_4213) );
CLKBUF_X2 inst_5086 ( .A(net_4405), .Z(net_5072) );
OAI21_X2 inst_533 ( .B1(net_3195), .B2(net_2967), .ZN(net_2900), .A(net_2410) );
INV_X4 inst_2478 ( .A(net_3081), .ZN(net_468) );
CLKBUF_X2 inst_5299 ( .A(net_5284), .Z(net_5285) );
CLKBUF_X2 inst_4972 ( .A(net_4400), .Z(net_4958) );
INV_X2 inst_2751 ( .A(net_1330), .ZN(net_1077) );
NAND2_X2 inst_1874 ( .A2(net_3959), .ZN(net_508), .A1(net_276) );
NAND2_X2 inst_1760 ( .A2(net_1394), .ZN(net_1239), .A1(net_37) );
INV_X4 inst_2291 ( .ZN(net_1694), .A(net_868) );
INV_X4 inst_2343 ( .ZN(net_611), .A(net_610) );
INV_X4 inst_2538 ( .ZN(net_3379), .A(net_3378) );
NAND2_X2 inst_2022 ( .ZN(net_3704), .A1(net_2357), .A2(net_1889) );
CLKBUF_X2 inst_4822 ( .A(net_4363), .Z(net_4808) );
INV_X2 inst_2821 ( .A(net_658), .ZN(net_539) );
DFF_X2 inst_3132 ( .D(net_2631), .QN(net_987), .CK(net_4812) );
AOI21_X2 inst_3960 ( .ZN(net_1711), .A(net_1561), .B1(net_433), .B2(net_168) );
NOR2_X2 inst_1095 ( .A2(net_4131), .ZN(net_360), .A1(net_178) );
OR3_X4 inst_176 ( .ZN(net_1274), .A2(net_312), .A1(net_266), .A3(net_263) );
INV_X4 inst_2439 ( .A(net_2988), .ZN(net_197) );
CLKBUF_X2 inst_4999 ( .A(net_4984), .Z(net_4985) );
INV_X2 inst_2826 ( .A(net_3941), .ZN(net_599) );
AOI221_X2 inst_3910 ( .B2(net_3998), .A(net_3325), .ZN(net_783), .C1(net_655), .B1(net_528), .C2(net_377) );
NAND3_X2 inst_1336 ( .A2(net_1401), .ZN(net_1126), .A1(net_406), .A3(net_263) );
NAND3_X2 inst_1332 ( .ZN(net_504), .A1(net_405), .A3(net_374), .A2(net_310) );
CLKBUF_X2 inst_4404 ( .A(net_4389), .Z(net_4390) );
NAND2_X2 inst_1841 ( .A2(net_3590), .ZN(net_843), .A1(net_788) );
CLKBUF_X2 inst_4500 ( .A(net_4485), .Z(net_4486) );
NAND2_X2 inst_1665 ( .ZN(net_2097), .A1(net_2096), .A2(net_195) );
DFF_X1 inst_3345 ( .D(net_2744), .QN(net_115), .CK(net_4448) );
CLKBUF_X2 inst_4763 ( .A(net_4748), .Z(net_4749) );
DFF_X1 inst_3264 ( .QN(net_3072), .D(net_2932), .CK(net_4721) );
CLKBUF_X2 inst_5169 ( .A(net_5154), .Z(net_5155) );
CLKBUF_X2 inst_4945 ( .A(net_4338), .Z(net_4931) );
OAI211_X2 inst_780 ( .C2(net_3348), .ZN(net_2841), .C1(net_2828), .B(net_2614), .A(net_2566) );
INV_X4 inst_2332 ( .A(net_3955), .ZN(net_674) );
AOI21_X2 inst_3967 ( .A(net_2525), .ZN(net_1364), .B1(net_1179), .B2(net_1175) );
INV_X4 inst_2310 ( .ZN(net_966), .A(net_791) );
NOR2_X2 inst_1089 ( .A1(net_3756), .ZN(net_424), .A2(net_373) );
AOI211_X2 inst_4018 ( .A(net_4185), .B(net_4083), .ZN(net_1810), .C1(net_1567), .C2(net_1045) );
NAND2_X2 inst_1767 ( .ZN(net_1627), .A2(net_1386), .A1(net_1232) );
AOI22_X2 inst_3669 ( .B1(net_570), .ZN(net_556), .A1(net_555), .B2(net_217), .A2(net_159) );
INV_X4 inst_2219 ( .ZN(net_2227), .A(net_2190) );
NAND3_X2 inst_1284 ( .A3(net_3127), .ZN(net_2297), .A1(net_2296), .A2(net_248) );
OAI21_X2 inst_546 ( .B2(net_2915), .B1(net_2887), .ZN(net_2885), .A(net_2438) );
INV_X4 inst_2465 ( .A(net_3092), .ZN(net_833) );
CLKBUF_X2 inst_5017 ( .A(net_4198), .Z(net_5003) );
INV_X4 inst_2361 ( .A(net_2514), .ZN(x475) );
NAND3_X2 inst_1290 ( .ZN(net_2257), .A1(net_2205), .A3(net_1951), .A2(net_1924) );
OAI21_X2 inst_704 ( .B2(net_3974), .ZN(net_893), .B1(net_754), .A(net_640) );
CLKBUF_X2 inst_5038 ( .A(net_5023), .Z(net_5024) );
CLKBUF_X2 inst_4542 ( .A(net_4527), .Z(net_4528) );
CLKBUF_X2 inst_5142 ( .A(net_5127), .Z(net_5128) );
INV_X4 inst_2226 ( .A(net_3428), .ZN(net_2049) );
OAI21_X2 inst_694 ( .B2(net_3123), .ZN(net_1330), .B1(net_822), .A(net_814) );
CLKBUF_X2 inst_4899 ( .A(net_4884), .Z(net_4885) );
NAND2_X2 inst_2046 ( .A1(net_3875), .A2(net_3859), .ZN(net_3850) );
CLKBUF_X2 inst_5079 ( .A(net_5064), .Z(net_5065) );
AND2_X4 inst_4129 ( .ZN(net_4056), .A2(net_3339), .A1(net_1247) );
INV_X4 inst_2498 ( .A(net_3164), .ZN(net_223) );
DFF_X2 inst_3154 ( .D(net_2260), .QN(net_46), .CK(net_4629) );
AOI221_X2 inst_3861 ( .B2(net_3120), .ZN(net_2021), .B1(net_2020), .C1(net_2019), .A(net_1899), .C2(x285) );
CLKBUF_X2 inst_4399 ( .A(net_4384), .Z(net_4385) );
CLKBUF_X2 inst_5211 ( .A(net_5196), .Z(net_5197) );
NAND3_X2 inst_1342 ( .A1(net_3782), .ZN(net_3407), .A3(net_3406), .A2(net_1376) );
INV_X2 inst_2971 ( .A(net_3043), .ZN(net_163) );
AND2_X2 inst_4196 ( .A2(net_2222), .ZN(net_1870), .A1(net_1862) );
AOI22_X2 inst_3524 ( .A2(net_3132), .A1(net_1923), .B1(net_1921), .ZN(net_1920), .B2(net_218) );
CLKBUF_X2 inst_4479 ( .A(net_4389), .Z(net_4465) );
CLKBUF_X2 inst_4396 ( .A(net_4293), .Z(net_4382) );
NOR2_X2 inst_1014 ( .A1(net_3486), .ZN(net_1867), .A2(net_1738) );
OAI211_X2 inst_787 ( .ZN(net_2760), .C2(net_2709), .B(net_2649), .A(net_2635), .C1(net_2603) );
INV_X4 inst_2531 ( .A(net_3618), .ZN(net_3290) );
CLKBUF_X2 inst_4549 ( .A(net_4534), .Z(net_4535) );
CLKBUF_X2 inst_4782 ( .A(net_4767), .Z(net_4768) );
AOI21_X2 inst_3933 ( .B2(net_3111), .ZN(net_2796), .B1(net_2792), .A(net_2745) );
NAND3_X2 inst_1347 ( .ZN(net_3476), .A3(net_3475), .A2(net_3474), .A1(net_3473) );
OAI211_X2 inst_825 ( .ZN(net_1464), .C2(net_1463), .A(net_1228), .C1(net_1036), .B(net_593) );
NAND2_X2 inst_1656 ( .A1(net_3200), .ZN(net_2112), .A2(net_1981) );
OAI21_X2 inst_509 ( .B1(net_3274), .B2(net_2965), .ZN(net_2933), .A(net_2443) );
INV_X4 inst_2586 ( .ZN(net_3655), .A(net_3653) );
INV_X2 inst_2687 ( .ZN(net_1788), .A(net_1708) );
NAND2_X2 inst_1680 ( .A1(net_3281), .ZN(net_2028), .A2(net_214) );
NAND2_X2 inst_1881 ( .ZN(net_891), .A1(net_413), .A2(net_335) );
NAND2_X2 inst_1626 ( .ZN(net_2601), .A2(net_2596), .A1(net_2389) );
INV_X4 inst_2622 ( .ZN(net_3953), .A(net_3913) );
SDFF_X2 inst_153 ( .SE(net_2218), .D(net_1610), .SI(net_211), .QN(net_55), .CK(net_4785) );
CLKBUF_X2 inst_4856 ( .A(net_4706), .Z(net_4842) );
NAND2_X2 inst_1892 ( .ZN(net_421), .A1(net_394), .A2(net_393) );
INV_X2 inst_3034 ( .A(net_3660), .ZN(net_3571) );
NAND2_X4 inst_1459 ( .A1(net_4152), .ZN(net_3858), .A2(net_1266) );
OAI21_X2 inst_726 ( .B1(net_3657), .A(net_3215), .ZN(net_602), .B2(net_320) );
OAI22_X2 inst_295 ( .A2(net_4034), .ZN(net_1704), .A1(net_1653), .B1(net_1165), .B2(net_1090) );
AND2_X4 inst_4094 ( .ZN(net_1955), .A2(net_1828), .A1(net_1827) );
OR2_X4 inst_209 ( .ZN(net_2327), .A1(net_2303), .A2(net_2214) );
AOI221_X2 inst_3894 ( .C2(net_4028), .A(net_2525), .C1(net_1394), .B1(net_1393), .ZN(net_1348), .B2(net_1326) );
CLKBUF_X2 inst_4726 ( .A(net_4711), .Z(net_4712) );
NOR2_X2 inst_1087 ( .ZN(net_584), .A1(net_394), .A2(net_393) );
NAND2_X2 inst_1781 ( .ZN(net_1300), .A2(net_1064), .A1(net_1063) );
OAI22_X2 inst_320 ( .B1(net_1614), .ZN(net_1070), .A1(net_1069), .A2(net_729), .B2(net_260) );
OAI21_X2 inst_607 ( .A(net_3886), .B1(net_3883), .B2(net_3516), .ZN(net_2329) );
INV_X2 inst_2769 ( .A(net_3573), .ZN(net_888) );
INV_X4 inst_2432 ( .A(net_2993), .ZN(net_181) );
NAND3_X2 inst_1375 ( .ZN(net_4192), .A2(net_3383), .A1(net_3382), .A3(net_1291) );
CLKBUF_X2 inst_4263 ( .A(net_4248), .Z(net_4249) );
CLKBUF_X2 inst_5061 ( .A(net_5046), .Z(net_5047) );
XOR2_X2 inst_1 ( .Z(net_2304), .A(net_2152), .B(net_1736) );
NAND2_X2 inst_1891 ( .A2(net_3590), .ZN(net_411), .A1(net_398) );
AOI21_X2 inst_3982 ( .B2(net_4144), .B1(net_3627), .ZN(net_946), .A(net_885) );
CLKBUF_X2 inst_4343 ( .A(net_4328), .Z(net_4329) );
CLKBUF_X2 inst_4564 ( .A(net_4549), .Z(net_4550) );
CLKBUF_X2 inst_4558 ( .A(net_4543), .Z(net_4544) );
CLKBUF_X2 inst_5258 ( .A(net_5243), .Z(net_5244) );
DFF_X2 inst_3215 ( .QN(net_3152), .D(net_803), .CK(net_4663) );
OR2_X4 inst_235 ( .ZN(net_3207), .A1(net_3206), .A2(net_2354) );
INV_X16 inst_3063 ( .A(net_3293), .ZN(net_1973) );
INV_X4 inst_2564 ( .ZN(net_3519), .A(net_2094) );
NAND2_X2 inst_1812 ( .A2(net_4120), .ZN(net_914), .A1(net_747) );
NOR2_X2 inst_1082 ( .ZN(net_585), .A2(net_584), .A1(net_422) );
AND2_X4 inst_4167 ( .ZN(net_4121), .A1(net_3160), .A2(net_3159) );
INV_X2 inst_2677 ( .ZN(net_1887), .A(net_1842) );
CLKBUF_X2 inst_4374 ( .A(net_4359), .Z(net_4360) );
NAND2_X2 inst_1995 ( .ZN(net_3480), .A1(net_2563), .A2(net_2003) );
XNOR2_X2 inst_105 ( .ZN(net_616), .A(net_309), .B(net_48) );
CLKBUF_X2 inst_4338 ( .A(net_4248), .Z(net_4324) );
AOI22_X2 inst_3518 ( .B1(net_4045), .B2(net_2051), .A1(net_1955), .ZN(net_1952), .A2(net_280) );
INV_X8 inst_2161 ( .ZN(net_3647), .A(net_3645) );
OAI21_X2 inst_625 ( .B2(net_4061), .ZN(net_2243), .A(net_2142), .B1(net_2127) );
CLKBUF_X2 inst_4721 ( .A(net_4706), .Z(net_4707) );
DFF_X1 inst_3367 ( .D(net_3697), .CK(net_4445), .Q(x256) );
INV_X2 inst_2835 ( .ZN(net_422), .A(net_421) );
OAI21_X2 inst_568 ( .B2(net_2907), .B1(net_2849), .ZN(net_2844), .A(net_2486) );
NAND2_X4 inst_1483 ( .ZN(net_3992), .A1(net_3991), .A2(net_3987) );
OAI21_X2 inst_523 ( .B2(net_2969), .B1(net_2923), .ZN(net_2914), .A(net_2412) );
INV_X2 inst_2731 ( .ZN(net_1396), .A(net_1348) );
INV_X4 inst_2207 ( .ZN(net_2252), .A(net_2224) );
NAND2_X2 inst_1492 ( .A1(net_3499), .ZN(net_2858), .A2(net_2630) );
OR3_X2 inst_181 ( .ZN(net_1721), .A3(net_1617), .A1(net_1587), .A2(net_1586) );
CLKBUF_X2 inst_5215 ( .A(net_4937), .Z(net_5201) );
CLKBUF_X2 inst_4234 ( .A(net_4219), .Z(net_4220) );
CLKBUF_X2 inst_4813 ( .A(net_4678), .Z(net_4799) );
AOI221_X2 inst_3892 ( .B2(net_2051), .C2(net_1394), .B1(net_1393), .ZN(net_1355), .A(net_1173), .C1(net_36) );
OAI21_X2 inst_713 ( .B2(net_874), .ZN(net_816), .A(net_815), .B1(net_616) );
AOI21_X4 inst_3930 ( .B2(net_3889), .B1(net_3838), .ZN(net_3700), .A(net_3567) );
INV_X2 inst_2867 ( .A(net_393), .ZN(net_329) );
INV_X2 inst_2898 ( .ZN(net_182), .A(net_114) );
OAI21_X2 inst_477 ( .ZN(net_2973), .B2(net_2972), .B1(net_2970), .A(net_2430) );
DFF_X1 inst_3398 ( .Q(net_3121), .D(net_1546), .CK(net_4306) );
NAND3_X2 inst_1368 ( .ZN(net_3989), .A3(net_3988), .A1(net_640), .A2(net_432) );
AOI22_X2 inst_3576 ( .A1(net_4060), .B1(net_4055), .ZN(net_1474), .B2(net_834), .A2(net_833) );
OAI221_X2 inst_423 ( .B1(net_3963), .B2(net_3338), .C2(net_3162), .ZN(net_1157), .A(net_1031), .C1(x475) );
OAI211_X2 inst_835 ( .C2(net_2637), .C1(net_1359), .ZN(net_1356), .A(net_1236), .B(net_593) );
NAND2_X1 inst_2088 ( .A2(net_4017), .A1(net_2969), .ZN(net_2419) );
DFF_X1 inst_3305 ( .QN(net_3019), .D(net_2869), .CK(net_5080) );
INV_X1 inst_3082 ( .ZN(net_3549), .A(net_3548) );
AND2_X4 inst_4137 ( .ZN(net_4066), .A1(net_2596), .A2(net_1032) );
DFF_X2 inst_3208 ( .QN(net_3162), .D(net_1157), .CK(net_5088) );
AND2_X4 inst_4134 ( .ZN(net_4063), .A2(net_1192), .A1(net_1136) );
NOR2_X2 inst_1112 ( .ZN(net_3327), .A2(net_3319), .A1(net_605) );
AOI22_X2 inst_3507 ( .B1(net_3676), .B2(net_3141), .A1(net_2012), .ZN(net_2010), .A2(net_379) );
OAI21_X2 inst_710 ( .ZN(net_1013), .A(net_750), .B1(net_725), .B2(net_526) );
AND3_X4 inst_4081 ( .ZN(net_4185), .A2(net_3571), .A1(net_618), .A3(net_594) );
NAND3_X1 inst_1379 ( .ZN(net_3350), .A2(net_3349), .A1(net_2550), .A3(net_1737) );
NOR2_X4 inst_941 ( .A1(net_3550), .ZN(net_3276), .A2(net_1457) );
OR2_X2 inst_271 ( .ZN(net_3771), .A2(net_2053), .A1(net_1808) );
DFF_X1 inst_3350 ( .D(net_2702), .QN(net_70), .CK(net_4267) );
NAND2_X2 inst_1817 ( .ZN(net_831), .A2(net_819), .A1(net_204) );
XNOR2_X2 inst_56 ( .B(net_3240), .ZN(net_2193), .A(net_2121) );
OAI22_X2 inst_308 ( .A2(net_1975), .A1(net_1461), .ZN(net_1333), .B1(net_1332), .B2(net_1200) );
NAND2_X2 inst_1546 ( .A2(net_4023), .A1(net_2961), .ZN(net_2476) );
NAND4_X2 inst_1230 ( .ZN(net_2222), .A4(net_565), .A1(net_546), .A2(net_500), .A3(net_482) );
OAI21_X4 inst_455 ( .B1(net_3673), .A(net_3430), .ZN(net_1457), .B2(net_1272) );
AOI22_X2 inst_3535 ( .A2(net_1908), .ZN(net_1770), .A1(net_1676), .B2(net_749), .B1(net_103) );
NAND2_X2 inst_1694 ( .A1(net_3293), .ZN(net_1976), .A2(net_202) );
INV_X2 inst_2871 ( .ZN(net_284), .A(net_109) );
INV_X4 inst_2540 ( .ZN(net_3397), .A(net_3109) );
AOI22_X2 inst_3497 ( .B1(net_3219), .ZN(net_2176), .A1(net_2134), .A2(net_597), .B2(net_596) );
NOR2_X2 inst_1064 ( .A2(net_3627), .ZN(net_885), .A1(net_511) );
AOI22_X2 inst_3629 ( .ZN(net_1638), .B1(net_931), .A1(net_800), .A2(net_401), .B2(net_267) );
AOI22_X2 inst_3599 ( .A1(net_4063), .B1(net_4058), .ZN(net_1418), .A2(net_237), .B2(net_157) );
INV_X2 inst_3024 ( .ZN(net_3459), .A(net_3458) );
OAI21_X2 inst_583 ( .B1(net_4036), .B2(net_2815), .ZN(net_2777), .A(net_1576) );
NAND2_X2 inst_1904 ( .A2(net_3166), .ZN(net_374), .A1(net_309) );
CLKBUF_X2 inst_5208 ( .A(net_5193), .Z(net_5194) );
AOI22_X2 inst_3581 ( .A1(net_4059), .B1(net_4056), .A2(net_4019), .B2(net_4017), .ZN(net_1469) );
CLKBUF_X2 inst_4414 ( .A(net_4399), .Z(net_4400) );
CLKBUF_X2 inst_4325 ( .A(net_4310), .Z(net_4311) );
CLKBUF_X2 inst_4833 ( .A(net_4818), .Z(net_4819) );
NAND2_X2 inst_2065 ( .ZN(net_3946), .A2(net_3124), .A1(net_3107) );
INV_X4 inst_2251 ( .A(net_4192), .ZN(net_1502) );
INV_X1 inst_3085 ( .ZN(net_3981), .A(net_3980) );
AOI21_X2 inst_3987 ( .A(net_4185), .B2(net_923), .ZN(net_792), .B1(net_692) );
AOI21_X2 inst_3951 ( .B1(net_3736), .ZN(net_1990), .A(net_1856), .B2(net_1439) );
CLKBUF_X2 inst_5124 ( .A(net_5109), .Z(net_5110) );
CLKBUF_X2 inst_4282 ( .A(net_4234), .Z(net_4268) );
CLKBUF_X2 inst_4863 ( .A(net_4848), .Z(net_4849) );
CLKBUF_X2 inst_4910 ( .A(net_4895), .Z(net_4896) );
NAND2_X2 inst_1899 ( .ZN(net_365), .A1(net_291), .A2(net_288) );
INV_X2 inst_2943 ( .A(net_3017), .ZN(net_140) );
NAND2_X2 inst_1593 ( .A1(net_2925), .ZN(net_2425), .A2(net_174) );
INV_X4 inst_2569 ( .ZN(net_3540), .A(net_3129) );
OAI21_X2 inst_724 ( .B2(net_1217), .ZN(net_620), .A(net_619), .B1(net_406) );
CLKBUF_X2 inst_4292 ( .A(net_4277), .Z(net_4278) );
INV_X2 inst_2716 ( .A(net_3802), .ZN(net_1772) );
INV_X4 inst_2449 ( .ZN(net_2623), .A(net_66) );
DFF_X1 inst_3228 ( .QN(net_3069), .D(net_2973), .CK(net_4882) );
NOR2_X4 inst_975 ( .A2(net_3997), .ZN(net_3932), .A1(net_3668) );
INV_X8 inst_2124 ( .A(net_3606), .ZN(net_399) );
INV_X2 inst_2789 ( .ZN(net_1253), .A(net_1131) );
DFF_X2 inst_3191 ( .QN(net_3163), .D(net_1697), .CK(net_5092) );
INV_X4 inst_2289 ( .ZN(net_1100), .A(net_880) );
NAND2_X4 inst_1435 ( .ZN(net_3674), .A1(net_3541), .A2(net_3270) );
NAND2_X4 inst_1431 ( .ZN(net_3660), .A1(net_3603), .A2(net_3243) );
AOI222_X1 inst_3760 ( .A2(net_3466), .C1(net_3119), .A1(net_2055), .B1(net_2054), .C2(net_2053), .ZN(net_2002), .B2(net_1468) );
NAND2_X4 inst_1398 ( .A1(net_3228), .ZN(net_1307), .A2(net_231) );
AOI222_X1 inst_3746 ( .C1(net_3504), .B1(net_3472), .A1(net_3469), .A2(net_3134), .ZN(net_2278), .B2(net_2051), .C2(net_874) );
NAND2_X2 inst_1804 ( .A1(net_4082), .ZN(net_1069), .A2(net_847) );
INV_X2 inst_2750 ( .A(net_2384), .ZN(net_1319) );
INV_X2 inst_2849 ( .ZN(net_375), .A(net_356) );
INV_X4 inst_2440 ( .A(net_3163), .ZN(net_144) );
AND2_X4 inst_4121 ( .ZN(net_4044), .A1(net_1875), .A2(net_1874) );
NAND2_X4 inst_1467 ( .ZN(net_3892), .A2(net_3716), .A1(net_3276) );
INV_X2 inst_2640 ( .ZN(net_2731), .A(net_2581) );
INV_X4 inst_2183 ( .ZN(net_2722), .A(net_2565) );
DFF_X1 inst_3327 ( .Q(net_3115), .D(net_2810), .CK(net_4371) );
CLKBUF_X2 inst_5068 ( .A(net_4589), .Z(net_5054) );
CLKBUF_X2 inst_4448 ( .A(net_4304), .Z(net_4434) );
INV_X2 inst_2659 ( .ZN(net_2113), .A(net_2039) );
INV_X8 inst_2134 ( .A(net_283), .ZN(net_279) );
NAND2_X2 inst_1744 ( .A2(net_1507), .A1(net_1441), .ZN(net_1436) );
CLKBUF_X2 inst_5018 ( .A(net_5003), .Z(net_5004) );
CLKBUF_X2 inst_4805 ( .A(net_4790), .Z(net_4791) );
INV_X2 inst_2834 ( .A(net_3156), .ZN(net_2514) );
CLKBUF_X2 inst_4784 ( .A(net_4769), .Z(net_4770) );
AND2_X4 inst_4117 ( .ZN(net_4035), .A1(net_2735), .A2(net_2694) );
NAND2_X2 inst_1513 ( .A2(net_4066), .ZN(net_2718), .A1(net_2612) );
NOR2_X2 inst_1155 ( .ZN(net_4057), .A2(net_1192), .A1(net_1191) );
OR2_X4 inst_207 ( .A1(net_3816), .ZN(net_2925), .A2(net_2354) );
DFF_X1 inst_3321 ( .QN(net_3000), .D(net_2846), .CK(net_5111) );
AND3_X4 inst_4080 ( .ZN(net_4162), .A1(net_3662), .A2(net_3642), .A3(net_3108) );
NAND2_X2 inst_1545 ( .A2(net_3402), .A1(net_3207), .ZN(net_2477) );
OAI22_X2 inst_333 ( .ZN(net_714), .A1(net_344), .B2(net_263), .B1(net_48), .A2(net_46) );
DFF_X1 inst_3338 ( .D(net_2763), .CK(net_4362), .Q(x0) );
OAI21_X2 inst_712 ( .ZN(net_1064), .B1(net_843), .A(net_842), .B2(net_669) );
NAND4_X2 inst_1215 ( .A1(net_2596), .ZN(net_1275), .A4(net_1126), .A2(net_960), .A3(net_406) );
CLKBUF_X2 inst_5279 ( .A(net_5264), .Z(net_5265) );
SDFF_X2 inst_131 ( .D(net_3483), .SI(net_3025), .Q(net_3025), .SE(net_2919), .CK(net_4892) );
OAI221_X2 inst_406 ( .ZN(net_2553), .A(net_1728), .B1(net_1614), .C1(net_1613), .B2(net_327), .C2(net_192) );
CLKBUF_X2 inst_4579 ( .A(net_4337), .Z(net_4565) );
OAI22_X2 inst_328 ( .ZN(net_880), .B2(net_721), .A1(net_641), .A2(net_329), .B1(net_42) );
DFF_X2 inst_3111 ( .QN(net_2992), .D(net_2800), .CK(net_5244) );
NAND2_X2 inst_2035 ( .ZN(net_3773), .A2(net_1845), .A1(net_1806) );
XNOR2_X2 inst_47 ( .B(net_3175), .ZN(net_2688), .A(net_2372) );
CLKBUF_X2 inst_4217 ( .A(net_4202), .Z(net_4203) );
INV_X2 inst_2764 ( .ZN(net_2131), .A(net_952) );
OAI211_X2 inst_818 ( .A(net_3487), .ZN(net_1799), .B(net_935), .C1(net_433), .C2(net_287) );
CLKBUF_X2 inst_5231 ( .A(net_4986), .Z(net_5217) );
NAND2_X2 inst_1984 ( .A1(net_3782), .ZN(net_3408), .A2(net_1376) );
AND2_X4 inst_4101 ( .A1(net_4081), .ZN(net_1155), .A2(net_686) );
DFF_X2 inst_3178 ( .QN(net_3166), .D(net_1830), .CK(net_4677) );
DFF_X1 inst_3274 ( .QN(net_3101), .D(net_2921), .CK(net_5086) );
AND2_X2 inst_4203 ( .A2(net_3344), .ZN(net_3269), .A1(net_3268) );
CLKBUF_X2 inst_4792 ( .A(net_4664), .Z(net_4778) );
INV_X2 inst_2840 ( .A(net_3395), .ZN(net_400) );
OAI21_X2 inst_525 ( .B2(net_2967), .B1(net_2923), .ZN(net_2911), .A(net_2404) );
INV_X2 inst_2781 ( .ZN(net_805), .A(net_759) );
OAI221_X2 inst_434 ( .C2(net_3468), .A(net_629), .B1(net_628), .C1(net_627), .ZN(net_625), .B2(net_402) );
NOR2_X2 inst_1032 ( .ZN(net_1505), .A1(net_1440), .A2(net_1439) );
NOR3_X2 inst_906 ( .A2(net_3984), .ZN(net_684), .A1(net_658), .A3(net_528) );
CLKBUF_X2 inst_4276 ( .A(net_4261), .Z(net_4262) );
CLKBUF_X2 inst_5222 ( .A(net_5207), .Z(net_5208) );
CLKBUF_X2 inst_5098 ( .A(net_4886), .Z(net_5084) );
NAND4_X2 inst_1248 ( .ZN(net_3611), .A4(net_3610), .A3(net_3609), .A2(net_3608), .A1(net_3607) );
INV_X4 inst_2598 ( .ZN(net_3746), .A(net_2876) );
INV_X4 inst_2402 ( .ZN(net_655), .A(net_359) );
NAND2_X4 inst_1392 ( .A1(net_3187), .ZN(net_2106), .A2(net_165) );
INV_X4 inst_2616 ( .A(net_3896), .ZN(net_3868) );
AND4_X4 inst_4044 ( .ZN(net_4050), .A1(net_1375), .A3(net_1209), .A2(net_1187), .A4(net_1019) );
NAND2_X4 inst_1476 ( .ZN(net_3939), .A1(net_3167), .A2(net_3109) );
INV_X4 inst_2249 ( .A(net_1459), .ZN(net_1378) );
AOI21_X2 inst_3998 ( .B1(net_3620), .ZN(net_3598), .B2(net_1636), .A(net_441) );
CLKBUF_X2 inst_4300 ( .A(net_4243), .Z(net_4286) );
MUX2_X2 inst_2113 ( .B(net_3133), .A(net_2222), .S(net_1071), .Z(net_868) );
CLKBUF_X2 inst_5249 ( .A(net_5234), .Z(net_5235) );
NAND2_X2 inst_1820 ( .A1(net_4098), .ZN(net_860), .A2(net_594) );
INV_X4 inst_2269 ( .ZN(net_1691), .A(net_1021) );
NAND2_X2 inst_1780 ( .A2(net_4109), .A1(net_1202), .ZN(net_1065) );
INV_X4 inst_2390 ( .ZN(net_366), .A(net_365) );
NAND2_X4 inst_1436 ( .A2(net_3819), .ZN(net_3679), .A1(net_3667) );
OR3_X2 inst_183 ( .A3(net_3968), .A2(net_3621), .A1(net_1058), .ZN(net_858) );
OAI211_X2 inst_852 ( .ZN(net_3321), .C1(net_3318), .A(net_3246), .B(net_1299), .C2(net_359) );
AOI221_X2 inst_3871 ( .B2(net_3113), .B1(net_2020), .C1(net_2019), .ZN(net_1933), .A(net_1858), .C2(x142) );
CLKBUF_X2 inst_4306 ( .A(net_4291), .Z(net_4292) );
CLKBUF_X2 inst_4729 ( .A(net_4655), .Z(net_4715) );
CLKBUF_X2 inst_4449 ( .A(net_4434), .Z(net_4435) );
NAND2_X4 inst_1474 ( .A1(net_3944), .ZN(net_3928), .A2(net_392) );
INV_X4 inst_2271 ( .ZN(net_1257), .A(net_1203) );
NAND2_X2 inst_2045 ( .ZN(net_3854), .A2(net_3853), .A1(net_3850) );
NAND2_X2 inst_1920 ( .A2(net_3161), .ZN(net_269), .A1(net_84) );
AOI222_X1 inst_3779 ( .ZN(net_1796), .A1(net_1795), .B1(net_1794), .C1(net_1793), .A2(net_641), .C2(net_379), .B2(net_284) );
NAND2_X2 inst_1848 ( .A2(net_838), .ZN(net_699), .A1(net_535) );
CLKBUF_X2 inst_4451 ( .A(net_4436), .Z(net_4437) );
NAND3_X2 inst_1311 ( .A1(net_2596), .A3(net_1717), .ZN(net_1030), .A2(net_921) );
OAI21_X2 inst_697 ( .A(net_1011), .ZN(net_953), .B1(net_789), .B2(net_614) );
DFF_X1 inst_3415 ( .Q(net_4032), .D(net_1352), .CK(net_4703) );
OAI21_X2 inst_487 ( .B1(net_3394), .B2(net_2972), .ZN(net_2955), .A(net_2428) );
CLKBUF_X2 inst_5159 ( .A(net_5144), .Z(net_5145) );
CLKBUF_X2 inst_4654 ( .A(net_4639), .Z(net_4640) );
NAND2_X2 inst_1640 ( .A1(net_4148), .ZN(net_3212), .A2(net_2105) );
AND2_X4 inst_4143 ( .ZN(net_4079), .A2(net_923), .A1(net_723) );
DFF_X1 inst_3234 ( .QN(net_3062), .D(net_2962), .CK(net_4872) );
CLKBUF_X2 inst_4747 ( .A(net_4438), .Z(net_4733) );
INV_X2 inst_2639 ( .ZN(net_2381), .A(net_2380) );
INV_X8 inst_2133 ( .A(net_3167), .ZN(net_268) );
CLKBUF_X2 inst_4630 ( .A(net_4615), .Z(net_4616) );
INV_X8 inst_2163 ( .ZN(net_3664), .A(net_3663) );
INV_X4 inst_2509 ( .ZN(net_619), .A(net_270) );
INV_X4 inst_2542 ( .ZN(net_3416), .A(net_2718) );
HA_X1 inst_3091 ( .S(net_1571), .CO(net_1570), .A(net_1342), .B(net_238) );
AND2_X2 inst_4197 ( .ZN(net_1601), .A1(net_1600), .A2(net_1514) );
CLKBUF_X2 inst_4668 ( .A(net_4653), .Z(net_4654) );
OAI221_X2 inst_417 ( .B1(net_3982), .ZN(net_1296), .C1(net_1295), .A(net_1098), .B2(net_717), .C2(net_259) );
NAND2_X2 inst_1861 ( .A1(net_3900), .A2(net_3441), .ZN(net_716) );
OAI21_X2 inst_671 ( .ZN(net_1593), .B1(net_1388), .A(net_1279), .B2(net_1103) );
XOR2_X2 inst_21 ( .Z(net_4071), .A(net_815), .B(net_617) );
AOI22_X2 inst_3570 ( .A1(net_4060), .B1(net_4055), .B2(net_3029), .A2(net_3028), .ZN(net_1480) );
CLKBUF_X2 inst_4524 ( .A(net_4361), .Z(net_4510) );
CLKBUF_X2 inst_4871 ( .A(net_4335), .Z(net_4857) );
CLKBUF_X2 inst_4835 ( .A(net_4601), .Z(net_4821) );
NAND2_X2 inst_2004 ( .A1(net_3550), .ZN(net_3527), .A2(net_3490) );
CLKBUF_X2 inst_4586 ( .A(net_4571), .Z(net_4572) );
CLKBUF_X2 inst_4257 ( .A(net_4242), .Z(net_4243) );
INV_X4 inst_2311 ( .A(net_1129), .ZN(net_790) );
AOI221_X2 inst_3885 ( .ZN(net_1658), .C1(net_1657), .C2(net_1656), .A(net_1251), .B1(net_1205), .B2(net_984) );
INV_X2 inst_2857 ( .A(net_4007), .ZN(net_377) );
OR2_X4 inst_220 ( .A1(net_4081), .ZN(net_1081), .A2(net_686) );
NAND2_X2 inst_1585 ( .A1(net_2915), .ZN(net_2435), .A2(net_163) );
NAND3_X2 inst_1317 ( .A3(net_3662), .A1(net_3523), .ZN(net_955), .A2(net_403) );
AOI22_X2 inst_3683 ( .B1(net_4123), .ZN(net_500), .A1(net_458), .B2(net_193), .A2(net_169) );
INV_X2 inst_2941 ( .A(net_3149), .ZN(net_282) );
OR2_X4 inst_245 ( .ZN(net_4133), .A1(net_3959), .A2(net_3952) );
NAND2_X2 inst_1873 ( .A2(net_4003), .ZN(net_658), .A1(net_517) );
AND2_X4 inst_4111 ( .A1(net_3654), .ZN(net_3243), .A2(net_283) );
OAI21_X2 inst_624 ( .B1(net_2235), .ZN(net_2157), .A(net_2045), .B2(net_106) );
SDFF_X2 inst_147 ( .D(net_3884), .SE(net_2625), .SI(net_93), .Q(net_93), .CK(net_4944) );
OAI22_X2 inst_313 ( .ZN(net_1164), .B1(net_641), .A1(net_533), .B2(net_529), .A2(net_523) );
NAND2_X2 inst_1676 ( .A1(net_2134), .ZN(net_2081), .A2(net_568) );
AND2_X4 inst_4170 ( .ZN(net_4124), .A2(net_3163), .A1(net_338) );
NOR2_X2 inst_1041 ( .A1(net_3964), .ZN(net_1328), .A2(net_1173) );
CLKBUF_X2 inst_5263 ( .A(net_5120), .Z(net_5249) );
NAND2_X1 inst_2086 ( .A2(net_4009), .A1(net_2972), .ZN(net_2433) );
DFF_X2 inst_3114 ( .D(net_2817), .QN(net_118), .CK(net_4597) );
AOI22_X2 inst_3577 ( .A1(net_4059), .B1(net_4056), .ZN(net_1473), .A2(net_195), .B2(net_194) );
INV_X2 inst_2637 ( .A(net_3693), .ZN(net_2511) );
AOI22_X2 inst_3624 ( .B2(net_3627), .ZN(net_1109), .A2(net_1011), .B1(net_948), .A1(net_888) );
OR2_X4 inst_236 ( .ZN(net_3208), .A1(net_3206), .A2(net_2352) );
CLKBUF_X2 inst_4539 ( .A(net_4524), .Z(net_4525) );
CLKBUF_X2 inst_4754 ( .A(net_4739), .Z(net_4740) );
OAI21_X2 inst_553 ( .B2(net_2925), .ZN(net_2873), .B1(net_2871), .A(net_2423) );
AOI221_X2 inst_3878 ( .B1(net_2020), .C1(net_2019), .ZN(net_1855), .A(net_1854), .B2(net_272), .C2(x409) );
DFF_X1 inst_3331 ( .D(net_2818), .QN(net_331), .CK(net_4323) );
CLKBUF_X2 inst_4532 ( .A(net_4517), .Z(net_4518) );
OR2_X4 inst_242 ( .ZN(net_3781), .A1(net_2212), .A2(net_1521) );
NOR2_X2 inst_986 ( .A1(net_3813), .ZN(net_2530), .A2(net_2529) );
DFF_X2 inst_3172 ( .D(net_1885), .QN(net_270), .CK(net_4849) );
CLKBUF_X2 inst_4983 ( .A(net_4422), .Z(net_4969) );
CLKBUF_X2 inst_4680 ( .A(net_4665), .Z(net_4666) );
NAND2_X4 inst_1422 ( .A2(net_3600), .ZN(net_3579), .A1(net_3238) );
AOI22_X2 inst_3508 ( .B1(net_3676), .B2(net_3136), .A1(net_2012), .ZN(net_2009), .A2(net_1797) );
CLKBUF_X2 inst_5132 ( .A(net_5117), .Z(net_5118) );
NAND4_X2 inst_1186 ( .ZN(net_1911), .A2(net_1757), .A1(net_1725), .A3(net_1721), .A4(net_1056) );
NAND2_X2 inst_1753 ( .ZN(net_1724), .A2(net_1300), .A1(net_1181) );
NAND2_X2 inst_1727 ( .ZN(net_1566), .A1(net_1565), .A2(net_1454) );
NAND4_X2 inst_1221 ( .ZN(net_952), .A4(net_736), .A3(net_569), .A2(net_489), .A1(net_476) );
NOR2_X1 inst_1166 ( .A1(net_2127), .ZN(net_1190), .A2(net_1189) );
NAND2_X2 inst_1739 ( .A2(net_3751), .ZN(net_1559), .A1(net_1437) );
XNOR2_X2 inst_116 ( .A(net_3875), .B(net_3858), .ZN(net_3224) );
NOR2_X2 inst_1133 ( .ZN(net_3656), .A1(net_3655), .A2(net_3477) );
OAI21_X2 inst_471 ( .B1(net_3509), .ZN(net_2979), .B2(net_2967), .A(net_2409) );
AND3_X2 inst_4087 ( .A2(net_4087), .ZN(net_1012), .A3(net_1011), .A1(net_145) );
CLKBUF_X2 inst_4580 ( .A(net_4565), .Z(net_4566) );
MUX2_X2 inst_2103 ( .S(net_2925), .Z(net_2575), .A(net_2573), .B(net_175) );
CLKBUF_X2 inst_4956 ( .A(net_4941), .Z(net_4942) );
AOI22_X2 inst_3609 ( .A1(net_4063), .B1(net_4058), .ZN(net_1408), .A2(net_597), .B2(net_596) );
CLKBUF_X2 inst_5139 ( .A(net_5124), .Z(net_5125) );
NOR3_X2 inst_896 ( .A2(net_3982), .A1(net_3781), .ZN(net_1702), .A3(net_56) );
CLKBUF_X2 inst_4750 ( .A(net_4735), .Z(net_4736) );
OAI22_X2 inst_339 ( .B1(net_3871), .A1(net_3556), .ZN(net_3217), .A2(net_2995), .B2(net_2994) );
INV_X2 inst_2664 ( .ZN(net_2351), .A(net_2099) );
OAI222_X2 inst_351 ( .C1(net_3784), .B2(net_3152), .A2(net_2189), .ZN(net_1934), .A1(net_1815), .B1(net_1814), .C2(net_119) );
INV_X4 inst_2608 ( .A(net_3817), .ZN(net_3816) );
INV_X4 inst_2557 ( .ZN(net_3497), .A(net_3494) );
INV_X4 inst_2521 ( .A(net_3370), .ZN(net_3252) );
OAI221_X2 inst_385 ( .B2(net_2699), .C2(net_2698), .ZN(net_2627), .B1(net_2626), .A(net_2532), .C1(net_2324) );
DFF_X1 inst_3319 ( .QN(net_3002), .D(net_2843), .CK(net_5071) );
INV_X2 inst_2653 ( .A(net_3827), .ZN(net_2630) );
CLKBUF_X2 inst_4621 ( .A(net_4606), .Z(net_4607) );
INV_X4 inst_2550 ( .ZN(net_3455), .A(net_2986) );
NAND2_X2 inst_1560 ( .A1(net_2912), .ZN(net_2462), .A2(net_227) );
AOI21_X2 inst_3932 ( .A(net_3465), .B2(net_3115), .ZN(net_2864), .B1(net_2822) );
CLKBUF_X2 inst_4281 ( .A(net_4266), .Z(net_4267) );
OAI21_X2 inst_596 ( .ZN(net_2624), .B1(net_2531), .A(net_1600), .B2(net_1443) );
INV_X2 inst_2771 ( .A(net_955), .ZN(net_883) );
CLKBUF_X2 inst_4687 ( .A(net_4287), .Z(net_4673) );
INV_X8 inst_2142 ( .A(net_3780), .ZN(net_3186) );
NAND2_X2 inst_1705 ( .ZN(net_1759), .A1(net_1758), .A2(net_53) );
CLKBUF_X2 inst_5110 ( .A(net_4702), .Z(net_5096) );
CLKBUF_X2 inst_4664 ( .A(net_4489), .Z(net_4650) );
OAI211_X2 inst_847 ( .C1(net_1274), .C2(net_988), .B(net_891), .ZN(net_704), .A(net_615) );
INV_X2 inst_2720 ( .ZN(net_1513), .A(net_1512) );
CLKBUF_X2 inst_5003 ( .A(net_4399), .Z(net_4989) );
CLKBUF_X2 inst_4458 ( .A(net_4443), .Z(net_4444) );
NAND2_X2 inst_1942 ( .ZN(net_3235), .A1(net_3187), .A2(net_221) );
NAND2_X2 inst_1716 ( .A1(net_3492), .A2(net_3364), .ZN(net_1690) );
DFF_X1 inst_3253 ( .QN(net_3088), .D(net_2944), .CK(net_4727) );
INV_X2 inst_2648 ( .A(net_3884), .ZN(net_2626) );
CLKBUF_X2 inst_5184 ( .A(net_5169), .Z(net_5170) );
CLKBUF_X2 inst_4596 ( .A(net_4573), .Z(net_4582) );
NOR2_X2 inst_1146 ( .ZN(net_3913), .A1(net_3489), .A2(net_3488) );
OAI21_X2 inst_637 ( .B2(net_2076), .ZN(net_2073), .A(net_1964), .B1(net_1677) );
AOI22_X2 inst_3708 ( .B1(net_4124), .A1(net_509), .ZN(net_456), .B2(net_236), .A2(net_151) );
OAI21_X2 inst_547 ( .B2(net_2912), .B1(net_2887), .ZN(net_2884), .A(net_2452) );
AOI211_X2 inst_4023 ( .ZN(net_1298), .B(net_1106), .C2(net_1094), .C1(net_840), .A(net_811) );
DFF_X2 inst_3105 ( .D(net_2827), .QN(net_245), .CK(net_4330) );
AOI22_X2 inst_3673 ( .ZN(net_548), .A1(net_458), .B1(net_457), .B2(net_221), .A2(net_155) );
AOI222_X1 inst_3781 ( .C1(net_4065), .B2(net_3789), .ZN(net_1725), .B1(net_1724), .A2(net_1581), .A1(net_1180), .C2(net_1113) );
CLKBUF_X2 inst_5162 ( .A(net_5147), .Z(net_5148) );
CLKBUF_X2 inst_4519 ( .A(net_4367), .Z(net_4505) );
AOI22_X2 inst_3539 ( .B1(net_1840), .A1(net_1698), .ZN(net_1669), .B2(net_179), .A2(net_77) );
INV_X4 inst_2457 ( .A(net_3078), .ZN(net_467) );
AOI22_X2 inst_3552 ( .A1(net_4060), .B1(net_4055), .ZN(net_1498), .A2(net_186), .B2(net_162) );
NAND2_X2 inst_1702 ( .ZN(net_1786), .A2(net_1785), .A1(net_1688) );
OAI33_X1 inst_274 ( .A1(net_1701), .B2(net_1606), .ZN(net_1556), .B1(net_1232), .B3(net_1173), .A3(net_444), .A2(net_143) );
NAND2_X2 inst_1607 ( .A1(net_2967), .ZN(net_2409), .A2(net_475) );
NAND3_X2 inst_1277 ( .ZN(net_2703), .A3(net_2691), .A1(net_2647), .A2(net_2593) );
INV_X2 inst_2817 ( .A(net_714), .ZN(net_604) );
AND3_X4 inst_4076 ( .ZN(net_4090), .A2(net_3959), .A3(net_3948), .A1(net_710) );
NAND2_X1 inst_2092 ( .A2(net_3968), .ZN(net_540), .A1(net_356) );
CLKBUF_X2 inst_4762 ( .A(net_4245), .Z(net_4748) );
OR3_X4 inst_164 ( .A2(net_2596), .ZN(net_2215), .A1(net_2214), .A3(net_2213) );
DFF_X2 inst_3207 ( .Q(net_3158), .D(net_1166), .CK(net_4824) );
DFF_X2 inst_3143 ( .QN(net_3103), .D(net_2542), .CK(net_4633) );
NAND2_X2 inst_1854 ( .A1(net_3243), .ZN(net_652), .A2(net_418) );
INV_X2 inst_2696 ( .ZN(net_1688), .A(net_1687) );
NAND2_X2 inst_1710 ( .A2(net_1772), .ZN(net_1734), .A1(net_1703) );
INV_X4 inst_2407 ( .ZN(net_528), .A(net_357) );
NAND2_X2 inst_1771 ( .ZN(net_1277), .A1(net_1158), .A2(net_973) );
INV_X2 inst_2880 ( .A(net_344), .ZN(net_263) );
CLKBUF_X2 inst_4884 ( .A(net_4869), .Z(net_4870) );
NAND2_X4 inst_1440 ( .ZN(net_3720), .A1(net_3678), .A2(net_3540) );
INV_X2 inst_2660 ( .ZN(net_2109), .A(net_2038) );
DFF_X2 inst_3142 ( .QN(net_2983), .D(net_2572), .CK(net_5228) );
INV_X4 inst_2305 ( .A(net_3924), .ZN(net_848) );
DFF_X1 inst_3355 ( .D(net_3695), .CK(net_4257), .Q(x142) );
OAI21_X2 inst_753 ( .ZN(net_3536), .B1(net_3533), .B2(net_3516), .A(net_3458) );
INV_X8 inst_2150 ( .ZN(net_3302), .A(net_3301) );
INV_X4 inst_2389 ( .A(net_826), .ZN(net_775) );
DFF_X1 inst_3427 ( .Q(net_4015), .D(net_4014), .CK(net_4910) );
NOR2_X4 inst_946 ( .ZN(net_3526), .A2(net_3168), .A1(net_268) );
NAND2_X2 inst_1954 ( .ZN(net_3285), .A1(net_3284), .A2(net_3182) );
INV_X4 inst_2260 ( .ZN(net_2141), .A(net_1172) );
CLKBUF_X2 inst_4946 ( .A(net_4643), .Z(net_4932) );
INV_X8 inst_2148 ( .A(net_3800), .ZN(net_3281) );
AOI21_X2 inst_3941 ( .ZN(net_2242), .B1(net_2238), .A(net_2188), .B2(net_1874) );
INV_X2 inst_2900 ( .A(net_3116), .ZN(net_1532) );
NAND2_X2 inst_1591 ( .A1(net_2972), .ZN(net_2427), .A2(net_834) );
DFF_X1 inst_3247 ( .QN(net_3091), .D(net_2948), .CK(net_4550) );
AOI22_X2 inst_3697 ( .B1(net_4124), .A1(net_509), .ZN(net_477), .A2(net_214), .B2(net_202) );
AOI221_X2 inst_3858 ( .B1(net_3736), .A(net_3362), .C2(net_3117), .C1(net_2115), .ZN(net_2046), .B2(net_239) );
OAI221_X2 inst_379 ( .B1(net_2670), .C1(net_2668), .ZN(net_2662), .B2(net_2661), .A(net_1386), .C2(net_331) );
CLKBUF_X2 inst_4625 ( .A(net_4610), .Z(net_4611) );
NOR2_X4 inst_926 ( .A2(net_3831), .A1(net_3266), .ZN(net_2210) );
AOI21_X4 inst_3922 ( .B2(net_3600), .ZN(net_2887), .B1(net_2878), .A(net_2124) );
NAND2_X2 inst_2053 ( .ZN(net_3895), .A2(net_3892), .A1(net_3347) );
NAND3_X2 inst_1325 ( .A2(net_3913), .ZN(net_1016), .A3(net_838), .A1(net_666) );
INV_X4 inst_2570 ( .ZN(net_3544), .A(net_3543) );
AND2_X4 inst_4153 ( .ZN(net_4102), .A2(net_3662), .A1(net_440) );
CLKBUF_X2 inst_4960 ( .A(net_4363), .Z(net_4946) );
CLKBUF_X2 inst_5105 ( .A(net_5090), .Z(net_5091) );
DFF_X1 inst_3312 ( .Q(net_3140), .D(net_2854), .CK(net_4519) );
AOI22_X2 inst_3646 ( .A1(net_4142), .B1(net_4112), .B2(net_2033), .ZN(net_756), .A2(x916) );
AOI22_X2 inst_3719 ( .A1(net_3815), .ZN(net_3607), .B1(net_3186), .A2(net_732), .B2(net_731) );
NOR3_X2 inst_891 ( .A3(net_3158), .ZN(net_2386), .A2(net_2384), .A1(net_2327) );
AND2_X4 inst_4095 ( .ZN(net_1741), .A1(net_1740), .A2(net_1705) );
XNOR2_X2 inst_74 ( .ZN(net_1462), .B(net_1461), .A(net_1329) );
NAND4_X2 inst_1235 ( .A2(net_3900), .A3(net_3243), .A4(net_721), .ZN(net_685), .A1(net_376) );
INV_X4 inst_2244 ( .A(net_1816), .ZN(net_1793) );
AOI22_X2 inst_3561 ( .B1(net_4062), .A1(net_4056), .ZN(net_1489), .A2(net_214), .B2(net_141) );
OAI22_X2 inst_288 ( .B1(net_1891), .ZN(net_1881), .A1(net_1880), .B2(net_508), .A2(net_276) );
DFF_X1 inst_3284 ( .QN(net_3052), .D(net_2896), .CK(net_4777) );
INV_X2 inst_3046 ( .ZN(net_3708), .A(net_1855) );
AOI22_X2 inst_3626 ( .A1(net_4115), .B1(net_1882), .ZN(net_940), .A2(net_773), .B2(net_210) );
AND4_X4 inst_4036 ( .ZN(net_2145), .A4(net_2144), .A1(net_2120), .A2(net_1867), .A3(net_1866) );
CLKBUF_X2 inst_4644 ( .A(net_4415), .Z(net_4630) );
CLKBUF_X2 inst_5244 ( .A(net_5229), .Z(net_5230) );
CLKBUF_X2 inst_4844 ( .A(net_4829), .Z(net_4830) );
CLKBUF_X2 inst_4512 ( .A(net_4497), .Z(net_4498) );
NAND3_X2 inst_1298 ( .A2(net_1636), .ZN(net_1563), .A1(net_1562), .A3(net_593) );
AOI222_X1 inst_3757 ( .A1(net_3676), .B1(net_2055), .C1(net_2054), .ZN(net_2035), .C2(net_425), .B2(net_379), .A2(net_295) );
NOR3_X2 inst_917 ( .ZN(net_4045), .A3(net_3447), .A1(net_1790), .A2(net_1772) );
AOI22_X2 inst_3712 ( .ZN(net_3205), .A1(net_3198), .A2(net_3023), .B2(net_3022), .B1(net_1982) );
NAND2_X2 inst_1743 ( .ZN(net_1503), .A1(net_1309), .A2(net_271) );
OAI221_X2 inst_372 ( .ZN(net_2685), .B2(net_2684), .B1(net_2670), .C1(net_2668), .A(net_1386), .C2(net_292) );
NAND2_X2 inst_1600 ( .A1(net_2969), .ZN(net_2417), .A2(net_488) );
CLKBUF_X2 inst_5022 ( .A(net_5007), .Z(net_5008) );
OR2_X4 inst_215 ( .A1(net_1445), .ZN(net_1374), .A2(net_300) );
INV_X2 inst_2850 ( .A(net_3526), .ZN(net_373) );
CLKBUF_X2 inst_5163 ( .A(net_5148), .Z(net_5149) );
INV_X4 inst_2624 ( .ZN(net_3968), .A(net_3967) );
OAI211_X2 inst_849 ( .B(net_3243), .ZN(net_719), .C1(net_666), .A(net_517), .C2(net_418) );
NAND2_X2 inst_1775 ( .A1(net_2213), .ZN(net_1359), .A2(net_1107) );
INV_X4 inst_2397 ( .A(net_3391), .ZN(net_1636) );
XOR2_X2 inst_3 ( .B(net_3255), .Z(net_1996), .A(net_1713) );
NOR2_X1 inst_1172 ( .ZN(net_4141), .A1(net_4081), .A2(net_1381) );
NOR2_X2 inst_1090 ( .A1(net_3391), .ZN(net_586), .A2(x974) );
INV_X2 inst_3060 ( .ZN(net_4172), .A(net_1994) );
AOI221_X2 inst_3903 ( .A(net_4078), .ZN(net_1112), .B2(net_990), .B1(net_911), .C1(net_892), .C2(net_361) );
INV_X4 inst_2372 ( .A(net_3900), .ZN(net_526) );
INV_X4 inst_2575 ( .ZN(net_3585), .A(net_3583) );
CLKBUF_X2 inst_5007 ( .A(net_4992), .Z(net_4993) );
OAI21_X2 inst_566 ( .B2(net_2912), .B1(net_2849), .ZN(net_2846), .A(net_2453) );
NAND2_X4 inst_1399 ( .ZN(net_796), .A2(net_672), .A1(net_665) );
NAND4_X2 inst_1239 ( .A1(net_3448), .ZN(net_3230), .A2(net_2597), .A4(net_2596), .A3(net_1295) );
CLKBUF_X2 inst_4357 ( .A(net_4342), .Z(net_4343) );
CLKBUF_X2 inst_4819 ( .A(net_4804), .Z(net_4805) );
DFF_X2 inst_3126 ( .QN(net_3142), .D(net_2687), .CK(net_4573) );
CLKBUF_X2 inst_4327 ( .A(net_4312), .Z(net_4313) );
OAI21_X2 inst_503 ( .B1(net_3394), .B2(net_3208), .ZN(net_2939), .A(net_2491) );
CLKBUF_X2 inst_4774 ( .A(net_4759), .Z(net_4760) );
INV_X4 inst_2333 ( .A(net_1071), .ZN(net_1036) );
NAND2_X2 inst_1936 ( .ZN(net_3203), .A1(net_3198), .A2(net_203) );
DFF_X2 inst_3193 ( .Q(net_3759), .D(net_3758), .QN(net_3168), .CK(net_5272) );
CLKBUF_X2 inst_5088 ( .A(net_5073), .Z(net_5074) );
AND2_X2 inst_4193 ( .A1(net_3448), .ZN(net_2710), .A2(net_1052) );
NAND2_X1 inst_2099 ( .ZN(net_3692), .A1(net_3688), .A2(net_2691) );
AND3_X4 inst_4069 ( .A1(net_4077), .ZN(net_1142), .A2(net_965), .A3(net_850) );
CLKBUF_X2 inst_5056 ( .A(net_5041), .Z(net_5042) );
NOR2_X2 inst_1097 ( .A1(net_3167), .A2(net_3109), .ZN(net_304) );
OAI21_X2 inst_686 ( .B1(net_3228), .B2(net_2037), .ZN(net_1308), .A(net_1259) );
AOI211_X2 inst_4016 ( .C1(net_4065), .ZN(net_1820), .B(net_1724), .C2(net_1663), .A(net_1043) );
CLKBUF_X2 inst_4892 ( .A(net_4877), .Z(net_4878) );
NAND2_X2 inst_1732 ( .A1(net_1556), .ZN(net_1553), .A2(x717) );
INV_X2 inst_2914 ( .A(net_3036), .ZN(net_172) );
INV_X2 inst_2888 ( .A(net_3044), .ZN(net_234) );
DFF_X1 inst_3294 ( .QN(net_3010), .D(net_2881), .CK(net_5121) );
INV_X2 inst_2741 ( .A(net_3966), .ZN(net_1267) );
AOI22_X2 inst_3643 ( .A1(net_4142), .B1(net_4112), .B2(net_1797), .ZN(net_759), .A2(x762) );
NOR2_X4 inst_967 ( .ZN(net_3857), .A2(net_3856), .A1(net_3855) );
INV_X8 inst_2119 ( .A(net_3556), .ZN(net_2134) );
NAND2_X2 inst_1929 ( .ZN(net_3192), .A1(net_3186), .A2(net_734) );
NAND2_X2 inst_1522 ( .A1(net_2959), .ZN(net_2500), .A2(net_737) );
DFF_X1 inst_3391 ( .D(net_1716), .QN(net_78), .CK(net_4246) );
NAND2_X2 inst_1794 ( .A1(net_1013), .ZN(net_1005), .A2(net_521) );
NAND4_X2 inst_1227 ( .ZN(net_800), .A4(net_634), .A3(net_566), .A2(net_483), .A1(net_466) );
INV_X4 inst_2324 ( .A(net_1024), .ZN(net_709) );
INV_X16 inst_3069 ( .A(net_4000), .ZN(net_3900) );
AOI22_X2 inst_3631 ( .ZN(net_879), .A2(net_458), .B2(net_457), .B1(net_190), .A1(net_161) );
NOR2_X2 inst_1101 ( .A2(net_3154), .A1(net_3108), .ZN(net_275) );
INV_X2 inst_3047 ( .ZN(net_3729), .A(net_3728) );
INV_X2 inst_2950 ( .A(net_3039), .ZN(net_205) );
AOI221_X2 inst_3847 ( .B1(net_3736), .ZN(net_2138), .C1(net_2137), .A(net_1941), .B2(net_330), .C2(net_216) );
INV_X2 inst_2897 ( .A(net_3008), .ZN(net_202) );
NOR4_X2 inst_861 ( .A1(net_1718), .ZN(net_1659), .A2(net_1657), .A3(net_1522), .A4(net_1149) );
INV_X4 inst_2529 ( .A(net_3283), .ZN(net_3280) );
NAND2_X2 inst_1787 ( .A1(net_3963), .A2(net_1837), .ZN(net_1031) );
INV_X2 inst_2990 ( .A(net_3152), .ZN(net_378) );
NAND3_X2 inst_1283 ( .ZN(net_2733), .A2(net_2377), .A1(net_2375), .A3(net_2374) );
INV_X4 inst_2451 ( .ZN(net_1874), .A(net_118) );
NAND4_X2 inst_1202 ( .ZN(net_2196), .A3(net_1473), .A4(net_1472), .A1(net_1407), .A2(net_1406) );
CLKBUF_X2 inst_4290 ( .A(net_4275), .Z(net_4276) );
NAND2_X2 inst_1540 ( .A1(net_2907), .ZN(net_2482), .A2(net_234) );
INV_X4 inst_2227 ( .ZN(net_2684), .A(net_2583) );
NAND2_X2 inst_1660 ( .ZN(net_2103), .A1(net_1982), .A2(net_193) );
INV_X2 inst_2742 ( .ZN(net_1227), .A(net_1226) );
AOI22_X2 inst_3536 ( .A2(net_1908), .ZN(net_1768), .A1(net_1767), .B2(net_749), .B1(net_96) );
OAI21_X2 inst_660 ( .ZN(net_2583), .B2(net_1975), .B1(net_1765), .A(net_1452) );
CLKBUF_X2 inst_5243 ( .A(net_4364), .Z(net_5229) );
CLKBUF_X2 inst_4375 ( .A(net_4238), .Z(net_4361) );
INV_X4 inst_2490 ( .A(net_3074), .ZN(net_558) );
OAI21_X2 inst_517 ( .B2(net_2959), .ZN(net_2924), .B1(net_2923), .A(net_2497) );
CLKBUF_X2 inst_5195 ( .A(net_4696), .Z(net_5181) );
NAND2_X2 inst_1576 ( .A1(net_2965), .ZN(net_2444), .A2(net_244) );
INV_X4 inst_2346 ( .ZN(net_722), .A(net_603) );
NAND4_X1 inst_1261 ( .ZN(net_4187), .A4(net_3530), .A2(net_3513), .A3(net_2679), .A1(net_2541) );
AOI22_X4 inst_3462 ( .ZN(net_3264), .A1(net_3263), .B1(net_1445), .A2(net_1374), .B2(net_300) );
CLKBUF_X2 inst_4254 ( .A(x1012), .Z(net_4240) );
CLKBUF_X2 inst_4330 ( .A(net_4315), .Z(net_4316) );
OAI22_X2 inst_310 ( .B1(net_3132), .ZN(net_1242), .A1(net_1099), .A2(net_1071), .B2(net_1036) );
CLKBUF_X2 inst_4368 ( .A(net_4353), .Z(net_4354) );
OAI211_X2 inst_794 ( .ZN(net_2636), .C1(net_2549), .A(net_2548), .C2(net_2547), .B(net_1740) );
INV_X2 inst_2754 ( .A(net_1183), .ZN(net_1004) );
NOR2_X2 inst_1005 ( .A2(net_3505), .ZN(net_1969), .A1(net_1833) );
INV_X2 inst_2759 ( .A(net_1137), .ZN(net_982) );
NOR2_X2 inst_1147 ( .ZN(net_3916), .A2(net_3914), .A1(net_525) );
NAND2_X2 inst_1768 ( .A1(net_4185), .ZN(net_1225), .A2(net_1011) );
NAND2_X2 inst_1580 ( .A1(net_2965), .ZN(net_2440), .A2(net_232) );
NAND2_X2 inst_1842 ( .ZN(net_844), .A2(net_775), .A1(net_435) );
INV_X2 inst_2688 ( .ZN(net_1756), .A(net_1722) );
INV_X2 inst_2917 ( .ZN(net_2307), .A(net_71) );
INV_X4 inst_2423 ( .ZN(net_347), .A(net_225) );
NAND2_X4 inst_1408 ( .A2(net_4135), .ZN(net_3301), .A1(net_3300) );
NOR2_X2 inst_996 ( .A1(net_2732), .ZN(net_2311), .A2(net_1905) );
INV_X4 inst_2351 ( .ZN(net_2525), .A(net_593) );
CLKBUF_X2 inst_5125 ( .A(net_5110), .Z(net_5111) );
NAND2_X2 inst_1853 ( .ZN(net_660), .A2(net_659), .A1(net_589) );
NAND2_X2 inst_1889 ( .A1(net_1636), .ZN(net_511), .A2(x974) );
NAND2_X2 inst_1527 ( .A1(net_3208), .ZN(net_2495), .A2(net_171) );
NAND2_X2 inst_2011 ( .ZN(net_3584), .A2(net_3583), .A1(net_2382) );
NAND2_X2 inst_1761 ( .A1(net_4031), .A2(net_1394), .ZN(net_1238) );
OAI21_X2 inst_740 ( .B1(net_3588), .ZN(net_3267), .B2(net_3208), .A(net_2490) );
OR2_X2 inst_264 ( .A1(net_4132), .A2(net_402), .ZN(net_395) );
AOI22_X2 inst_3703 ( .ZN(net_465), .A1(net_458), .B1(net_457), .B2(net_197), .A2(net_175) );
AND2_X4 inst_4189 ( .ZN(net_4186), .A2(net_591), .A1(net_583) );
XNOR2_X2 inst_84 ( .ZN(net_1222), .B(net_987), .A(net_875) );
NAND3_X2 inst_1333 ( .A3(net_3662), .A2(net_3613), .ZN(net_531), .A1(net_424) );
NAND2_X2 inst_1937 ( .A1(net_3769), .ZN(net_3214), .A2(net_368) );
OR3_X4 inst_173 ( .A1(net_4113), .A3(net_3387), .ZN(net_814), .A2(net_632) );
AOI22_X2 inst_3710 ( .B1(net_4123), .A1(net_571), .ZN(net_443), .B2(net_177), .A2(net_153) );
CLKBUF_X2 inst_4405 ( .A(net_4220), .Z(net_4391) );
OAI21_X2 inst_611 ( .ZN(net_2354), .A(net_2299), .B1(net_2298), .B2(net_2181) );
AOI21_X2 inst_3953 ( .ZN(net_1753), .A(net_1702), .B1(net_1651), .B2(net_231) );
INV_X4 inst_2487 ( .A(net_3013), .ZN(net_155) );
NAND2_X2 inst_1551 ( .A1(net_2961), .ZN(net_2471), .A2(net_467) );
NAND4_X1 inst_1260 ( .ZN(net_506), .A4(net_505), .A1(net_327), .A2(net_289), .A3(net_260) );
NOR2_X2 inst_1088 ( .A1(net_4127), .ZN(net_449), .A2(net_42) );
NAND2_X2 inst_1943 ( .A1(net_4182), .ZN(net_3245), .A2(net_3244) );
OAI21_X2 inst_490 ( .B1(net_3588), .B2(net_2969), .ZN(net_2952), .A(net_2413) );
DFF_X1 inst_3332 ( .Q(net_3151), .D(net_2821), .CK(net_4366) );
CLKBUF_X2 inst_4898 ( .A(net_4883), .Z(net_4884) );
INV_X2 inst_2717 ( .A(net_3515), .ZN(net_2323) );
INV_X4 inst_2218 ( .A(net_3556), .ZN(net_2082) );
AND2_X4 inst_4176 ( .ZN(net_4130), .A2(net_3388), .A1(net_3127) );
SDFF_X2 inst_129 ( .D(net_3483), .SI(net_3028), .Q(net_3028), .SE(net_2907), .CK(net_5061) );
NAND3_X2 inst_1309 ( .A1(net_4069), .ZN(net_1114), .A2(net_409), .A3(net_207) );
INV_X2 inst_2740 ( .ZN(net_1270), .A(net_1218) );
NAND2_X2 inst_1754 ( .ZN(net_1294), .A2(net_1293), .A1(net_1172) );
NAND2_X2 inst_1531 ( .A1(net_3208), .ZN(net_2491), .A2(net_551) );
INV_X2 inst_2931 ( .A(net_3000), .ZN(net_236) );
CLKBUF_X2 inst_4768 ( .A(net_4753), .Z(net_4754) );
CLKBUF_X2 inst_4938 ( .A(net_4322), .Z(net_4924) );
INV_X4 inst_2530 ( .ZN(net_3283), .A(net_3281) );
INV_X2 inst_2727 ( .ZN(net_1451), .A(net_1450) );
INV_X2 inst_2922 ( .A(net_3159), .ZN(net_220) );
AOI221_X2 inst_3803 ( .C1(net_2781), .B1(net_2775), .ZN(net_2772), .A(net_2671), .B2(net_318), .C2(net_77) );
DFF_X2 inst_3183 ( .D(net_1749), .QN(net_106), .CK(net_4528) );
NAND2_X2 inst_1503 ( .ZN(net_2794), .A1(net_2730), .A2(net_2695) );
OAI21_X1 inst_777 ( .A(net_3858), .B2(net_3827), .B1(net_3405), .ZN(net_3329) );
CLKBUF_X2 inst_4312 ( .A(net_4297), .Z(net_4298) );
AOI221_X2 inst_3802 ( .C1(net_2781), .B1(net_2775), .ZN(net_2773), .A(net_2662), .B2(net_331), .C2(net_255) );
CLKBUF_X2 inst_5016 ( .A(net_5001), .Z(net_5002) );
NOR2_X2 inst_1037 ( .ZN(net_1284), .A1(net_1283), .A2(net_586) );
NOR2_X4 inst_933 ( .A2(net_3641), .A1(net_3576), .ZN(net_1272) );
OAI22_X2 inst_300 ( .ZN(net_1546), .B2(net_1545), .A1(net_1543), .B1(net_1542), .A2(net_318) );
AOI22_X2 inst_3596 ( .A1(net_4062), .B1(net_4057), .ZN(net_1421), .A2(net_519), .B2(net_478) );
AOI22_X2 inst_3724 ( .ZN(net_3651), .B1(net_3647), .A1(net_3185), .A2(net_462), .B2(net_461) );
NAND4_X2 inst_1250 ( .ZN(net_3826), .A1(net_3825), .A4(net_3767), .A3(net_3766), .A2(net_3590) );
NAND4_X2 inst_1226 ( .A3(net_2717), .A2(net_1274), .A4(net_1126), .ZN(net_793), .A1(net_686) );
NOR2_X2 inst_1013 ( .A2(net_3321), .ZN(net_1838), .A1(net_1739) );
OAI221_X2 inst_446 ( .B1(net_4161), .ZN(net_3749), .B2(net_3407), .C1(net_2328), .A(net_2021), .C2(net_67) );
CLKBUF_X2 inst_4965 ( .A(net_4950), .Z(net_4951) );
NAND2_X2 inst_1979 ( .ZN(net_3382), .A1(net_3377), .A2(net_3376) );
OAI221_X2 inst_364 ( .ZN(net_2742), .B1(net_2733), .C1(net_2731), .C2(net_2663), .A(net_2644), .B2(net_1818) );
AOI22_X2 inst_3613 ( .A1(net_4063), .B1(net_4058), .ZN(net_1404), .B2(net_235), .A2(net_232) );
INV_X4 inst_2354 ( .ZN(net_1606), .A(net_947) );
CLKBUF_X2 inst_4923 ( .A(net_4908), .Z(net_4909) );
OAI211_X2 inst_824 ( .C1(net_3964), .ZN(net_1816), .A(net_1450), .C2(net_1324), .B(net_671) );
INV_X2 inst_2997 ( .A(net_3003), .ZN(net_219) );
AOI22_X2 inst_3533 ( .ZN(net_1822), .B2(net_1821), .A1(net_1758), .B1(net_1169), .A2(net_54) );
CLKBUF_X2 inst_4712 ( .A(net_4697), .Z(net_4698) );
OAI221_X2 inst_411 ( .B2(net_3789), .ZN(net_1547), .A(net_1390), .B1(net_1343), .C2(net_1089), .C1(net_1040) );
XNOR2_X2 inst_124 ( .ZN(net_4154), .B(net_3459), .A(net_3457) );
AOI22_X2 inst_3515 ( .B1(net_4045), .B2(net_3466), .ZN(net_1956), .A1(net_1955), .A2(net_256) );
AOI222_X1 inst_3750 ( .C1(net_3116), .A2(net_3115), .ZN(net_2056), .A1(net_2055), .B2(net_2054), .C2(net_2053), .B1(net_1910) );
AOI211_X2 inst_4026 ( .B(net_4070), .C2(net_1636), .ZN(net_1226), .A(net_1173), .C1(net_883) );
AND4_X2 inst_4056 ( .ZN(net_1516), .A1(net_1327), .A4(net_1274), .A2(net_1268), .A3(net_1030) );
CLKBUF_X2 inst_4382 ( .A(net_4367), .Z(net_4368) );
CLKBUF_X2 inst_4401 ( .A(net_4386), .Z(net_4387) );
DFF_X1 inst_3430 ( .Q(net_4021), .D(net_4020), .CK(net_4899) );
AOI221_X2 inst_3869 ( .A(net_3362), .B2(net_3117), .B1(net_2020), .C1(net_2019), .ZN(net_1936), .C2(x204) );
AOI22_X2 inst_3488 ( .B1(net_2752), .ZN(net_2605), .A2(net_2520), .A1(net_2275), .B2(net_51) );
NAND3_X4 inst_1270 ( .ZN(net_3954), .A1(net_3927), .A3(net_3451), .A2(net_3450) );
CLKBUF_X2 inst_4563 ( .A(net_4548), .Z(net_4549) );
XNOR2_X2 inst_61 ( .A(net_3256), .ZN(net_2163), .B(net_1644) );
OR2_X4 inst_203 ( .ZN(net_2912), .A2(net_2354), .A1(net_2351) );
NOR2_X2 inst_1139 ( .ZN(net_3786), .A2(net_3266), .A1(net_2209) );
NAND2_X2 inst_1519 ( .A1(net_2959), .ZN(net_2503), .A2(net_150) );
INV_X8 inst_2156 ( .A(net_3939), .ZN(net_3612) );
CLKBUF_X2 inst_4989 ( .A(net_4974), .Z(net_4975) );
CLKBUF_X2 inst_4507 ( .A(net_4492), .Z(net_4493) );
NAND2_X2 inst_1571 ( .A1(net_2912), .ZN(net_2450), .A2(net_215) );
CLKBUF_X2 inst_4324 ( .A(net_4296), .Z(net_4310) );
OAI21_X4 inst_456 ( .A(net_3945), .ZN(net_392), .B1(net_313), .B2(net_275) );
OAI211_X2 inst_832 ( .ZN(net_1360), .C1(net_1359), .A(net_1241), .B(net_593), .C2(net_315) );
INV_X4 inst_2515 ( .A(net_3283), .ZN(net_3178) );
NAND2_X2 inst_1491 ( .A1(net_3368), .A2(net_3296), .ZN(net_2859) );
NAND2_X4 inst_1402 ( .A2(net_3662), .ZN(net_434), .A1(net_407) );
OAI33_X1 inst_275 ( .ZN(net_3796), .A3(net_3792), .B3(net_2717), .A1(net_1297), .A2(net_1288), .B1(net_730), .B2(net_631) );
XNOR2_X2 inst_117 ( .B(net_3859), .ZN(net_3592), .A(net_3511) );
INV_X2 inst_2676 ( .ZN(net_1896), .A(net_1895) );
CLKBUF_X2 inst_5172 ( .A(net_4970), .Z(net_5158) );
DFF_X2 inst_3106 ( .QN(net_3131), .D(net_2830), .CK(net_4490) );
AOI22_X2 inst_3728 ( .ZN(net_3864), .A1(net_3178), .B1(net_2099), .A2(net_226), .B2(net_167) );
SDFF_X2 inst_154 ( .SE(net_2514), .D(net_1886), .SI(net_86), .Q(net_86), .CK(net_4980) );
INV_X4 inst_2416 ( .A(net_3106), .ZN(net_257) );
AND2_X4 inst_4106 ( .A2(net_3163), .ZN(net_458), .A1(net_345) );
AOI221_X2 inst_3812 ( .B2(net_3134), .ZN(net_2592), .B1(net_2591), .C1(net_2590), .C2(net_2589), .A(net_1090) );
OAI21_X4 inst_465 ( .ZN(net_3770), .B1(net_3634), .A(net_1602), .B2(net_923) );
INV_X4 inst_2304 ( .ZN(net_2053), .A(net_1845) );
AOI21_X2 inst_3959 ( .B1(net_1797), .ZN(net_1639), .A(net_1561), .B2(net_433) );
INV_X4 inst_2503 ( .A(net_3155), .ZN(net_207) );
CLKBUF_X2 inst_4877 ( .A(net_4862), .Z(net_4863) );
CLKBUF_X2 inst_4518 ( .A(net_4503), .Z(net_4504) );
CLKBUF_X2 inst_4240 ( .A(net_4225), .Z(net_4226) );
INV_X4 inst_2173 ( .ZN(net_2871), .A(net_2837) );
NAND2_X2 inst_1790 ( .ZN(net_1587), .A2(net_958), .A1(net_937) );
XNOR2_X2 inst_94 ( .ZN(net_715), .A(net_714), .B(net_43) );
DFF_X2 inst_3214 ( .QN(net_3153), .D(net_806), .CK(net_4666) );
NAND2_X2 inst_1905 ( .A2(net_3127), .ZN(net_343), .A1(net_299) );
INV_X4 inst_2264 ( .ZN(net_1518), .A(net_1151) );
NAND3_X1 inst_1378 ( .A2(net_3530), .A1(net_3513), .ZN(net_3295), .A3(net_2679) );
OR2_X4 inst_243 ( .A2(net_4000), .ZN(net_3907), .A1(net_719) );
CLKBUF_X2 inst_4345 ( .A(net_4278), .Z(net_4331) );
OAI221_X2 inst_424 ( .B1(net_3839), .C2(net_3681), .ZN(net_1271), .C1(net_1152), .B2(net_877), .A(net_860) );
OAI21_X2 inst_591 ( .B1(net_3693), .A(net_3229), .ZN(net_2647), .B2(net_71) );
INV_X2 inst_2697 ( .ZN(net_1778), .A(net_1686) );
DFF_X2 inst_3166 ( .D(net_1997), .QN(net_108), .CK(net_4533) );
XOR2_X2 inst_15 ( .A(net_1100), .B(net_1092), .Z(net_1087) );
AOI222_X1 inst_3747 ( .C1(net_3504), .B1(net_3472), .A1(net_3469), .A2(net_3136), .B2(net_3115), .ZN(net_2277), .C2(net_261) );
AOI22_X2 inst_3656 ( .ZN(net_598), .A1(net_597), .B1(net_596), .A2(net_571), .B2(net_570) );
INV_X4 inst_2237 ( .A(net_2144), .ZN(net_1779) );
CLKBUF_X2 inst_4417 ( .A(net_4402), .Z(net_4403) );
AOI22_X2 inst_3496 ( .A1(net_2249), .ZN(net_2211), .B1(net_2153), .A2(net_2141), .B2(net_297) );
INV_X8 inst_2123 ( .ZN(net_570), .A(net_367) );
DFF_X1 inst_3229 ( .QN(net_3066), .D(net_2958), .CK(net_4880) );
CLKBUF_X2 inst_4918 ( .A(net_4367), .Z(net_4904) );
INV_X2 inst_2706 ( .ZN(net_1665), .A(net_1664) );
AND2_X4 inst_4135 ( .ZN(net_4064), .A2(net_2522), .A1(net_2518) );
OAI21_X2 inst_476 ( .B1(net_3509), .B2(net_3208), .ZN(net_2974), .A(net_2494) );
AOI222_X1 inst_3742 ( .A1(net_4189), .C1(net_3504), .B1(net_3472), .ZN(net_2319), .A2(net_2037), .C2(net_393), .B2(net_228) );
INV_X4 inst_2499 ( .ZN(net_1439), .A(net_62) );
INV_X2 inst_2827 ( .A(net_3614), .ZN(net_522) );
XOR2_X2 inst_20 ( .Z(net_4037), .A(net_2379), .B(net_1782) );
INV_X4 inst_2448 ( .A(net_3082), .ZN(net_551) );
NAND3_X2 inst_1369 ( .A3(net_4004), .ZN(net_3987), .A2(net_3986), .A1(net_3395) );
AOI21_X2 inst_3988 ( .B2(net_923), .ZN(net_741), .A(net_740), .B1(net_655) );
OAI222_X2 inst_349 ( .C1(net_3784), .A2(net_2131), .ZN(net_1939), .A1(net_1815), .B1(net_1814), .B2(net_505), .C2(net_115) );
CLKBUF_X2 inst_4994 ( .A(net_4979), .Z(net_4980) );
INV_X4 inst_2541 ( .ZN(net_3399), .A(net_3102) );
OAI21_X2 inst_576 ( .B2(net_2917), .B1(net_2803), .ZN(net_2802), .A(net_2403) );
NAND2_X2 inst_1693 ( .A1(net_3293), .ZN(net_1977), .A2(net_227) );
CLKBUF_X2 inst_4249 ( .A(net_4217), .Z(net_4235) );
CLKBUF_X2 inst_4235 ( .A(net_4220), .Z(net_4221) );
INV_X4 inst_2561 ( .A(net_3858), .ZN(net_3514) );
DFF_X1 inst_3306 ( .QN(net_3018), .D(net_2865), .CK(net_5075) );
NOR2_X2 inst_1020 ( .A2(net_4089), .ZN(net_1854), .A1(net_1815) );
INV_X2 inst_2876 ( .A(net_3270), .ZN(net_262) );
INV_X2 inst_3055 ( .A(net_3943), .ZN(net_3929) );
NOR2_X4 inst_976 ( .A1(net_3997), .ZN(net_3935), .A2(net_3789) );
AOI21_X2 inst_3952 ( .B2(net_4086), .A(net_3963), .B1(net_1844), .ZN(net_1843) );
CLKBUF_X2 inst_4226 ( .A(net_4211), .Z(net_4212) );
NAND3_X2 inst_1279 ( .ZN(net_2748), .A1(net_2680), .A2(net_1518), .A3(net_1213) );
INV_X4 inst_2252 ( .ZN(net_1306), .A(net_1305) );
AOI22_X2 inst_3588 ( .A1(net_4062), .B1(net_4057), .ZN(net_1429), .B2(net_177), .A2(net_159) );
NOR2_X2 inst_1096 ( .A2(net_3164), .A1(net_3162), .ZN(net_338) );
CLKBUF_X2 inst_4229 ( .A(net_4214), .Z(net_4215) );
CLKBUF_X2 inst_4552 ( .A(net_4366), .Z(net_4538) );
INV_X4 inst_2238 ( .ZN(net_1862), .A(net_1815) );
CLKBUF_X2 inst_5207 ( .A(net_5192), .Z(net_5193) );
INV_X2 inst_2763 ( .ZN(net_1068), .A(net_962) );
CLKBUF_X2 inst_5072 ( .A(net_4791), .Z(net_5058) );
CLKBUF_X2 inst_4543 ( .A(net_4199), .Z(net_4529) );
NAND2_X2 inst_1839 ( .A1(net_4106), .ZN(net_1152), .A2(net_326) );
DFF_X2 inst_3151 ( .D(net_2257), .QN(net_192), .CK(net_4464) );
OAI21_X2 inst_761 ( .A(net_3989), .ZN(net_3783), .B2(net_3681), .B1(net_867) );
CLKBUF_X2 inst_4867 ( .A(net_4395), .Z(net_4853) );
DFF_X1 inst_3399 ( .Q(net_3118), .D(net_1534), .CK(net_4303) );
DFF_X1 inst_3414 ( .D(net_1361), .Q(net_30), .CK(net_4295) );
CLKBUF_X2 inst_4436 ( .A(net_4421), .Z(net_4422) );
CLKBUF_X2 inst_4495 ( .A(net_4480), .Z(net_4481) );
INV_X2 inst_2803 ( .A(net_844), .ZN(net_726) );
NAND2_X4 inst_1432 ( .A1(net_3769), .ZN(net_3663), .A2(net_3590) );
OAI21_X2 inst_725 ( .ZN(net_1400), .A(net_363), .B2(net_322), .B1(net_164) );
AND2_X4 inst_4120 ( .ZN(net_4043), .A1(net_2114), .A2(net_1611) );
INV_X1 inst_3084 ( .ZN(net_3689), .A(net_3688) );
CLKBUF_X2 inst_5097 ( .A(net_5082), .Z(net_5083) );
INV_X4 inst_2259 ( .ZN(net_1181), .A(net_1180) );
NAND3_X2 inst_1337 ( .ZN(net_3260), .A1(net_3257), .A2(net_2892), .A3(net_2890) );
INV_X4 inst_2464 ( .A(net_3070), .ZN(net_492) );
INV_X2 inst_2641 ( .ZN(net_2340), .A(net_2320) );
HA_X1 inst_3096 ( .B(net_3103), .S(net_1154), .CO(net_822), .A(net_688) );
INV_X2 inst_3015 ( .ZN(net_3402), .A(net_3010) );
AOI21_X2 inst_4010 ( .ZN(net_4161), .B1(net_2243), .A(net_2123), .B2(net_182) );
NAND2_X2 inst_1638 ( .ZN(net_2186), .A1(net_2185), .A2(net_1771) );
DFF_X1 inst_3328 ( .D(net_2807), .QN(net_292), .CK(net_4487) );
INV_X4 inst_2441 ( .A(net_3154), .ZN(net_218) );
NOR2_X2 inst_1111 ( .ZN(net_3314), .A1(net_3313), .A2(net_1509) );
DFF_X1 inst_3220 ( .QN(net_3060), .D(net_2975), .CK(net_4608) );
INV_X2 inst_2658 ( .ZN(net_2249), .A(net_2153) );
NOR3_X4 inst_878 ( .A3(net_3760), .A2(net_3754), .ZN(net_3603), .A1(net_268) );
CLKBUF_X2 inst_4959 ( .A(net_4363), .Z(net_4945) );
OAI21_X2 inst_480 ( .B1(net_2970), .ZN(net_2966), .B2(net_2965), .A(net_2444) );
NAND2_X2 inst_1926 ( .ZN(net_3189), .A1(net_3186), .A2(net_150) );
CLKBUF_X2 inst_4631 ( .A(net_4306), .Z(net_4617) );
CLKBUF_X2 inst_4351 ( .A(net_4336), .Z(net_4337) );
OAI21_X2 inst_564 ( .B2(net_2917), .B1(net_2849), .ZN(net_2848), .A(net_2396) );
INV_X2 inst_2986 ( .ZN(net_128), .A(net_74) );
CLKBUF_X2 inst_4783 ( .A(net_4768), .Z(net_4769) );
INV_X4 inst_2206 ( .ZN(net_2253), .A(net_2232) );
INV_X2 inst_2792 ( .A(net_965), .ZN(net_787) );
OAI21_X2 inst_739 ( .ZN(net_3241), .B1(net_3240), .B2(net_1975), .A(net_1720) );
AOI221_X2 inst_3862 ( .C2(net_3543), .ZN(net_2018), .B1(net_2017), .C1(net_2016), .A(net_1892), .B2(net_364) );
XNOR2_X2 inst_46 ( .A(net_3692), .ZN(net_2587), .B(net_1449) );
NOR2_X4 inst_934 ( .A2(net_4186), .ZN(net_915), .A1(net_796) );
INV_X4 inst_2537 ( .ZN(net_3349), .A(net_3348) );
NOR2_X2 inst_1000 ( .ZN(net_2031), .A1(net_1973), .A2(net_126) );
NOR2_X2 inst_1126 ( .ZN(net_3472), .A1(net_3471), .A2(net_1835) );
AOI22_X2 inst_3470 ( .B2(net_3120), .A1(net_2724), .B1(net_2722), .ZN(net_2720), .A2(net_31) );
CLKBUF_X2 inst_5304 ( .A(net_4742), .Z(net_5290) );
OAI211_X2 inst_796 ( .ZN(net_2273), .C2(net_2272), .B(net_2237), .C1(net_2190), .A(net_2006) );
INV_X4 inst_2585 ( .ZN(net_3653), .A(net_3169) );
OAI21_X2 inst_633 ( .ZN(net_2078), .B2(net_2076), .A(net_1967), .B1(net_1668) );
INV_X4 inst_2364 ( .ZN(net_691), .A(net_442) );
CLKBUF_X2 inst_4299 ( .A(net_4256), .Z(net_4285) );
OAI21_X2 inst_524 ( .B1(net_3302), .ZN(net_2913), .B2(net_2912), .A(net_2450) );
NAND2_X2 inst_1882 ( .A2(net_2037), .ZN(net_426), .A1(net_401) );
XNOR2_X2 inst_104 ( .B(net_3418), .ZN(net_452), .A(net_366) );
AND3_X4 inst_4060 ( .A1(net_4042), .A2(net_3506), .ZN(net_2534), .A3(net_2125) );
INV_X4 inst_2285 ( .A(net_1332), .ZN(net_1118) );
INV_X4 inst_2331 ( .A(net_2717), .ZN(net_847) );
CLKBUF_X2 inst_4478 ( .A(net_4463), .Z(net_4464) );
DFF_X1 inst_3344 ( .D(net_2779), .CK(net_4350), .Q(x90) );
NAND2_X2 inst_1499 ( .ZN(net_2818), .A1(net_2773), .A2(net_2716) );
INV_X4 inst_2377 ( .ZN(net_2737), .A(net_409) );
INV_X4 inst_2522 ( .ZN(net_3255), .A(net_3254) );
INV_X2 inst_2972 ( .ZN(net_238), .A(net_116) );
CLKBUF_X2 inst_4862 ( .A(net_4847), .Z(net_4848) );
OAI21_X2 inst_727 ( .B2(net_3662), .ZN(net_693), .A(net_424), .B1(net_368) );
CLKBUF_X2 inst_4663 ( .A(net_4648), .Z(net_4649) );
CLKBUF_X2 inst_4804 ( .A(net_4254), .Z(net_4790) );
NOR3_X2 inst_882 ( .ZN(net_2835), .A1(net_2786), .A2(net_2765), .A3(net_2712) );
INV_X2 inst_2874 ( .ZN(net_1173), .A(x1023) );
CLKBUF_X2 inst_4607 ( .A(net_4592), .Z(net_4593) );
INV_X4 inst_2431 ( .ZN(net_225), .A(net_44) );
DFF_X1 inst_3297 ( .QN(net_3007), .D(net_2886), .CK(net_5259) );
CLKBUF_X2 inst_5216 ( .A(net_4810), .Z(net_5202) );
INV_X2 inst_2938 ( .ZN(net_1507), .A(net_63) );
CLKBUF_X2 inst_5257 ( .A(net_5242), .Z(net_5243) );
CLKBUF_X2 inst_4423 ( .A(net_4334), .Z(net_4409) );
CLKBUF_X2 inst_5083 ( .A(net_5068), .Z(net_5069) );
NAND3_X2 inst_1346 ( .A3(net_3634), .A2(net_3620), .ZN(net_3431), .A1(net_1267) );
OAI21_X2 inst_708 ( .B2(net_4186), .A(net_3627), .B1(net_986), .ZN(net_971) );
AOI22_X2 inst_3523 ( .A2(net_3136), .B2(net_3111), .A1(net_1923), .ZN(net_1922), .B1(net_1921) );
CLKBUF_X2 inst_4855 ( .A(net_4840), .Z(net_4841) );
NAND3_X2 inst_1374 ( .ZN(net_4191), .A1(net_1290), .A3(net_593), .A2(net_178) );
NOR2_X4 inst_953 ( .A1(net_4157), .A2(net_3917), .ZN(net_3675) );
CLKBUF_X2 inst_5108 ( .A(net_4596), .Z(net_5094) );
CLKBUF_X2 inst_4342 ( .A(net_4327), .Z(net_4328) );
INV_X4 inst_2510 ( .A(net_3058), .ZN(net_567) );
AOI22_X2 inst_3510 ( .B1(net_3676), .B2(net_3134), .A1(net_2012), .ZN(net_2007), .A2(net_378) );
CLKBUF_X2 inst_4277 ( .A(net_4254), .Z(net_4263) );
NOR2_X2 inst_1071 ( .ZN(net_1176), .A1(net_750), .A2(net_399) );
CLKBUF_X2 inst_5060 ( .A(net_5045), .Z(net_5046) );
CLKBUF_X2 inst_4339 ( .A(net_4324), .Z(net_4325) );
CLKBUF_X2 inst_5291 ( .A(net_4543), .Z(net_5277) );
NAND2_X4 inst_1421 ( .ZN(net_3580), .A1(net_3579), .A2(net_2312) );
DFF_X1 inst_3373 ( .QN(net_3122), .D(net_2256), .CK(net_4481) );
NAND2_X2 inst_1994 ( .ZN(net_3481), .A2(net_3480), .A1(net_3479) );
CLKBUF_X2 inst_4902 ( .A(net_4355), .Z(net_4888) );
CLKBUF_X2 inst_4262 ( .A(net_4247), .Z(net_4248) );
CLKBUF_X2 inst_5298 ( .A(net_4298), .Z(net_5284) );
AOI22_X2 inst_3664 ( .A1(net_571), .B1(net_570), .ZN(net_563), .A2(net_219), .B2(net_160) );
CLKBUF_X2 inst_4720 ( .A(net_4705), .Z(net_4706) );
AOI22_X2 inst_3486 ( .A1(net_4038), .A2(net_3385), .B1(net_2657), .ZN(net_2650), .B2(net_361) );
INV_X8 inst_2162 ( .ZN(net_3654), .A(net_3653) );
CLKBUF_X2 inst_4986 ( .A(net_4545), .Z(net_4972) );
OAI221_X2 inst_392 ( .C2(net_3408), .B1(net_2361), .ZN(net_2360), .C1(net_2219), .A(net_1930), .B2(net_108) );
XNOR2_X2 inst_120 ( .ZN(net_4132), .B(net_290), .A(net_46) );
OAI22_X2 inst_294 ( .A1(net_3781), .B1(net_1884), .ZN(net_1742), .A2(net_1590), .B2(net_266) );
CLKBUF_X2 inst_4398 ( .A(net_4383), .Z(net_4384) );
AND2_X4 inst_4165 ( .ZN(net_4119), .A1(net_401), .A2(net_260) );
NAND2_X2 inst_1514 ( .ZN(net_2550), .A1(net_2549), .A2(net_2548) );
DFF_X1 inst_3384 ( .D(net_1897), .Q(net_83), .CK(net_4474) );
INV_X4 inst_2272 ( .ZN(net_1023), .A(net_972) );
NAND2_X2 inst_1608 ( .A1(net_2967), .ZN(net_2408), .A2(net_519) );
OAI21_X2 inst_567 ( .B2(net_2909), .B1(net_2849), .ZN(net_2845), .A(net_2467) );
DFF_X2 inst_3200 ( .QN(net_3108), .D(net_1629), .CK(net_4828) );
OAI211_X2 inst_810 ( .ZN(net_1630), .B(net_1628), .C1(net_1627), .A(net_1557), .C2(net_1124) );
OR2_X4 inst_230 ( .ZN(net_1826), .A1(net_412), .A2(net_389) );
NAND2_X2 inst_1601 ( .A1(net_2969), .ZN(net_2416), .A2(net_479) );
NAND2_X4 inst_1484 ( .ZN(net_4000), .A1(net_3999), .A2(net_3171) );
INV_X2 inst_3035 ( .ZN(net_3575), .A(net_3574) );
AOI22_X2 inst_3526 ( .A2(net_3138), .A1(net_1923), .B1(net_1921), .ZN(net_1918), .B2(net_1326) );
OAI211_X2 inst_856 ( .ZN(net_3758), .B(net_1628), .C1(net_1627), .A(net_1552), .C2(net_385) );
NAND2_X2 inst_1893 ( .ZN(net_533), .A2(net_385), .A1(net_334) );

endmodule
