module s510 (
cnt509,
pcnt12,
cnt283,
cnt44,
cnt13,
pcnt241,
blif_clk_net,
pcnt6,
cnt261,
john,
pcnt17,
cnt511,
cnt272,
cnt21,
cnt567,
cnt10,
cnt45,
pcnt27,
cnt284,
cnt591,
blif_reset_net,
cclr,
vsync,
cblank,
csync,
pc,
csm,
pclr);

// Start PIs
input cnt509;
input pcnt12;
input cnt283;
input cnt44;
input cnt13;
input pcnt241;
input blif_clk_net;
input pcnt6;
input cnt261;
input john;
input pcnt17;
input cnt511;
input cnt272;
input cnt21;
input cnt567;
input cnt10;
input cnt45;
input pcnt27;
input cnt284;
input cnt591;
input blif_reset_net;

// Start POs
output cclr;
output vsync;
output cblank;
output csync;
output pc;
output csm;
output pclr;

// Start wires
wire net_47;
wire net_176;
wire net_215;
wire net_137;
wire net_132;
wire net_54;
wire net_237;
wire net_105;
wire vsync;
wire net_129;
wire net_119;
wire net_98;
wire net_12;
wire net_151;
wire net_53;
wire net_93;
wire net_210;
wire net_168;
wire net_259;
wire net_269;
wire net_127;
wire pclr;
wire net_76;
wire net_101;
wire net_187;
wire net_111;
wire net_264;
wire net_90;
wire net_225;
wire net_283;
wire net_100;
wire net_85;
wire net_263;
wire net_252;
wire net_124;
wire net_240;
wire net_160;
wire net_221;
wire net_115;
wire net_4;
wire net_17;
wire net_164;
wire cnt13;
wire pcnt241;
wire net_87;
wire net_0;
wire net_35;
wire net_16;
wire net_239;
wire net_193;
wire net_157;
wire net_257;
wire net_233;
wire net_42;
wire net_120;
wire net_201;
wire net_109;
wire net_80;
wire net_65;
wire blif_reset_net;
wire net_50;
wire net_234;
wire net_96;
wire net_66;
wire net_38;
wire net_167;
wire net_207;
wire net_136;
wire net_280;
wire net_19;
wire net_126;
wire net_278;
wire net_34;
wire net_108;
wire net_270;
wire net_183;
wire net_150;
wire net_63;
wire net_274;
wire pcnt12;
wire net_30;
wire net_189;
wire net_24;
wire net_99;
wire net_186;
wire net_46;
wire net_118;
wire net_216;
wire net_146;
wire pcnt27;
wire net_122;
wire net_7;
wire net_224;
wire net_172;
wire net_52;
wire net_165;
wire pc;
wire net_13;
wire net_246;
wire net_94;
wire net_219;
wire net_18;
wire net_131;
wire net_114;
wire net_196;
wire net_29;
wire net_149;
wire net_142;
wire net_248;
wire net_31;
wire net_36;
wire net_158;
wire net_41;
wire net_198;
wire net_253;
wire net_276;
wire net_209;
wire net_3;
wire net_154;
wire john;
wire net_213;
wire net_238;
wire net_260;
wire net_28;
wire net_97;
wire net_182;
wire net_192;
wire net_60;
wire net_267;
wire net_273;
wire net_256;
wire net_58;
wire net_82;
wire net_64;
wire cnt567;
wire net_121;
wire cnt45;
wire net_73;
wire net_200;
wire net_177;
wire net_75;
wire net_86;
wire net_206;
wire net_195;
wire net_125;
wire net_107;
wire net_166;
wire net_223;
wire net_179;
wire net_235;
wire net_159;
wire net_61;
wire net_62;
wire net_6;
wire net_217;
wire net_271;
wire net_23;
wire cnt10;
wire net_117;
wire net_74;
wire net_250;
wire net_205;
wire net_135;
wire net_265;
wire net_242;
wire net_130;
wire cclr;
wire net_147;
wire net_14;
wire net_220;
wire net_26;
wire net_113;
wire blif_clk_net;
wire net_32;
wire csm;
wire net_40;
wire net_282;
wire net_69;
wire cblank;
wire cnt284;
wire net_161;
wire net_141;
wire net_83;
wire net_95;
wire net_173;
wire net_78;
wire net_27;
wire cnt44;
wire net_56;
wire net_155;
wire net_261;
wire net_191;
wire net_22;
wire net_181;
wire net_39;
wire net_245;
wire net_2;
wire net_102;
wire net_144;
wire net_227;
wire net_9;
wire net_59;
wire net_162;
wire net_230;
wire net_44;
wire net_277;
wire net_134;
wire net_199;
wire net_45;
wire net_89;
wire cnt272;
wire net_185;
wire net_272;
wire net_178;
wire net_236;
wire net_208;
wire net_212;
wire net_243;
wire cnt283;
wire net_222;
wire net_152;
wire net_116;
wire net_175;
wire net_91;
wire net_55;
wire net_106;
wire net_258;
wire net_255;
wire net_140;
wire net_266;
wire net_247;
wire pcnt17;
wire net_279;
wire net_104;
wire net_148;
wire net_72;
wire net_25;
wire net_229;
wire net_70;
wire net_251;
wire net_194;
wire net_241;
wire net_5;
wire net_244;
wire net_128;
wire net_138;
wire pcnt6;
wire net_184;
wire net_11;
wire net_123;
wire csync;
wire net_262;
wire net_170;
wire net_68;
wire net_77;
wire net_214;
wire net_249;
wire net_20;
wire net_49;
wire net_15;
wire net_275;
wire net_57;
wire net_71;
wire net_153;
wire net_156;
wire net_84;
wire net_218;
wire cnt261;
wire net_174;
wire net_231;
wire net_92;
wire net_1;
wire net_112;
wire net_103;
wire net_139;
wire net_226;
wire net_43;
wire net_228;
wire net_10;
wire net_180;
wire net_21;
wire net_169;
wire net_51;
wire net_79;
wire net_171;
wire net_143;
wire cnt509;
wire net_190;
wire net_88;
wire net_145;
wire net_281;
wire net_197;
wire net_204;
wire net_81;
wire net_232;
wire net_163;
wire net_254;
wire net_67;
wire net_37;
wire net_202;
wire net_268;
wire cnt511;
wire cnt21;
wire net_188;
wire net_110;
wire net_48;
wire net_33;
wire net_8;
wire net_211;
wire cnt591;
wire net_133;
wire net_203;

// Start cells
DFFR_X2 inst_257 ( .QN(net_238), .RN(net_235), .D(net_232), .CK(net_275) );
CLKBUF_X2 inst_290 ( .A(net_282), .Z(net_283) );
NAND2_X2 inst_145 ( .ZN(net_188), .A1(net_110), .A2(net_34) );
CLKBUF_X2 inst_272 ( .A(net_264), .Z(net_265) );
NAND2_X2 inst_103 ( .ZN(net_254), .A1(net_23), .A2(net_0) );
INV_X2 inst_248 ( .ZN(net_246), .A(net_142) );
INV_X2 inst_228 ( .A(net_79), .ZN(net_12) );
NAND2_X2 inst_125 ( .ZN(net_108), .A1(net_96), .A2(net_71) );
INV_X4 inst_207 ( .ZN(net_192), .A(net_149) );
NAND2_X2 inst_138 ( .ZN(net_160), .A1(net_159), .A2(net_157) );
NAND2_X2 inst_159 ( .ZN(net_228), .A1(net_211), .A2(net_209) );
NAND2_X2 inst_134 ( .A2(net_225), .ZN(net_146), .A1(net_127) );
INV_X2 inst_244 ( .ZN(net_125), .A(net_111) );
NAND2_X2 inst_131 ( .ZN(net_128), .A1(net_127), .A2(net_89) );
INV_X4 inst_214 ( .ZN(net_159), .A(net_115) );
INV_X4 inst_180 ( .A(net_238), .ZN(net_104) );
NAND2_X1 inst_160 ( .ZN(net_9), .A1(pcnt17), .A2(cnt284) );
NOR2_X2 inst_33 ( .ZN(net_88), .A2(net_43), .A1(net_23) );
NOR2_X2 inst_47 ( .ZN(net_135), .A2(net_81), .A1(net_18) );
NOR3_X2 inst_19 ( .ZN(net_239), .A1(net_231), .A3(net_230), .A2(net_228) );
OR2_X2 inst_8 ( .ZN(net_171), .A2(net_170), .A1(net_67) );
INV_X2 inst_232 ( .A(net_199), .ZN(net_34) );
INV_X2 inst_247 ( .ZN(net_212), .A(net_113) );
NOR2_X4 inst_27 ( .A2(net_253), .ZN(net_148), .A1(net_142) );
NAND2_X2 inst_100 ( .ZN(net_15), .A2(net_6), .A1(cnt44) );
CLKBUF_X2 inst_279 ( .A(net_271), .Z(net_272) );
INV_X1 inst_253 ( .ZN(net_235), .A(blif_reset_net) );
INV_X4 inst_211 ( .ZN(net_115), .A(net_86) );
INV_X8 inst_162 ( .ZN(net_60), .A(net_11) );
NAND2_X4 inst_93 ( .A2(net_245), .ZN(net_78), .A1(net_57) );
NAND3_X2 inst_81 ( .ZN(net_208), .A2(net_207), .A3(net_122), .A1(net_55) );
NAND2_X2 inst_139 ( .ZN(net_165), .A1(net_106), .A2(net_83) );
NAND2_X2 inst_155 ( .ZN(net_206), .A2(net_155), .A1(net_149) );
NOR2_X2 inst_59 ( .ZN(net_223), .A2(net_217), .A1(net_150) );
NAND2_X2 inst_135 ( .A1(net_207), .ZN(net_151), .A2(net_93) );
INV_X4 inst_196 ( .A(net_173), .ZN(net_49) );
NOR2_X2 inst_55 ( .ZN(net_191), .A2(net_147), .A1(net_97) );
NOR2_X2 inst_37 ( .A2(net_199), .A1(net_100), .ZN(net_61) );
INV_X2 inst_237 ( .ZN(net_63), .A(net_62) );
NAND2_X2 inst_148 ( .ZN(net_194), .A1(net_141), .A2(net_103) );
AND2_X4 inst_264 ( .A2(net_261), .ZN(net_40), .A1(net_10) );
INV_X4 inst_191 ( .ZN(net_102), .A(net_74) );
NAND3_X2 inst_84 ( .ZN(net_218), .A3(net_197), .A1(net_161), .A2(net_158) );
NOR2_X2 inst_51 ( .ZN(net_147), .A2(net_118), .A1(cnt284) );
NAND2_X2 inst_142 ( .ZN(net_177), .A2(net_154), .A1(net_140) );
NAND3_X2 inst_80 ( .A3(net_252), .A1(net_251), .ZN(net_204), .A2(net_73) );
INV_X4 inst_173 ( .ZN(net_23), .A(net_13) );
INV_X2 inst_224 ( .ZN(net_4), .A(cnt511) );
INV_X4 inst_216 ( .ZN(net_141), .A(net_140) );
NAND3_X2 inst_78 ( .ZN(net_193), .A2(net_192), .A1(net_168), .A3(net_153) );
CLKBUF_X2 inst_287 ( .A(net_273), .Z(net_280) );
NOR2_X2 inst_42 ( .ZN(net_120), .A1(net_62), .A2(net_24) );
INV_X2 inst_241 ( .A(net_105), .ZN(net_77) );
INV_X4 inst_177 ( .ZN(net_14), .A(net_13) );
INV_X2 inst_231 ( .A(net_40), .ZN(net_32) );
CLKBUF_X2 inst_270 ( .A(blif_clk_net), .Z(net_263) );
INV_X4 inst_183 ( .ZN(net_52), .A(net_24) );
NOR2_X4 inst_26 ( .ZN(net_249), .A1(net_65), .A2(net_60) );
NAND2_X2 inst_151 ( .ZN(net_197), .A2(net_128), .A1(net_33) );
NOR2_X1 inst_64 ( .ZN(net_182), .A1(net_181), .A2(net_167) );
NAND2_X2 inst_107 ( .A1(net_98), .ZN(net_64), .A2(net_40) );
NAND4_X2 inst_70 ( .ZN(net_233), .A2(net_225), .A4(net_224), .A1(net_223), .A3(net_179) );
NAND2_X2 inst_129 ( .ZN(net_124), .A2(net_123), .A1(net_96) );
NAND2_X4 inst_92 ( .A2(net_244), .ZN(net_65), .A1(net_38) );
INV_X4 inst_189 ( .A(net_57), .ZN(net_47) );
INV_X2 inst_223 ( .ZN(net_3), .A(cnt591) );
NOR4_X2 inst_11 ( .ZN(net_215), .A4(net_183), .A1(net_176), .A2(net_145), .A3(net_119) );
INV_X4 inst_188 ( .ZN(net_75), .A(net_23) );
NOR3_X2 inst_14 ( .A2(net_173), .ZN(net_132), .A1(net_131), .A3(net_98) );
NOR2_X2 inst_31 ( .A2(net_262), .ZN(net_41), .A1(net_23) );
INV_X2 inst_252 ( .ZN(net_176), .A(net_175) );
NAND2_X2 inst_158 ( .A1(net_257), .ZN(net_227), .A2(net_199) );
NAND2_X2 inst_141 ( .ZN(net_174), .A2(net_172), .A1(net_149) );
NOR2_X1 inst_62 ( .A1(net_238), .ZN(net_53), .A2(net_27) );
INV_X4 inst_200 ( .A(net_49), .ZN(net_48) );
INV_X2 inst_251 ( .ZN(net_175), .A(net_159) );
CLKBUF_X2 inst_286 ( .A(net_278), .Z(net_279) );
NOR2_X2 inst_57 ( .ZN(net_210), .A2(net_195), .A1(net_152) );
NAND2_X2 inst_102 ( .A2(net_261), .A1(net_260), .ZN(net_44) );
NOR2_X2 inst_32 ( .ZN(net_30), .A2(net_29), .A1(john) );
NAND2_X2 inst_144 ( .ZN(net_184), .A2(net_183), .A1(net_159) );
INV_X4 inst_195 ( .A(net_44), .ZN(net_35) );
NOR2_X4 inst_21 ( .A1(net_261), .A2(net_260), .ZN(net_38) );
CLKBUF_X2 inst_281 ( .A(net_272), .Z(net_274) );
NAND2_X4 inst_97 ( .ZN(net_255), .A1(net_120), .A2(net_96) );
NAND2_X2 inst_124 ( .ZN(net_256), .A1(net_104), .A2(net_63) );
NOR3_X2 inst_18 ( .ZN(net_243), .A1(net_164), .A3(net_162), .A2(net_61) );
INV_X4 inst_208 ( .ZN(net_87), .A(net_78) );
NAND3_X2 inst_88 ( .A3(net_240), .A1(net_239), .ZN(net_236), .A2(net_210) );
INV_X2 inst_220 ( .ZN(net_0), .A(cnt21) );
OR2_X2 inst_9 ( .ZN(net_179), .A1(net_178), .A2(net_170) );
NAND2_X2 inst_113 ( .A2(net_173), .A1(net_102), .ZN(net_72) );
INV_X4 inst_198 ( .ZN(net_207), .A(net_49) );
NOR2_X2 inst_50 ( .A1(net_149), .ZN(net_145), .A2(net_144) );
NAND2_X2 inst_137 ( .ZN(net_158), .A2(net_157), .A1(net_96) );
INV_X2 inst_245 ( .A(net_225), .ZN(net_103) );
NAND2_X2 inst_130 ( .A2(net_186), .ZN(net_126), .A1(net_125) );
INV_X2 inst_227 ( .ZN(net_6), .A(pcnt12) );
INV_X2 inst_226 ( .ZN(net_5), .A(pcnt17) );
DFFR_X2 inst_260 ( .QN(net_259), .D(net_236), .RN(net_235), .CK(net_273) );
INV_X4 inst_176 ( .A(net_13), .ZN(net_10) );
NOR2_X2 inst_58 ( .ZN(net_217), .A1(net_192), .A2(net_191) );
NAND2_X2 inst_147 ( .ZN(net_190), .A2(net_146), .A1(net_144) );
NAND3_X2 inst_87 ( .ZN(net_232), .A3(net_221), .A1(net_203), .A2(net_134) );
NOR2_X2 inst_61 ( .A1(net_241), .ZN(net_230), .A2(net_96) );
INV_X4 inst_203 ( .ZN(net_137), .A(net_75) );
INV_X4 inst_212 ( .ZN(net_131), .A(net_87) );
INV_X2 inst_234 ( .ZN(net_51), .A(net_50) );
OR3_X2 inst_0 ( .ZN(net_219), .A1(net_207), .A2(net_175), .A3(net_125) );
INV_X4 inst_184 ( .ZN(net_37), .A(net_26) );
INV_X2 inst_236 ( .A(net_68), .ZN(net_56) );
NOR4_X2 inst_10 ( .A3(net_199), .ZN(net_195), .A2(net_163), .A4(net_45), .A1(net_30) );
OR2_X2 inst_4 ( .ZN(net_91), .A2(net_90), .A1(net_52) );
NOR2_X1 inst_65 ( .A2(net_219), .A1(net_186), .ZN(csm) );
NOR2_X2 inst_28 ( .ZN(net_17), .A1(net_4), .A2(pcnt241) );
INV_X2 inst_242 ( .ZN(net_81), .A(net_80) );
CLKBUF_X2 inst_275 ( .A(net_267), .Z(net_268) );
NAND2_X2 inst_117 ( .ZN(net_89), .A2(net_88), .A1(net_16) );
NAND2_X4 inst_98 ( .ZN(net_251), .A1(net_249), .A2(cnt10) );
AND3_X2 inst_263 ( .ZN(net_117), .A1(net_116), .A2(net_96), .A3(net_88) );
INV_X4 inst_190 ( .ZN(net_100), .A(net_31) );
INV_X4 inst_204 ( .ZN(net_149), .A(net_75) );
INV_X4 inst_185 ( .ZN(net_25), .A(net_24) );
NOR2_X2 inst_49 ( .ZN(net_200), .A1(net_84), .A2(net_75) );
NAND2_X2 inst_154 ( .ZN(net_203), .A2(net_180), .A1(net_49) );
NOR3_X2 inst_13 ( .ZN(net_157), .A3(net_78), .A1(net_29), .A2(net_19) );
NAND3_X2 inst_75 ( .ZN(net_106), .A1(net_105), .A3(net_104), .A2(cnt509) );
INV_X4 inst_166 ( .ZN(net_253), .A(cnt45) );
NAND2_X2 inst_116 ( .ZN(net_129), .A2(net_53), .A1(net_52) );
INV_X8 inst_163 ( .A(net_261), .ZN(net_26) );
NOR2_X2 inst_54 ( .A2(net_172), .ZN(net_166), .A1(net_133) );
NAND3_X2 inst_79 ( .A1(net_246), .ZN(net_198), .A2(pcnt6), .A3(cnt284) );
NAND2_X2 inst_109 ( .ZN(net_127), .A1(net_52), .A2(net_41) );
NAND2_X2 inst_106 ( .A1(net_238), .ZN(net_39), .A2(net_38) );
INV_X2 inst_219 ( .A(net_249), .ZN(net_248) );
INV_X4 inst_201 ( .ZN(net_168), .A(net_49) );
NOR2_X2 inst_43 ( .A2(net_258), .ZN(net_95), .A1(net_64) );
DFFR_X2 inst_255 ( .QN(net_262), .RN(net_235), .D(net_222), .CK(net_283) );
NAND2_X2 inst_128 ( .ZN(net_114), .A2(net_80), .A1(cnt567) );
NAND3_X2 inst_73 ( .ZN(net_73), .A3(net_40), .A1(net_25), .A2(cnt21) );
DFFR_X2 inst_256 ( .QN(net_237), .RN(net_235), .D(net_229), .CK(net_279) );
NOR2_X4 inst_23 ( .ZN(net_70), .A1(net_44), .A2(net_43) );
NAND2_X4 inst_94 ( .ZN(net_225), .A1(net_178), .A2(net_47) );
AND3_X4 inst_262 ( .ZN(net_226), .A2(net_225), .A3(net_206), .A1(net_201) );
INV_X2 inst_243 ( .ZN(net_93), .A(net_92) );
CLKBUF_X2 inst_285 ( .A(net_277), .Z(net_278) );
NOR3_X2 inst_15 ( .ZN(net_150), .A2(net_149), .A3(net_116), .A1(net_48) );
INV_X4 inst_218 ( .ZN(net_231), .A(net_227) );
INV_X4 inst_197 ( .A(net_49), .ZN(net_42) );
INV_X2 inst_250 ( .A(net_172), .ZN(net_122) );
INV_X4 inst_179 ( .A(net_238), .ZN(net_29) );
NOR2_X4 inst_24 ( .ZN(net_46), .A1(net_37), .A2(net_11) );
OR2_X2 inst_6 ( .ZN(net_155), .A1(net_154), .A2(net_153) );
NAND2_X2 inst_114 ( .ZN(net_92), .A1(net_75), .A2(net_74) );
INV_X4 inst_194 ( .A(net_98), .ZN(net_54) );
NAND3_X2 inst_76 ( .A2(net_192), .ZN(net_134), .A1(net_133), .A3(net_111) );
NAND2_X2 inst_150 ( .A2(net_256), .A1(net_255), .ZN(net_247) );
INV_X4 inst_172 ( .A(net_79), .ZN(net_8) );
CLKBUF_X2 inst_277 ( .A(net_269), .Z(net_270) );
NAND3_X2 inst_83 ( .ZN(net_214), .A3(net_213), .A1(net_174), .A2(net_102) );
NAND2_X2 inst_121 ( .ZN(net_101), .A2(net_100), .A1(net_86) );
NAND2_X2 inst_123 ( .ZN(net_163), .A2(net_107), .A1(net_52) );
OR3_X1 inst_2 ( .A1(net_216), .A3(net_212), .A2(net_143), .ZN(cclr) );
NAND3_X2 inst_86 ( .A2(net_219), .A1(net_194), .A3(net_171), .ZN(cblank) );
NAND2_X2 inst_118 ( .ZN(net_113), .A2(net_70), .A1(net_7) );
NOR2_X4 inst_20 ( .A1(net_260), .ZN(net_98), .A2(net_21) );
NAND2_X2 inst_153 ( .ZN(net_202), .A2(net_200), .A1(net_42) );
NOR2_X2 inst_38 ( .ZN(net_154), .A1(net_74), .A2(net_36) );
NOR2_X2 inst_52 ( .A2(net_248), .ZN(net_162), .A1(net_17) );
NAND2_X4 inst_90 ( .A1(net_250), .A2(net_238), .ZN(net_43) );
AND2_X4 inst_267 ( .ZN(net_59), .A1(net_57), .A2(net_3) );
NAND2_X2 inst_140 ( .ZN(net_213), .A1(net_173), .A2(net_172) );
INV_X4 inst_209 ( .ZN(net_111), .A(net_76) );
DFFR_X2 inst_259 ( .QN(net_260), .RN(net_235), .D(net_234), .CK(net_270) );
INV_X2 inst_221 ( .ZN(net_1), .A(cnt567) );
NOR2_X2 inst_40 ( .ZN(net_123), .A2(net_39), .A1(net_23) );
INV_X4 inst_167 ( .A(net_262), .ZN(net_79) );
INV_X2 inst_246 ( .A(net_131), .ZN(net_110) );
CLKBUF_X2 inst_289 ( .A(net_281), .Z(net_282) );
NAND2_X4 inst_95 ( .A2(net_186), .ZN(net_142), .A1(net_46) );
OR3_X1 inst_1 ( .A3(net_212), .A2(net_182), .A1(net_166), .ZN(pc) );
CLKBUF_X2 inst_282 ( .A(net_274), .Z(net_275) );
NAND4_X2 inst_72 ( .A4(net_243), .A1(net_242), .ZN(net_234), .A2(net_205), .A3(net_112) );
NOR2_X2 inst_44 ( .ZN(net_97), .A2(net_96), .A1(net_76) );
CLKBUF_X2 inst_274 ( .A(net_266), .Z(net_267) );
INV_X4 inst_174 ( .ZN(net_244), .A(net_13) );
NAND2_X2 inst_115 ( .A1(net_96), .ZN(net_82), .A2(net_56) );
INV_X2 inst_235 ( .ZN(net_55), .A(net_54) );
INV_X4 inst_210 ( .A(net_86), .ZN(net_84) );
INV_X8 inst_164 ( .ZN(net_57), .A(net_26) );
OR2_X2 inst_5 ( .A2(net_127), .ZN(net_94), .A1(net_68) );
CLKBUF_X2 inst_278 ( .A(net_264), .Z(net_271) );
NAND2_X2 inst_157 ( .A2(net_208), .A1(net_94), .ZN(pclr) );
INV_X2 inst_239 ( .A(net_127), .ZN(net_69) );
NAND2_X2 inst_105 ( .ZN(net_62), .A2(net_37), .A1(net_31) );
NAND4_X2 inst_68 ( .ZN(net_222), .A4(net_193), .A2(net_169), .A1(net_160), .A3(net_156) );
INV_X4 inst_213 ( .ZN(net_172), .A(net_99) );
NOR2_X2 inst_53 ( .ZN(net_164), .A2(net_163), .A1(cnt13) );
INV_X4 inst_175 ( .ZN(net_96), .A(net_79) );
INV_X4 inst_205 ( .ZN(net_80), .A(net_64) );
INV_X1 inst_254 ( .ZN(net_107), .A(net_65) );
INV_X2 inst_225 ( .ZN(net_258), .A(cnt283) );
NAND2_X2 inst_133 ( .A2(net_249), .ZN(net_136), .A1(cnt511) );
NAND2_X2 inst_112 ( .ZN(net_116), .A1(net_68), .A2(net_44) );
NAND4_X2 inst_67 ( .ZN(net_221), .A3(net_213), .A4(net_189), .A2(net_115), .A1(net_72) );
INV_X4 inst_181 ( .ZN(net_245), .A(net_23) );
NAND2_X2 inst_127 ( .ZN(net_112), .A1(net_111), .A2(net_69) );
NOR2_X2 inst_29 ( .ZN(net_18), .A1(net_1), .A2(pcnt27) );
INV_X4 inst_186 ( .ZN(net_173), .A(net_29) );
NOR3_X2 inst_17 ( .ZN(net_205), .A2(net_138), .A3(net_135), .A1(net_132) );
NAND2_X2 inst_146 ( .ZN(net_189), .A2(net_139), .A1(net_100) );
INV_X2 inst_249 ( .ZN(net_119), .A(net_118) );
INV_X4 inst_202 ( .ZN(net_144), .A(net_102) );
INV_X4 inst_187 ( .ZN(net_27), .A(net_26) );
INV_X4 inst_206 ( .ZN(net_86), .A(net_52) );
NAND2_X2 inst_122 ( .ZN(net_170), .A1(net_102), .A2(net_87) );
NAND2_X2 inst_126 ( .ZN(net_109), .A2(net_107), .A1(net_28) );
NOR2_X4 inst_25 ( .ZN(net_105), .A2(net_60), .A1(net_50) );
INV_X2 inst_240 ( .ZN(net_71), .A(net_70) );
NAND2_X2 inst_110 ( .A1(net_260), .ZN(net_90), .A2(net_41) );
NAND3_X2 inst_74 ( .ZN(net_83), .A1(net_66), .A3(net_35), .A2(cnt45) );
CLKBUF_X2 inst_288 ( .A(net_280), .Z(net_281) );
INV_X2 inst_229 ( .A(net_260), .ZN(net_19) );
NAND2_X4 inst_99 ( .A1(net_247), .ZN(net_211), .A2(cnt44) );
NOR2_X2 inst_35 ( .ZN(net_178), .A2(net_79), .A1(net_52) );
NAND4_X2 inst_69 ( .ZN(net_229), .A4(net_214), .A2(net_202), .A3(net_190), .A1(net_184) );
NOR2_X2 inst_48 ( .A2(net_225), .ZN(net_138), .A1(net_137) );
NAND3_X2 inst_82 ( .ZN(net_257), .A1(net_198), .A2(net_136), .A3(net_114) );
NOR2_X2 inst_46 ( .ZN(net_153), .A2(net_116), .A1(net_79) );
NOR2_X2 inst_30 ( .ZN(net_20), .A2(net_12), .A1(net_2) );
NAND2_X2 inst_136 ( .ZN(net_156), .A1(net_149), .A2(net_108) );
NAND2_X2 inst_108 ( .A1(net_238), .ZN(net_66), .A2(net_22) );
INV_X2 inst_233 ( .A(net_43), .ZN(net_36) );
INV_X4 inst_165 ( .A(net_259), .ZN(net_13) );
CLKBUF_X2 inst_271 ( .A(net_263), .Z(net_264) );
CLKBUF_X2 inst_283 ( .A(net_272), .Z(net_276) );
NOR2_X4 inst_22 ( .A1(net_260), .ZN(net_31), .A2(net_13) );
NOR2_X2 inst_34 ( .ZN(net_45), .A2(net_20), .A1(cnt10) );
NOR3_X4 inst_12 ( .ZN(net_241), .A1(net_204), .A3(net_148), .A2(net_95) );
NAND4_X2 inst_71 ( .A2(net_226), .A4(net_188), .A1(net_124), .A3(net_90), .ZN(csync) );
NOR2_X2 inst_56 ( .ZN(net_240), .A2(net_187), .A1(net_117) );
NAND2_X2 inst_104 ( .A2(net_238), .ZN(net_28), .A1(cnt13) );
NOR2_X2 inst_60 ( .ZN(net_242), .A2(net_220), .A1(net_121) );
INV_X4 inst_168 ( .A(net_237), .ZN(net_11) );
INV_X4 inst_169 ( .ZN(net_250), .A(net_11) );
INV_X4 inst_215 ( .A(net_149), .ZN(net_140) );
NAND2_X1 inst_161 ( .ZN(net_139), .A2(net_99), .A1(net_74) );
NOR3_X2 inst_16 ( .ZN(net_152), .A3(net_129), .A1(net_92), .A2(cnt261) );
CLKBUF_X2 inst_276 ( .A(net_268), .Z(net_269) );
OR2_X4 inst_3 ( .A2(net_262), .ZN(net_22), .A1(net_21) );
NAND2_X2 inst_156 ( .ZN(net_209), .A2(net_165), .A1(net_137) );
INV_X4 inst_170 ( .A(net_79), .ZN(net_7) );
DFFR_X2 inst_258 ( .QN(net_261), .RN(net_235), .D(net_233), .CK(net_265) );
NOR2_X2 inst_41 ( .ZN(net_85), .A2(net_59), .A1(net_58) );
INV_X4 inst_199 ( .ZN(net_76), .A(net_47) );
NAND2_X4 inst_91 ( .A2(net_260), .ZN(net_50), .A1(net_26) );
NAND2_X2 inst_132 ( .ZN(net_130), .A1(net_129), .A2(net_113) );
NAND2_X2 inst_143 ( .ZN(net_180), .A2(net_101), .A1(net_32) );
NOR2_X2 inst_36 ( .ZN(net_58), .A1(net_57), .A2(cnt272) );
NAND2_X2 inst_152 ( .ZN(net_201), .A1(net_200), .A2(net_199) );
AND2_X4 inst_265 ( .A2(net_260), .ZN(net_186), .A1(net_14) );
NAND2_X4 inst_96 ( .A2(net_254), .ZN(net_252), .A1(net_105) );
NOR2_X2 inst_45 ( .A2(net_199), .ZN(net_183), .A1(net_111) );
NAND2_X2 inst_101 ( .ZN(net_16), .A2(net_5), .A1(cnt284) );
AND2_X2 inst_269 ( .ZN(net_161), .A2(net_109), .A1(net_77) );
INV_X2 inst_238 ( .ZN(net_67), .A(net_66) );
AND4_X2 inst_261 ( .ZN(net_187), .A3(net_186), .A2(net_178), .A1(net_173), .A4(net_85) );
INV_X4 inst_178 ( .A(net_60), .ZN(net_24) );
NAND3_X1 inst_89 ( .A1(net_215), .A3(net_126), .A2(net_82), .ZN(vsync) );
NAND2_X2 inst_111 ( .A1(net_173), .ZN(net_133), .A2(net_54) );
NAND4_X2 inst_66 ( .ZN(net_216), .A3(net_181), .A2(net_177), .A1(net_151), .A4(net_131) );
AND2_X2 inst_268 ( .ZN(net_121), .A2(net_120), .A1(net_15) );
OR2_X2 inst_7 ( .ZN(net_169), .A1(net_168), .A2(net_167) );
NOR2_X1 inst_63 ( .A1(net_207), .ZN(net_143), .A2(net_142) );
INV_X4 inst_182 ( .ZN(net_74), .A(net_19) );
CLKBUF_X2 inst_273 ( .A(net_265), .Z(net_266) );
NAND2_X2 inst_120 ( .ZN(net_167), .A1(net_111), .A2(net_98) );
NAND2_X2 inst_119 ( .A1(net_238), .ZN(net_118), .A2(net_51) );
CLKBUF_X2 inst_284 ( .A(net_276), .Z(net_277) );
INV_X2 inst_222 ( .ZN(net_2), .A(john) );
INV_X4 inst_192 ( .A(net_74), .ZN(net_33) );
CLKBUF_X2 inst_280 ( .A(net_272), .Z(net_273) );
NAND3_X2 inst_85 ( .ZN(net_220), .A3(net_196), .A2(net_185), .A1(net_91) );
AND2_X4 inst_266 ( .A2(net_238), .ZN(net_199), .A1(net_8) );
NAND2_X2 inst_149 ( .ZN(net_196), .A2(net_130), .A1(net_23) );
INV_X4 inst_193 ( .ZN(net_181), .A(net_41) );
NOR2_X2 inst_39 ( .ZN(net_99), .A1(net_79), .A2(net_78) );
INV_X2 inst_230 ( .ZN(net_68), .A(net_38) );
INV_X4 inst_217 ( .ZN(net_224), .A(net_218) );
NAND3_X2 inst_77 ( .ZN(net_185), .A3(net_123), .A2(net_52), .A1(net_9) );
INV_X4 inst_171 ( .ZN(net_21), .A(net_11) );

endmodule
