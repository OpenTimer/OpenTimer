module c7552_slack (
n94,
n18,
n172,
n61,
n188,
n133,
n53,
n178,
n55,
n213,
n63,
n239,
n220,
n65,
n231,
n208,
n113,
n162,
n184,
n74,
n1,
n3749,
n2230,
n160,
n80,
n4394,
n226,
n210,
n150,
n78,
n109,
n89,
n114,
n176,
n3711,
n180,
n2239,
n141,
n153,
n83,
n2224,
n3729,
n3723,
n124,
n2247,
n103,
n216,
n223,
n157,
n196,
n155,
n69,
n197,
n81,
n4420,
n32,
n202,
n4405,
n190,
n76,
n240,
n4526,
n57,
n9,
n111,
n1486,
n1492,
n151,
n12,
n2236,
n2211,
n205,
n191,
n29,
n234,
n206,
n97,
n177,
n147,
n232,
n47,
n50,
n4437,
n2208,
n159,
n73,
n173,
n62,
n4400,
n228,
n87,
n23,
n193,
n130,
n38,
n4410,
n127,
n2204,
n219,
n4432,
n179,
n227,
n118,
n1469,
n4528,
n238,
n161,
n201,
n88,
n54,
n237,
n169,
n2218,
n75,
n64,
n60,
n82,
n3743,
n1480,
n189,
n1197,
n171,
n134,
n221,
n230,
n175,
n212,
n4427,
n112,
n167,
n35,
n166,
n135,
n154,
n164,
n85,
n4415,
n222,
n1462,
n185,
n203,
n152,
n170,
n199,
n2256,
n181,
n187,
n214,
n3698,
n100,
n211,
n3737,
n1496,
n115,
n207,
n1459,
n217,
n168,
n26,
n195,
n209,
n163,
n198,
n2253,
n183,
n182,
n215,
n218,
n3701,
n86,
n59,
n5,
n4393,
n165,
n110,
n158,
n1455,
n121,
n84,
n58,
n15,
n144,
n79,
n41,
n3705,
n229,
n138,
n66,
n56,
n192,
n194,
n186,
n77,
n3717,
n106,
n235,
n204,
n70,
n224,
n233,
n156,
n174,
n225,
n44,
n236,
n200,
n408,
n399,
n278,
n2,
n370,
n350,
n319,
n522,
n307,
n368,
n556,
n406,
n471,
n436,
n540,
n412,
n304,
n292,
n532,
n528,
n480,
n422,
n404,
n432,
n444,
n333,
n488,
n391,
n276,
n558,
n486,
n258,
n560,
n362,
n281,
n546,
n330,
n448,
n289,
n341,
n324,
n554,
n526,
n264,
n496,
n442,
n410,
n524,
n416,
n538,
n3,
n552,
n469,
n382,
n492,
n414,
n246,
n286,
n295,
n394,
n536,
n249,
n327,
n365,
n453,
n313,
n279,
n379,
n548,
n298,
n356,
n373,
n252,
n446,
n321,
n438,
n284,
n530,
n450,
n550,
n359,
n336,
n534,
n301,
n344,
n397,
n338,
n418,
n490,
n542,
n440,
n388,
n484,
n270,
n385,
n482,
n478,
n347,
n544,
n316,
n310,
n402,
n494,
n419,
n273,
n353,
n376);

// Start PIs
input n94;
input n18;
input n172;
input n61;
input n188;
input n133;
input n53;
input n178;
input n55;
input n213;
input n63;
input n239;
input n220;
input n65;
input n231;
input n208;
input n113;
input n162;
input n184;
input n74;
input n1;
input n3749;
input n2230;
input n160;
input n80;
input n4394;
input n226;
input n210;
input n150;
input n78;
input n109;
input n89;
input n114;
input n176;
input n3711;
input n180;
input n2239;
input n141;
input n153;
input n83;
input n2224;
input n3729;
input n3723;
input n124;
input n2247;
input n103;
input n216;
input n223;
input n157;
input n196;
input n155;
input n69;
input n197;
input n81;
input n4420;
input n32;
input n202;
input n4405;
input n190;
input n76;
input n240;
input n4526;
input n57;
input n9;
input n111;
input n1486;
input n1492;
input n151;
input n12;
input n2236;
input n2211;
input n205;
input n191;
input n29;
input n234;
input n206;
input n97;
input n177;
input n147;
input n232;
input n47;
input n50;
input n4437;
input n2208;
input n159;
input n73;
input n173;
input n62;
input n4400;
input n228;
input n87;
input n23;
input n193;
input n130;
input n38;
input n4410;
input n127;
input n2204;
input n219;
input n4432;
input n179;
input n227;
input n118;
input n1469;
input n4528;
input n238;
input n161;
input n201;
input n88;
input n54;
input n237;
input n169;
input n2218;
input n75;
input n64;
input n60;
input n82;
input n3743;
input n1480;
input n189;
input n1197;
input n171;
input n134;
input n221;
input n230;
input n175;
input n212;
input n4427;
input n112;
input n167;
input n35;
input n166;
input n135;
input n154;
input n164;
input n85;
input n4415;
input n222;
input n1462;
input n185;
input n203;
input n152;
input n170;
input n199;
input n2256;
input n181;
input n187;
input n214;
input n3698;
input n100;
input n211;
input n3737;
input n1496;
input n115;
input n207;
input n1459;
input n217;
input n168;
input n26;
input n195;
input n209;
input n163;
input n198;
input n2253;
input n183;
input n182;
input n215;
input n218;
input n3701;
input n86;
input n59;
input n5;
input n4393;
input n165;
input n110;
input n158;
input n1455;
input n121;
input n84;
input n58;
input n15;
input n144;
input n79;
input n41;
input n3705;
input n229;
input n138;
input n66;
input n56;
input n192;
input n194;
input n186;
input n77;
input n3717;
input n106;
input n235;
input n204;
input n70;
input n224;
input n233;
input n156;
input n174;
input n225;
input n44;
input n236;
input n200;

// Start POs
output n408;
output n399;
output n278;
output n2;
output n370;
output n350;
output n319;
output n522;
output n307;
output n368;
output n556;
output n406;
output n471;
output n436;
output n540;
output n412;
output n304;
output n292;
output n532;
output n528;
output n480;
output n422;
output n404;
output n432;
output n444;
output n333;
output n488;
output n391;
output n276;
output n558;
output n486;
output n258;
output n560;
output n362;
output n281;
output n546;
output n330;
output n448;
output n289;
output n341;
output n324;
output n554;
output n526;
output n264;
output n496;
output n442;
output n410;
output n524;
output n416;
output n538;
output n3;
output n552;
output n469;
output n382;
output n492;
output n414;
output n246;
output n286;
output n295;
output n394;
output n536;
output n249;
output n327;
output n365;
output n453;
output n313;
output n279;
output n379;
output n548;
output n298;
output n356;
output n373;
output n252;
output n446;
output n321;
output n438;
output n284;
output n530;
output n450;
output n550;
output n359;
output n336;
output n534;
output n301;
output n344;
output n397;
output n338;
output n418;
output n490;
output n542;
output n440;
output n388;
output n484;
output n270;
output n385;
output n482;
output n478;
output n347;
output n544;
output n316;
output n310;
output n402;
output n494;
output n419;
output n273;
output n353;
output n376;

// Start wires
wire n408;
wire n319;
wire net_796;
wire net_416;
wire net_215;
wire net_933;
wire net_54;
wire net_526;
wire net_943;
wire n436;
wire net_834;
wire net_429;
wire net_694;
wire net_129;
wire net_648;
wire net_373;
wire net_98;
wire net_739;
wire net_980;
wire net_151;
wire net_356;
wire net_53;
wire net_452;
wire n63;
wire net_974;
wire net_545;
wire net_284;
wire net_560;
wire net_774;
wire net_923;
wire net_826;
wire net_439;
wire net_259;
wire net_548;
wire n333;
wire net_501;
wire n560;
wire n2230;
wire net_187;
wire net_111;
wire net_264;
wire net_225;
wire n150;
wire net_636;
wire n78;
wire net_263;
wire net_252;
wire net_124;
wire net_343;
wire net_160;
wire n141;
wire net_832;
wire net_322;
wire net_511;
wire n3723;
wire net_815;
wire net_901;
wire net_420;
wire net_665;
wire net_447;
wire net_871;
wire net_410;
wire net_508;
wire net_390;
wire n536;
wire net_35;
wire n365;
wire net_586;
wire n453;
wire n313;
wire net_703;
wire net_239;
wire net_193;
wire net_310;
wire n1486;
wire net_120;
wire net_292;
wire net_201;
wire net_109;
wire net_80;
wire n234;
wire n206;
wire net_96;
wire net_167;
wire net_651;
wire net_682;
wire net_989;
wire net_280;
wire net_744;
wire n159;
wire net_495;
wire net_34;
wire net_458;
wire net_108;
wire net_598;
wire net_685;
wire n478;
wire n87;
wire n130;
wire net_789;
wire n38;
wire net_971;
wire n4410;
wire n310;
wire net_593;
wire net_617;
wire net_672;
wire net_777;
wire net_1007;
wire net_554;
wire net_490;
wire net_742;
wire net_1014;
wire net_46;
wire n60;
wire net_584;
wire net_969;
wire n175;
wire net_632;
wire net_538;
wire net_165;
wire net_883;
wire net_843;
wire net_821;
wire net_464;
wire net_366;
wire net_13;
wire n448;
wire net_747;
wire net_446;
wire n554;
wire n1462;
wire n410;
wire n170;
wire n2256;
wire net_248;
wire net_384;
wire n3;
wire net_964;
wire n1496;
wire net_198;
wire n26;
wire n195;
wire net_209;
wire net_3;
wire n163;
wire net_634;
wire net_294;
wire net_802;
wire net_371;
wire n110;
wire n58;
wire n15;
wire net_1004;
wire net_848;
wire net_485;
wire net_997;
wire n194;
wire net_1031;
wire n336;
wire net_503;
wire net_256;
wire net_850;
wire n3717;
wire net_82;
wire net_64;
wire net_996;
wire net_726;
wire net_679;
wire net_1028;
wire net_308;
wire net_75;
wire n347;
wire net_959;
wire net_515;
wire net_600;
wire net_757;
wire net_701;
wire net_206;
wire net_125;
wire net_397;
wire net_808;
wire net_223;
wire net_1009;
wire net_715;
wire net_235;
wire net_890;
wire net_606;
wire net_623;
wire n188;
wire net_663;
wire net_320;
wire net_579;
wire net_250;
wire net_769;
wire n65;
wire net_312;
wire net_986;
wire net_130;
wire net_572;
wire n208;
wire n231;
wire net_286;
wire net_147;
wire net_787;
wire net_481;
wire net_369;
wire n486;
wire net_403;
wire net_32;
wire net_1025;
wire n80;
wire n330;
wire net_935;
wire net_282;
wire net_645;
wire net_426;
wire net_780;
wire net_841;
wire net_609;
wire net_541;
wire net_414;
wire n2224;
wire n83;
wire net_794;
wire n2247;
wire net_799;
wire net_528;
wire n197;
wire n69;
wire net_1012;
wire net_456;
wire net_155;
wire net_705;
wire net_335;
wire net_907;
wire net_506;
wire net_181;
wire n76;
wire net_349;
wire net_39;
wire net_1036;
wire net_245;
wire n446;
wire net_395;
wire net_331;
wire n530;
wire net_493;
wire n2236;
wire net_816;
wire net_386;
wire net_987;
wire net_641;
wire net_277;
wire n50;
wire n344;
wire net_919;
wire n418;
wire net_89;
wire n4437;
wire net_290;
wire net_680;
wire n23;
wire net_931;
wire net_338;
wire net_1039;
wire net_721;
wire net_243;
wire net_400;
wire n399;
wire n179;
wire net_759;
wire net_1018;
wire net_602;
wire net_175;
wire net_657;
wire n2218;
wire net_823;
wire net_106;
wire net_140;
wire net_740;
wire net_247;
wire n1480;
wire net_329;
wire net_279;
wire net_698;
wire net_897;
wire net_25;
wire net_70;
wire net_691;
wire n112;
wire net_194;
wire net_962;
wire net_730;
wire net_615;
wire net_478;
wire net_441;
wire net_596;
wire net_138;
wire net_749;
wire net_1019;
wire net_804;
wire net_333;
wire net_639;
wire net_728;
wire n289;
wire n324;
wire net_957;
wire net_1006;
wire net_719;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_77;
wire net_20;
wire n214;
wire n181;
wire net_878;
wire net_1033;
wire net_49;
wire net_518;
wire net_861;
wire net_15;
wire net_57;
wire net_71;
wire net_771;
wire net_929;
wire n3701;
wire net_1;
wire net_708;
wire n5;
wire net_696;
wire n165;
wire net_537;
wire net_180;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire net_432;
wire net_513;
wire net_204;
wire net_232;
wire n338;
wire net_604;
wire net_163;
wire net_967;
wire n542;
wire net_67;
wire n224;
wire net_268;
wire n174;
wire net_459;
wire net_483;
wire net_48;
wire net_8;
wire net_737;
wire net_203;
wire net_505;
wire net_176;
wire net_296;
wire net_137;
wire net_992;
wire net_613;
wire net_237;
wire n172;
wire n94;
wire net_782;
wire n53;
wire net_614;
wire net_532;
wire net_93;
wire net_578;
wire n220;
wire net_786;
wire net_302;
wire net_889;
wire n184;
wire net_127;
wire net_984;
wire net_348;
wire net_753;
wire n1;
wire net_626;
wire net_101;
wire net_906;
wire net_388;
wire net_326;
wire net_707;
wire net_589;
wire net_100;
wire net_655;
wire n526;
wire net_686;
wire net_652;
wire net_536;
wire net_455;
wire net_221;
wire net_115;
wire net_689;
wire net_751;
wire net_393;
wire net_442;
wire net_830;
wire net_542;
wire n216;
wire n246;
wire net_575;
wire net_877;
wire net_595;
wire net_378;
wire n223;
wire net_408;
wire net_724;
wire net_1026;
wire net_423;
wire n190;
wire net_328;
wire net_157;
wire net_42;
wire n2211;
wire n191;
wire net_874;
wire net_66;
wire net_466;
wire net_868;
wire net_765;
wire n359;
wire net_675;
wire net_818;
wire net_938;
wire net_443;
wire net_922;
wire net_522;
wire net_270;
wire n385;
wire net_183;
wire net_668;
wire net_150;
wire net_304;
wire net_1011;
wire n278;
wire net_811;
wire net_352;
wire n1469;
wire n350;
wire net_800;
wire n238;
wire net_977;
wire net_644;
wire n307;
wire net_30;
wire net_643;
wire net_852;
wire net_436;
wire n540;
wire net_24;
wire net_622;
wire n304;
wire net_186;
wire net_812;
wire n1197;
wire n167;
wire net_792;
wire n432;
wire net_1000;
wire n488;
wire net_1035;
wire net_1016;
wire net_767;
wire n85;
wire net_825;
wire net_219;
wire net_18;
wire net_309;
wire net_659;
wire net_131;
wire net_196;
wire net_913;
wire net_29;
wire net_358;
wire n203;
wire net_837;
wire n152;
wire net_899;
wire net_1010;
wire net_516;
wire net_31;
wire net_927;
wire n115;
wire n3737;
wire net_956;
wire n1459;
wire net_713;
wire n2253;
wire net_693;
wire net_360;
wire net_213;
wire net_729;
wire n4393;
wire net_863;
wire net_260;
wire net_947;
wire net_438;
wire n321;
wire n284;
wire net_732;
wire net_580;
wire n450;
wire n229;
wire net_314;
wire net_904;
wire net_341;
wire net_952;
wire n397;
wire net_468;
wire net_58;
wire n484;
wire net_970;
wire net_798;
wire net_488;
wire n44;
wire net_73;
wire net_807;
wire net_86;
wire net_945;
wire net_179;
wire net_159;
wire net_61;
wire net_449;
wire net_383;
wire n133;
wire n471;
wire net_62;
wire n178;
wire net_6;
wire net_553;
wire net_534;
wire net_217;
wire n55;
wire net_733;
wire net_887;
wire net_903;
wire n213;
wire net_763;
wire net_427;
wire net_486;
wire net_135;
wire net_915;
wire net_473;
wire net_406;
wire n422;
wire net_633;
wire net_324;
wire net_113;
wire net_710;
wire net_497;
wire n546;
wire net_454;
wire net_462;
wire net_418;
wire net_40;
wire net_872;
wire n264;
wire net_709;
wire n109;
wire net_161;
wire n442;
wire n2239;
wire net_300;
wire n538;
wire net_748;
wire net_677;
wire net_95;
wire n103;
wire net_173;
wire net_78;
wire net_990;
wire net_950;
wire net_1003;
wire net_514;
wire net_376;
wire net_22;
wire net_354;
wire net_524;
wire net_646;
wire net_363;
wire net_445;
wire net_573;
wire n205;
wire net_776;
wire net_866;
wire net_44;
wire net_784;
wire net_520;
wire net_422;
wire n301;
wire net_1032;
wire net_561;
wire net_567;
wire n2208;
wire net_45;
wire net_381;
wire net_591;
wire net_746;
wire n62;
wire net_981;
wire n4400;
wire net_272;
wire n193;
wire net_178;
wire net_845;
wire n127;
wire net_1024;
wire n219;
wire n544;
wire net_762;
wire n227;
wire net_695;
wire net_839;
wire net_814;
wire n88;
wire net_556;
wire net_941;
wire n169;
wire net_893;
wire net_809;
wire net_629;
wire net_55;
wire net_559;
wire net_635;
wire net_255;
wire net_266;
wire net_1037;
wire net_345;
wire net_859;
wire net_620;
wire net_619;
wire net_350;
wire net_398;
wire net_306;
wire net_954;
wire n528;
wire n444;
wire net_500;
wire n276;
wire n154;
wire n164;
wire net_631;
wire net_11;
wire net_123;
wire net_994;
wire net_527;
wire net_362;
wire net_262;
wire net_318;
wire net_68;
wire n211;
wire n469;
wire net_976;
wire n394;
wire net_316;
wire net_865;
wire net_84;
wire net_670;
wire net_611;
wire net_231;
wire n379;
wire net_103;
wire net_226;
wire net_1021;
wire net_228;
wire n252;
wire net_926;
wire n41;
wire n3705;
wire net_966;
wire net_143;
wire n56;
wire net_190;
wire net_391;
wire net_1002;
wire net_533;
wire net_145;
wire net_911;
wire net_37;
wire n233;
wire n156;
wire net_582;
wire net_188;
wire net_755;
wire net_509;
wire n482;
wire net_661;
wire net_881;
wire net_211;
wire net_133;
wire net_568;
wire n2;
wire net_47;
wire net_1008;
wire n522;
wire n556;
wire n61;
wire net_557;
wire net_119;
wire net_210;
wire net_168;
wire net_916;
wire n532;
wire net_741;
wire net_477;
wire net_940;
wire n404;
wire net_385;
wire net_851;
wire net_269;
wire net_469;
wire n160;
wire net_847;
wire net_727;
wire net_90;
wire net_671;
wire net_283;
wire net_85;
wire net_778;
wire net_770;
wire n176;
wire net_404;
wire net_1005;
wire n180;
wire net_240;
wire n124;
wire net_4;
wire net_895;
wire net_295;
wire n196;
wire n81;
wire n32;
wire n4420;
wire net_307;
wire net_344;
wire net_16;
wire n279;
wire net_884;
wire net_712;
wire net_257;
wire n57;
wire net_233;
wire net_474;
wire net_472;
wire net_958;
wire net_65;
wire n550;
wire net_995;
wire net_896;
wire net_484;
wire net_136;
wire net_207;
wire net_944;
wire net_700;
wire net_961;
wire net_126;
wire n173;
wire n73;
wire net_278;
wire net_571;
wire net_63;
wire n494;
wire n4432;
wire net_274;
wire net_601;
wire n118;
wire net_321;
wire net_425;
wire n4528;
wire net_287;
wire net_189;
wire net_930;
wire net_833;
wire net_829;
wire net_720;
wire net_99;
wire n64;
wire net_480;
wire net_216;
wire net_934;
wire net_433;
wire net_836;
wire net_900;
wire net_717;
wire n4427;
wire net_544;
wire net_368;
wire n480;
wire net_224;
wire net_684;
wire net_52;
wire n166;
wire net_608;
wire n258;
wire net_370;
wire net_510;
wire net_413;
wire net_1020;
wire net_716;
wire net_114;
wire net_973;
wire net_1034;
wire net_860;
wire net_36;
wire net_870;
wire n207;
wire net_253;
wire net_637;
wire net_276;
wire net_311;
wire net_760;
wire net_494;
wire net_547;
wire net_873;
wire net_154;
wire net_666;
wire n86;
wire net_507;
wire net_616;
wire n158;
wire net_238;
wire net_817;
wire net_28;
wire net_529;
wire net_704;
wire n79;
wire net_587;
wire net_97;
wire n186;
wire net_192;
wire net_793;
wire net_649;
wire net_460;
wire n204;
wire n235;
wire net_650;
wire net_291;
wire net_457;
wire net_735;
wire net_772;
wire net_857;
wire net_867;
wire net_121;
wire net_200;
wire net_597;
wire net_743;
wire n200;
wire net_396;
wire n316;
wire net_195;
wire net_107;
wire net_166;
wire net_530;
wire n406;
wire net_849;
wire net_594;
wire net_603;
wire net_23;
wire net_271;
wire net_117;
wire net_74;
wire net_673;
wire net_401;
wire net_642;
wire net_205;
wire net_699;
wire net_242;
wire net_359;
wire net_440;
wire n162;
wire net_758;
wire net_26;
wire net_470;
wire net_920;
wire net_334;
wire net_430;
wire net_882;
wire net_718;
wire net_365;
wire net_820;
wire net_380;
wire n496;
wire net_141;
wire n3711;
wire net_467;
wire n524;
wire net_83;
wire net_879;
wire n416;
wire net_372;
wire net_437;
wire n295;
wire net_56;
wire n249;
wire net_566;
wire net_968;
wire n4405;
wire net_336;
wire net_803;
wire n240;
wire net_624;
wire net_555;
wire net_2;
wire net_9;
wire n111;
wire n438;
wire n151;
wire n12;
wire net_298;
wire net_790;
wire net_688;
wire net_697;
wire net_998;
wire net_475;
wire net_563;
wire net_605;
wire net_199;
wire net_502;
wire net_431;
wire net_835;
wire net_924;
wire net_898;
wire net_638;
wire net_909;
wire n370;
wire net_222;
wire net_932;
wire net_152;
wire net_313;
wire n368;
wire net_489;
wire net_714;
wire n237;
wire n75;
wire net_683;
wire net_258;
wire net_607;
wire net_148;
wire net_419;
wire net_251;
wire net_972;
wire net_244;
wire net_664;
wire net_936;
wire net_128;
wire net_585;
wire net_840;
wire net_819;
wire n362;
wire net_827;
wire net_549;
wire net_785;
wire net_374;
wire net_411;
wire net_854;
wire net_788;
wire net_214;
wire n187;
wire net_249;
wire n100;
wire n552;
wire n382;
wire net_979;
wire n168;
wire net_706;
wire n209;
wire net_156;
wire net_1013;
wire net_842;
wire net_810;
wire net_92;
wire net_112;
wire net_394;
wire n59;
wire net_139;
wire net_551;
wire n1455;
wire net_332;
wire net_409;
wire n84;
wire n138;
wire net_463;
wire net_492;
wire net_656;
wire net_88;
wire n77;
wire net_197;
wire net_766;
wire n106;
wire net_81;
wire n388;
wire n440;
wire net_402;
wire net_202;
wire n270;
wire n225;
wire net_110;
wire net_722;
wire net_379;
wire net_33;
wire net_988;
wire net_918;
wire net_949;
wire net_289;
wire net_450;
wire net_621;
wire net_435;
wire net_132;
wire n18;
wire net_105;
wire net_12;
wire net_978;
wire n239;
wire n113;
wire net_569;
wire net_768;
wire net_1017;
wire net_955;
wire n74;
wire net_327;
wire net_357;
wire n391;
wire net_960;
wire net_630;
wire net_999;
wire net_76;
wire net_1029;
wire net_908;
wire n4394;
wire net_353;
wire net_822;
wire net_801;
wire net_519;
wire net_412;
wire net_838;
wire n153;
wire n3729;
wire net_17;
wire net_319;
wire net_453;
wire n286;
wire net_581;
wire net_164;
wire n155;
wire net_731;
wire net_377;
wire net_87;
wire net_0;
wire net_288;
wire net_1038;
wire net_912;
wire n202;
wire net_658;
wire net_805;
wire net_734;
wire n4526;
wire net_540;
wire net_512;
wire net_779;
wire n1492;
wire net_662;
wire net_862;
wire net_951;
wire net_891;
wire net_50;
wire net_806;
wire n97;
wire net_234;
wire net_38;
wire n177;
wire n147;
wire net_342;
wire n47;
wire net_975;
wire net_612;
wire net_19;
wire n490;
wire net_738;
wire net_946;
wire net_892;
wire net_504;
wire net_855;
wire n228;
wire net_674;
wire net_618;
wire n2204;
wire net_303;
wire n273;
wire n161;
wire net_491;
wire net_965;
wire net_681;
wire net_948;
wire net_783;
wire net_392;
wire net_118;
wire n82;
wire n3743;
wire net_754;
wire n189;
wire net_421;
wire net_146;
wire n171;
wire net_921;
wire net_764;
wire net_550;
wire net_876;
wire net_122;
wire net_417;
wire n230;
wire net_7;
wire n35;
wire net_172;
wire n281;
wire net_428;
wire net_94;
wire net_246;
wire net_461;
wire net_640;
wire net_482;
wire n222;
wire net_991;
wire net_905;
wire net_775;
wire net_149;
wire net_142;
wire net_752;
wire n199;
wire net_387;
wire net_654;
wire net_858;
wire net_330;
wire net_888;
wire net_498;
wire net_535;
wire net_158;
wire n414;
wire net_676;
wire net_41;
wire n327;
wire n198;
wire net_577;
wire n183;
wire net_570;
wire n182;
wire n215;
wire net_444;
wire net_525;
wire net_1023;
wire net_844;
wire n548;
wire net_325;
wire net_797;
wire n356;
wire net_301;
wire n121;
wire net_299;
wire n144;
wire net_985;
wire n66;
wire net_182;
wire net_60;
wire net_521;
wire net_337;
wire net_590;
wire net_267;
wire net_273;
wire net_424;
wire net_576;
wire net_690;
wire net_465;
wire n236;
wire net_177;
wire net_523;
wire net_407;
wire net_476;
wire net_564;
wire n376;
wire net_382;
wire net_725;
wire net_583;
wire net_813;
wire net_953;
wire net_351;
wire net_1027;
wire net_894;
wire net_340;
wire net_265;
wire net_517;
wire net_434;
wire net_628;
wire net_791;
wire net_939;
wire net_824;
wire net_14;
wire net_220;
wire n558;
wire net_293;
wire n3749;
wire net_942;
wire n226;
wire n210;
wire n341;
wire net_69;
wire net_543;
wire n114;
wire n89;
wire net_925;
wire net_625;
wire net_339;
wire net_993;
wire n492;
wire net_361;
wire net_864;
wire net_27;
wire n157;
wire net_317;
wire net_856;
wire net_305;
wire net_880;
wire net_191;
wire net_261;
wire net_558;
wire net_660;
wire net_144;
wire net_102;
wire net_227;
wire net_59;
wire n9;
wire net_162;
wire n29;
wire net_1001;
wire net_781;
wire net_230;
wire net_910;
wire n232;
wire net_653;
wire n534;
wire net_134;
wire net_1022;
wire net_678;
wire net_546;
wire net_185;
wire net_702;
wire net_588;
wire net_928;
wire net_667;
wire net_853;
wire n402;
wire net_208;
wire net_236;
wire net_1015;
wire net_212;
wire net_315;
wire net_487;
wire net_552;
wire net_914;
wire net_415;
wire net_116;
wire n201;
wire n54;
wire net_347;
wire net_756;
wire net_91;
wire net_297;
wire net_346;
wire n412;
wire net_875;
wire net_104;
wire net_448;
wire n134;
wire net_72;
wire net_886;
wire n221;
wire n292;
wire net_229;
wire n212;
wire net_627;
wire net_917;
wire net_241;
wire net_687;
wire net_5;
wire net_405;
wire n135;
wire net_983;
wire net_355;
wire net_184;
wire net_711;
wire net_599;
wire net_610;
wire n4415;
wire net_723;
wire n185;
wire net_389;
wire net_831;
wire net_902;
wire net_451;
wire n3698;
wire net_323;
wire net_963;
wire net_846;
wire net_750;
wire net_736;
wire net_275;
wire net_399;
wire net_539;
wire n217;
wire net_692;
wire net_153;
wire net_218;
wire net_174;
wire n218;
wire net_375;
wire net_562;
wire n298;
wire net_364;
wire net_43;
wire n373;
wire net_10;
wire net_592;
wire net_21;
wire net_79;
wire net_647;
wire net_885;
wire net_1030;
wire n192;
wire net_773;
wire net_285;
wire net_281;
wire net_828;
wire net_869;
wire net_669;
wire net_937;
wire net_254;
wire n70;
wire net_761;
wire net_496;
wire net_479;
wire net_574;
wire net_795;
wire net_982;
wire n419;
wire net_745;
wire n353;

// Start cells
NAND2_X1 inst_696 ( .ZN(net_190), .A2(net_146), .A1(net_39) );
NOR2_X1 inst_481 ( .ZN(net_875), .A1(net_768), .A2(net_711) );
XNOR2_X1 inst_228 ( .ZN(net_844), .B(net_842), .A(net_781) );
XNOR2_X1 inst_125 ( .ZN(net_603), .A(net_333), .B(n2211) );
NOR2_X1 inst_486 ( .A2(net_856), .ZN(net_789), .A1(net_602) );
INV_X1 inst_1025 ( .ZN(net_491), .A(net_490) );
NAND2_X1 inst_707 ( .ZN(net_280), .A2(net_154), .A1(net_56) );
NAND2_X1 inst_779 ( .ZN(net_559), .A1(net_533), .A2(net_491) );
NOR2_X1 inst_395 ( .A1(net_164), .ZN(net_158), .A2(net_91) );
NAND2_X1 inst_841 ( .ZN(net_971), .A2(net_936), .A1(net_879) );
XNOR2_X1 inst_244 ( .ZN(net_943), .B(net_854), .A(net_514) );
NOR2_X1 inst_452 ( .A2(net_999), .ZN(net_502), .A1(net_501) );
NAND2_X1 inst_689 ( .ZN(net_265), .A2(net_131), .A1(net_77) );
NOR2_X1 inst_430 ( .ZN(net_433), .A2(net_179), .A1(n4427) );
XNOR2_X1 inst_214 ( .ZN(net_781), .B(net_733), .A(net_732) );
NAND4_X1 inst_548 ( .A4(net_741), .A1(net_706), .A2(net_705), .A3(net_704), .ZN(n412) );
NOR2_X1 inst_515 ( .ZN(net_1011), .A2(net_1007), .A1(net_729) );
NAND2_X1 inst_772 ( .ZN(net_544), .A2(net_422), .A1(net_386) );
NAND2_X1 inst_728 ( .ZN(net_167), .A2(net_132), .A1(net_33) );
INV_X1 inst_944 ( .ZN(net_15), .A(n3705) );
NAND2_X1 inst_642 ( .ZN(net_74), .A2(n238), .A1(n18) );
NOR2_X1 inst_459 ( .ZN(net_805), .A1(net_531), .A2(net_399) );
INV_X1 inst_1018 ( .ZN(net_720), .A(net_432) );
NOR2_X1 inst_445 ( .A2(net_1012), .ZN(net_615), .A1(net_498) );
NAND2_X1 inst_850 ( .ZN(net_988), .A2(net_970), .A1(net_776) );
NAND2_X1 inst_709 ( .ZN(net_157), .A1(net_156), .A2(net_93) );
XNOR2_X1 inst_93 ( .A(net_266), .ZN(net_227), .B(net_114) );
NAND2_X1 inst_700 ( .ZN(net_271), .A2(net_140), .A1(net_48) );
INV_X2 inst_920 ( .A(net_373), .ZN(net_164) );
NAND2_X1 inst_606 ( .ZN(net_39), .A2(n198), .A1(n18) );
NOR2_X1 inst_367 ( .A1(net_191), .ZN(net_91), .A2(n170) );
INV_X1 inst_957 ( .ZN(net_26), .A(n82) );
INV_X1 inst_979 ( .A(net_331), .ZN(net_236) );
NAND2_X1 inst_853 ( .ZN(net_1003), .A2(net_985), .A1(net_766) );
INV_X1 inst_1008 ( .ZN(net_1025), .A(net_623) );
XNOR2_X1 inst_139 ( .ZN(net_422), .A(net_290), .B(n4437) );
NAND2_X1 inst_657 ( .A2(net_191), .ZN(net_145), .A1(n94) );
NAND3_X1 inst_559 ( .ZN(net_477), .A3(net_476), .A1(net_305), .A2(net_304) );
NAND3_X1 inst_584 ( .ZN(net_750), .A1(net_658), .A3(net_657), .A2(net_484) );
NAND4_X1 inst_521 ( .ZN(n404), .A4(n240), .A3(n228), .A2(n184), .A1(n150) );
NOR2_X1 inst_470 ( .A2(net_808), .ZN(net_708), .A1(net_677) );
NAND4_X1 inst_535 ( .A1(net_722), .ZN(net_674), .A3(net_592), .A4(net_591), .A2(net_389) );
NOR2_X1 inst_450 ( .A2(net_956), .A1(net_728), .ZN(net_496) );
NAND2_X1 inst_745 ( .ZN(net_506), .A2(net_352), .A1(net_108) );
NAND4_X1 inst_520 ( .ZN(n410), .A4(n199), .A3(n188), .A2(n172), .A1(n162) );
XNOR2_X1 inst_237 ( .ZN(net_874), .A(net_827), .B(net_774) );
XNOR2_X1 inst_148 ( .ZN(net_597), .A(net_406), .B(net_309) );
NAND4_X1 inst_554 ( .A3(net_986), .A4(net_935), .A1(net_891), .A2(net_836), .ZN(n270) );
XNOR2_X1 inst_191 ( .ZN(net_707), .B(net_636), .A(net_508) );
CLKBUF_X1 inst_1063 ( .Z(n530), .A(n4420) );
NAND2_X1 inst_813 ( .ZN(net_754), .A2(net_753), .A1(n4526) );
XOR2_X1 inst_51 ( .Z(net_344), .A(net_343), .B(net_342) );
OR2_X4 inst_315 ( .ZN(net_677), .A1(net_536), .A2(net_231) );
XOR2_X1 inst_80 ( .Z(net_780), .A(net_779), .B(net_778) );
NAND2_X1 inst_836 ( .ZN(net_962), .A1(net_907), .A2(net_899) );
CLKBUF_X1 inst_1066 ( .Z(n524), .A(n4437) );
INV_X1 inst_974 ( .A(net_333), .ZN(net_240) );
XNOR2_X1 inst_216 ( .ZN(net_788), .A(net_715), .B(net_241) );
CLKBUF_X1 inst_1059 ( .Z(n538), .A(n4400) );
XNOR2_X1 inst_241 ( .ZN(net_930), .A(net_884), .B(net_844) );
CLKBUF_X1 inst_1075 ( .Z(n482), .A(n2253) );
MUX2_X2 inst_862 ( .Z(net_214), .S(net_191), .A(net_8), .B(n62) );
AND2_X4 inst_1116 ( .ZN(net_561), .A1(net_480), .A2(net_467) );
XNOR2_X1 inst_151 ( .ZN(net_445), .A(net_330), .B(net_294) );
XOR2_X1 inst_64 ( .Z(net_377), .A(net_376), .B(net_375) );
INV_X1 inst_1001 ( .ZN(net_1016), .A(net_442) );
NAND2_X1 inst_743 ( .A2(net_293), .ZN(net_201), .A1(net_115) );
NOR2_X1 inst_415 ( .ZN(net_245), .A2(net_172), .A1(n4415) );
NAND2_X1 inst_828 ( .ZN(net_871), .A1(net_867), .A2(net_850) );
AND3_X4 inst_1104 ( .A3(net_608), .ZN(net_602), .A1(net_601), .A2(net_592) );
MUX2_X2 inst_892 ( .S(net_987), .Z(net_830), .A(net_829), .B(net_828) );
XNOR2_X1 inst_223 ( .ZN(net_837), .A(net_788), .B(net_661) );
AND2_X4 inst_1132 ( .ZN(net_550), .A2(net_549), .A1(net_432) );
NOR2_X1 inst_402 ( .ZN(net_351), .A1(net_164), .A2(net_104) );
INV_X1 inst_968 ( .A(net_262), .ZN(net_172) );
NAND2_X1 inst_819 ( .A2(net_987), .ZN(net_809), .A1(net_808) );
OR2_X2 inst_340 ( .A1(net_570), .ZN(net_541), .A2(net_540) );
NOR2_X1 inst_494 ( .A1(net_1020), .ZN(net_986), .A2(net_807) );
OR2_X4 inst_329 ( .ZN(net_685), .A1(net_628), .A2(net_538) );
INV_X1 inst_938 ( .ZN(net_115), .A(n3749) );
NAND3_X1 inst_574 ( .ZN(net_612), .A1(net_611), .A3(net_598), .A2(net_487) );
NOR2_X1 inst_386 ( .A2(net_162), .ZN(net_129), .A1(net_128) );
XNOR2_X1 inst_158 ( .A(net_485), .ZN(net_453), .B(net_452) );
XNOR2_X1 inst_141 ( .ZN(net_535), .B(net_392), .A(net_232) );
INV_X1 inst_936 ( .ZN(net_12), .A(n1496) );
NOR2_X1 inst_507 ( .ZN(net_917), .A2(net_916), .A1(net_747) );
NAND3_X1 inst_571 ( .ZN(net_649), .A3(net_578), .A1(net_519), .A2(net_467) );
MUX2_X2 inst_884 ( .S(net_191), .Z(net_119), .B(net_10), .A(n1459) );
NAND2_X1 inst_711 ( .ZN(net_328), .A2(net_126), .A1(net_54) );
NAND2_X1 inst_827 ( .ZN(net_890), .A1(net_867), .A2(net_834) );
NAND4_X1 inst_552 ( .ZN(net_921), .A1(net_920), .A2(net_895), .A4(net_813), .A3(net_767) );
NAND2_X1 inst_599 ( .ZN(net_373), .A2(n9), .A1(n12) );
INV_X1 inst_1033 ( .A(net_893), .ZN(net_675) );
NOR2_X1 inst_469 ( .ZN(net_692), .A1(net_590), .A2(net_516) );
XOR2_X1 inst_18 ( .Z(net_564), .A(net_259), .B(net_258) );
MUX2_X2 inst_915 ( .Z(net_1036), .B(net_1032), .A(net_1026), .S(n4526) );
NAND2_X1 inst_811 ( .A1(net_762), .ZN(net_755), .A2(net_735) );
NAND4_X1 inst_541 ( .ZN(net_699), .A1(net_579), .A2(net_562), .A4(net_481), .A3(net_194) );
XNOR2_X1 inst_208 ( .ZN(net_770), .B(net_680), .A(net_405) );
XOR2_X1 inst_9 ( .A(net_314), .Z(net_217), .B(net_216) );
XNOR2_X1 inst_113 ( .ZN(net_371), .A(net_157), .B(net_110) );
NOR2_X1 inst_505 ( .ZN(net_936), .A1(net_913), .A2(net_886) );
NOR3_X1 inst_356 ( .ZN(net_977), .A1(net_934), .A3(net_900), .A2(net_825) );
CLKBUF_X1 inst_1058 ( .Z(n540), .A(n4393) );
XNOR2_X1 inst_198 ( .ZN(net_738), .B(net_637), .A(net_509) );
INV_X1 inst_952 ( .ZN(net_22), .A(n1492) );
MUX2_X2 inst_897 ( .Z(net_866), .A(net_865), .B(net_864), .S(net_785) );
NAND2_X1 inst_784 ( .ZN(net_633), .A2(net_526), .A1(net_429) );
NAND2_X1 inst_721 ( .A1(net_191), .ZN(net_168), .A2(net_156) );
MUX2_X2 inst_902 ( .Z(net_949), .B(net_947), .A(net_946), .S(net_907) );
XNOR2_X1 inst_293 ( .B(net_1014), .A(net_1001), .ZN(n310) );
NAND2_X1 inst_778 ( .A1(net_751), .ZN(net_658), .A2(net_551) );
NAND2_X1 inst_636 ( .ZN(net_68), .A2(n206), .A1(n18) );
NAND2_X1 inst_632 ( .ZN(net_64), .A2(n189), .A1(n18) );
XOR2_X1 inst_0 ( .Z(net_381), .B(net_182), .A(n38) );
XNOR2_X1 inst_184 ( .ZN(net_795), .A(net_673), .B(net_659) );
NAND2_X1 inst_690 ( .ZN(net_320), .A2(net_139), .A1(net_60) );
NOR2_X1 inst_433 ( .ZN(net_569), .A2(net_418), .A1(net_366) );
NAND2_X1 inst_781 ( .ZN(net_731), .A2(net_627), .A1(net_524) );
NAND2_X1 inst_732 ( .A1(net_264), .A2(net_211), .ZN(net_192) );
XNOR2_X1 inst_98 ( .A(net_283), .B(net_280), .ZN(net_255) );
XNOR2_X1 inst_263 ( .B(net_962), .A(net_596), .ZN(n356) );
XNOR2_X1 inst_185 ( .ZN(net_701), .B(net_586), .A(net_395) );
INV_X1 inst_959 ( .ZN(net_80), .A(n5) );
XOR2_X1 inst_75 ( .Z(net_803), .A(net_720), .B(net_662) );
OR2_X4 inst_332 ( .ZN(net_824), .A1(net_756), .A2(net_755) );
XNOR2_X1 inst_166 ( .ZN(net_510), .B(net_370), .A(net_357) );
MUX2_X2 inst_868 ( .Z(net_285), .S(net_191), .A(net_112), .B(n75) );
XNOR2_X1 inst_163 ( .ZN(net_507), .B(net_324), .A(net_252) );
NOR2_X1 inst_394 ( .ZN(net_362), .A1(net_164), .A2(net_102) );
XOR2_X1 inst_79 ( .B(net_1025), .A(net_686), .Z(n391) );
XNOR2_X1 inst_106 ( .ZN(net_334), .A(net_333), .B(net_141) );
NOR2_X1 inst_422 ( .ZN(net_248), .A2(net_180), .A1(n2256) );
XNOR2_X1 inst_201 ( .ZN(net_741), .B(net_640), .A(net_445) );
INV_X1 inst_927 ( .ZN(net_4), .A(n3737) );
NAND2_X1 inst_605 ( .ZN(net_38), .A2(n226), .A1(n18) );
CLKBUF_X1 inst_1084 ( .Z(n440), .A(n1492) );
OR4_X1 inst_304 ( .ZN(net_851), .A2(n416), .A4(n414), .A3(n412), .A1(n404) );
NAND2_X1 inst_752 ( .ZN(net_244), .A2(net_240), .A1(n2211) );
INV_X1 inst_1027 ( .A(net_591), .ZN(net_537) );
XOR2_X1 inst_73 ( .Z(net_829), .A(net_536), .B(net_534) );
AND2_X4 inst_1143 ( .ZN(net_991), .A2(net_974), .A1(net_551) );
NOR2_X1 inst_378 ( .A1(net_191), .ZN(net_103), .A2(n167) );
MUX2_X2 inst_890 ( .Z(net_341), .S(net_191), .A(net_122), .B(n112) );
NOR2_X1 inst_361 ( .A1(net_191), .ZN(net_85), .A2(n169) );
INV_X1 inst_1024 ( .ZN(net_594), .A(net_522) );
INV_X1 inst_1016 ( .ZN(net_1004), .A(net_414) );
NAND2_X1 inst_659 ( .A2(net_191), .ZN(net_154), .A1(n29) );
XNOR2_X1 inst_250 ( .B(net_905), .A(net_898), .ZN(n344) );
NAND2_X1 inst_848 ( .ZN(net_985), .A2(net_958), .A1(net_743) );
NAND2_X1 inst_786 ( .ZN(net_660), .A2(net_659), .A1(net_540) );
NOR2_X1 inst_397 ( .ZN(net_358), .A1(net_164), .A2(net_100) );
NOR2_X1 inst_504 ( .ZN(net_906), .A2(net_896), .A1(net_764) );
CLKBUF_X1 inst_1048 ( .Z(n560), .A(n3698) );
NOR2_X1 inst_440 ( .A1(net_1027), .A2(net_963), .ZN(net_608) );
XOR2_X1 inst_2 ( .A(net_341), .Z(net_205), .B(net_204) );
NAND2_X1 inst_644 ( .ZN(net_76), .A2(n220), .A1(n18) );
MUX2_X2 inst_918 ( .Z(net_1039), .B(net_1034), .A(net_1030), .S(net_931) );
CLKBUF_X1 inst_1091 ( .A(n341), .Z(n286) );
NAND3_X1 inst_578 ( .ZN(net_729), .A1(net_620), .A3(net_619), .A2(net_506) );
MUX2_X2 inst_888 ( .Z(net_220), .S(net_191), .A(net_14), .B(n64) );
XOR2_X1 inst_52 ( .Z(net_347), .A(net_346), .B(net_345) );
NAND2_X1 inst_668 ( .A2(net_191), .ZN(net_147), .A1(n32) );
XNOR2_X1 inst_221 ( .ZN(net_826), .A(net_770), .B(net_672) );
NAND3_X1 inst_556 ( .A1(net_80), .ZN(n292), .A3(n134), .A2(n133) );
NAND2_X1 inst_650 ( .A2(net_191), .ZN(net_149), .A1(n103) );
XNOR2_X1 inst_289 ( .ZN(net_1024), .A(net_1012), .B(net_1002) );
INV_X1 inst_987 ( .A(net_277), .ZN(net_186) );
NOR2_X1 inst_432 ( .A1(net_406), .ZN(net_405), .A2(net_404) );
NAND2_X1 inst_679 ( .ZN(net_325), .A2(net_125), .A1(net_57) );
NOR2_X1 inst_420 ( .ZN(net_533), .A2(net_183), .A1(n2247) );
XNOR2_X1 inst_282 ( .ZN(net_1015), .A(net_1004), .B(net_998) );
NOR2_X1 inst_513 ( .ZN(net_994), .A2(net_991), .A1(net_750) );
NAND2_X1 inst_754 ( .ZN(net_460), .A2(net_242), .A1(n2239) );
XOR2_X1 inst_44 ( .Z(net_478), .B(net_320), .A(net_314) );
NOR2_X1 inst_371 ( .ZN(net_182), .A1(net_96), .A2(n2204) );
OR2_X4 inst_314 ( .A1(net_321), .A2(net_216), .ZN(net_196) );
NOR2_X1 inst_435 ( .A2(net_967), .ZN(net_427), .A1(net_426) );
NAND2_X1 inst_597 ( .ZN(net_31), .A2(n18), .A1(n160) );
NAND2_X1 inst_687 ( .ZN(net_323), .A2(net_140), .A1(net_62) );
NAND2_X1 inst_774 ( .ZN(net_668), .A2(net_597), .A1(net_415) );
NAND2_X1 inst_621 ( .ZN(net_124), .A1(n4528), .A2(n1492) );
NAND2_X1 inst_838 ( .A2(net_923), .ZN(net_922), .A1(net_678) );
INV_X1 inst_985 ( .ZN(net_392), .A(net_231) );
NAND2_X1 inst_628 ( .ZN(net_60), .A2(n18), .A1(n179) );
NAND2_X1 inst_815 ( .ZN(net_785), .A2(net_784), .A1(net_736) );
NOR2_X1 inst_472 ( .ZN(net_710), .A1(net_676), .A2(net_653) );
NOR2_X1 inst_447 ( .A1(net_1016), .ZN(net_617), .A2(net_503) );
NOR2_X1 inst_457 ( .ZN(net_709), .A1(net_524), .A2(net_490) );
MUX2_X2 inst_875 ( .Z(net_259), .S(net_191), .A(net_4), .B(n54) );
NAND2_X1 inst_665 ( .ZN(net_406), .A2(net_191), .A1(n3701) );
CLKBUF_X1 inst_1073 ( .Z(n486), .A(n2239) );
AND2_X4 inst_1117 ( .ZN(net_576), .A2(net_412), .A1(net_303) );
AND2_X4 inst_1130 ( .A1(net_603), .A2(net_551), .ZN(net_543) );
XNOR2_X1 inst_127 ( .ZN(net_462), .A(net_367), .B(n2247) );
MUX2_X2 inst_855 ( .S(net_191), .Z(net_107), .A(net_22), .B(n1455) );
NOR2_X1 inst_413 ( .ZN(net_751), .A2(net_240), .A1(n2211) );
XNOR2_X1 inst_146 ( .ZN(net_397), .B(net_229), .A(net_205) );
OR2_X4 inst_334 ( .ZN(net_894), .A2(net_833), .A1(net_757) );
MUX2_X2 inst_859 ( .Z(net_284), .S(net_191), .A(net_109), .B(n76) );
XNOR2_X1 inst_187 ( .ZN(net_703), .B(net_588), .A(net_230) );
XNOR2_X1 inst_206 ( .ZN(net_769), .A(net_683), .B(net_243) );
NAND2_X1 inst_805 ( .ZN(net_889), .A1(net_709), .A2(net_648) );
XNOR2_X1 inst_122 ( .ZN(net_463), .A(net_346), .B(n2253) );
XOR2_X1 inst_25 ( .Z(net_276), .A(net_275), .B(net_274) );
NOR3_X1 inst_354 ( .ZN(net_716), .A1(net_550), .A3(net_434), .A2(net_401) );
NOR2_X1 inst_405 ( .ZN(net_200), .A1(net_164), .A2(net_106) );
AND2_X4 inst_1145 ( .ZN(net_1008), .A2(net_1007), .A1(net_696) );
NOR2_X1 inst_492 ( .ZN(net_825), .A1(net_824), .A2(net_823) );
INV_X1 inst_1042 ( .ZN(net_822), .A(net_821) );
NAND2_X1 inst_817 ( .ZN(net_786), .A2(net_782), .A1(net_719) );
OR2_X4 inst_326 ( .ZN(net_526), .A2(net_525), .A1(net_483) );
NAND4_X1 inst_518 ( .ZN(n408), .A4(n186), .A3(n185), .A1(n183), .A2(n182) );
XOR2_X1 inst_69 ( .Z(net_799), .B(net_596), .A(net_485) );
NOR2_X1 inst_373 ( .A1(net_191), .ZN(net_98), .A2(n212) );
XOR2_X1 inst_82 ( .Z(net_804), .A(net_803), .B(net_802) );
XNOR2_X1 inst_108 ( .ZN(net_418), .A(net_358), .B(net_354) );
NAND2_X1 inst_844 ( .ZN(net_997), .A1(net_950), .A2(net_922) );
NAND3_X1 inst_595 ( .ZN(net_953), .A1(net_951), .A3(net_930), .A2(net_819) );
XOR2_X1 inst_22 ( .Z(net_268), .A(net_267), .B(net_266) );
AND2_X4 inst_1121 ( .A2(net_469), .ZN(net_421), .A1(net_295) );
AND3_X4 inst_1102 ( .ZN(net_679), .A3(net_611), .A2(net_598), .A1(net_597) );
NOR2_X1 inst_460 ( .ZN(net_532), .A2(net_441), .A1(net_248) );
INV_X1 inst_970 ( .A(net_318), .ZN(net_174) );
OR3_X4 inst_307 ( .A2(net_720), .A3(net_596), .ZN(net_520), .A1(net_485) );
NAND2_X1 inst_767 ( .ZN(net_655), .A2(net_592), .A1(net_556) );
NAND2_X1 inst_638 ( .ZN(net_70), .A2(n194), .A1(n18) );
XNOR2_X1 inst_161 ( .ZN(net_457), .A(net_337), .B(net_260) );
NAND3_X1 inst_560 ( .ZN(net_479), .A3(net_471), .A1(net_363), .A2(net_362) );
NAND2_X1 inst_749 ( .ZN(net_241), .A2(net_236), .A1(n4394) );
NAND3_X1 inst_586 ( .ZN(net_840), .A1(net_697), .A3(net_557), .A2(net_504) );
NAND2_X1 inst_702 ( .ZN(net_267), .A2(net_150), .A1(net_53) );
XOR2_X1 inst_16 ( .Z(net_252), .A(net_190), .B(net_167) );
NAND2_X1 inst_717 ( .ZN(net_264), .A2(net_143), .A1(net_58) );
XNOR2_X1 inst_276 ( .ZN(net_1002), .A(net_1001), .B(net_966) );
INV_X1 inst_1030 ( .ZN(net_650), .A(net_649) );
NAND2_X1 inst_718 ( .ZN(net_283), .A2(net_155), .A1(net_68) );
INV_X1 inst_1029 ( .ZN(net_648), .A(net_647) );
XNOR2_X1 inst_156 ( .ZN(net_450), .B(net_374), .A(net_350) );
INV_X1 inst_950 ( .ZN(net_20), .A(n69) );
CLKBUF_X1 inst_1068 ( .Z(n496), .A(n2208) );
MUX2_X2 inst_886 ( .Z(net_378), .S(net_191), .A(net_23), .B(n79) );
NAND2_X1 inst_802 ( .ZN(net_694), .A1(net_625), .A2(net_618) );
XNOR2_X1 inst_296 ( .ZN(net_1034), .B(net_1029), .A(net_1024) );
XNOR2_X1 inst_91 ( .A(net_315), .ZN(net_221), .B(net_220) );
MUX2_X2 inst_905 ( .S(net_962), .B(net_858), .A(net_802), .Z(n347) );
XNOR2_X1 inst_132 ( .ZN(net_673), .A(net_292), .B(n3743) );
OR2_X2 inst_342 ( .A2(net_921), .A1(net_915), .ZN(n264) );
NAND4_X1 inst_526 ( .A2(net_578), .ZN(net_562), .A4(net_561), .A1(net_518), .A3(net_391) );
INV_X1 inst_1006 ( .A(net_911), .ZN(net_882) );
NOR2_X1 inst_463 ( .ZN(net_555), .A2(net_554), .A1(net_498) );
XNOR2_X1 inst_96 ( .ZN(net_253), .A(net_159), .B(net_134) );
XNOR2_X1 inst_101 ( .ZN(net_311), .A(net_310), .B(net_264) );
OR2_X4 inst_319 ( .A2(net_1029), .ZN(net_554), .A1(net_484) );
NOR2_X1 inst_400 ( .ZN(net_360), .A1(net_164), .A2(net_95) );
NAND2_X1 inst_614 ( .ZN(net_47), .A2(n187), .A1(n18) );
NAND2_X1 inst_649 ( .A2(net_191), .ZN(net_148), .A1(n66) );
NAND2_X1 inst_821 ( .A2(net_950), .ZN(net_821), .A1(net_647) );
XNOR2_X1 inst_261 ( .ZN(net_957), .A(net_956), .B(net_912) );
INV_X1 inst_1031 ( .ZN(net_652), .A(net_651) );
INV_X1 inst_980 ( .A(net_345), .ZN(net_180) );
NOR2_X1 inst_500 ( .A2(net_904), .ZN(net_886), .A1(net_768) );
INV_X1 inst_945 ( .ZN(net_16), .A(n1486) );
NOR2_X1 inst_510 ( .ZN(net_961), .A2(net_959), .A1(net_746) );
XNOR2_X1 inst_268 ( .A(net_999), .ZN(net_979), .B(net_940) );
NOR2_X1 inst_369 ( .A1(net_191), .ZN(net_94), .A2(n214) );
INV_X1 inst_995 ( .ZN(net_925), .A(net_415) );
NAND4_X1 inst_550 ( .ZN(net_869), .A4(net_817), .A1(net_584), .A3(net_479), .A2(net_473) );
NAND2_X1 inst_830 ( .ZN(net_878), .A2(net_877), .A1(net_710) );
NAND2_X1 inst_603 ( .ZN(net_36), .A2(n196), .A1(n18) );
OR2_X4 inst_327 ( .A1(net_728), .ZN(net_620), .A2(net_529) );
XOR2_X1 inst_85 ( .B(net_1027), .A(net_961), .Z(n362) );
XNOR2_X1 inst_291 ( .ZN(net_1028), .B(net_1027), .A(net_1010) );
CLKBUF_X1 inst_1060 ( .Z(n536), .A(n4405) );
XNOR2_X1 inst_266 ( .ZN(net_968), .A(net_967), .B(net_926) );
NAND2_X1 inst_776 ( .ZN(net_920), .A2(net_420), .A1(n38) );
MUX2_X2 inst_900 ( .Z(net_945), .B(net_943), .A(net_942), .S(net_761) );
MUX2_X2 inst_866 ( .Z(net_308), .S(net_191), .A(net_111), .B(n59) );
XOR2_X1 inst_77 ( .Z(net_794), .A(net_745), .B(net_713) );
XNOR2_X1 inst_171 ( .ZN(net_586), .B(net_394), .A(net_222) );
NAND3_X1 inst_558 ( .A3(net_567), .ZN(net_475), .A2(net_355), .A1(net_341) );
NAND3_X1 inst_594 ( .ZN(net_952), .A1(net_951), .A2(net_950), .A3(net_928) );
XNOR2_X1 inst_145 ( .ZN(net_396), .B(net_227), .A(net_221) );
XNOR2_X1 inst_290 ( .ZN(net_1026), .B(net_1025), .A(net_1005) );
NOR2_X1 inst_374 ( .A1(net_191), .ZN(net_99), .A2(n173) );
XNOR2_X1 inst_272 ( .B(net_1012), .A(net_954), .ZN(n316) );
NOR2_X1 inst_502 ( .ZN(net_900), .A2(net_890), .A1(net_889) );
XNOR2_X1 inst_103 ( .ZN(net_319), .A(net_318), .B(net_317) );
NAND2_X1 inst_814 ( .ZN(net_767), .A1(net_766), .A2(net_742) );
XNOR2_X1 inst_248 ( .ZN(net_947), .B(net_860), .A(net_452) );
NOR2_X1 inst_389 ( .ZN(net_365), .A1(net_164), .A2(net_85) );
INV_X1 inst_925 ( .ZN(net_112), .A(n3717) );
NAND2_X1 inst_789 ( .A2(net_776), .ZN(net_664), .A1(net_522) );
NOR2_X1 inst_357 ( .A1(net_191), .ZN(net_81), .A2(n177) );
AND2_X4 inst_1120 ( .ZN(net_566), .A2(net_476), .A1(net_417) );
AND2_X4 inst_1141 ( .ZN(net_959), .A2(net_916), .A1(net_548) );
NAND2_X1 inst_809 ( .ZN(net_723), .A1(net_722), .A2(net_666) );
MUX2_X2 inst_881 ( .Z(net_314), .S(net_191), .A(net_117), .B(n84) );
INV_X1 inst_932 ( .ZN(net_8), .A(n4437) );
NAND2_X1 inst_822 ( .ZN(net_816), .A2(net_812), .A1(n89) );
MUX2_X2 inst_913 ( .A(net_1020), .B(net_1019), .S(net_993), .Z(n276) );
XNOR2_X1 inst_180 ( .ZN(net_640), .B(net_444), .A(net_276) );
AND2_X4 inst_1125 ( .A2(net_673), .ZN(net_436), .A1(net_435) );
INV_X1 inst_947 ( .ZN(net_18), .A(n2256) );
MUX2_X2 inst_912 ( .S(net_1018), .A(net_535), .B(net_534), .Z(n469) );
NAND2_X1 inst_731 ( .ZN(net_390), .A1(net_191), .A2(net_190) );
NAND2_X1 inst_609 ( .ZN(net_42), .A2(n217), .A1(n18) );
INV_X1 inst_1022 ( .A(net_630), .ZN(net_487) );
NAND2_X1 inst_795 ( .A2(net_684), .ZN(net_680), .A1(net_539) );
XNOR2_X1 inst_301 ( .B(net_1038), .A(net_984), .ZN(n370) );
NOR2_X1 inst_363 ( .A1(net_191), .ZN(net_87), .A2(n153) );
XOR2_X1 inst_27 ( .Z(net_518), .A(net_281), .B(net_280) );
XNOR2_X1 inst_247 ( .ZN(net_946), .B(net_859), .A(net_454) );
NOR2_X1 inst_403 ( .ZN(net_349), .A1(net_164), .A2(net_92) );
XNOR2_X1 inst_302 ( .A(net_1039), .B(net_981), .ZN(n321) );
OR2_X4 inst_322 ( .A2(net_1027), .ZN(net_552), .A1(net_497) );
NAND2_X1 inst_673 ( .A2(net_191), .ZN(net_151), .A1(n138) );
XNOR2_X1 inst_211 ( .ZN(net_858), .B(net_749), .A(net_717) );
NAND2_X1 inst_619 ( .ZN(net_52), .A2(n190), .A1(n18) );
NAND2_X1 inst_681 ( .ZN(net_258), .A2(net_127), .A1(net_40) );
NAND3_X1 inst_561 ( .ZN(net_481), .A3(net_480), .A2(net_323), .A1(net_285) );
NOR2_X1 inst_412 ( .ZN(net_452), .A2(net_239), .A1(n4420) );
NOR2_X1 inst_449 ( .A2(net_963), .ZN(net_495), .A1(net_383) );
NAND2_X1 inst_639 ( .ZN(net_71), .A2(n201), .A1(n18) );
MUX2_X2 inst_877 ( .Z(net_209), .S(net_191), .A(net_115), .B(n56) );
XNOR2_X1 inst_155 ( .ZN(net_449), .A(net_369), .B(net_347) );
NOR2_X1 inst_464 ( .ZN(net_659), .A2(net_546), .A1(net_435) );
MUX2_X2 inst_871 ( .Z(net_300), .S(net_191), .A(net_113), .B(n81) );
OR2_X2 inst_341 ( .ZN(net_545), .A2(net_544), .A1(net_486) );
INV_X1 inst_962 ( .ZN(net_28), .A(n2211) );
XNOR2_X1 inst_196 ( .A(net_925), .B(net_631), .ZN(n397) );
NAND4_X1 inst_532 ( .ZN(net_580), .A1(net_576), .A4(net_564), .A3(net_376), .A2(net_375) );
XOR2_X1 inst_55 ( .Z(net_357), .A(net_356), .B(net_355) );
NAND2_X1 inst_641 ( .ZN(net_73), .A2(n18), .A1(n158) );
NOR2_X1 inst_498 ( .A1(net_892), .ZN(net_870), .A2(net_849) );
NAND2_X1 inst_684 ( .ZN(net_136), .A2(net_135), .A1(net_43) );
XNOR2_X1 inst_298 ( .B(net_1023), .A(net_989), .ZN(n327) );
AND2_X4 inst_1137 ( .ZN(net_686), .A1(net_685), .A2(net_684) );
XOR2_X1 inst_42 ( .Z(net_413), .A(net_308), .B(net_307) );
OR2_X4 inst_323 ( .A2(net_1031), .ZN(net_557), .A1(net_506) );
NAND3_X1 inst_588 ( .ZN(net_856), .A1(net_723), .A3(net_552), .A2(net_501) );
NOR3_X1 inst_350 ( .ZN(net_766), .A3(net_381), .A2(net_163), .A1(net_129) );
XNOR2_X1 inst_231 ( .ZN(net_855), .A(net_796), .B(net_791) );
AND2_X4 inst_1138 ( .ZN(net_700), .A2(net_646), .A1(net_198) );
AND2_X4 inst_1119 ( .A1(net_572), .A2(net_469), .ZN(net_416) );
INV_X1 inst_1038 ( .ZN(net_743), .A(net_742) );
NAND2_X1 inst_793 ( .A1(net_692), .ZN(net_672), .A2(net_668) );
NAND2_X1 inst_715 ( .ZN(net_379), .A2(net_125), .A1(net_55) );
NOR2_X1 inst_437 ( .ZN(net_546), .A2(net_511), .A1(net_483) );
INV_X1 inst_940 ( .ZN(net_14), .A(n2236) );
INV_X1 inst_1004 ( .ZN(net_733), .A(net_463) );
XNOR2_X1 inst_189 ( .ZN(net_705), .B(net_642), .A(net_449) );
XOR2_X1 inst_14 ( .A(net_373), .B(net_228), .Z(net_225) );
NOR2_X1 inst_475 ( .A1(net_1025), .ZN(net_687), .A2(net_685) );
XOR2_X1 inst_31 ( .B(net_304), .Z(net_287), .A(net_286) );
INV_X1 inst_1045 ( .A(net_898), .ZN(net_872) );
NAND4_X1 inst_528 ( .ZN(net_670), .A1(net_573), .A3(net_572), .A2(net_469), .A4(net_270) );
MUX2_X2 inst_865 ( .Z(net_204), .S(net_191), .A(net_16), .B(n88) );
XNOR2_X1 inst_252 ( .ZN(net_912), .A(net_911), .B(net_874) );
MUX2_X2 inst_903 ( .S(net_962), .B(net_455), .A(net_453), .Z(n353) );
XOR2_X1 inst_62 ( .Z(net_596), .B(net_325), .A(n4420) );
INV_X1 inst_956 ( .ZN(net_25), .A(n4415) );
XNOR2_X1 inst_251 ( .ZN(net_910), .B(net_880), .A(net_873) );
NOR3_X1 inst_352 ( .ZN(net_681), .A1(net_528), .A2(net_440), .A3(net_438) );
NAND3_X1 inst_575 ( .A2(net_747), .ZN(net_614), .A1(net_613), .A3(net_608) );
CLKBUF_X1 inst_1074 ( .Z(n484), .A(n2247) );
NAND2_X1 inst_846 ( .A2(net_971), .ZN(net_970), .A1(net_594) );
XNOR2_X1 inst_286 ( .B(net_1016), .A(net_988), .ZN(n333) );
MUX2_X2 inst_879 ( .Z(net_363), .S(net_191), .A(net_11), .B(n109) );
NOR2_X1 inst_484 ( .A2(net_840), .ZN(net_774), .A1(net_605) );
NAND2_X1 inst_627 ( .ZN(net_59), .A2(n232), .A1(n18) );
XOR2_X1 inst_32 ( .B(net_302), .Z(net_288), .A(net_265) );
NOR4_X1 inst_344 ( .A2(net_1025), .A3(net_1004), .A1(net_967), .ZN(net_735), .A4(net_668) );
NOR2_X1 inst_428 ( .ZN(net_435), .A2(net_184), .A1(n3737) );
INV_X1 inst_969 ( .A(net_351), .ZN(net_173) );
NAND2_X1 inst_629 ( .ZN(net_61), .A2(n229), .A1(n18) );
AND3_X4 inst_1100 ( .ZN(net_644), .A3(net_478), .A1(net_197), .A2(net_196) );
NOR2_X1 inst_407 ( .ZN(net_372), .A1(net_164), .A2(net_82) );
NAND2_X1 inst_791 ( .ZN(net_667), .A2(net_658), .A1(net_657) );
NAND2_X1 inst_623 ( .ZN(net_55), .A2(n192), .A1(n18) );
CLKBUF_X1 inst_1072 ( .Z(n488), .A(n2236) );
INV_X1 inst_1044 ( .ZN(net_983), .A(net_866) );
XNOR2_X1 inst_97 ( .ZN(net_254), .A(net_166), .B(net_130) );
NAND2_X1 inst_616 ( .ZN(net_49), .A2(n239), .A1(n18) );
MUX2_X2 inst_898 ( .Z(net_898), .A(net_865), .B(net_864), .S(net_852) );
NAND2_X1 inst_775 ( .ZN(net_628), .A2(net_597), .A1(n4526) );
NAND4_X1 inst_533 ( .A1(net_645), .ZN(net_582), .A4(net_478), .A3(net_321), .A2(net_216) );
NAND2_X1 inst_620 ( .ZN(net_53), .A2(n18), .A1(n171) );
AND3_X4 inst_1107 ( .ZN(net_607), .A3(net_606), .A2(net_603), .A1(net_437) );
NAND2_X1 inst_652 ( .A2(net_191), .ZN(net_156), .A1(n70) );
XNOR2_X1 inst_137 ( .ZN(net_432), .A(net_289), .B(n4432) );
NAND2_X1 inst_677 ( .ZN(net_121), .A2(net_120), .A1(n38) );
NOR2_X1 inst_425 ( .ZN(net_249), .A2(net_178), .A1(n1486) );
XNOR2_X1 inst_130 ( .ZN(net_389), .A(net_262), .B(n4415) );
NAND2_X1 inst_722 ( .ZN(net_282), .A2(net_149), .A1(net_72) );
XNOR2_X1 inst_227 ( .ZN(net_843), .B(net_842), .A(net_780) );
CLKBUF_X1 inst_1095 ( .A(n264), .Z(n258) );
NAND2_X1 inst_760 ( .ZN(net_538), .A1(net_415), .A2(net_414) );
NAND2_X1 inst_746 ( .ZN(net_309), .A2(net_224), .A1(net_191) );
XNOR2_X1 inst_176 ( .ZN(net_636), .B(net_451), .A(net_257) );
XOR2_X1 inst_58 ( .Z(net_471), .B(net_338), .A(net_202) );
XOR2_X1 inst_87 ( .B(net_1029), .A(net_994), .Z(n313) );
CLKBUF_X1 inst_1054 ( .Z(n548), .A(n3737) );
INV_X1 inst_972 ( .A(net_272), .ZN(net_175) );
INV_X1 inst_983 ( .A(net_367), .ZN(net_183) );
NAND2_X1 inst_800 ( .ZN(net_691), .A1(net_622), .A2(net_616) );
NAND2_X1 inst_780 ( .A2(net_805), .ZN(net_626), .A1(net_492) );
XOR2_X1 inst_10 ( .B(net_361), .Z(net_218), .A(net_199) );
XOR2_X1 inst_4 ( .A(net_375), .B(net_259), .Z(net_208) );
AND2_X4 inst_1110 ( .ZN(net_163), .A2(net_162), .A1(net_128) );
NAND3_X1 inst_581 ( .ZN(net_624), .A1(net_623), .A3(net_611), .A2(net_590) );
NAND2_X1 inst_600 ( .ZN(net_33), .A2(n208), .A1(n18) );
XOR2_X1 inst_28 ( .Z(net_480), .B(net_282), .A(net_206) );
CLKBUF_X1 inst_1089 ( .A(n471), .Z(n419) );
XOR2_X1 inst_49 ( .A(net_360), .Z(net_340), .B(net_200) );
XNOR2_X1 inst_204 ( .ZN(net_800), .B(net_720), .A(net_663) );
NAND3_X1 inst_592 ( .ZN(net_932), .A1(net_931), .A3(net_930), .A2(net_821) );
NAND4_X1 inst_546 ( .A1(net_739), .A2(net_738), .A4(net_737), .A3(net_707), .ZN(n416) );
INV_X1 inst_993 ( .A(net_512), .ZN(net_483) );
MUX2_X2 inst_910 ( .S(net_997), .A(net_779), .B(net_734), .Z(n301) );
NAND2_X1 inst_704 ( .ZN(net_152), .A2(net_137), .A1(net_41) );
NAND2_X1 inst_693 ( .ZN(net_310), .A2(net_144), .A1(net_70) );
NOR2_X1 inst_390 ( .ZN(net_343), .A1(net_164), .A2(net_84) );
CLKBUF_X1 inst_1062 ( .Z(n532), .A(n4415) );
NOR2_X1 inst_359 ( .A1(net_191), .ZN(net_83), .A2(n154) );
CLKBUF_X1 inst_1055 ( .Z(n546), .A(n3743) );
NAND2_X1 inst_765 ( .ZN(net_529), .A2(net_442), .A1(net_411) );
XNOR2_X1 inst_256 ( .B(net_956), .ZN(net_927), .A(net_883) );
NAND2_X1 inst_694 ( .ZN(net_307), .A2(net_145), .A1(net_44) );
NAND2_X1 inst_630 ( .ZN(net_62), .A2(n205), .A1(n18) );
INV_X1 inst_937 ( .ZN(net_111), .A(n4405) );
NOR2_X1 inst_401 ( .ZN(net_346), .A1(net_164), .A2(net_83) );
INV_X1 inst_923 ( .ZN(net_2), .A(n1469) );
NOR2_X1 inst_512 ( .ZN(net_976), .A2(net_960), .A1(net_856) );
MUX2_X2 inst_908 ( .Z(net_984), .S(net_983), .B(net_949), .A(net_948) );
NOR3_X1 inst_355 ( .ZN(net_914), .A1(net_870), .A3(net_869), .A2(net_187) );
NAND2_X1 inst_782 ( .ZN(net_631), .A1(net_630), .A2(net_628) );
XNOR2_X1 inst_218 ( .ZN(net_798), .A(net_797), .B(net_748) );
NAND2_X1 inst_647 ( .ZN(net_78), .A2(n224), .A1(n18) );
XOR2_X1 inst_6 ( .B(net_300), .Z(net_212), .A(net_211) );
XNOR2_X1 inst_194 ( .ZN(net_732), .B(net_731), .A(net_460) );
INV_X1 inst_1014 ( .ZN(net_1027), .A(net_722) );
NAND2_X1 inst_787 ( .A2(net_797), .ZN(net_661), .A1(net_537) );
NAND2_X1 inst_825 ( .ZN(net_877), .A2(net_847), .A1(net_754) );
NAND2_X1 inst_833 ( .ZN(net_899), .A2(net_898), .A1(net_654) );
XNOR2_X1 inst_123 ( .ZN(net_387), .A(net_329), .B(n3737) );
NOR2_X1 inst_509 ( .ZN(net_974), .A1(net_939), .A2(net_909) );
INV_X1 inst_930 ( .ZN(net_6), .A(n4432) );
NAND2_X1 inst_699 ( .ZN(net_286), .A2(net_148), .A1(net_64) );
INV_X1 inst_960 ( .ZN(net_27), .A(n58) );
XNOR2_X1 inst_118 ( .ZN(net_1001), .A(net_343), .B(n2236) );
INV_X1 inst_935 ( .ZN(net_11), .A(n2253) );
XNOR2_X1 inst_153 ( .ZN(net_447), .A(net_327), .B(net_291) );
NOR2_X1 inst_442 ( .A2(net_963), .A1(net_905), .ZN(net_591) );
XOR2_X1 inst_38 ( .Z(net_303), .A(net_302), .B(net_301) );
NOR2_X1 inst_381 ( .ZN(net_162), .A1(net_96), .A2(n1455) );
NAND2_X1 inst_726 ( .ZN(net_292), .A2(net_165), .A1(net_59) );
XNOR2_X1 inst_295 ( .ZN(net_1033), .B(net_1031), .A(net_1017) );
MUX2_X2 inst_883 ( .S(net_191), .Z(net_118), .B(net_27), .A(n4393) );
XNOR2_X1 inst_209 ( .ZN(net_884), .B(net_726), .A(net_682) );
INV_X1 inst_964 ( .ZN(net_169), .A(net_168) );
CLKBUF_X1 inst_1087 ( .Z(n432), .A(n1) );
XOR2_X1 inst_40 ( .Z(net_476), .B(net_286), .A(net_214) );
OR2_X4 inst_320 ( .A1(net_571), .ZN(net_540), .A2(net_511) );
XNOR2_X1 inst_167 ( .ZN(net_513), .A(net_512), .B(net_511) );
NAND2_X1 inst_607 ( .ZN(net_40), .A2(n202), .A1(n18) );
INV_X1 inst_1026 ( .ZN(net_595), .A(net_492) );
NAND2_X1 inst_756 ( .ZN(net_609), .A1(net_590), .A2(net_414) );
XNOR2_X1 inst_95 ( .ZN(net_230), .A(net_123), .B(net_107) );
XOR2_X1 inst_1 ( .A(net_363), .Z(net_203), .B(net_202) );
NOR2_X1 inst_439 ( .A1(net_1031), .A2(net_956), .ZN(net_604) );
OR2_X4 inst_331 ( .A1(net_814), .ZN(net_757), .A2(net_670) );
CLKBUF_X1 inst_1070 ( .Z(n492), .A(n2224) );
XNOR2_X1 inst_235 ( .ZN(net_862), .A(net_861), .B(net_806) );
NAND2_X1 inst_750 ( .ZN(net_243), .A2(net_235), .A1(n1462) );
OR2_X4 inst_317 ( .ZN(net_382), .A2(net_381), .A1(net_162) );
AND2_X4 inst_1123 ( .ZN(net_425), .A2(net_424), .A1(net_379) );
CLKBUF_X1 inst_1082 ( .Z(n444), .A(n1480) );
NAND2_X1 inst_667 ( .A2(net_191), .ZN(net_131), .A1(n100) );
XNOR2_X1 inst_278 ( .A(net_1016), .ZN(net_1006), .B(net_972) );
NOR2_X1 inst_467 ( .ZN(net_558), .A2(net_557), .A1(net_503) );
INV_X1 inst_992 ( .ZN(net_728), .A(net_384) );
XNOR2_X1 inst_105 ( .ZN(net_324), .A(net_323), .B(net_282) );
NOR2_X1 inst_488 ( .A2(net_987), .ZN(net_807), .A1(net_677) );
NOR2_X1 inst_387 ( .A1(net_164), .ZN(net_130), .A2(net_98) );
INV_X1 inst_997 ( .A(net_965), .ZN(net_489) );
MUX2_X2 inst_857 ( .Z(net_228), .S(net_191), .A(net_24), .B(n113) );
XNOR2_X1 inst_254 ( .B(net_939), .ZN(net_919), .A(net_888) );
NAND2_X1 inst_654 ( .A2(net_191), .ZN(net_139), .A1(n144) );
NAND2_X1 inst_625 ( .ZN(net_57), .A2(n222), .A1(n18) );
XNOR2_X1 inst_225 ( .ZN(net_839), .B(net_775), .A(net_772) );
NOR2_X1 inst_508 ( .ZN(net_938), .A2(net_906), .A1(net_814) );
NAND3_X1 inst_568 ( .ZN(net_584), .A3(net_563), .A2(net_361), .A1(net_360) );
NAND4_X1 inst_523 ( .A2(net_568), .A4(net_567), .ZN(net_466), .A1(net_358), .A3(net_354) );
NOR2_X1 inst_365 ( .A1(net_191), .ZN(net_89), .A2(n211) );
XOR2_X1 inst_67 ( .Z(net_967), .B(net_272), .A(n3723) );
INV_X1 inst_954 ( .ZN(net_23), .A(n4420) );
XNOR2_X1 inst_181 ( .ZN(net_641), .B(net_446), .A(net_279) );
AND2_X4 inst_1135 ( .ZN(net_671), .A2(net_574), .A1(net_192) );
NOR2_X1 inst_391 ( .ZN(net_356), .A1(net_164), .A2(net_101) );
NAND2_X1 inst_661 ( .A2(net_191), .ZN(net_144), .A1(n121) );
NAND3_X1 inst_590 ( .ZN(net_813), .A1(net_812), .A3(net_675), .A2(n89) );
NAND2_X1 inst_713 ( .ZN(net_275), .A2(net_154), .A1(net_74) );
XNOR2_X1 inst_202 ( .ZN(net_792), .A(net_660), .B(net_570) );
NAND2_X1 inst_634 ( .ZN(net_66), .A2(n225), .A1(n18) );
NOR2_X1 inst_419 ( .ZN(net_247), .A2(net_171), .A1(n2236) );
AND3_X4 inst_1105 ( .ZN(net_678), .A2(net_615), .A3(net_606), .A1(net_603) );
INV_X1 inst_981 ( .A(net_275), .ZN(net_181) );
NOR2_X1 inst_477 ( .A2(net_750), .ZN(net_718), .A1(net_543) );
NOR2_X1 inst_423 ( .ZN(net_531), .A2(net_174), .A1(n2218) );
CLKBUF_X1 inst_1069 ( .Z(n494), .A(n2218) );
NAND2_X1 inst_835 ( .ZN(net_931), .A1(net_904), .A2(net_871) );
XNOR2_X1 inst_136 ( .ZN(net_696), .A(net_348), .B(n1480) );
XOR2_X1 inst_30 ( .Z(net_467), .B(net_323), .A(net_285) );
OR2_X4 inst_330 ( .A1(net_756), .A2(net_668), .ZN(net_629) );
NAND2_X1 inst_610 ( .ZN(net_43), .A2(n181), .A1(n18) );
AND2_X4 inst_1112 ( .A2(net_965), .A1(net_751), .ZN(net_399) );
INV_X1 inst_1036 ( .ZN(net_845), .A(net_712) );
XNOR2_X1 inst_233 ( .ZN(net_859), .B(net_858), .A(net_801) );
NAND2_X1 inst_710 ( .ZN(net_290), .A2(net_148), .A1(net_37) );
XNOR2_X1 inst_165 ( .ZN(net_509), .B(net_340), .A(net_339) );
INV_X1 inst_941 ( .ZN(net_756), .A(n4526) );
XNOR2_X1 inst_271 ( .ZN(net_990), .A(net_989), .B(net_957) );
XOR2_X1 inst_34 ( .Z(net_294), .A(net_293), .B(net_292) );
XOR2_X1 inst_12 ( .B(net_308), .A(net_297), .Z(net_222) );
INV_X1 inst_1047 ( .ZN(net_951), .A(net_931) );
NAND4_X1 inst_529 ( .ZN(net_574), .A2(net_573), .A4(net_572), .A1(net_421), .A3(net_269) );
XOR2_X1 inst_56 ( .Z(net_567), .B(net_356), .A(net_204) );
XOR2_X1 inst_71 ( .A(net_462), .Z(net_461), .B(net_460) );
OR3_X4 inst_308 ( .A2(net_720), .ZN(net_676), .A1(net_596), .A3(net_544) );
XOR2_X1 inst_60 ( .Z(net_369), .A(net_368), .B(net_367) );
NOR2_X1 inst_455 ( .A2(net_925), .A1(net_630), .ZN(net_516) );
CLKBUF_X1 inst_1064 ( .Z(n528), .A(n4427) );
NAND2_X1 inst_675 ( .A2(net_80), .ZN(n289), .A1(n1197) );
NAND2_X1 inst_758 ( .A1(net_911), .ZN(net_522), .A2(net_411) );
NOR2_X1 inst_496 ( .ZN(net_849), .A1(net_848), .A2(net_815) );
MUX2_X2 inst_860 ( .S(net_191), .Z(net_110), .B(net_20), .A(n3698) );
OR2_X4 inst_336 ( .ZN(net_934), .A1(net_913), .A2(net_885) );
NAND3_X1 inst_563 ( .ZN(net_758), .A3(net_576), .A2(net_564), .A1(net_377) );
NAND3_X1 inst_583 ( .ZN(net_746), .A1(net_656), .A3(net_655), .A2(net_497) );
INV_X1 inst_943 ( .ZN(net_108), .A(n106) );
XNOR2_X1 inst_258 ( .A(net_965), .ZN(net_941), .B(net_903) );
NOR2_X1 inst_376 ( .A1(net_191), .ZN(net_101), .A2(n166) );
XNOR2_X1 inst_143 ( .ZN(net_394), .B(net_226), .A(net_212) );
XNOR2_X1 inst_265 ( .ZN(net_966), .A(net_965), .B(net_919) );
NOR2_X1 inst_482 ( .A2(net_772), .ZN(net_771), .A1(net_599) );
INV_X1 inst_1040 ( .ZN(net_765), .A(net_764) );
NAND2_X1 inst_682 ( .ZN(net_293), .A2(net_131), .A1(net_35) );
NAND2_X1 inst_736 ( .A1(net_321), .A2(net_216), .ZN(net_197) );
NAND4_X1 inst_544 ( .ZN(net_764), .A4(net_671), .A2(net_565), .A1(net_470), .A3(net_408) );
XNOR2_X1 inst_238 ( .ZN(net_881), .B(net_880), .A(net_839) );
CLKBUF_X1 inst_1093 ( .A(n292), .Z(n281) );
NAND4_X1 inst_539 ( .ZN(net_848), .A4(net_581), .A2(net_575), .A3(net_477), .A1(net_195) );
NAND2_X1 inst_724 ( .ZN(net_277), .A2(net_142), .A1(net_38) );
MUX2_X2 inst_895 ( .B(net_853), .S(net_852), .A(net_794), .Z(n376) );
XNOR2_X1 inst_178 ( .ZN(net_638), .B(net_510), .A(net_359) );
XNOR2_X1 inst_111 ( .ZN(net_366), .A(net_365), .B(net_364) );
INV_X1 inst_975 ( .A(net_289), .ZN(net_177) );
NAND2_X1 inst_734 ( .A1(net_282), .A2(net_206), .ZN(net_194) );
CLKBUF_X1 inst_1077 ( .Z(n478), .A(n2211) );
XNOR2_X1 inst_222 ( .ZN(net_827), .A(net_769), .B(net_664) );
XNOR2_X1 inst_284 ( .B(net_1018), .A(net_536), .ZN(n471) );
NAND2_X1 inst_806 ( .ZN(net_714), .A2(net_713), .A1(net_541) );
XNOR2_X1 inst_280 ( .ZN(net_1010), .B(net_1009), .A(net_979) );
NAND2_X1 inst_763 ( .ZN(net_524), .A2(net_462), .A1(net_388) );
NOR4_X1 inst_346 ( .ZN(net_907), .A2(net_690), .A1(net_553), .A4(net_502), .A3(net_245) );
NOR2_X1 inst_491 ( .A1(net_865), .ZN(net_847), .A2(net_763) );
CLKBUF_X1 inst_1052 ( .Z(n552), .A(n3723) );
INV_X1 inst_978 ( .A(net_325), .ZN(net_239) );
CLKBUF_X1 inst_1079 ( .Z(n450), .A(n1459) );
NAND2_X1 inst_842 ( .ZN(net_954), .A2(net_924), .A1(net_805) );
NAND4_X1 inst_537 ( .ZN(net_646), .A1(net_645), .A2(net_644), .A3(net_267), .A4(net_266) );
NAND2_X1 inst_826 ( .ZN(net_850), .A2(net_847), .A1(net_824) );
NAND4_X1 inst_551 ( .ZN(net_913), .A4(net_820), .A3(net_559), .A1(net_532), .A2(net_465) );
CLKBUF_X1 inst_1051 ( .Z(n554), .A(n3717) );
XNOR2_X1 inst_207 ( .B(net_1004), .A(net_693), .ZN(n394) );
NOR3_X1 inst_353 ( .ZN(net_713), .A1(net_547), .A3(net_436), .A2(net_430) );
NOR2_X1 inst_495 ( .A2(net_847), .ZN(net_846), .A1(net_845) );
NOR2_X1 inst_506 ( .ZN(net_915), .A2(net_914), .A1(net_893) );
XNOR2_X1 inst_159 ( .A(net_485), .ZN(net_455), .B(net_454) );
MUX2_X2 inst_872 ( .Z(net_306), .S(net_191), .A(net_29), .B(n60) );
INV_X1 inst_951 ( .ZN(net_21), .A(n3743) );
XNOR2_X1 inst_134 ( .ZN(net_601), .A(net_331), .B(n4394) );
CLKBUF_X1 inst_1085 ( .Z(n438), .A(n1496) );
OR2_X4 inst_333 ( .A2(net_865), .ZN(net_864), .A1(net_762) );
NAND2_X1 inst_712 ( .ZN(net_342), .A2(net_160), .A1(net_73) );
XNOR2_X1 inst_131 ( .ZN(net_592), .A(net_278), .B(n4405) );
NOR2_X1 inst_406 ( .ZN(net_355), .A1(net_164), .A2(net_103) );
XNOR2_X1 inst_160 ( .ZN(net_456), .B(net_288), .A(net_256) );
NOR2_X1 inst_462 ( .A1(net_999), .ZN(net_553), .A2(net_552) );
OR2_X4 inst_328 ( .A1(net_880), .ZN(net_539), .A2(net_538) );
MUX2_X2 inst_869 ( .Z(net_281), .S(net_191), .A(net_15), .B(n74) );
XOR2_X1 inst_19 ( .Z(net_263), .A(net_262), .B(net_261) );
XOR2_X1 inst_47 ( .Z(net_332), .B(net_331), .A(net_138) );
XOR2_X1 inst_8 ( .B(net_305), .Z(net_215), .A(net_214) );
NAND2_X1 inst_818 ( .A2(net_867), .ZN(net_823), .A1(net_744) );
NOR2_X1 inst_370 ( .A1(net_191), .ZN(net_95), .A2(n175) );
NAND2_X1 inst_762 ( .ZN(net_420), .A2(net_382), .A1(net_182) );
NAND3_X1 inst_573 ( .ZN(net_653), .A3(net_613), .A2(net_608), .A1(net_601) );
XNOR2_X1 inst_100 ( .A(net_267), .ZN(net_260), .B(net_136) );
INV_X1 inst_965 ( .A(net_290), .ZN(net_170) );
INV_X1 inst_921 ( .ZN(net_0), .A(n4400) );
XNOR2_X1 inst_279 ( .B(net_975), .A(net_965), .ZN(n319) );
XOR2_X1 inst_81 ( .Z(net_796), .A(net_795), .B(net_794) );
NAND2_X1 inst_612 ( .ZN(net_45), .A2(n18), .A1(n159) );
NAND4_X1 inst_525 ( .ZN(net_473), .A3(net_472), .A4(net_471), .A2(net_400), .A1(net_238) );
INV_X1 inst_1012 ( .ZN(net_1009), .A(net_592) );
MUX2_X2 inst_901 ( .Z(net_948), .A(net_947), .B(net_946), .S(net_811) );
NOR2_X1 inst_434 ( .ZN(net_645), .A2(net_409), .A1(net_316) );
NAND2_X1 inst_790 ( .ZN(net_666), .A2(net_656), .A1(net_655) );
INV_X1 inst_1032 ( .ZN(net_654), .A(net_653) );
INV_X1 inst_1009 ( .ZN(net_956), .A(net_411) );
NAND2_X1 inst_751 ( .ZN(net_514), .A2(net_234), .A1(n3729) );
MUX2_X2 inst_906 ( .Z(net_978), .S(net_977), .A(net_863), .B(net_830) );
NAND2_X1 inst_845 ( .A2(net_971), .ZN(net_969), .A1(net_652) );
NAND2_X1 inst_733 ( .A1(net_356), .A2(net_204), .ZN(net_193) );
NOR2_X1 inst_377 ( .A1(net_191), .ZN(net_102), .A2(n174) );
XNOR2_X1 inst_142 ( .ZN(net_393), .B(net_210), .A(net_208) );
XOR2_X1 inst_78 ( .Z(net_802), .A(net_749), .B(net_716) );
XNOR2_X1 inst_177 ( .ZN(net_637), .B(net_457), .A(net_322) );
NAND2_X1 inst_783 ( .ZN(net_632), .A2(net_610), .A1(net_609) );
MUX2_X2 inst_885 ( .Z(net_216), .S(net_191), .A(net_9), .B(n83) );
XNOR2_X1 inst_183 ( .ZN(net_643), .B(net_450), .A(net_353) );
NAND2_X1 inst_852 ( .ZN(net_996), .A2(net_995), .A1(net_728) );
AND2_X4 inst_1142 ( .ZN(net_960), .A2(net_959), .A1(net_722) );
INV_X1 inst_928 ( .ZN(n341), .A(n15) );
INV_X1 inst_1028 ( .A(net_758), .ZN(net_600) );
XNOR2_X1 inst_107 ( .ZN(net_337), .A(net_336), .B(net_335) );
NOR2_X1 inst_393 ( .ZN(net_336), .A1(net_164), .A2(net_81) );
NAND2_X1 inst_615 ( .ZN(net_48), .A2(n236), .A1(n18) );
INV_X1 inst_990 ( .ZN(net_486), .A(net_452) );
XNOR2_X1 inst_92 ( .A(net_269), .ZN(net_226), .B(net_118) );
NOR4_X1 inst_345 ( .ZN(net_950), .A2(net_691), .A1(net_555), .A4(net_500), .A3(net_247) );
CLKBUF_X1 inst_1050 ( .Z(n556), .A(n3711) );
NAND2_X1 inst_643 ( .ZN(net_75), .A2(n235), .A1(n18) );
NAND2_X1 inst_697 ( .ZN(net_312), .A2(net_147), .A1(net_79) );
NOR2_X1 inst_487 ( .A2(net_861), .ZN(net_790), .A1(net_607) );
XNOR2_X1 inst_200 ( .ZN(net_740), .B(net_639), .A(net_393) );
XOR2_X1 inst_57 ( .Z(net_472), .A(net_361), .B(net_360) );
OR2_X4 inst_338 ( .A2(net_977), .ZN(net_973), .A1(net_808) );
NOR2_X1 inst_417 ( .ZN(net_401), .A2(net_177), .A1(n4432) );
NAND2_X1 inst_671 ( .A2(net_191), .ZN(net_135), .A1(n141) );
INV_X1 inst_1017 ( .ZN(net_1031), .A(net_696) );
XOR2_X1 inst_21 ( .Z(net_412), .B(net_265), .A(net_209) );
NAND3_X1 inst_579 ( .A1(net_722), .ZN(net_621), .A3(net_613), .A2(net_556) );
XNOR2_X1 inst_281 ( .ZN(net_1013), .A(net_1012), .B(net_980) );
CLKBUF_X1 inst_1094 ( .A(n341), .Z(n279) );
NAND3_X1 inst_585 ( .ZN(net_772), .A1(net_689), .A3(net_494), .A2(net_426) );
NAND2_X1 inst_698 ( .ZN(net_261), .A2(net_144), .A1(net_78) );
MUX2_X2 inst_893 ( .S(net_852), .B(net_515), .A(net_513), .Z(n382) );
XOR2_X1 inst_88 ( .B(net_1031), .A(net_1011), .Z(n330) );
NOR2_X1 inst_410 ( .ZN(net_384), .A2(net_235), .A1(n1462) );
OR2_X4 inst_316 ( .ZN(net_233), .A1(net_232), .A2(net_231) );
XNOR2_X1 inst_220 ( .ZN(net_806), .A(net_805), .B(net_752) );
NAND2_X1 inst_851 ( .ZN(net_993), .A1(net_987), .A2(net_973) );
NAND2_X1 inst_831 ( .ZN(net_879), .A2(net_877), .A1(net_875) );
NOR2_X1 inst_360 ( .A1(net_191), .ZN(net_84), .A2(n157) );
NOR2_X1 inst_383 ( .A2(net_124), .ZN(net_116), .A1(n38) );
INV_X1 inst_1023 ( .ZN(net_880), .A(net_597) );
XOR2_X1 inst_50 ( .Z(net_568), .B(net_355), .A(net_341) );
NAND2_X1 inst_773 ( .ZN(net_1019), .A2(net_677), .A1(net_443) );
XNOR2_X1 inst_245 ( .ZN(net_942), .B(net_855), .A(net_512) );
NAND3_X1 inst_569 ( .ZN(net_808), .A2(net_696), .A1(net_617), .A3(net_594) );
CLKBUF_X1 inst_1080 ( .Z(n448), .A(n1469) );
AND2_X4 inst_1124 ( .ZN(net_434), .A1(net_433), .A2(net_432) );
NAND2_X1 inst_678 ( .ZN(net_232), .A2(net_124), .A1(n38) );
NAND2_X1 inst_624 ( .ZN(net_56), .A2(n207), .A1(n18) );
AND3_X4 inst_1103 ( .ZN(net_599), .A3(net_598), .A1(net_597), .A2(net_414) );
XNOR2_X1 inst_260 ( .ZN(net_955), .B(net_925), .A(net_910) );
AND2_X4 inst_1129 ( .A1(net_601), .A2(net_548), .ZN(net_542) );
NAND2_X1 inst_854 ( .A2(net_1003), .A1(net_920), .ZN(n249) );
XNOR2_X1 inst_147 ( .ZN(net_398), .A(net_218), .B(net_203) );
NAND2_X1 inst_837 ( .ZN(net_908), .A2(net_897), .A1(net_797) );
OR2_X4 inst_313 ( .A1(net_200), .A2(net_199), .ZN(net_188) );
NAND2_X1 inst_744 ( .ZN(net_504), .A2(net_348), .A1(net_122) );
NAND4_X1 inst_549 ( .A4(net_875), .ZN(net_818), .A3(net_753), .A2(net_712), .A1(n4526) );
INV_X1 inst_1041 ( .A(net_950), .ZN(net_819) );
XNOR2_X1 inst_234 ( .ZN(net_860), .A(net_804), .B(net_799) );
NAND4_X1 inst_522 ( .ZN(net_465), .A1(net_464), .A3(net_463), .A4(net_462), .A2(net_439) );
XNOR2_X1 inst_236 ( .ZN(net_873), .A(net_826), .B(net_771) );
INV_X1 inst_1002 ( .ZN(net_745), .A(net_428) );
NOR2_X1 inst_478 ( .ZN(net_721), .A1(net_720), .A2(net_665) );
NAND4_X1 inst_553 ( .ZN(net_981), .A3(net_953), .A2(net_952), .A1(net_932), .A4(net_929) );
XOR2_X1 inst_65 ( .Z(net_380), .A(net_379), .B(net_378) );
NAND4_X1 inst_536 ( .ZN(net_593), .A4(net_568), .A1(net_488), .A3(net_365), .A2(net_364) );
XNOR2_X1 inst_242 ( .ZN(net_887), .A(net_837), .B(net_789) );
INV_X1 inst_986 ( .A(net_346), .ZN(net_185) );
NAND2_X1 inst_688 ( .ZN(net_141), .A2(net_135), .A1(net_34) );
NOR2_X1 inst_516 ( .ZN(net_1014), .A2(net_992), .A1(net_861) );
NAND2_X1 inst_804 ( .ZN(net_697), .A1(net_696), .A2(net_634) );
XNOR2_X1 inst_190 ( .ZN(net_706), .B(net_643), .A(net_254) );
XOR2_X1 inst_13 ( .B(net_284), .A(net_281), .Z(net_223) );
INV_X8 inst_919 ( .ZN(net_191), .A(n18) );
XNOR2_X1 inst_116 ( .ZN(net_374), .A(net_373), .B(net_372) );
NOR2_X1 inst_416 ( .ZN(net_556), .A2(net_186), .A1(n4400) );
NAND2_X1 inst_598 ( .ZN(net_32), .A2(n227), .A1(n18) );
AND2_X4 inst_1133 ( .ZN(net_585), .A2(net_475), .A1(net_193) );
NOR2_X1 inst_471 ( .ZN(net_867), .A1(net_676), .A2(net_674) );
NAND2_X1 inst_799 ( .ZN(net_690), .A1(net_621), .A2(net_614) );
XNOR2_X1 inst_219 ( .ZN(net_801), .A(net_800), .B(net_799) );
NAND2_X1 inst_738 ( .ZN(net_237), .A1(net_200), .A2(net_199) );
NAND2_X1 inst_719 ( .ZN(net_289), .A2(net_161), .A1(net_76) );
NAND2_X1 inst_840 ( .ZN(net_935), .A2(net_934), .A1(net_708) );
XNOR2_X1 inst_255 ( .ZN(net_926), .B(net_925), .A(net_881) );
NAND4_X1 inst_542 ( .ZN(net_761), .A3(net_624), .A4(net_612), .A2(net_530), .A1(net_474) );
XNOR2_X1 inst_128 ( .ZN(net_411), .A(net_351), .B(n1469) );
NOR2_X1 inst_453 ( .ZN(net_505), .A1(net_504), .A2(net_503) );
AND2_X4 inst_1134 ( .ZN(net_665), .A2(net_545), .A1(net_423) );
NOR2_X1 inst_493 ( .ZN(net_833), .A1(net_832), .A2(net_783) );
XOR2_X1 inst_23 ( .A(net_295), .Z(net_270), .B(net_269) );
MUX2_X2 inst_896 ( .Z(net_863), .B(net_829), .A(net_828), .S(net_809) );
OR2_X2 inst_339 ( .ZN(n402), .A2(n57), .A1(n5) );
AND2_X4 inst_1113 ( .ZN(net_563), .A2(net_471), .A1(net_400) );
NOR3_X1 inst_351 ( .ZN(net_762), .A1(net_571), .A2(net_570), .A3(net_525) );
NOR2_X1 inst_408 ( .ZN(net_166), .A1(net_164), .A2(net_89) );
INV_X1 inst_973 ( .A(net_292), .ZN(net_176) );
AND2_X4 inst_1144 ( .ZN(net_992), .A2(net_991), .A1(net_724) );
OR2_X4 inst_325 ( .A1(net_630), .ZN(net_610), .A2(net_538) );
NOR2_X1 inst_461 ( .ZN(net_627), .A1(net_533), .A2(net_527) );
NOR2_X1 inst_385 ( .ZN(net_367), .A1(net_164), .A2(net_97) );
NAND2_X1 inst_829 ( .ZN(net_876), .A1(net_875), .A2(net_846) );
NAND2_X1 inst_812 ( .ZN(net_736), .A2(net_735), .A1(n4526) );
XNOR2_X1 inst_197 ( .ZN(net_737), .B(net_635), .A(net_456) );
XNOR2_X1 inst_179 ( .ZN(net_639), .B(net_458), .A(net_223) );
XOR2_X1 inst_24 ( .Z(net_273), .A(net_272), .B(net_271) );
INV_X1 inst_955 ( .ZN(net_24), .A(n1462) );
XNOR2_X1 inst_114 ( .ZN(net_989), .A(net_349), .B(n1486) );
AND2_X4 inst_1122 ( .ZN(net_527), .A1(net_464), .A2(net_462) );
XOR2_X1 inst_76 ( .Z(net_778), .A(net_726), .B(net_681) );
NAND2_X1 inst_617 ( .ZN(net_50), .A2(n237), .A1(n18) );
AND2_X4 inst_1127 ( .ZN(net_441), .A1(net_440), .A2(net_439) );
XNOR2_X1 inst_150 ( .ZN(net_444), .B(net_273), .A(net_251) );
XNOR2_X1 inst_172 ( .ZN(net_587), .B(net_396), .A(net_217) );
NOR2_X1 inst_362 ( .A1(net_191), .ZN(net_86), .A2(n165) );
XNOR2_X1 inst_277 ( .ZN(net_1005), .A(net_1004), .B(net_968) );
XOR2_X1 inst_83 ( .B(net_967), .A(net_773), .Z(n388) );
XNOR2_X1 inst_121 ( .ZN(net_439), .A(net_345), .B(n2256) );
MUX2_X2 inst_887 ( .Z(net_364), .S(net_191), .A(net_2), .B(n111) );
OR3_X4 inst_306 ( .A1(net_1025), .A3(net_967), .A2(net_493), .ZN(net_474) );
NAND4_X1 inst_534 ( .ZN(net_589), .A4(net_569), .A2(net_567), .A3(net_403), .A1(net_228) );
CLKBUF_X1 inst_1065 ( .Z(n526), .A(n4432) );
CLKBUF_X1 inst_1057 ( .Z(n542), .A(n3701) );
NAND2_X1 inst_596 ( .ZN(net_30), .A2(n18), .A1(n178) );
XNOR2_X1 inst_90 ( .ZN(net_536), .A(net_124), .B(n38) );
XNOR2_X1 inst_140 ( .ZN(net_534), .B(net_392), .A(net_116) );
XNOR2_X1 inst_267 ( .A(net_989), .ZN(net_972), .B(net_927) );
NAND2_X1 inst_847 ( .ZN(net_995), .A2(net_971), .A1(net_911) );
NAND2_X1 inst_748 ( .ZN(net_484), .A2(net_317), .A1(net_117) );
AND2_X2 inst_1146 ( .ZN(n278), .A1(n163), .A2(n1) );
NAND2_X1 inst_716 ( .ZN(net_318), .A2(net_151), .A1(net_31) );
NAND2_X1 inst_637 ( .ZN(net_69), .A2(n233), .A1(n18) );
NAND4_X1 inst_530 ( .ZN(net_575), .A2(net_476), .A1(net_425), .A4(net_417), .A3(net_378) );
NAND4_X1 inst_547 ( .A4(net_740), .A1(net_703), .A2(net_702), .A3(net_701), .ZN(n414) );
NAND2_X1 inst_792 ( .ZN(net_893), .A1(net_766), .A2(net_669) );
NAND2_X1 inst_720 ( .ZN(net_329), .A2(net_127), .A1(net_69) );
INV_X1 inst_958 ( .ZN(net_122), .A(n1480) );
NOR2_X1 inst_368 ( .A1(net_191), .ZN(net_92), .A2(n213) );
INV_X1 inst_1010 ( .ZN(net_517), .A(net_388) );
NAND2_X1 inst_803 ( .ZN(net_695), .A1(net_673), .A2(net_633) );
NAND2_X1 inst_769 ( .ZN(net_431), .A1(net_430), .A2(net_428) );
XNOR2_X1 inst_174 ( .B(net_756), .A(net_597), .ZN(n373) );
XNOR2_X1 inst_274 ( .ZN(net_998), .A(net_967), .B(net_955) );
NAND2_X1 inst_662 ( .A2(net_191), .ZN(net_160), .A1(n135) );
NAND2_X1 inst_701 ( .ZN(net_272), .A2(net_149), .A1(net_75) );
XNOR2_X1 inst_164 ( .ZN(net_508), .B(net_313), .A(net_287) );
MUX2_X2 inst_867 ( .Z(net_206), .S(net_191), .A(net_5), .B(n73) );
NAND2_X1 inst_820 ( .A2(net_907), .ZN(net_811), .A1(net_674) );
XOR2_X1 inst_5 ( .B(net_301), .Z(net_210), .A(net_209) );
XNOR2_X1 inst_157 ( .ZN(net_451), .B(net_311), .A(net_296) );
NAND2_X1 inst_729 ( .ZN(net_302), .A2(net_165), .A1(net_71) );
XNOR2_X1 inst_213 ( .ZN(net_777), .A(net_776), .B(net_730) );
XOR2_X1 inst_68 ( .Z(net_571), .B(net_328), .A(n3729) );
NAND2_X1 inst_604 ( .ZN(net_37), .A2(n219), .A1(n18) );
XOR2_X1 inst_53 ( .Z(net_350), .A(net_349), .B(net_348) );
INV_X1 inst_1007 ( .ZN(net_939), .A(net_603) );
XNOR2_X1 inst_205 ( .ZN(net_752), .A(net_751), .B(net_750) );
NAND2_X1 inst_753 ( .ZN(net_454), .A2(net_239), .A1(n4420) );
NOR2_X1 inst_380 ( .A1(net_191), .ZN(net_105), .A2(n164) );
INV_X1 inst_946 ( .ZN(net_17), .A(n85) );
NAND2_X1 inst_651 ( .A2(net_191), .ZN(net_140), .A1(n23) );
XNOR2_X1 inst_292 ( .ZN(net_1030), .B(net_1029), .A(net_1013) );
INV_X1 inst_999 ( .A(net_1001), .ZN(net_498) );
NOR2_X1 inst_379 ( .A1(net_191), .ZN(net_104), .A2(n216) );
INV_X1 inst_926 ( .ZN(net_113), .A(n4410) );
XNOR2_X1 inst_186 ( .ZN(net_702), .B(net_587), .A(net_398) );
XOR2_X1 inst_17 ( .A(net_376), .B(net_258), .Z(net_256) );
NAND2_X1 inst_706 ( .ZN(net_295), .A2(net_153), .A1(net_47) );
NAND2_X1 inst_759 ( .ZN(net_490), .A1(net_463), .A2(net_439) );
XNOR2_X1 inst_249 ( .B(net_939), .ZN(net_903), .A(net_862) );
MUX2_X2 inst_863 ( .Z(net_269), .S(net_191), .A(net_19), .B(n77) );
NAND2_X1 inst_839 ( .ZN(net_924), .A2(net_923), .A1(net_595) );
INV_X1 inst_1015 ( .ZN(net_905), .A(net_601) );
XNOR2_X1 inst_240 ( .ZN(net_928), .B(net_843), .A(net_464) );
XNOR2_X1 inst_110 ( .B(net_365), .ZN(net_359), .A(net_358) );
MUX2_X2 inst_891 ( .S(net_191), .Z(net_123), .A(net_12), .B(n2204) );
XOR2_X1 inst_74 ( .Z(net_779), .A(net_733), .B(net_627) );
XNOR2_X1 inst_288 ( .ZN(net_1022), .B(net_1009), .A(net_1000) );
XNOR2_X1 inst_229 ( .B(net_852), .A(net_571), .ZN(n385) );
NOR2_X1 inst_396 ( .A1(net_164), .ZN(net_159), .A2(net_86) );
XNOR2_X1 inst_99 ( .A(net_307), .B(net_298), .ZN(net_257) );
NAND2_X1 inst_669 ( .A2(net_191), .ZN(net_146), .A1(n41) );
NAND2_X1 inst_664 ( .A2(net_191), .ZN(net_127), .A1(n127) );
XNOR2_X1 inst_283 ( .ZN(net_1017), .A(net_1016), .B(net_990) );
OR3_X2 inst_311 ( .ZN(net_891), .A1(net_890), .A3(net_889), .A2(net_835) );
MUX2_X2 inst_917 ( .Z(net_1038), .A(net_1035), .B(net_1028), .S(net_983) );
NOR2_X1 inst_372 ( .A1(net_191), .ZN(net_97), .A2(n155) );
INV_X1 inst_988 ( .ZN(net_238), .A(net_237) );
XNOR2_X1 inst_215 ( .ZN(net_787), .A(net_718), .B(net_244) );
XNOR2_X1 inst_169 ( .ZN(net_842), .A(net_517), .B(net_462) );
NOR2_X1 inst_421 ( .ZN(net_440), .A2(net_185), .A1(n2253) );
CLKBUF_X1 inst_1092 ( .A(n289), .Z(n284) );
NAND4_X1 inst_555 ( .A3(net_986), .A4(net_937), .A2(net_876), .A1(net_818), .ZN(n246) );
NAND2_X1 inst_849 ( .ZN(net_1018), .A1(net_987), .A2(net_969) );
NAND2_X1 inst_816 ( .ZN(net_852), .A2(net_784), .A1(net_688) );
NOR2_X1 inst_431 ( .ZN(net_391), .A2(net_390), .A1(net_169) );
XOR2_X1 inst_3 ( .B(net_285), .Z(net_207), .A(net_206) );
NOR4_X1 inst_348 ( .A4(net_892), .ZN(net_812), .A1(net_758), .A3(net_757), .A2(net_649) );
CLKBUF_X1 inst_1090 ( .Z(n3), .A(n1) );
MUX2_X2 inst_889 ( .Z(net_375), .S(net_191), .A(net_1), .B(n53) );
NAND3_X1 inst_577 ( .ZN(net_618), .A1(net_617), .A3(net_604), .A2(net_384) );
NAND3_X1 inst_566 ( .ZN(net_581), .A3(net_566), .A2(net_312), .A1(net_306) );
XOR2_X1 inst_36 ( .Z(net_299), .A(net_298), .B(net_297) );
NAND2_X1 inst_656 ( .A2(net_191), .ZN(net_126), .A1(n130) );
NAND2_X1 inst_645 ( .ZN(net_77), .A2(n200), .A1(n18) );
XOR2_X1 inst_45 ( .Z(net_327), .A(net_326), .B(net_325) );
NOR2_X1 inst_503 ( .ZN(net_916), .A1(net_905), .A2(net_872) );
NOR2_X1 inst_451 ( .ZN(net_500), .A1(net_499), .A2(net_498) );
AND3_X4 inst_1108 ( .ZN(net_684), .A1(net_610), .A3(net_609), .A2(net_493) );
XNOR2_X1 inst_269 ( .A(net_1001), .ZN(net_980), .B(net_941) );
NOR2_X1 inst_458 ( .ZN(net_530), .A2(net_427), .A1(net_250) );
NOR2_X1 inst_444 ( .A1(net_1029), .ZN(net_606), .A2(net_489) );
NAND2_X1 inst_797 ( .ZN(net_688), .A2(net_679), .A1(n4526) );
AND4_X1 inst_1097 ( .A2(net_480), .ZN(net_468), .A4(net_467), .A3(net_284), .A1(net_283) );
NAND2_X1 inst_686 ( .ZN(net_317), .A2(net_139), .A1(net_45) );
NAND2_X1 inst_741 ( .ZN(net_497), .A2(net_278), .A1(net_111) );
NOR2_X1 inst_514 ( .ZN(net_1007), .A2(net_995), .A1(net_529) );
INV_X1 inst_967 ( .A(net_372), .ZN(net_235) );
NAND2_X1 inst_685 ( .ZN(net_138), .A2(net_137), .A1(net_32) );
XOR2_X1 inst_63 ( .Z(net_485), .B(net_326), .A(n4427) );
XNOR2_X1 inst_119 ( .ZN(net_442), .A(net_352), .B(n106) );
INV_X1 inst_939 ( .ZN(net_13), .A(n2239) );
NAND2_X1 inst_676 ( .A2(net_191), .ZN(net_125), .A1(n35) );
AND2_X4 inst_1118 ( .ZN(net_573), .A2(net_413), .A1(net_299) );
AND2_X4 inst_1115 ( .A2(net_568), .ZN(net_403), .A1(net_373) );
MUX2_X2 inst_874 ( .S(net_191), .Z(net_114), .B(net_26), .A(n2208) );
INV_X1 inst_1019 ( .ZN(net_1029), .A(net_724) );
INV_X1 inst_1021 ( .A(net_1020), .ZN(net_443) );
NOR2_X1 inst_473 ( .ZN(net_712), .A1(net_677), .A2(net_651) );
AND2_X4 inst_1131 ( .A1(net_673), .ZN(net_547), .A2(net_546) );
CLKBUF_X1 inst_1076 ( .Z(n480), .A(n2256) );
XNOR2_X1 inst_217 ( .ZN(net_793), .A(net_792), .B(net_791) );
NAND3_X1 inst_572 ( .A1(net_911), .ZN(net_651), .A3(net_617), .A2(net_604) );
NAND2_X1 inst_742 ( .ZN(net_426), .A2(net_271), .A1(net_112) );
NAND2_X1 inst_691 ( .ZN(net_298), .A2(net_142), .A1(net_36) );
AND3_X4 inst_1101 ( .ZN(net_519), .A3(net_518), .A2(net_480), .A1(net_407) );
NOR2_X1 inst_427 ( .ZN(net_250), .A2(net_175), .A1(n3723) );
XNOR2_X1 inst_257 ( .A(net_963), .ZN(net_940), .B(net_902) );
NOR2_X1 inst_485 ( .ZN(net_783), .A2(net_782), .A1(net_758) );
NAND2_X1 inst_770 ( .ZN(net_657), .A1(net_531), .A2(net_437) );
NAND3_X1 inst_565 ( .ZN(net_577), .A3(net_576), .A1(net_259), .A2(net_258) );
MUX2_X2 inst_861 ( .Z(net_315), .S(net_191), .B(net_17), .A(n2230) );
NAND2_X1 inst_672 ( .A2(net_191), .ZN(net_150), .A1(n147) );
XNOR2_X1 inst_138 ( .ZN(net_724), .A(net_342), .B(n2230) );
NAND2_X1 inst_622 ( .ZN(net_54), .A2(n234), .A1(n18) );
NOR2_X1 inst_409 ( .ZN(net_512), .A2(net_234), .A1(n3729) );
MUX2_X2 inst_899 ( .Z(net_944), .A(net_943), .B(net_942), .S(net_760) );
XOR2_X1 inst_33 ( .Z(net_291), .A(net_290), .B(net_289) );
NAND2_X1 inst_703 ( .ZN(net_321), .A2(net_151), .A1(net_67) );
OR2_X4 inst_312 ( .A1(net_191), .ZN(net_93), .A2(n3701) );
NAND2_X1 inst_660 ( .A2(net_191), .ZN(net_142), .A1(n97) );
INV_X1 inst_977 ( .A(net_326), .ZN(net_179) );
NOR2_X1 inst_517 ( .ZN(net_1023), .A2(net_1008), .A1(net_840) );
OR3_X4 inst_309 ( .ZN(net_895), .A1(net_894), .A2(net_893), .A3(net_892) );
XNOR2_X1 inst_232 ( .ZN(net_857), .A(net_856), .B(net_798) );
NOR4_X1 inst_347 ( .ZN(net_987), .A2(net_694), .A1(net_558), .A4(net_505), .A3(net_249) );
NAND2_X1 inst_768 ( .A1(net_435), .ZN(net_429), .A2(net_428) );
NAND2_X1 inst_663 ( .A2(net_191), .ZN(net_155), .A1(n26) );
XNOR2_X1 inst_297 ( .ZN(net_1035), .B(net_1027), .A(net_1022) );
NAND2_X1 inst_755 ( .ZN(net_1020), .A2(net_233), .A1(net_121) );
CLKBUF_X1 inst_1067 ( .Z(n522), .A(n4394) );
OR3_X2 inst_310 ( .ZN(net_410), .A1(net_409), .A2(net_335), .A3(net_315) );
INV_X1 inst_1043 ( .A(net_847), .ZN(net_834) );
XNOR2_X1 inst_253 ( .ZN(net_918), .B(net_905), .A(net_887) );
INV_X1 inst_971 ( .A(net_368), .ZN(net_242) );
XNOR2_X1 inst_162 ( .ZN(net_458), .B(net_371), .A(net_207) );
NAND3_X1 inst_589 ( .ZN(net_861), .A1(net_725), .A3(net_554), .A2(net_499) );
NAND2_X1 inst_794 ( .ZN(net_768), .A1(net_709), .A2(net_678) );
INV_X1 inst_1005 ( .ZN(net_511), .A(net_387) );
NAND2_X1 inst_602 ( .ZN(net_35), .A2(n231), .A1(n18) );
XOR2_X1 inst_59 ( .Z(net_400), .A(net_363), .B(net_362) );
XNOR2_X1 inst_135 ( .ZN(net_414), .A(net_274), .B(n3711) );
INV_X1 inst_996 ( .A(net_989), .ZN(net_503) );
XOR2_X1 inst_37 ( .Z(net_469), .B(net_310), .A(net_300) );
AND4_X1 inst_1098 ( .ZN(net_698), .A4(net_563), .A3(net_472), .A1(net_237), .A2(net_188) );
NAND2_X1 inst_740 ( .ZN(net_501), .A2(net_261), .A1(net_113) );
XNOR2_X1 inst_264 ( .ZN(net_964), .A(net_963), .B(net_918) );
XOR2_X1 inst_84 ( .B(net_963), .A(net_917), .Z(n368) );
INV_X1 inst_924 ( .ZN(net_3), .A(n2230) );
OR4_X1 inst_303 ( .ZN(net_836), .A2(net_835), .A4(net_823), .A1(net_756), .A3(net_755) );
XNOR2_X1 inst_173 ( .ZN(net_588), .B(net_397), .A(net_219) );
NAND2_X1 inst_723 ( .ZN(net_304), .A2(net_161), .A1(net_52) );
XNOR2_X1 inst_224 ( .ZN(net_838), .A(net_787), .B(net_626) );
NAND2_X1 inst_611 ( .ZN(net_44), .A2(n195), .A1(n18) );
XNOR2_X1 inst_287 ( .B(net_1031), .ZN(net_1021), .A(net_1006) );
NOR2_X1 inst_426 ( .ZN(net_590), .A2(net_181), .A1(n3705) );
NAND2_X1 inst_618 ( .ZN(net_51), .A2(n221), .A1(n18) );
NAND2_X1 inst_648 ( .ZN(net_79), .A2(n191), .A1(n18) );
CLKBUF_X1 inst_1088 ( .A(n469), .Z(n422) );
XNOR2_X1 inst_270 ( .B(net_971), .A(net_882), .ZN(n324) );
NOR2_X1 inst_474 ( .A2(net_729), .ZN(net_683), .A1(net_523) );
XOR2_X1 inst_26 ( .Z(net_279), .A(net_278), .B(net_277) );
NAND2_X1 inst_766 ( .A1(net_433), .ZN(net_423), .A2(net_422) );
NOR2_X1 inst_490 ( .ZN(net_815), .A1(net_814), .A2(net_765) );
INV_X1 inst_984 ( .A(net_329), .ZN(net_184) );
NAND2_X1 inst_801 ( .ZN(net_693), .A1(net_692), .A2(net_629) );
NAND2_X1 inst_626 ( .ZN(net_58), .A2(n193), .A1(n18) );
NAND2_X1 inst_692 ( .ZN(net_262), .A2(net_143), .A1(net_63) );
XOR2_X1 inst_70 ( .B(net_464), .A(net_462), .Z(net_459) );
XNOR2_X1 inst_129 ( .ZN(net_388), .A(net_368), .B(n2239) );
MUX2_X2 inst_870 ( .Z(net_301), .S(net_191), .A(net_21), .B(n55) );
XOR2_X1 inst_11 ( .B(net_364), .A(net_354), .Z(net_219) );
NAND2_X1 inst_631 ( .ZN(net_63), .A2(n223), .A1(n18) );
CLKBUF_X1 inst_1056 ( .Z(n544), .A(n3749) );
XNOR2_X1 inst_188 ( .ZN(net_704), .B(net_641), .A(net_447) );
NOR2_X1 inst_441 ( .ZN(net_488), .A2(net_418), .A1(net_385) );
NAND2_X1 inst_798 ( .ZN(net_689), .A2(net_632), .A1(net_623) );
NAND2_X1 inst_808 ( .ZN(net_719), .A2(net_650), .A1(n89) );
NAND3_X1 inst_557 ( .A1(net_572), .ZN(net_408), .A2(net_310), .A3(net_300) );
NAND2_X1 inst_777 ( .A1(net_747), .ZN(net_656), .A2(net_548) );
NOR2_X1 inst_398 ( .ZN(net_345), .A1(net_164), .A2(net_87) );
AND2_X4 inst_1128 ( .ZN(net_528), .A2(net_527), .A1(net_463) );
NOR2_X1 inst_436 ( .A1(net_1004), .A2(net_967), .ZN(net_611) );
INV_X1 inst_1037 ( .ZN(net_784), .A(net_761) );
NAND2_X1 inst_823 ( .ZN(net_817), .A2(net_759), .A1(net_698) );
INV_X1 inst_933 ( .ZN(net_9), .A(n2218) );
XNOR2_X1 inst_300 ( .B(net_1037), .A(net_978), .ZN(n338) );
XNOR2_X1 inst_102 ( .A(net_335), .ZN(net_316), .B(net_315) );
INV_X1 inst_1013 ( .A(net_673), .ZN(net_570) );
NOR2_X1 inst_446 ( .A2(net_1009), .A1(net_963), .ZN(net_548) );
NOR2_X1 inst_364 ( .A1(net_191), .ZN(net_88), .A2(n156) );
XNOR2_X1 inst_144 ( .ZN(net_395), .B(net_215), .A(net_213) );
XNOR2_X1 inst_195 ( .ZN(net_734), .B(net_733), .A(net_731) );
NAND2_X1 inst_824 ( .ZN(net_820), .A2(net_819), .A1(net_709) );
NOR2_X1 inst_411 ( .ZN(net_747), .A2(net_236), .A1(n4394) );
XNOR2_X1 inst_124 ( .ZN(net_911), .A(net_372), .B(n1462) );
MUX2_X2 inst_880 ( .Z(net_361), .S(net_191), .A(net_7), .B(n86) );
NAND2_X1 inst_680 ( .ZN(net_376), .A2(net_126), .A1(net_65) );
NAND2_X1 inst_785 ( .ZN(net_634), .A2(net_620), .A1(net_619) );
NAND2_X1 inst_737 ( .A1(net_336), .A2(net_220), .ZN(net_198) );
INV_X1 inst_961 ( .ZN(net_109), .A(n3711) );
MUX2_X2 inst_876 ( .Z(net_305), .S(net_191), .A(net_6), .B(n61) );
NAND4_X1 inst_545 ( .ZN(net_759), .A4(net_700), .A1(net_583), .A2(net_582), .A3(net_410) );
NOR2_X1 inst_399 ( .ZN(net_338), .A1(net_164), .A2(net_99) );
NAND4_X1 inst_527 ( .ZN(net_565), .A1(net_416), .A4(net_413), .A3(net_298), .A2(net_297) );
XNOR2_X1 inst_226 ( .ZN(net_841), .A(net_840), .B(net_777) );
NOR2_X1 inst_414 ( .ZN(net_464), .A2(net_242), .A1(n2239) );
XOR2_X1 inst_61 ( .A(net_373), .Z(net_370), .B(net_158) );
XNOR2_X1 inst_203 ( .ZN(net_748), .A(net_747), .B(net_746) );
NAND4_X1 inst_531 ( .ZN(net_579), .A4(net_578), .A1(net_561), .A2(net_281), .A3(net_280) );
NAND3_X1 inst_562 ( .ZN(net_482), .A3(net_412), .A2(net_302), .A1(net_301) );
XNOR2_X1 inst_212 ( .ZN(net_775), .B(net_727), .A(net_692) );
AND2_X4 inst_1139 ( .ZN(net_763), .A1(net_762), .A2(net_761) );
NOR2_X1 inst_499 ( .A2(net_904), .A1(net_889), .ZN(net_885) );
OR2_X4 inst_335 ( .ZN(net_901), .A2(net_894), .A1(net_892) );
NAND2_X1 inst_674 ( .A2(net_191), .ZN(net_143), .A1(n47) );
NOR2_X1 inst_466 ( .ZN(net_662), .A2(net_549), .A1(net_433) );
NAND2_X1 inst_658 ( .A2(net_191), .ZN(net_153), .A1(n118) );
INV_X1 inst_989 ( .ZN(net_404), .A(net_309) );
NOR2_X1 inst_456 ( .A1(net_1016), .ZN(net_523), .A2(net_522) );
NAND2_X1 inst_832 ( .A2(net_898), .ZN(net_897), .A1(net_591) );
XNOR2_X1 inst_275 ( .ZN(net_1000), .A(net_999), .B(net_964) );
XNOR2_X1 inst_117 ( .ZN(net_437), .A(net_317), .B(n2224) );
MUX2_X2 inst_858 ( .Z(net_354), .S(net_191), .A(net_108), .B(n87) );
NOR2_X1 inst_438 ( .ZN(net_549), .A1(net_486), .A2(net_485) );
AND2_X4 inst_1109 ( .ZN(net_335), .A2(net_160), .A1(net_30) );
NOR2_X1 inst_501 ( .ZN(net_896), .A2(net_868), .A1(net_670) );
NAND3_X1 inst_587 ( .ZN(net_865), .A3(net_695), .A1(net_431), .A2(net_201) );
CLKBUF_X1 inst_1081 ( .Z(n446), .A(n106) );
XNOR2_X1 inst_154 ( .ZN(net_448), .A(net_344), .B(net_334) );
NAND2_X1 inst_666 ( .A2(net_191), .ZN(net_161), .A1(n50) );
OR2_X4 inst_324 ( .A1(net_733), .A2(net_524), .ZN(net_521) );
NOR2_X1 inst_465 ( .ZN(net_797), .A1(net_556), .A2(net_495) );
XOR2_X1 inst_54 ( .Z(net_353), .A(net_352), .B(net_351) );
XNOR2_X1 inst_109 ( .ZN(net_409), .A(net_336), .B(net_220) );
NAND3_X1 inst_570 ( .A2(net_724), .ZN(net_647), .A1(net_615), .A3(net_595) );
NAND2_X1 inst_640 ( .ZN(net_72), .A2(n204), .A1(n18) );
XOR2_X1 inst_43 ( .A(net_379), .Z(net_313), .B(net_312) );
XNOR2_X1 inst_94 ( .ZN(net_229), .A(net_228), .B(net_119) );
AND2_X4 inst_1114 ( .A2(net_422), .ZN(net_402), .A1(net_401) );
NOR2_X1 inst_454 ( .A2(net_1012), .ZN(net_551), .A1(net_489) );
NOR2_X1 inst_375 ( .A1(net_191), .ZN(net_100), .A2(n168) );
INV_X1 inst_942 ( .ZN(net_128), .A(n38) );
MUX2_X2 inst_904 ( .S(net_962), .A(net_803), .B(net_800), .Z(n350) );
XNOR2_X1 inst_262 ( .B(net_1009), .A(net_908), .ZN(n365) );
XNOR2_X1 inst_243 ( .ZN(net_888), .A(net_838), .B(net_790) );
XNOR2_X1 inst_285 ( .A(net_996), .B(net_956), .ZN(n336) );
NOR2_X1 inst_424 ( .ZN(net_560), .A2(net_173), .A1(n1469) );
NAND3_X1 inst_591 ( .A1(net_931), .ZN(net_929), .A3(net_928), .A2(net_822) );
NOR2_X1 inst_497 ( .ZN(net_868), .A1(net_832), .A2(net_831) );
XOR2_X1 inst_15 ( .Z(net_251), .B(net_224), .A(net_133) );
NAND2_X1 inst_757 ( .ZN(net_630), .A1(net_406), .A2(net_404) );
OR2_X2 inst_343 ( .A2(net_938), .A1(net_848), .ZN(n252) );
INV_X1 inst_1035 ( .ZN(net_711), .A(net_710) );
AND3_X4 inst_1106 ( .A2(net_911), .ZN(net_605), .A3(net_604), .A1(net_442) );
OR2_X4 inst_337 ( .ZN(net_937), .A2(net_936), .A1(net_845) );
NAND4_X1 inst_543 ( .ZN(net_742), .A2(net_593), .A4(net_589), .A3(net_585), .A1(net_466) );
INV_X1 inst_929 ( .ZN(net_5), .A(n3723) );
INV_X1 inst_982 ( .A(net_328), .ZN(net_234) );
CLKBUF_X1 inst_1078 ( .Z(n453), .A(n1) );
NAND2_X1 inst_670 ( .A2(net_191), .ZN(net_132), .A1(n44) );
XNOR2_X1 inst_299 ( .B(net_1036), .A(net_982), .ZN(n399) );
INV_X1 inst_1034 ( .ZN(net_835), .A(net_708) );
NOR2_X1 inst_476 ( .A2(net_746), .ZN(net_715), .A1(net_542) );
NOR2_X1 inst_418 ( .ZN(net_246), .A2(net_170), .A1(n4437) );
MUX2_X2 inst_864 ( .Z(net_211), .S(net_191), .A(net_25), .B(n80) );
XOR2_X1 inst_86 ( .B(net_999), .A(net_976), .Z(n359) );
INV_X1 inst_949 ( .ZN(net_19), .A(n4394) );
XOR2_X1 inst_20 ( .Z(net_572), .B(net_264), .A(net_211) );
NAND2_X1 inst_613 ( .ZN(net_46), .A2(n18), .A1(n151) );
INV_X1 inst_1039 ( .A(net_889), .ZN(net_744) );
NAND2_X1 inst_714 ( .ZN(net_326), .A2(net_147), .A1(net_51) );
NOR4_X1 inst_349 ( .ZN(net_904), .A1(net_810), .A2(net_721), .A4(net_402), .A3(net_246) );
NOR2_X1 inst_483 ( .ZN(net_773), .A2(net_772), .A1(net_687) );
NAND3_X1 inst_576 ( .A2(net_751), .ZN(net_616), .A1(net_615), .A3(net_606) );
XNOR2_X1 inst_259 ( .A(net_939), .B(net_923), .ZN(n295) );
INV_X1 inst_1046 ( .A(net_923), .ZN(net_909) );
XNOR2_X1 inst_246 ( .B(net_905), .ZN(net_902), .A(net_857) );
INV_X1 inst_1020 ( .ZN(net_749), .A(net_422) );
CLKBUF_X1 inst_1061 ( .Z(n534), .A(n4410) );
NAND2_X1 inst_635 ( .ZN(net_67), .A2(n180), .A1(n18) );
NAND2_X1 inst_807 ( .ZN(net_717), .A2(net_716), .A1(net_520) );
NAND2_X1 inst_705 ( .ZN(net_333), .A2(net_150), .A1(net_46) );
XOR2_X1 inst_72 ( .Z(net_791), .B(net_571), .A(net_511) );
MUX2_X2 inst_911 ( .S(net_997), .B(net_884), .A(net_778), .Z(n298) );
INV_X1 inst_976 ( .A(net_349), .ZN(net_178) );
NAND4_X1 inst_519 ( .ZN(n406), .A4(n230), .A3(n218), .A1(n210), .A2(n152) );
MUX2_X2 inst_909 ( .S(net_997), .B(net_461), .A(net_459), .Z(n304) );
INV_X1 inst_1003 ( .ZN(net_726), .A(net_439) );
NAND3_X1 inst_582 ( .A1(net_696), .ZN(net_625), .A3(net_617), .A2(net_560) );
CLKBUF_X1 inst_1096 ( .Z(n2), .A(n1) );
NAND2_X1 inst_683 ( .ZN(net_133), .A2(net_132), .A1(net_49) );
NAND2_X1 inst_735 ( .A1(net_286), .A2(net_214), .ZN(net_195) );
CLKBUF_X1 inst_1053 ( .Z(n550), .A(n3729) );
XNOR2_X1 inst_115 ( .ZN(net_965), .A(net_318), .B(n2218) );
XNOR2_X1 inst_210 ( .ZN(net_853), .B(net_745), .A(net_714) );
MUX2_X2 inst_894 ( .S(net_852), .A(net_795), .B(net_792), .Z(n379) );
INV_X1 inst_994 ( .A(net_567), .ZN(net_385) );
NAND2_X1 inst_761 ( .ZN(net_525), .A2(net_428), .A1(net_387) );
XNOR2_X1 inst_239 ( .ZN(net_883), .B(net_882), .A(net_841) );
XNOR2_X1 inst_175 ( .ZN(net_635), .B(net_507), .A(net_255) );
NAND3_X1 inst_593 ( .ZN(net_933), .A1(net_914), .A3(net_901), .A2(net_816) );
NAND2_X1 inst_725 ( .ZN(net_224), .A2(net_146), .A1(net_61) );
NAND2_X1 inst_747 ( .ZN(net_499), .A2(net_342), .A1(net_3) );
NAND2_X1 inst_843 ( .ZN(net_958), .A2(net_933), .A1(net_669) );
NAND2_X1 inst_601 ( .ZN(net_34), .A2(n18), .A1(n161) );
XNOR2_X1 inst_133 ( .ZN(net_722), .A(net_261), .B(n4410) );
XNOR2_X1 inst_112 ( .ZN(net_415), .A(net_275), .B(n3705) );
MUX2_X2 inst_916 ( .Z(net_1037), .A(net_1033), .B(net_1021), .S(net_977) );
NAND2_X1 inst_764 ( .A2(net_965), .A1(net_603), .ZN(net_492) );
NOR2_X1 inst_479 ( .ZN(net_782), .A2(net_699), .A1(net_468) );
OR4_X1 inst_305 ( .A4(net_851), .ZN(n418), .A3(n410), .A2(n408), .A1(n406) );
AND2_X4 inst_1111 ( .A1(net_338), .A2(net_202), .ZN(net_187) );
XOR2_X1 inst_29 ( .Z(net_578), .A(net_284), .B(net_283) );
NAND2_X1 inst_771 ( .ZN(net_619), .A1(net_560), .A2(net_442) );
MUX2_X2 inst_878 ( .Z(net_199), .S(net_191), .A(net_13), .B(n63) );
XNOR2_X1 inst_126 ( .ZN(net_623), .A(net_271), .B(n3717) );
NOR2_X1 inst_480 ( .A2(net_761), .ZN(net_760), .A1(net_735) );
NAND4_X1 inst_538 ( .ZN(net_832), .A2(net_580), .A4(net_577), .A3(net_482), .A1(net_189) );
NAND3_X1 inst_564 ( .ZN(net_814), .A3(net_566), .A2(net_424), .A1(net_380) );
NAND2_X1 inst_646 ( .ZN(net_120), .A1(n4528), .A2(n1496) );
INV_X1 inst_963 ( .ZN(net_29), .A(n4427) );
AND2_X4 inst_1140 ( .ZN(net_831), .A2(net_786), .A1(net_600) );
NOR2_X1 inst_382 ( .A1(net_191), .ZN(net_106), .A2(n176) );
XOR2_X1 inst_35 ( .Z(net_296), .B(net_295), .A(net_152) );
NAND2_X1 inst_739 ( .ZN(net_493), .A2(net_274), .A1(net_109) );
INV_X1 inst_948 ( .ZN(net_117), .A(n2224) );
CLKBUF_X1 inst_1086 ( .Z(n436), .A(n1462) );
NOR2_X1 inst_358 ( .A1(net_191), .ZN(net_82), .A2(n209) );
XOR2_X1 inst_48 ( .B(net_362), .Z(net_339), .A(net_338) );
MUX2_X2 inst_907 ( .Z(net_982), .A(net_945), .B(net_944), .S(n4526) );
XOR2_X1 inst_46 ( .Z(net_330), .A(net_329), .B(net_328) );
INV_X1 inst_934 ( .ZN(net_10), .A(n114) );
INV_X1 inst_922 ( .ZN(net_1), .A(n3729) );
INV_X1 inst_1000 ( .A(net_485), .ZN(net_386) );
AND2_X4 inst_1126 ( .A1(net_533), .A2(net_463), .ZN(net_438) );
NOR2_X1 inst_443 ( .A1(net_1025), .A2(net_925), .ZN(net_598) );
NAND2_X1 inst_796 ( .ZN(net_682), .A2(net_681), .A1(net_521) );
NAND2_X1 inst_633 ( .ZN(net_65), .A2(n203), .A1(n18) );
NAND4_X1 inst_524 ( .A4(net_572), .ZN(net_470), .A2(net_469), .A3(net_308), .A1(net_307) );
NAND2_X1 inst_655 ( .A2(net_191), .ZN(net_137), .A1(n115) );
XNOR2_X1 inst_104 ( .ZN(net_322), .A(net_321), .B(net_320) );
NOR2_X1 inst_448 ( .A1(net_1009), .A2(net_999), .ZN(net_613) );
CLKBUF_X1 inst_1049 ( .Z(n558), .A(n3705) );
XNOR2_X1 inst_168 ( .ZN(net_515), .A(net_514), .B(net_511) );
MUX2_X2 inst_914 ( .A(net_1020), .B(net_1019), .S(net_1018), .Z(n273) );
NAND2_X1 inst_695 ( .ZN(net_278), .A2(net_145), .A1(net_66) );
NAND2_X1 inst_730 ( .A1(net_265), .A2(net_209), .ZN(net_189) );
NOR2_X1 inst_384 ( .ZN(net_368), .A1(net_164), .A2(net_88) );
NAND2_X1 inst_727 ( .ZN(net_331), .A2(net_153), .A1(net_42) );
MUX2_X2 inst_873 ( .Z(net_202), .S(net_191), .A(net_18), .B(n110) );
OR2_X4 inst_321 ( .A2(net_1025), .ZN(net_494), .A1(net_493) );
NAND2_X1 inst_653 ( .A2(net_191), .ZN(net_165), .A1(n124) );
INV_X1 inst_991 ( .A(net_747), .ZN(net_383) );
NAND2_X1 inst_608 ( .ZN(net_41), .A2(n197), .A1(n18) );
NAND2_X1 inst_834 ( .ZN(net_923), .A1(net_904), .A2(net_878) );
MUX2_X2 inst_882 ( .Z(net_266), .S(net_191), .A(net_28), .B(n65) );
XNOR2_X1 inst_170 ( .ZN(net_828), .A(net_536), .B(net_535) );
NAND3_X1 inst_580 ( .A1(net_724), .ZN(net_622), .A3(net_615), .A2(net_531) );
INV_X1 inst_966 ( .A(net_343), .ZN(net_171) );
NOR2_X1 inst_511 ( .ZN(net_975), .A2(net_974), .A1(net_751) );
XOR2_X1 inst_41 ( .Z(net_424), .B(net_312), .A(net_306) );
XNOR2_X1 inst_199 ( .ZN(net_739), .B(net_638), .A(net_253) );
NAND2_X1 inst_708 ( .ZN(net_274), .A2(net_155), .A1(net_50) );
XNOR2_X1 inst_152 ( .ZN(net_446), .B(net_332), .A(net_263) );
INV_X1 inst_953 ( .ZN(net_96), .A(n4528) );
CLKBUF_X1 inst_1071 ( .Z(n490), .A(n2230) );
AND4_X1 inst_1099 ( .ZN(net_669), .A1(net_569), .A2(net_568), .A4(net_567), .A3(net_225) );
NOR2_X1 inst_468 ( .ZN(net_776), .A1(net_560), .A2(net_496) );
INV_X1 inst_1011 ( .ZN(net_999), .A(net_389) );
NOR2_X1 inst_429 ( .ZN(net_430), .A2(net_176), .A1(n3743) );
NAND4_X1 inst_540 ( .ZN(net_892), .A4(net_698), .A2(net_645), .A3(net_644), .A1(net_268) );
NOR2_X1 inst_404 ( .ZN(net_348), .A1(net_164), .A2(net_94) );
INV_X1 inst_998 ( .ZN(net_1012), .A(net_437) );
XNOR2_X1 inst_89 ( .ZN(net_231), .A(net_120), .B(n38) );
NOR2_X1 inst_388 ( .A1(net_164), .ZN(net_134), .A2(net_105) );
XOR2_X1 inst_66 ( .Z(net_963), .B(net_277), .A(n4400) );
XOR2_X1 inst_7 ( .A(net_378), .B(net_306), .Z(net_213) );
NOR2_X1 inst_392 ( .ZN(net_352), .A1(net_164), .A2(net_90) );
XNOR2_X1 inst_182 ( .ZN(net_642), .B(net_448), .A(net_319) );
XNOR2_X1 inst_273 ( .B(net_997), .A(net_517), .ZN(n307) );
XNOR2_X1 inst_120 ( .ZN(net_428), .A(net_293), .B(n3749) );
XNOR2_X1 inst_294 ( .ZN(net_1032), .B(net_1025), .A(net_1015) );
NAND2_X1 inst_788 ( .ZN(net_663), .A2(net_662), .A1(net_419) );
NOR2_X1 inst_489 ( .A2(net_907), .ZN(net_810), .A1(net_676) );
INV_X1 inst_931 ( .ZN(net_7), .A(n2247) );
XNOR2_X1 inst_192 ( .ZN(net_727), .B(net_684), .A(net_630) );
NOR2_X1 inst_366 ( .A1(net_191), .ZN(net_90), .A2(n215) );
CLKBUF_X1 inst_1083 ( .Z(n442), .A(n1486) );
NAND3_X1 inst_567 ( .A3(net_645), .ZN(net_583), .A1(net_320), .A2(net_314) );
XNOR2_X1 inst_149 ( .ZN(net_407), .B(net_390), .A(net_168) );
XNOR2_X1 inst_193 ( .ZN(net_730), .A(net_729), .B(net_728) );
OR2_X4 inst_318 ( .A1(net_596), .A2(net_485), .ZN(net_419) );
NAND2_X1 inst_810 ( .ZN(net_725), .A1(net_724), .A2(net_667) );
AND2_X4 inst_1136 ( .A1(net_762), .ZN(net_753), .A2(net_679) );
XOR2_X1 inst_39 ( .Z(net_417), .A(net_305), .B(net_304) );
XNOR2_X1 inst_230 ( .ZN(net_854), .B(net_853), .A(net_793) );
MUX2_X2 inst_856 ( .Z(net_297), .S(net_191), .A(net_0), .B(n78) );

endmodule
