module s1494 (
v4,
v3,
CLR,
v5,
v1,
v0,
blif_clk_net,
v2,
v6,
blif_reset_net,
v13_D_7,
v13_D_15,
v13_D_11,
v13_D_23,
v13_D_17,
v13_D_9,
v13_D_22,
v13_D_20,
v13_D_19,
v13_D_12,
v13_D_18,
v13_D_8,
v13_D_21,
v13_D_6,
v13_D_13,
v13_D_10,
v13_D_24,
v13_D_14,
v13_D_16);

// Start PIs
input v4;
input v3;
input CLR;
input v5;
input v1;
input v0;
input blif_clk_net;
input v2;
input v6;
input blif_reset_net;

// Start POs
output v13_D_7;
output v13_D_15;
output v13_D_11;
output v13_D_23;
output v13_D_17;
output v13_D_9;
output v13_D_22;
output v13_D_20;
output v13_D_19;
output v13_D_12;
output v13_D_18;
output v13_D_8;
output v13_D_21;
output v13_D_6;
output v13_D_13;
output v13_D_10;
output v13_D_24;
output v13_D_14;
output v13_D_16;

// Start wires
wire net_568;
wire net_47;
wire net_416;
wire net_215;
wire net_54;
wire net_526;
wire net_429;
wire net_694;
wire net_557;
wire net_129;
wire net_648;
wire net_373;
wire net_119;
wire net_98;
wire net_739;
wire v13_D_19;
wire net_151;
wire net_356;
wire net_53;
wire net_452;
wire net_210;
wire net_545;
wire net_284;
wire net_168;
wire net_560;
wire net_774;
wire net_741;
wire net_477;
wire net_439;
wire net_385;
wire net_259;
wire net_269;
wire net_548;
wire net_469;
wire net_501;
wire net_187;
wire net_111;
wire net_727;
wire net_264;
wire net_90;
wire net_671;
wire net_225;
wire net_283;
wire net_636;
wire net_85;
wire net_263;
wire net_252;
wire net_124;
wire net_778;
wire net_343;
wire net_770;
wire net_404;
wire net_240;
wire net_160;
wire net_322;
wire net_511;
wire net_4;
wire net_420;
wire net_665;
wire net_447;
wire net_295;
wire net_410;
wire net_508;
wire net_390;
wire net_307;
wire net_35;
wire net_586;
wire net_344;
wire v6;
wire net_16;
wire net_703;
wire v13_D_20;
wire net_712;
wire net_239;
wire net_193;
wire net_257;
wire net_310;
wire net_233;
wire net_474;
wire net_120;
wire net_292;
wire net_201;
wire net_472;
wire net_109;
wire net_80;
wire net_65;
wire net_96;
wire net_484;
wire net_167;
wire net_207;
wire net_136;
wire net_651;
wire net_700;
wire net_682;
wire net_280;
wire net_126;
wire net_744;
wire net_495;
wire net_278;
wire net_34;
wire net_458;
wire net_108;
wire net_598;
wire net_685;
wire net_571;
wire net_63;
wire net_593;
wire net_617;
wire net_601;
wire net_274;
wire net_672;
wire net_777;
wire net_554;
wire net_425;
wire net_321;
wire net_287;
wire net_189;
wire v13_D_23;
wire net_490;
wire net_742;
wire net_720;
wire net_99;
wire net_46;
wire net_480;
wire net_216;
wire net_433;
wire net_584;
wire net_717;
wire net_544;
wire net_368;
wire net_224;
wire net_684;
wire net_632;
wire net_52;
wire net_538;
wire net_165;
wire net_608;
wire net_510;
wire net_370;
wire net_464;
wire net_366;
wire net_13;
wire net_413;
wire net_747;
wire net_446;
wire net_716;
wire net_114;
wire v13_D_10;
wire net_248;
wire net_384;
wire net_36;
wire net_198;
wire net_637;
wire net_253;
wire net_311;
wire net_276;
wire net_760;
wire net_494;
wire net_209;
wire net_3;
wire net_547;
wire net_634;
wire net_294;
wire net_154;
wire net_666;
wire net_507;
wire net_616;
wire net_371;
wire net_238;
wire net_529;
wire net_28;
wire net_704;
wire v13_D_24;
wire net_587;
wire net_485;
wire net_97;
wire net_192;
wire net_649;
wire net_503;
wire net_256;
wire net_460;
wire net_82;
wire net_650;
wire net_64;
wire net_457;
wire net_291;
wire net_735;
wire net_726;
wire net_772;
wire net_679;
wire net_121;
wire net_597;
wire net_200;
wire net_308;
wire net_75;
wire net_515;
wire net_743;
wire net_600;
wire net_396;
wire net_757;
wire net_701;
wire net_206;
wire net_195;
wire net_125;
wire net_397;
wire net_107;
wire net_166;
wire net_223;
wire net_715;
wire net_235;
wire v13_D_7;
wire net_530;
wire net_606;
wire net_623;
wire net_663;
wire net_603;
wire net_594;
wire net_320;
wire net_271;
wire net_23;
wire net_117;
wire net_74;
wire net_673;
wire net_642;
wire net_579;
wire net_401;
wire net_250;
wire net_205;
wire net_769;
wire net_699;
wire net_242;
wire net_312;
wire net_130;
wire net_572;
wire net_359;
wire net_440;
wire net_286;
wire net_147;
wire net_481;
wire net_369;
wire net_758;
wire net_470;
wire net_26;
wire net_403;
wire net_334;
wire blif_clk_net;
wire net_32;
wire net_430;
wire net_718;
wire net_365;
wire net_282;
wire net_645;
wire net_426;
wire net_380;
wire net_141;
wire net_780;
wire net_467;
wire v1;
wire net_83;
wire net_609;
wire net_541;
wire net_414;
wire net_372;
wire net_437;
wire net_528;
wire net_56;
wire net_566;
wire net_456;
wire net_155;
wire net_705;
wire net_335;
wire net_506;
wire net_181;
wire net_336;
wire net_624;
wire net_349;
wire net_39;
wire net_555;
wire net_245;
wire net_2;
wire v3;
wire net_9;
wire net_395;
wire net_331;
wire net_298;
wire net_493;
wire net_688;
wire net_697;
wire net_475;
wire net_563;
wire net_386;
wire net_641;
wire net_605;
wire net_277;
wire net_199;
wire net_502;
wire net_431;
wire net_89;
wire net_290;
wire net_680;
wire net_338;
wire net_721;
wire net_638;
wire v13_D_14;
wire net_243;
wire net_400;
wire net_759;
wire net_222;
wire net_602;
wire net_313;
wire net_152;
wire net_489;
wire net_714;
wire net_175;
wire net_657;
wire net_106;
wire net_683;
wire net_607;
wire net_258;
wire net_140;
wire net_740;
wire net_247;
wire net_329;
wire net_279;
wire net_148;
wire net_698;
wire v13_D_8;
wire net_419;
wire net_25;
wire v13_D_13;
wire net_70;
wire net_691;
wire net_251;
wire net_194;
wire net_730;
wire net_615;
wire net_478;
wire net_244;
wire net_664;
wire net_585;
wire net_441;
wire net_128;
wire net_596;
wire v5;
wire net_138;
wire net_749;
wire net_333;
wire net_639;
wire net_728;
wire net_549;
wire net_374;
wire net_719;
wire net_411;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_77;
wire net_214;
wire net_249;
wire net_20;
wire net_49;
wire net_518;
wire v4;
wire net_15;
wire net_57;
wire net_706;
wire net_71;
wire net_771;
wire net_156;
wire net_394;
wire net_92;
wire net_1;
wire net_112;
wire net_708;
wire net_139;
wire net_696;
wire net_551;
wire net_537;
wire net_332;
wire net_180;
wire net_409;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire net_492;
wire net_463;
wire net_656;
wire net_432;
wire net_88;
wire net_197;
wire net_513;
wire net_204;
wire net_766;
wire net_81;
wire net_232;
wire net_604;
wire net_163;
wire net_402;
wire net_67;
wire v13_D_9;
wire net_202;
wire net_268;
wire net_110;
wire net_722;
wire net_379;
wire net_459;
wire net_483;
wire net_48;
wire net_33;
wire net_8;
wire net_737;
wire net_203;
wire net_450;
wire net_289;
wire net_505;
wire net_621;
wire net_435;
wire net_176;
wire net_137;
wire net_296;
wire net_132;
wire net_613;
wire net_237;
wire net_105;
wire net_782;
wire net_614;
wire net_532;
wire net_12;
wire net_93;
wire net_578;
wire net_302;
wire net_569;
wire v13_D_16;
wire net_768;
wire net_127;
wire net_327;
wire net_357;
wire net_348;
wire net_753;
wire net_630;
wire net_76;
wire net_626;
wire net_101;
wire net_388;
wire net_326;
wire net_353;
wire net_707;
wire net_589;
wire net_519;
wire net_100;
wire net_412;
wire net_655;
wire net_686;
wire net_652;
wire net_536;
wire CLR;
wire net_455;
wire net_221;
wire net_115;
wire net_689;
wire v2;
wire net_751;
wire net_393;
wire net_442;
wire net_17;
wire net_319;
wire net_542;
wire net_453;
wire net_575;
wire net_595;
wire net_581;
wire net_378;
wire net_164;
wire net_408;
wire net_724;
wire net_731;
wire net_377;
wire net_87;
wire net_0;
wire net_288;
wire net_423;
wire net_658;
wire net_328;
wire net_734;
wire net_157;
wire net_540;
wire net_512;
wire net_42;
wire net_779;
wire net_662;
wire blif_reset_net;
wire net_50;
wire net_234;
wire net_38;
wire net_66;
wire net_466;
wire net_765;
wire net_675;
wire net_342;
wire net_612;
wire net_19;
wire net_738;
wire net_443;
wire net_504;
wire net_522;
wire net_270;
wire net_674;
wire net_183;
wire net_668;
wire net_618;
wire v13_D_6;
wire net_150;
wire net_303;
wire net_304;
wire net_352;
wire net_491;
wire net_644;
wire net_30;
wire net_681;
wire net_643;
wire net_783;
wire net_436;
wire net_24;
wire net_392;
wire net_622;
wire net_186;
wire net_118;
wire net_754;
wire net_421;
wire net_146;
wire net_764;
wire net_550;
wire net_122;
wire net_417;
wire net_7;
wire v0;
wire net_172;
wire net_428;
wire net_94;
wire net_246;
wire net_461;
wire net_767;
wire net_219;
wire net_640;
wire net_18;
wire net_309;
wire net_482;
wire net_659;
wire net_131;
wire net_196;
wire net_29;
wire net_775;
wire net_358;
wire net_142;
wire net_149;
wire net_752;
wire net_516;
wire net_654;
wire net_31;
wire net_387;
wire net_330;
wire net_535;
wire net_498;
wire net_158;
wire net_676;
wire net_41;
wire v13_D_15;
wire net_713;
wire net_577;
wire net_693;
wire net_360;
wire net_570;
wire net_525;
wire net_444;
wire net_213;
wire net_325;
wire net_729;
wire net_301;
wire net_260;
wire net_299;
wire net_438;
wire net_732;
wire net_580;
wire net_314;
wire net_182;
wire net_521;
wire net_60;
wire net_590;
wire net_337;
wire net_341;
wire net_267;
wire net_273;
wire net_424;
wire net_468;
wire net_58;
wire net_690;
wire net_576;
wire net_488;
wire net_73;
wire net_465;
wire net_86;
wire net_177;
wire net_523;
wire net_407;
wire net_476;
wire net_564;
wire net_382;
wire net_179;
wire net_725;
wire net_159;
wire net_61;
wire net_583;
wire net_449;
wire net_383;
wire net_62;
wire net_6;
wire net_553;
wire net_534;
wire net_217;
wire net_351;
wire v13_D_12;
wire net_733;
wire net_763;
wire net_427;
wire net_486;
wire net_135;
wire net_340;
wire net_265;
wire net_517;
wire net_628;
wire net_434;
wire net_406;
wire net_473;
wire net_220;
wire net_14;
wire net_633;
wire net_293;
wire net_324;
wire net_113;
wire net_710;
wire net_497;
wire net_454;
wire net_418;
wire net_462;
wire net_40;
wire net_69;
wire net_543;
wire net_709;
wire net_161;
wire net_625;
wire net_300;
wire net_339;
wire net_748;
wire net_677;
wire net_95;
wire net_173;
wire net_361;
wire net_78;
wire net_27;
wire net_317;
wire net_305;
wire v13_D_11;
wire net_514;
wire net_191;
wire net_261;
wire net_22;
wire net_376;
wire net_558;
wire net_354;
wire net_660;
wire net_524;
wire net_144;
wire net_102;
wire net_227;
wire net_59;
wire net_646;
wire net_363;
wire net_445;
wire net_573;
wire net_162;
wire net_776;
wire net_781;
wire net_44;
wire net_230;
wire net_653;
wire net_784;
wire net_520;
wire net_422;
wire net_134;
wire net_678;
wire net_546;
wire net_561;
wire net_567;
wire net_45;
wire net_381;
wire net_702;
wire net_591;
wire net_185;
wire v13_D_22;
wire net_746;
wire net_588;
wire v13_D_18;
wire net_272;
wire net_178;
wire net_667;
wire net_208;
wire net_236;
wire net_487;
wire net_212;
wire net_315;
wire net_762;
wire net_552;
wire net_695;
wire net_415;
wire net_116;
wire net_556;
wire net_347;
wire net_756;
wire net_91;
wire net_297;
wire net_346;
wire net_629;
wire net_55;
wire net_559;
wire net_635;
wire net_255;
wire net_266;
wire net_345;
wire net_104;
wire net_620;
wire net_448;
wire net_619;
wire net_72;
wire net_350;
wire net_229;
wire net_398;
wire net_627;
wire net_306;
wire net_687;
wire net_241;
wire net_5;
wire net_405;
wire net_500;
wire net_355;
wire net_184;
wire net_711;
wire net_599;
wire net_631;
wire net_11;
wire net_610;
wire net_723;
wire net_123;
wire net_527;
wire net_262;
wire net_362;
wire net_389;
wire net_68;
wire net_318;
wire net_451;
wire net_323;
wire net_750;
wire net_736;
wire net_275;
wire net_539;
wire net_399;
wire net_692;
wire net_153;
wire v13_D_17;
wire net_316;
wire net_218;
wire net_84;
wire net_670;
wire net_174;
wire net_611;
wire net_231;
wire net_562;
wire net_103;
wire net_375;
wire net_226;
wire net_364;
wire net_43;
wire v13_D_21;
wire net_10;
wire net_228;
wire net_592;
wire net_21;
wire net_647;
wire net_79;
wire net_143;
wire net_190;
wire net_773;
wire net_391;
wire net_533;
wire net_145;
wire net_285;
wire net_281;
wire net_669;
wire net_254;
wire net_37;
wire net_582;
wire net_188;
wire net_761;
wire net_496;
wire net_755;
wire net_509;
wire net_574;
wire net_479;
wire net_661;
wire net_211;
wire net_133;
wire net_745;

// Start cells
INV_X4 inst_537 ( .A(net_190), .ZN(net_10) );
INV_X4 inst_696 ( .A(net_429), .ZN(net_372) );
NAND2_X2 inst_481 ( .A1(net_638), .A2(net_627), .ZN(v13_D_10) );
INV_X4 inst_551 ( .ZN(net_193), .A(net_48) );
NAND2_X4 inst_228 ( .A2(net_758), .A1(net_706), .ZN(net_606) );
NOR2_X1 inst_125 ( .A2(net_615), .A1(net_446), .ZN(v13_D_18) );
NAND2_X1 inst_486 ( .A1(net_760), .ZN(net_15), .A2(net_0) );
INV_X8 inst_506 ( .ZN(net_57), .A(net_48) );
NAND2_X1 inst_495 ( .ZN(net_475), .A1(net_400), .A2(net_354) );
NAND2_X2 inst_353 ( .ZN(net_400), .A2(net_399), .A1(net_296) );
NAND2_X4 inst_207 ( .A2(net_737), .A1(net_736), .ZN(net_182) );
NAND3_X2 inst_159 ( .A1(net_718), .A3(net_393), .ZN(net_289), .A2(net_148) );
INV_X4 inst_707 ( .ZN(net_458), .A(net_376) );
AND2_X2 inst_779 ( .A1(net_504), .ZN(net_221), .A2(net_220) );
NAND2_X2 inst_395 ( .ZN(net_496), .A1(net_385), .A2(net_285) );
NAND4_X2 inst_134 ( .ZN(net_503), .A1(net_502), .A3(net_501), .A4(net_112), .A2(net_66) );
NAND2_X2 inst_244 ( .A2(net_760), .ZN(net_97), .A1(net_31) );
NAND2_X2 inst_333 ( .ZN(net_345), .A1(net_344), .A2(net_185) );
INV_X4 inst_712 ( .ZN(net_522), .A(net_479) );
NAND2_X2 inst_452 ( .ZN(net_610), .A2(net_582), .A1(net_414) );
INV_X4 inst_689 ( .ZN(net_429), .A(net_390) );
NAND2_X2 inst_430 ( .ZN(net_566), .A1(net_491), .A2(net_485) );
NAND4_X2 inst_131 ( .ZN(net_411), .A2(net_226), .A4(net_222), .A3(net_219), .A1(net_164) );
NAND2_X2 inst_406 ( .ZN(net_521), .A1(net_520), .A2(net_452) );
NAND2_X4 inst_214 ( .ZN(net_719), .A1(net_225), .A2(net_110) );
NAND2_X2 inst_462 ( .ZN(net_623), .A2(net_589), .A1(net_551) );
NAND3_X2 inst_160 ( .ZN(net_291), .A2(net_255), .A1(net_174), .A3(net_105) );
NAND2_X2 inst_328 ( .ZN(net_332), .A2(net_251), .A1(net_139) );
NOR2_X4 inst_47 ( .A1(net_760), .ZN(net_79), .A2(net_1) );
OR2_X2 inst_19 ( .ZN(net_325), .A1(net_324), .A2(net_294) );
INV_X4 inst_548 ( .A(net_760), .ZN(net_58) );
INV_X8 inst_515 ( .ZN(net_363), .A(net_78) );
OR2_X4 inst_8 ( .A1(net_762), .ZN(net_716), .A2(v0) );
AND2_X4 inst_772 ( .ZN(net_216), .A1(net_54), .A2(net_17) );
INV_X2 inst_728 ( .A(net_131), .ZN(net_90) );
DFFR_X2 inst_762 ( .QN(net_762), .RN(net_657), .D(net_653), .CK(net_766) );
NAND2_X2 inst_370 ( .ZN(net_442), .A2(net_313), .A1(net_211) );
INV_X4 inst_573 ( .ZN(net_725), .A(net_40) );
NOR2_X2 inst_100 ( .ZN(net_437), .A1(net_326), .A2(net_312) );
INV_X4 inst_642 ( .A(net_253), .ZN(net_240) );
NAND2_X2 inst_459 ( .ZN(net_620), .A2(net_597), .A1(net_186) );
NAND2_X2 inst_279 ( .A1(net_756), .ZN(net_336), .A2(net_131) );
NAND2_X2 inst_445 ( .ZN(net_595), .A1(net_594), .A2(net_537) );
INV_X4 inst_709 ( .ZN(net_575), .A(net_491) );
NOR2_X2 inst_93 ( .ZN(net_374), .A1(net_257), .A2(net_221) );
INV_X4 inst_700 ( .A(net_603), .ZN(net_416) );
NOR2_X2 inst_81 ( .A1(net_211), .ZN(net_203), .A2(net_10) );
INV_X4 inst_612 ( .ZN(net_119), .A(net_91) );
INV_X4 inst_606 ( .A(net_125), .ZN(net_116) );
NAND2_X2 inst_367 ( .ZN(net_439), .A1(net_299), .A2(net_235) );
INV_X4 inst_525 ( .ZN(net_46), .A(v0) );
NAND4_X2 inst_139 ( .ZN(net_619), .A2(net_586), .A4(net_543), .A3(net_448), .A1(net_223) );
INV_X4 inst_657 ( .ZN(net_412), .A(net_268) );
INV_X4 inst_559 ( .ZN(net_23), .A(net_22) );
INV_X4 inst_584 ( .ZN(net_78), .A(net_31) );
INV_X8 inst_521 ( .ZN(net_316), .A(net_233) );
CLKBUF_X2 inst_790 ( .A(net_770), .Z(net_771) );
NAND2_X2 inst_434 ( .ZN(net_574), .A2(net_513), .A1(net_341) );
NAND2_X2 inst_470 ( .ZN(net_632), .A2(net_612), .A1(net_577) );
INV_X2 inst_751 ( .ZN(net_319), .A(net_249) );
INV_X4 inst_535 ( .A(net_46), .ZN(net_8) );
NAND2_X2 inst_450 ( .ZN(net_607), .A2(net_574), .A1(net_544) );
INV_X2 inst_745 ( .ZN(net_235), .A(net_234) );
INV_X8 inst_520 ( .A(net_535), .ZN(net_314) );
NAND2_X2 inst_237 ( .A1(net_762), .A2(net_761), .ZN(net_29) );
NAND3_X4 inst_148 ( .ZN(net_636), .A3(net_606), .A1(net_536), .A2(net_444) );
INV_X4 inst_554 ( .ZN(net_131), .A(net_58) );
INV_X2 inst_733 ( .ZN(net_110), .A(net_109) );
NAND2_X2 inst_377 ( .ZN(net_465), .A1(net_394), .A2(net_342) );
NAND3_X2 inst_191 ( .A3(net_667), .A1(net_666), .ZN(net_650), .A2(net_529) );
NOR2_X4 inst_51 ( .ZN(net_94), .A2(net_50), .A1(net_31) );
NAND3_X4 inst_142 ( .ZN(net_751), .A2(net_675), .A1(net_674), .A3(net_36) );
NAND2_X2 inst_315 ( .ZN(net_277), .A2(net_200), .A1(net_10) );
NOR2_X2 inst_80 ( .A2(net_747), .A1(net_746), .ZN(net_198) );
NAND2_X4 inst_216 ( .A1(net_710), .ZN(net_691), .A2(net_190) );
NOR2_X2 inst_78 ( .A1(net_425), .ZN(net_173), .A2(net_104) );
NAND2_X2 inst_241 ( .A2(net_760), .ZN(net_77), .A1(net_48) );
NAND3_X2 inst_177 ( .ZN(net_534), .A2(net_501), .A1(net_450), .A3(net_431) );
CLKBUF_X2 inst_783 ( .A(blif_clk_net), .Z(net_764) );
NAND3_X2 inst_183 ( .A2(net_753), .A1(net_752), .ZN(net_682), .A3(net_664) );
NAND3_X2 inst_151 ( .ZN(net_259), .A1(net_135), .A2(net_58), .A3(net_22) );
NOR2_X2 inst_64 ( .ZN(net_24), .A1(net_12), .A2(v1) );
INV_X2 inst_743 ( .A(net_340), .ZN(net_181) );
NAND2_X2 inst_415 ( .A1(net_596), .ZN(net_537), .A2(net_490) );
INV_X4 inst_615 ( .ZN(net_162), .A(net_95) );
NAND2_X2 inst_393 ( .A1(net_526), .ZN(net_493), .A2(net_373) );
NOR2_X2 inst_107 ( .ZN(net_530), .A1(net_455), .A2(net_293) );
NOR2_X2 inst_92 ( .ZN(net_317), .A2(net_303), .A1(net_238) );
NAND2_X2 inst_345 ( .ZN(net_371), .A1(net_275), .A2(net_250) );
NAND2_X4 inst_223 ( .A1(net_748), .ZN(net_700), .A2(net_169) );
NAND2_X2 inst_402 ( .ZN(net_515), .A2(net_441), .A1(net_129) );
NAND2_X2 inst_340 ( .ZN(net_366), .A1(net_349), .A2(net_273) );
INV_X4 inst_643 ( .ZN(net_272), .A(net_157) );
INV_X4 inst_697 ( .ZN(net_550), .A(net_377) );
NAND2_X1 inst_494 ( .ZN(net_452), .A2(net_451), .A1(net_316) );
NAND2_X1 inst_487 ( .A2(net_135), .ZN(net_98), .A1(net_14) );
NAND2_X2 inst_329 ( .ZN(net_335), .A2(net_334), .A1(net_316) );
INV_X4 inst_574 ( .A(net_79), .ZN(net_49) );
NAND2_X2 inst_386 ( .ZN(net_482), .A1(net_481), .A2(net_338) );
NAND3_X2 inst_158 ( .ZN(net_288), .A2(net_287), .A1(net_156), .A3(net_150) );
NAND4_X2 inst_141 ( .A1(net_720), .ZN(net_633), .A3(net_583), .A4(net_467), .A2(net_330) );
NAND2_X4 inst_200 ( .A1(net_725), .ZN(net_118), .A2(net_79) );
INV_X8 inst_507 ( .ZN(net_106), .A(net_31) );
INV_X4 inst_571 ( .A(net_758), .ZN(net_600) );
NOR2_X4 inst_57 ( .ZN(net_150), .A2(net_70), .A1(net_31) );
NAND2_X2 inst_338 ( .ZN(net_361), .A2(net_207), .A1(net_70) );
INV_X4 inst_711 ( .ZN(net_492), .A(net_491) );
INV_X4 inst_552 ( .ZN(net_68), .A(net_55) );
INV_X4 inst_599 ( .A(net_393), .ZN(net_104) );
NAND2_X2 inst_417 ( .ZN(net_539), .A2(net_477), .A1(net_260) );
INV_X4 inst_671 ( .ZN(net_404), .A(net_242) );
INV_X4 inst_579 ( .ZN(net_136), .A(net_30) );
OR2_X2 inst_21 ( .ZN(net_337), .A2(net_336), .A1(net_151) );
NAND2_X2 inst_469 ( .ZN(net_630), .A2(net_610), .A1(net_474) );
NAND2_X2 inst_281 ( .A2(net_245), .ZN(net_195), .A1(net_178) );
INV_X4 inst_585 ( .ZN(net_393), .A(net_84) );
INV_X4 inst_698 ( .ZN(net_489), .A(net_378) );
OR2_X2 inst_18 ( .A2(net_758), .A1(net_544), .ZN(net_307) );
INV_X4 inst_541 ( .ZN(net_542), .A(net_287) );
NAND2_X2 inst_410 ( .ZN(net_527), .A1(net_526), .A2(net_418) );
NAND2_X4 inst_208 ( .ZN(net_740), .A2(net_131), .A1(net_124) );
NOR2_X2 inst_88 ( .A1(net_347), .ZN(net_310), .A2(net_139) );
NAND2_X2 inst_316 ( .ZN(net_278), .A2(net_191), .A1(net_49) );
NAND2_X4 inst_220 ( .A1(net_729), .ZN(net_445), .A2(net_106) );
OR2_X4 inst_9 ( .ZN(net_586), .A1(net_44), .A2(v4) );
NOR2_X2 inst_113 ( .ZN(net_590), .A2(net_561), .A1(net_481) );
INV_X8 inst_505 ( .A(net_761), .ZN(net_48) );
NAND2_X2 inst_356 ( .ZN(net_407), .A2(net_291), .A1(net_126) );
NAND2_X2 inst_383 ( .ZN(net_471), .A2(net_398), .A1(net_114) );
NAND2_X2 inst_360 ( .ZN(net_418), .A2(net_397), .A1(net_381) );
AND2_X4 inst_773 ( .A1(net_762), .ZN(net_747), .A2(net_31) );
NAND2_X4 inst_198 ( .ZN(net_81), .A2(net_50), .A1(net_17) );
NOR2_X4 inst_50 ( .A1(net_193), .ZN(net_178), .A2(net_2) );
NAND2_X2 inst_245 ( .ZN(net_60), .A2(net_26), .A1(net_17) );
INV_X4 inst_569 ( .A(net_303), .ZN(net_37) );
INV_X4 inst_678 ( .ZN(net_385), .A(net_314) );
INV_X4 inst_624 ( .ZN(net_321), .A(net_281) );
NAND2_X2 inst_260 ( .A2(net_718), .A1(net_716), .ZN(net_707) );
CLKBUF_X2 inst_784 ( .A(net_764), .Z(net_765) );
INV_X2 inst_721 ( .ZN(net_28), .A(net_17) );
NAND3_X4 inst_147 ( .ZN(net_631), .A3(net_601), .A1(net_591), .A2(net_493) );
INV_X2 inst_744 ( .A(net_643), .ZN(net_186) );
NAND2_X2 inst_313 ( .ZN(net_275), .A2(net_274), .A1(net_237) );
NAND2_X2 inst_293 ( .A2(net_297), .ZN(net_219), .A1(net_206) );
AND2_X2 inst_778 ( .A2(net_211), .ZN(net_204), .A1(net_115) );
INV_X4 inst_636 ( .ZN(net_149), .A(net_148) );
INV_X4 inst_632 ( .ZN(net_197), .A(net_127) );
INV_X4 inst_549 ( .ZN(net_53), .A(net_48) );
NAND2_X2 inst_234 ( .A1(net_762), .ZN(net_40), .A2(net_17) );
XNOR2_X2 inst_0 ( .ZN(net_495), .A(net_316), .B(net_84) );
INV_X8 inst_522 ( .A(net_520), .ZN(net_456) );
NAND3_X2 inst_184 ( .ZN(net_706), .A3(net_669), .A1(net_668), .A2(net_478) );
INV_X4 inst_690 ( .ZN(net_402), .A(net_316) );
NAND2_X2 inst_236 ( .A2(net_287), .A1(net_54), .ZN(net_20) );
NAND2_X2 inst_433 ( .ZN(net_570), .A1(net_569), .A2(net_531) );
INV_X4 inst_553 ( .ZN(net_56), .A(net_22) );
NAND2_X2 inst_478 ( .ZN(net_645), .A1(net_643), .A2(net_626) );
NOR2_X2 inst_65 ( .A2(net_762), .ZN(net_27), .A1(net_4) );
INV_X4 inst_536 ( .A(net_54), .ZN(net_50) );
NAND2_X2 inst_242 ( .ZN(net_82), .A1(net_55), .A2(net_53) );
INV_X4 inst_688 ( .ZN(net_426), .A(net_306) );
AND2_X2 inst_781 ( .A1(net_451), .ZN(net_422), .A2(net_333) );
INV_X2 inst_732 ( .ZN(net_108), .A(net_107) );
INV_X8 inst_516 ( .ZN(net_686), .A(net_118) );
NOR2_X2 inst_98 ( .ZN(net_433), .A2(net_317), .A1(net_314) );
NAND2_X2 inst_263 ( .ZN(net_140), .A1(net_77), .A2(net_16) );
NAND3_X2 inst_190 ( .A1(net_645), .A3(net_635), .A2(net_599), .ZN(v13_D_24) );
NAND3_X2 inst_185 ( .ZN(net_599), .A1(net_562), .A3(net_443), .A2(net_34) );
OR2_X4 inst_13 ( .ZN(net_401), .A1(net_390), .A2(net_274) );
NOR2_X2 inst_75 ( .A1(net_762), .ZN(net_156), .A2(net_131) );
NAND2_X2 inst_332 ( .A2(net_346), .ZN(net_343), .A1(net_211) );
NAND3_X2 inst_166 ( .A2(net_751), .A1(net_750), .A3(net_698), .ZN(net_384) );
NOR2_X2 inst_116 ( .ZN(net_624), .A2(net_590), .A1(net_405) );
INV_X4 inst_598 ( .A(net_102), .ZN(net_76) );
NAND2_X2 inst_416 ( .ZN(net_538), .A2(net_487), .A1(net_385) );
NAND3_X2 inst_163 ( .A1(net_745), .ZN(net_376), .A2(net_102), .A3(net_31) );
NAND2_X2 inst_471 ( .ZN(net_635), .A2(net_623), .A1(net_603) );
NAND2_X2 inst_394 ( .ZN(net_494), .A2(net_380), .A1(v4) );
NOR2_X2 inst_79 ( .A1(net_730), .ZN(net_234), .A2(net_127) );
CLKBUF_X2 inst_799 ( .A(net_779), .Z(net_780) );
NOR2_X2 inst_106 ( .A2(net_697), .A1(net_696), .ZN(net_689) );
INV_X2 inst_738 ( .ZN(net_146), .A(net_145) );
NAND2_X2 inst_422 ( .ZN(net_553), .A1(net_552), .A2(net_466) );
NAND2_X4 inst_219 ( .A1(net_722), .ZN(net_396), .A2(net_106) );
INV_X2 inst_719 ( .A(net_760), .ZN(net_9) );
NAND2_X4 inst_201 ( .A2(net_542), .A1(net_161), .ZN(net_88) );
INV_X4 inst_605 ( .ZN(net_737), .A(net_82) );
NAND2_X2 inst_304 ( .A1(net_526), .ZN(net_462), .A2(net_255) );
INV_X2 inst_752 ( .A(net_446), .ZN(net_380) );
INV_X4 inst_542 ( .A(net_10), .ZN(net_7) );
NAND2_X2 inst_255 ( .A2(net_758), .ZN(net_114), .A1(net_113) );
NAND2_X2 inst_453 ( .ZN(net_612), .A1(net_611), .A2(net_585) );
NAND4_X2 inst_128 ( .A2(net_499), .A1(net_303), .ZN(net_282), .A4(net_281), .A3(net_253) );
NOR2_X2 inst_73 ( .ZN(net_746), .A1(net_287), .A2(net_128) );
NAND2_X1 inst_493 ( .A2(net_354), .ZN(net_309), .A1(net_308) );
NAND2_X2 inst_378 ( .A1(net_510), .ZN(net_466), .A2(net_170) );
OR2_X2 inst_23 ( .ZN(net_352), .A1(net_347), .A2(net_204) );
NAND2_X2 inst_339 ( .ZN(net_365), .A1(net_364), .A2(net_209) );
NAND2_X2 inst_351 ( .ZN(net_392), .A1(net_391), .A2(net_281) );
NAND2_X2 inst_361 ( .ZN(net_420), .A1(net_419), .A2(net_332) );
NAND2_X2 inst_408 ( .A1(net_542), .ZN(net_523), .A2(net_415) );
NAND2_X2 inst_325 ( .ZN(net_327), .A1(net_326), .A2(net_324) );
NAND2_X2 inst_461 ( .A2(net_758), .A1(net_711), .ZN(net_662) );
NAND2_X2 inst_385 ( .ZN(net_480), .A1(net_456), .A2(net_322) );
NAND2_X4 inst_197 ( .ZN(net_99), .A2(net_42), .A1(net_21) );
INV_X4 inst_659 ( .ZN(net_242), .A(net_240) );
NAND2_X2 inst_250 ( .A2(net_274), .ZN(net_92), .A1(net_28) );
NAND3_X2 inst_179 ( .ZN(net_549), .A2(net_457), .A3(net_451), .A1(net_309) );
OR2_X2 inst_24 ( .ZN(net_490), .A1(net_489), .A2(net_408) );
NOR2_X2 inst_114 ( .ZN(net_608), .A2(net_580), .A1(net_547) );
CLKBUF_X2 inst_786 ( .A(net_765), .Z(net_767) );
INV_X4 inst_617 ( .ZN(net_100), .A(net_99) );
NOR2_X2 inst_76 ( .ZN(net_399), .A2(net_134), .A1(net_131) );
NAND2_X2 inst_397 ( .ZN(net_506), .A2(net_473), .A1(net_306) );
INV_X8 inst_504 ( .ZN(net_17), .A(net_5) );
NAND3_X2 inst_150 ( .A3(net_761), .ZN(net_33), .A2(net_32), .A1(net_12) );
NAND3_X2 inst_172 ( .ZN(net_434), .A2(net_393), .A3(net_262), .A1(net_89) );
NAND2_X2 inst_362 ( .ZN(net_421), .A2(net_345), .A1(net_301) );
NAND2_X2 inst_277 ( .ZN(net_710), .A2(net_92), .A1(net_60) );
NOR2_X2 inst_83 ( .ZN(net_254), .A2(net_253), .A1(net_139) );
NOR2_X2 inst_121 ( .A1(net_690), .A2(net_654), .ZN(net_653) );
INV_X4 inst_534 ( .ZN(net_134), .A(net_54) );
NAND2_X2 inst_440 ( .ZN(net_585), .A1(net_533), .A2(net_523) );
NAND2_X2 inst_306 ( .ZN(net_735), .A2(net_259), .A1(net_155) );
OR3_X2 inst_2 ( .A1(net_368), .ZN(net_228), .A3(net_227), .A2(net_36) );
INV_X4 inst_644 ( .A(net_388), .ZN(net_265) );
INV_X4 inst_596 ( .ZN(net_425), .A(net_75) );
INV_X4 inst_578 ( .ZN(net_210), .A(net_52) );
NOR2_X4 inst_52 ( .ZN(net_176), .A2(net_93), .A1(net_31) );
NOR2_X2 inst_90 ( .A2(net_600), .A1(net_314), .ZN(net_312) );
NAND2_X2 inst_267 ( .ZN(net_155), .A2(net_154), .A1(net_96) );
NAND4_X2 inst_140 ( .ZN(net_621), .A1(net_584), .A3(net_558), .A4(net_519), .A2(net_483) );
INV_X4 inst_668 ( .ZN(net_238), .A(net_237) );
NAND2_X4 inst_221 ( .A1(net_708), .ZN(net_658), .A2(net_134) );
INV_X2 inst_748 ( .ZN(net_280), .A(net_279) );
INV_X2 inst_716 ( .ZN(net_0), .A(v3) );
INV_X4 inst_556 ( .ZN(net_303), .A(net_18) );
INV_X4 inst_650 ( .A(net_643), .ZN(net_594) );
INV_X4 inst_637 ( .ZN(net_196), .A(net_132) );
NAND2_X2 inst_289 ( .ZN(net_596), .A2(net_274), .A1(net_132) );
CLKBUF_X2 inst_792 ( .A(net_772), .Z(net_773) );
INV_X4 inst_547 ( .ZN(net_14), .A(net_13) );
INV_X4 inst_530 ( .ZN(net_190), .A(v3) );
INV_X2 inst_720 ( .ZN(net_62), .A(net_24) );
NAND2_X2 inst_432 ( .ZN(net_568), .A2(net_527), .A1(net_506) );
INV_X4 inst_679 ( .ZN(net_358), .A(net_341) );
NAND2_X2 inst_420 ( .ZN(net_551), .A1(net_550), .A2(net_495) );
NAND2_X2 inst_282 ( .A1(net_707), .ZN(net_705), .A2(net_197) );
NAND2_X2 inst_368 ( .ZN(net_440), .A1(net_316), .A2(net_184) );
INV_X8 inst_513 ( .ZN(net_124), .A(net_69) );
CLKBUF_X2 inst_803 ( .A(net_783), .Z(net_784) );
INV_X2 inst_754 ( .A(net_572), .ZN(net_469) );
AND2_X4 inst_769 ( .A2(net_761), .A1(net_759), .ZN(net_274) );
NOR3_X2 inst_44 ( .A1(net_494), .A3(net_374), .A2(net_67), .ZN(v13_D_15) );
NAND2_X2 inst_274 ( .ZN(net_177), .A2(net_176), .A1(net_59) );
NAND3_X2 inst_174 ( .A3(net_727), .A2(net_726), .ZN(net_680), .A1(net_288) );
NAND2_X2 inst_371 ( .ZN(net_444), .A2(net_443), .A1(net_378) );
INV_X4 inst_701 ( .ZN(net_755), .A(net_369) );
INV_X4 inst_662 ( .ZN(net_263), .A(net_209) );
NAND2_X2 inst_314 ( .A1(net_526), .ZN(net_276), .A2(net_216) );
NAND2_X2 inst_435 ( .ZN(net_576), .A1(net_575), .A2(net_516) );
NAND3_X2 inst_164 ( .ZN(net_382), .A3(net_381), .A1(net_362), .A2(net_210) );
OR2_X4 inst_5 ( .ZN(net_451), .A1(net_3), .A2(v4) );
INV_X4 inst_597 ( .ZN(net_674), .A(net_102) );
INV_X2 inst_729 ( .ZN(net_730), .A(net_95) );
NAND3_X2 inst_157 ( .ZN(net_249), .A3(net_248), .A1(net_121), .A2(net_56) );
INV_X4 inst_687 ( .ZN(net_520), .A(net_435) );
AND2_X4 inst_774 ( .A1(net_758), .ZN(net_340), .A2(net_31) );
INV_X4 inst_621 ( .ZN(net_388), .A(net_103) );
NOR2_X2 inst_68 ( .ZN(net_121), .A2(net_58), .A1(net_17) );
NAND2_X4 inst_213 ( .ZN(net_544), .A1(net_157), .A2(net_132) );
INV_X4 inst_604 ( .ZN(net_168), .A(net_142) );
NOR2_X4 inst_53 ( .A2(net_760), .ZN(net_225), .A1(net_87) );
INV_X4 inst_628 ( .ZN(net_148), .A(net_119) );
INV_X2 inst_753 ( .ZN(net_398), .A(net_397) );
NAND2_X4 inst_205 ( .ZN(net_138), .A2(net_137), .A1(net_136) );
NAND2_X2 inst_472 ( .A1(net_643), .ZN(net_637), .A2(net_621) );
NAND2_X2 inst_447 ( .ZN(net_695), .A2(net_563), .A1(net_548) );
NAND2_X2 inst_380 ( .ZN(net_467), .A2(net_401), .A1(net_358) );
NAND2_X2 inst_457 ( .A2(net_571), .A1(net_500), .ZN(v13_D_19) );
INV_X4 inst_651 ( .A(net_643), .ZN(net_183) );
INV_X4 inst_665 ( .ZN(net_347), .A(net_237) );
NAND2_X2 inst_292 ( .A2(net_542), .ZN(net_218), .A1(net_160) );
NAND2_X2 inst_379 ( .ZN(net_757), .A2(net_407), .A1(net_212) );
NAND4_X2 inst_127 ( .ZN(net_727), .A2(net_287), .A4(net_161), .A1(net_70), .A3(net_31) );
NAND3_X2 inst_186 ( .ZN(net_618), .A2(net_556), .A3(net_534), .A1(net_366) );
OR2_X2 inst_17 ( .A2(net_762), .ZN(net_756), .A1(net_178) );
INV_X4 inst_706 ( .ZN(net_457), .A(net_456) );
INV_X1 inst_759 ( .A(net_546), .ZN(net_508) );
NAND2_X2 inst_413 ( .ZN(net_532), .A2(net_423), .A1(net_419) );
NAND3_X4 inst_146 ( .ZN(net_541), .A3(net_445), .A2(net_410), .A1(net_396) );
NAND2_X2 inst_249 ( .ZN(net_736), .A1(net_704), .A2(net_84) );
NAND2_X2 inst_334 ( .ZN(net_449), .A1(net_347), .A2(net_346) );
NAND3_X2 inst_187 ( .ZN(net_723), .A3(net_663), .A1(net_662), .A2(net_282) );
NAND2_X4 inst_206 ( .ZN(net_175), .A1(net_76), .A2(net_31) );
NOR2_X2 inst_122 ( .A1(net_714), .ZN(net_655), .A2(net_654) );
OR2_X2 inst_25 ( .A1(net_758), .ZN(net_511), .A2(net_510) );
NAND2_X2 inst_354 ( .ZN(net_403), .A2(net_399), .A1(net_290) );
NAND2_X2 inst_405 ( .ZN(net_519), .A1(net_502), .A2(net_432) );
NAND2_X1 inst_492 ( .A1(net_542), .ZN(net_208), .A2(net_152) );
NAND2_X2 inst_240 ( .ZN(net_47), .A1(net_46), .A2(net_36) );
NAND2_X2 inst_326 ( .A2(net_526), .ZN(net_329), .A1(net_211) );
NOR2_X2 inst_110 ( .ZN(net_580), .A1(net_578), .A2(net_517) );
INV_X8 inst_518 ( .ZN(net_297), .A(net_124) );
NOR2_X2 inst_74 ( .A2(net_762), .A1(net_346), .ZN(net_130) );
NAND2_X2 inst_288 ( .ZN(net_212), .A1(net_211), .A2(net_210) );
NAND2_X2 inst_396 ( .A1(net_502), .ZN(net_497), .A2(net_379) );
NAND2_X4 inst_229 ( .ZN(net_744), .A1(net_715), .A2(net_600) );
NOR2_X2 inst_99 ( .ZN(net_436), .A1(net_435), .A2(net_310) );
NOR2_X2 inst_69 ( .A1(net_760), .ZN(net_294), .A2(net_55) );
NAND2_X2 inst_373 ( .A1(net_502), .ZN(net_448), .A2(net_336) );
NOR2_X2 inst_82 ( .A1(net_287), .ZN(net_239), .A2(net_167) );
INV_X4 inst_669 ( .ZN(net_391), .A(net_211) );
NOR2_X2 inst_108 ( .ZN(net_555), .A2(net_505), .A1(net_173) );
INV_X4 inst_664 ( .ZN(net_304), .A(net_215) );
INV_X4 inst_595 ( .A(net_453), .ZN(net_74) );
NAND2_X2 inst_283 ( .ZN(net_199), .A1(net_193), .A2(net_133) );
OR2_X2 inst_22 ( .ZN(net_339), .A2(net_338), .A1(net_227) );
NAND2_X2 inst_311 ( .ZN(net_271), .A2(net_188), .A1(net_7) );
NAND2_X2 inst_460 ( .ZN(net_622), .A2(net_604), .A1(net_565) );
NAND2_X2 inst_372 ( .ZN(net_447), .A2(net_446), .A1(net_128) );
NAND3_X2 inst_169 ( .A2(net_545), .ZN(net_427), .A1(net_426), .A3(net_425) );
NAND2_X4 inst_215 ( .ZN(net_731), .A1(net_665), .A2(net_99) );
NAND2_X2 inst_307 ( .ZN(net_261), .A2(net_260), .A1(net_240) );
AND3_X2 inst_767 ( .A2(net_564), .A3(net_542), .ZN(net_505), .A1(net_504) );
INV_X4 inst_638 ( .ZN(net_202), .A(net_150) );
NAND2_X2 inst_421 ( .ZN(net_667), .A1(net_526), .A2(net_509) );
NAND3_X2 inst_161 ( .ZN(net_664), .A1(net_375), .A3(net_213), .A2(net_137) );
INV_X4 inst_560 ( .A(net_137), .ZN(net_45) );
INV_X2 inst_749 ( .ZN(net_454), .A(net_431) );
INV_X4 inst_586 ( .ZN(net_229), .A(net_59) );
INV_X4 inst_702 ( .ZN(net_572), .A(net_456) );
INV_X4 inst_555 ( .ZN(net_375), .A(net_18) );
OR2_X2 inst_16 ( .ZN(net_128), .A1(net_68), .A2(net_31) );
INV_X2 inst_717 ( .ZN(net_12), .A(v6) );
NAND2_X2 inst_276 ( .ZN(net_185), .A1(net_184), .A2(net_101) );
INV_X2 inst_718 ( .ZN(net_3), .A(v5) );
NAND2_X2 inst_431 ( .ZN(net_567), .A2(net_532), .A1(net_402) );
NAND2_X2 inst_348 ( .A1(net_431), .ZN(net_379), .A2(net_280) );
OR3_X2 inst_3 ( .ZN(net_663), .A1(net_292), .A3(net_153), .A2(net_18) );
NAND3_X2 inst_156 ( .A2(net_762), .ZN(net_247), .A3(net_246), .A1(net_245) );
INV_X4 inst_577 ( .A(net_406), .ZN(net_91) );
CLKBUF_X2 inst_802 ( .A(net_782), .Z(net_783) );
INV_X4 inst_566 ( .ZN(net_206), .A(net_131) );
NAND2_X2 inst_296 ( .ZN(net_226), .A2(net_111), .A1(net_73) );
NOR2_X2 inst_91 ( .ZN(net_378), .A2(net_368), .A1(net_316) );
NAND4_X2 inst_132 ( .A2(net_721), .ZN(net_498), .A1(net_462), .A4(net_348), .A3(net_271) );
NAND2_X2 inst_342 ( .A1(net_735), .ZN(net_369), .A2(net_368) );
INV_X4 inst_526 ( .ZN(net_137), .A(v1) );
NOR3_X2 inst_36 ( .ZN(net_293), .A1(net_292), .A2(net_284), .A3(net_51) );
INV_X4 inst_656 ( .ZN(net_341), .A(net_139) );
INV_X4 inst_645 ( .ZN(net_233), .A(net_160) );
NAND2_X2 inst_463 ( .A2(net_592), .A1(net_424), .ZN(v13_D_22) );
INV_X8 inst_503 ( .ZN(net_31), .A(net_1) );
NOR2_X2 inst_96 ( .ZN(net_405), .A1(net_404), .A2(net_272) );
NOR3_X2 inst_45 ( .A2(net_594), .A3(net_555), .A1(net_460), .ZN(v13_D_21) );
NAND2_X2 inst_451 ( .ZN(net_609), .A2(net_579), .A1(net_549) );
NOR2_X2 inst_101 ( .ZN(net_472), .A2(net_395), .A1(net_350) );
NAND2_X2 inst_319 ( .ZN(net_377), .A2(net_211), .A1(net_11) );
NAND2_X2 inst_269 ( .ZN(net_163), .A1(net_162), .A2(net_161) );
NAND2_X2 inst_458 ( .A2(net_758), .A1(net_695), .ZN(net_688) );
NAND2_X2 inst_444 ( .ZN(net_593), .A2(net_566), .A1(net_550) );
NAND2_X2 inst_400 ( .ZN(net_512), .A2(net_439), .A1(net_263) );
CLKBUF_X2 inst_797 ( .A(net_777), .Z(net_778) );
INV_X4 inst_614 ( .ZN(net_107), .A(net_94) );
INV_X4 inst_686 ( .A(net_552), .ZN(net_300) );
INV_X4 inst_649 ( .ZN(net_174), .A(net_130) );
INV_X2 inst_741 ( .A(net_363), .ZN(net_158) );
NAND2_X2 inst_261 ( .ZN(net_703), .A2(net_125), .A1(net_6) );
INV_X8 inst_514 ( .ZN(net_255), .A(net_102) );
MUX2_X1 inst_500 ( .S(net_613), .A(net_609), .B(net_568), .Z(v13_D_7) );
INV_X8 inst_510 ( .ZN(net_93), .A(net_17) );
NAND2_X2 inst_268 ( .ZN(net_159), .A2(net_120), .A1(net_79) );
INV_X4 inst_685 ( .ZN(net_564), .A(net_552) );
NAND2_X2 inst_369 ( .ZN(net_441), .A1(net_360), .A2(net_298) );
INV_X4 inst_550 ( .ZN(net_44), .A(net_14) );
NOR2_X4 inst_63 ( .ZN(net_701), .A1(net_639), .A2(net_631) );
NOR2_X2 inst_119 ( .A1(net_709), .A2(net_654), .ZN(net_651) );
INV_X4 inst_603 ( .ZN(net_169), .A(net_81) );
NAND2_X2 inst_327 ( .A1(net_431), .ZN(net_331), .A2(net_330) );
INV_X4 inst_676 ( .A(net_316), .ZN(net_286) );
NOR2_X2 inst_85 ( .ZN(net_267), .A2(net_265), .A1(net_86) );
NAND2_X2 inst_291 ( .A1(net_762), .ZN(net_569), .A2(net_189) );
NAND2_X2 inst_266 ( .A2(net_758), .ZN(net_292), .A1(net_90) );
AND2_X4 inst_776 ( .ZN(net_724), .A1(net_550), .A2(net_371) );
NAND2_X2 inst_473 ( .ZN(net_638), .A2(net_622), .A1(net_575) );
NAND2_X4 inst_217 ( .ZN(net_729), .A1(net_719), .A2(net_259) );
INV_X4 inst_572 ( .ZN(net_39), .A(net_38) );
INV_X2 inst_742 ( .ZN(net_167), .A(net_166) );
NOR2_X2 inst_77 ( .A1(net_758), .ZN(net_356), .A2(net_70) );
NAND3_X2 inst_171 ( .ZN(net_432), .A2(net_431), .A1(net_352), .A3(net_297) );
INV_X4 inst_691 ( .ZN(net_502), .A(net_385) );
INV_X4 inst_558 ( .A(net_48), .ZN(net_21) );
NAND2_X2 inst_427 ( .ZN(net_558), .A2(net_468), .A1(net_300) );
NAND2_X2 inst_257 ( .ZN(net_659), .A2(net_294), .A1(net_189) );
INV_X4 inst_594 ( .A(net_102), .ZN(net_73) );
NAND3_X4 inst_145 ( .ZN(net_693), .A3(net_295), .A2(net_217), .A1(net_199) );
NAND2_X2 inst_290 ( .ZN(net_217), .A1(net_216), .A2(net_140) );
NAND2_X2 inst_374 ( .ZN(net_450), .A1(net_449), .A2(net_315) );
NAND2_X2 inst_272 ( .ZN(net_170), .A1(net_169), .A2(net_168) );
INV_X8 inst_502 ( .A(net_763), .ZN(net_5) );
NOR2_X2 inst_103 ( .ZN(net_514), .A2(net_436), .A1(net_402) );
NAND2_X2 inst_485 ( .A2(net_647), .A1(net_383), .ZN(v13_D_17) );
AND2_X4 inst_770 ( .A2(net_542), .ZN(net_141), .A1(net_42) );
INV_X4 inst_565 ( .ZN(net_52), .A(net_29) );
NAND2_X2 inst_248 ( .ZN(net_109), .A2(net_41), .A1(v3) );
INV_X4 inst_672 ( .A(net_338), .ZN(net_244) );
INV_X4 inst_622 ( .ZN(net_230), .A(net_104) );
NAND4_X2 inst_138 ( .ZN(net_711), .A4(net_671), .A1(net_670), .A2(net_569), .A3(net_528) );
NAND2_X2 inst_389 ( .ZN(net_486), .A2(net_367), .A1(net_356) );
CLKBUF_X2 inst_789 ( .A(net_769), .Z(net_770) );
NAND2_X2 inst_357 ( .ZN(net_748), .A2(net_258), .A1(net_202) );
NAND2_X2 inst_409 ( .A1(net_546), .ZN(net_525), .A2(net_429) );
NAND3_X2 inst_180 ( .A3(net_678), .A1(net_677), .ZN(net_661), .A2(net_302) );
INV_X4 inst_703 ( .ZN(net_546), .A(net_402) );
NOR3_X4 inst_33 ( .A3(net_724), .A1(net_723), .ZN(net_690), .A2(net_524) );
NAND2_X2 inst_312 ( .ZN(net_273), .A1(net_272), .A2(net_268) );
INV_X4 inst_660 ( .ZN(net_251), .A(net_202) );
INV_X2 inst_731 ( .ZN(net_355), .A(net_154) );
INV_X4 inst_609 ( .ZN(net_139), .A(net_131) );
INV_X8 inst_517 ( .ZN(net_643), .A(net_613) );
NAND2_X2 inst_309 ( .ZN(net_733), .A2(net_159), .A1(net_122) );
NAND2_X4 inst_232 ( .A2(net_758), .A1(net_694), .ZN(net_666) );
NAND2_X2 inst_347 ( .ZN(net_753), .A1(net_375), .A2(net_278) );
AND3_X2 inst_768 ( .ZN(net_587), .A1(net_586), .A2(net_552), .A3(net_475) );
CLKBUF_X2 inst_795 ( .A(net_775), .Z(net_776) );
INV_X4 inst_663 ( .ZN(net_214), .A(net_213) );
NAND2_X2 inst_301 ( .ZN(net_241), .A1(net_240), .A2(net_98) );
NAND2_X2 inst_363 ( .A1(net_758), .ZN(net_423), .A2(net_351) );
INV_X16 inst_755 ( .ZN(net_102), .A(net_93) );
NOR4_X2 inst_27 ( .ZN(net_696), .A1(net_391), .A3(net_375), .A2(net_292), .A4(net_198) );
NAND2_X2 inst_247 ( .A1(net_762), .A2(net_718), .ZN(net_69) );
NAND2_X2 inst_297 ( .A2(net_703), .ZN(net_702), .A1(net_187) );
NAND2_X2 inst_403 ( .ZN(net_516), .A2(net_438), .A1(net_339) );
NAND2_X2 inst_302 ( .A1(net_526), .A2(net_281), .ZN(net_250) );
NAND2_X2 inst_310 ( .ZN(net_270), .A1(net_269), .A2(net_268) );
NAND2_X2 inst_322 ( .A2(net_758), .ZN(net_446), .A1(net_211) );
INV_X4 inst_673 ( .ZN(net_306), .A(net_251) );
NAND2_X2 inst_253 ( .ZN(net_111), .A1(net_82), .A2(net_33) );
NAND2_X4 inst_211 ( .ZN(net_362), .A2(net_132), .A1(net_70) );
INV_X4 inst_619 ( .ZN(net_269), .A(net_128) );
INV_X4 inst_681 ( .ZN(net_435), .A(net_211) );
NAND3_X2 inst_162 ( .ZN(net_328), .A3(net_246), .A1(net_192), .A2(net_137) );
INV_X4 inst_589 ( .A(net_113), .ZN(net_75) );
INV_X4 inst_561 ( .A(net_303), .ZN(net_113) );
CLKBUF_X2 inst_794 ( .A(net_766), .Z(net_775) );
NAND2_X2 inst_412 ( .ZN(net_531), .A1(net_464), .A2(net_241) );
NAND2_X2 inst_449 ( .A1(net_643), .ZN(net_605), .A2(net_573) );
INV_X4 inst_639 ( .ZN(net_268), .A(net_260) );
NAND3_X2 inst_155 ( .ZN(net_243), .A3(net_145), .A2(net_78), .A1(net_63) );
NAND2_X2 inst_464 ( .ZN(net_625), .A2(net_616), .A1(net_611) );
INV_X4 inst_602 ( .A(net_94), .ZN(net_80) );
NOR2_X4 inst_59 ( .A1(net_762), .ZN(net_349), .A2(net_106) );
NAND4_X2 inst_135 ( .A2(net_643), .ZN(net_571), .A4(net_488), .A1(net_416), .A3(net_229) );
NAND2_X2 inst_341 ( .ZN(net_367), .A2(net_252), .A1(net_205) );
NAND2_X4 inst_196 ( .A1(net_55), .ZN(net_43), .A2(net_42) );
INV_X4 inst_532 ( .ZN(net_13), .A(net_3) );
NOR2_X4 inst_55 ( .A1(net_246), .ZN(net_157), .A2(net_131) );
NOR3_X2 inst_37 ( .A2(net_594), .A1(net_231), .A3(net_146), .ZN(v13_D_20) );
INV_X4 inst_641 ( .ZN(net_419), .A(net_156) );
MUX2_X2 inst_498 ( .S(net_762), .A(net_303), .Z(net_285), .B(net_284) );
INV_X2 inst_740 ( .A(net_363), .ZN(net_151) );
INV_X4 inst_684 ( .A(net_385), .ZN(net_299) );
NAND2_X2 inst_264 ( .ZN(net_692), .A1(net_142), .A2(net_141) );
NOR2_X2 inst_84 ( .ZN(net_256), .A1(net_234), .A2(net_131) );
INV_X2 inst_723 ( .A(net_762), .ZN(net_732) );
NAND3_X2 inst_173 ( .A3(net_758), .A1(net_685), .ZN(net_677), .A2(net_147) );
NAND2_X2 inst_298 ( .ZN(net_750), .A2(net_738), .A1(net_166) );
NAND2_X2 inst_303 ( .A1(net_526), .ZN(net_252), .A2(net_72) );
INV_X4 inst_611 ( .ZN(net_120), .A(net_99) );
NAND2_X4 inst_224 ( .A1(net_734), .ZN(net_669), .A2(net_535) );
NOR3_X2 inst_42 ( .ZN(net_547), .A2(net_546), .A3(net_545), .A1(net_472) );
NAND2_X2 inst_287 ( .A2(net_399), .ZN(net_308), .A1(net_269) );
NAND2_X2 inst_323 ( .ZN(net_742), .A1(net_321), .A2(net_320) );
INV_X4 inst_618 ( .ZN(net_326), .A(net_36) );
NAND2_X2 inst_426 ( .ZN(net_557), .A1(net_510), .A2(net_471) );
INV_X4 inst_588 ( .ZN(net_65), .A(net_64) );
INV_X4 inst_648 ( .ZN(net_215), .A(net_171) );
NAND2_X2 inst_350 ( .A2(net_717), .ZN(net_387), .A1(net_359) );
NAND2_X4 inst_231 ( .A2(net_689), .A1(net_688), .ZN(net_684) );
NAND2_X2 inst_270 ( .ZN(net_164), .A2(net_162), .A1(net_83) );
NAND2_X2 inst_474 ( .ZN(net_640), .A2(net_630), .A1(net_508) );
CLKBUF_X2 inst_793 ( .A(net_773), .Z(net_774) );
AND3_X4 inst_766 ( .ZN(net_681), .A3(net_248), .A2(net_154), .A1(net_35) );
INV_X4 inst_715 ( .ZN(net_714), .A(net_650) );
NOR4_X2 inst_26 ( .ZN(net_455), .A2(net_454), .A3(net_453), .A1(net_425), .A4(net_404) );
NAND2_X2 inst_437 ( .ZN(net_579), .A1(net_578), .A2(net_515) );
NAND2_X1 inst_490 ( .A1(net_346), .A2(net_135), .ZN(net_129) );
CLKBUF_X2 inst_801 ( .A(net_781), .Z(net_782) );
INV_X4 inst_626 ( .ZN(net_253), .A(net_116) );
INV_X4 inst_692 ( .ZN(net_578), .A(net_358) );
NOR2_X2 inst_70 ( .A1(net_732), .ZN(net_85), .A2(net_17) );
NAND4_X2 inst_129 ( .A4(net_340), .ZN(net_283), .A1(net_91), .A3(net_45), .A2(net_37) );
NAND3_X2 inst_189 ( .A3(net_637), .A1(net_595), .A2(net_459), .ZN(v13_D_8) );
OR2_X4 inst_11 ( .A1(net_721), .ZN(net_179), .A2(net_137) );
INV_X4 inst_631 ( .A(net_139), .ZN(net_126) );
NAND3_X2 inst_188 ( .A2(net_634), .A3(net_629), .A1(net_593), .ZN(v13_D_14) );
OR2_X2 inst_14 ( .A1(net_31), .ZN(net_25), .A2(net_24) );
NAND2_X2 inst_475 ( .A1(net_643), .ZN(net_641), .A2(net_632) );
NAND2_X2 inst_441 ( .ZN(net_588), .A1(net_525), .A2(net_484) );
NOR3_X4 inst_31 ( .ZN(net_728), .A3(net_683), .A1(net_682), .A2(net_225) );
INV_X4 inst_528 ( .A(net_759), .ZN(net_1) );
NAND2_X2 inst_252 ( .ZN(net_101), .A2(net_52), .A1(net_23) );
CLKBUF_X2 inst_798 ( .A(net_778), .Z(net_779) );
NOR2_X4 inst_62 ( .A1(net_728), .ZN(net_639), .A2(net_545) );
AND2_X4 inst_777 ( .ZN(net_536), .A2(net_486), .A1(net_307) );
INV_X4 inst_557 ( .A(net_115), .ZN(net_38) );
NAND2_X2 inst_251 ( .ZN(net_721), .A2(net_193), .A1(net_93) );
NAND2_X2 inst_352 ( .A1(net_552), .ZN(net_394), .A2(net_393) );
INV_X4 inst_575 ( .ZN(net_66), .A(net_44) );
NAND2_X2 inst_398 ( .ZN(net_507), .A2(net_382), .A1(net_158) );
NAND2_X2 inst_286 ( .ZN(net_207), .A1(net_206), .A2(net_144) );
NAND2_X2 inst_436 ( .A1(net_578), .ZN(net_577), .A2(net_512) );
NAND2_X2 inst_484 ( .A2(net_713), .A1(net_712), .ZN(net_648) );
INV_X4 inst_627 ( .ZN(net_245), .A(net_88) );
NAND2_X2 inst_300 ( .ZN(net_685), .A1(net_179), .A2(net_165) );
NOR2_X2 inst_102 ( .ZN(net_668), .A2(net_384), .A1(net_319) );
NOR3_X4 inst_32 ( .ZN(net_709), .A1(net_636), .A3(net_389), .A2(net_305) );
NAND2_X2 inst_344 ( .A2(net_692), .A1(net_691), .ZN(net_676) );
NAND2_X2 inst_428 ( .ZN(net_559), .A1(net_511), .A2(net_357) );
NAND2_X2 inst_446 ( .ZN(net_597), .A1(net_596), .A2(net_538) );
NAND2_X2 inst_364 ( .ZN(net_430), .A1(net_429), .A2(net_412) );
NAND3_X4 inst_144 ( .A1(net_731), .ZN(net_410), .A3(net_131), .A2(net_78) );
INV_X4 inst_629 ( .ZN(net_123), .A(net_106) );
NAND2_X4 inst_195 ( .ZN(net_287), .A2(v4), .A1(v5) );
NAND2_X2 inst_407 ( .A1(net_693), .ZN(net_670), .A2(net_106) );
CLKBUF_X2 inst_791 ( .A(net_767), .Z(net_772) );
INV_X4 inst_623 ( .A(net_162), .ZN(net_105) );
NAND2_X2 inst_411 ( .A1(net_550), .ZN(net_529), .A2(net_420) );
NOR2_X2 inst_97 ( .ZN(net_408), .A2(net_254), .A1(net_135) );
INV_X4 inst_616 ( .ZN(net_504), .A(net_97) );
AND2_X4 inst_775 ( .ZN(net_683), .A1(net_176), .A2(net_142) );
NOR2_X1 inst_124 ( .ZN(net_738), .A1(net_190), .A2(net_17) );
INV_X4 inst_533 ( .A(net_12), .ZN(net_6) );
INV_X4 inst_620 ( .ZN(net_613), .A(net_501) );
INV_X4 inst_652 ( .A(net_762), .ZN(net_237) );
INV_X4 inst_680 ( .A(net_431), .ZN(net_364) );
CLKBUF_X2 inst_785 ( .A(net_765), .Z(net_766) );
INV_X2 inst_737 ( .A(net_425), .ZN(net_143) );
NAND4_X2 inst_137 ( .A2(net_659), .A1(net_658), .ZN(net_581), .A4(net_328), .A3(net_247) );
INV_X4 inst_677 ( .A(net_347), .ZN(net_290) );
NAND2_X2 inst_425 ( .ZN(net_556), .A1(net_542), .A2(net_465) );
INV_X4 inst_545 ( .A(net_762), .ZN(net_55) );
NAND4_X2 inst_130 ( .A2(net_758), .ZN(net_409), .A4(net_406), .A3(net_368), .A1(net_203) );
INV_X2 inst_722 ( .A(net_38), .ZN(net_34) );
NAND2_X4 inst_227 ( .A1(net_660), .ZN(net_601), .A2(net_600) );
NAND2_X2 inst_399 ( .ZN(net_509), .A2(net_392), .A1(net_335) );
DFFR_X2 inst_760 ( .QN(net_763), .RN(net_657), .D(net_651), .CK(net_780) );
INV_X2 inst_746 ( .A(net_308), .ZN(net_257) );
INV_X4 inst_527 ( .ZN(net_54), .A(v2) );
NAND2_X4 inst_226 ( .A1(net_661), .ZN(net_591), .A2(net_113) );
NAND3_X2 inst_176 ( .ZN(net_533), .A1(net_440), .A3(net_269), .A2(net_75) );
NOR2_X4 inst_58 ( .A1(net_227), .ZN(net_180), .A2(net_109) );
NAND2_X2 inst_414 ( .ZN(net_634), .A1(net_492), .A2(net_482) );
NOR2_X2 inst_87 ( .ZN(net_305), .A2(net_304), .A1(net_80) );
NOR2_X4 inst_61 ( .A2(net_681), .A1(net_680), .ZN(net_560) );
INV_X4 inst_562 ( .ZN(net_84), .A(net_26) );
INV_X4 inst_531 ( .A(net_46), .ZN(net_2) );
NAND2_X4 inst_203 ( .A1(net_762), .ZN(net_152), .A2(net_106) );
NAND2_X4 inst_212 ( .ZN(net_745), .A1(net_171), .A2(net_138) );
MUX2_X2 inst_499 ( .A(net_388), .B(net_356), .Z(net_353), .S(net_211) );
NAND2_X2 inst_335 ( .ZN(net_726), .A1(net_705), .A2(net_504) );
INV_X4 inst_674 ( .ZN(net_359), .A(net_314) );
CLKBUF_X2 inst_800 ( .A(net_766), .Z(net_781) );
NAND2_X2 inst_466 ( .ZN(net_627), .A2(net_618), .A1(net_572) );
AND2_X2 inst_780 ( .ZN(net_350), .A2(net_349), .A1(net_38) );
INV_X4 inst_658 ( .ZN(net_460), .A(net_200) );
OR2_X4 inst_10 ( .A2(net_762), .ZN(net_224), .A1(net_115) );
OR3_X2 inst_4 ( .ZN(net_357), .A2(net_356), .A3(net_355), .A1(net_13) );
NAND2_X2 inst_456 ( .ZN(net_617), .A2(net_570), .A1(net_504) );
INV_X4 inst_581 ( .A(net_545), .ZN(net_453) );
INV_X4 inst_600 ( .ZN(net_281), .A(net_77) );
NOR3_X4 inst_28 ( .ZN(net_754), .A3(net_718), .A1(net_419), .A2(net_106) );
NAND2_X2 inst_275 ( .A1(net_504), .ZN(net_354), .A2(net_178) );
NOR2_X2 inst_117 ( .A2(net_608), .A1(net_469), .ZN(v13_D_9) );
NAND2_X2 inst_438 ( .ZN(net_582), .A2(net_518), .A1(net_386) );
MUX2_X1 inst_501 ( .A(net_646), .B(net_602), .S(net_385), .Z(v13_D_12) );
NOR2_X4 inst_49 ( .ZN(net_346), .A1(net_54), .A2(net_53) );
NAND2_X4 inst_204 ( .A2(net_760), .ZN(net_171), .A1(net_36) );
INV_X4 inst_587 ( .ZN(net_246), .A(net_70) );
INV_X4 inst_666 ( .ZN(net_431), .A(net_139) );
NAND3_X2 inst_154 ( .ZN(net_232), .A2(net_176), .A3(net_103), .A1(net_10) );
INV_X4 inst_592 ( .ZN(net_71), .A(net_70) );
INV_X4 inst_546 ( .A(net_758), .ZN(net_11) );
NAND2_X2 inst_324 ( .ZN(net_323), .A1(net_322), .A2(net_320) );
NAND2_X2 inst_465 ( .ZN(net_626), .A2(net_617), .A1(net_434) );
INV_X4 inst_704 ( .ZN(net_491), .A(net_385) );
NOR2_X2 inst_109 ( .ZN(net_561), .A2(net_476), .A1(net_311) );
NOR2_X4 inst_54 ( .A2(net_760), .ZN(net_154), .A1(net_93) );
INV_X4 inst_693 ( .ZN(net_414), .A(net_358) );
INV_X4 inst_570 ( .A(net_758), .ZN(net_545) );
NAND2_X2 inst_390 ( .ZN(net_752), .A2(net_411), .A1(net_363) );
INV_X4 inst_640 ( .ZN(net_200), .A(net_153) );
NOR3_X2 inst_43 ( .A2(net_755), .A1(net_754), .A3(net_679), .ZN(net_563) );
NAND2_X2 inst_359 ( .ZN(net_417), .A2(net_327), .A1(net_266) );
DFFR_X1 inst_765 ( .QN(net_758), .RN(net_657), .D(net_648), .CK(net_784) );
NAND2_X2 inst_256 ( .ZN(net_665), .A1(net_81), .A2(net_68) );
INV_X4 inst_694 ( .ZN(net_360), .A(net_359) );
NOR2_X2 inst_94 ( .ZN(net_473), .A2(net_390), .A1(net_236) );
NAND2_X2 inst_454 ( .ZN(net_614), .A1(net_613), .A2(net_588) );
INV_X4 inst_630 ( .ZN(net_368), .A(net_106) );
NAND2_X2 inst_375 ( .ZN(net_459), .A1(net_426), .A2(net_325) );
NAND2_X2 inst_401 ( .A1(net_569), .ZN(net_513), .A2(net_442) );
NAND2_X2 inst_262 ( .ZN(net_133), .A1(net_132), .A2(net_15) );
INV_X8 inst_512 ( .ZN(net_132), .A(net_43) );
NAND2_X2 inst_355 ( .A1(net_733), .ZN(net_671), .A2(net_406) );
NAND2_X2 inst_243 ( .ZN(net_284), .A1(net_56), .A2(net_10) );
NAND2_X2 inst_285 ( .A1(net_499), .ZN(net_302), .A2(net_121) );
INV_X4 inst_591 ( .ZN(net_673), .A(net_545) );
NAND2_X2 inst_424 ( .ZN(net_554), .A1(net_520), .A2(net_470) );
AND2_X2 inst_782 ( .ZN(net_463), .A1(net_462), .A2(net_323) );
NAND2_X1 inst_497 ( .ZN(net_602), .A2(net_553), .A1(net_377) );
NAND2_X4 inst_218 ( .ZN(net_510), .A1(net_286), .A2(net_121) );
OR2_X2 inst_15 ( .A1(net_758), .ZN(net_86), .A2(net_31) );
INV_X1 inst_757 ( .ZN(net_657), .A(blif_reset_net) );
INV_X4 inst_647 ( .ZN(net_213), .A(net_197) );
NAND2_X2 inst_343 ( .A1(net_435), .ZN(net_370), .A2(net_304) );
OR2_X4 inst_6 ( .A2(net_760), .ZN(net_227), .A1(net_42) );
NAND3_X1 inst_194 ( .A2(net_634), .A1(net_605), .A3(net_596), .ZN(v13_D_11) );
INV_X4 inst_543 ( .ZN(net_115), .A(net_8) );
NAND2_X2 inst_337 ( .A1(net_716), .ZN(net_351), .A2(net_201) );
CLKBUF_X2 inst_787 ( .A(net_767), .Z(net_768) );
INV_X4 inst_670 ( .ZN(net_390), .A(net_320) );
NOR2_X2 inst_123 ( .A1(net_687), .ZN(net_656), .A2(net_654) );
INV_X8 inst_509 ( .ZN(net_70), .A(net_57) );
NAND2_X2 inst_299 ( .ZN(net_722), .A1(net_197), .A2(net_172) );
INV_X4 inst_699 ( .ZN(net_481), .A(net_414) );
NAND2_X2 inst_418 ( .ZN(net_540), .A1(net_480), .A2(net_276) );
NAND2_X2 inst_476 ( .ZN(net_642), .A2(net_625), .A1(net_614) );
NOR2_X2 inst_118 ( .A2(net_624), .A1(net_181), .ZN(v13_D_23) );
NOR2_X2 inst_86 ( .ZN(net_697), .A1(net_303), .A2(net_302) );
NAND3_X2 inst_153 ( .ZN(net_231), .A1(net_230), .A2(net_229), .A3(net_62) );
OR2_X2 inst_20 ( .A1(net_399), .A2(net_349), .ZN(net_333) );
NAND2_X2 inst_442 ( .ZN(net_720), .A2(net_554), .A1(net_385) );
INV_X4 inst_613 ( .ZN(net_127), .A(net_61) );
NOR3_X2 inst_38 ( .ZN(net_679), .A1(net_354), .A2(net_287), .A3(net_196) );
INV_X4 inst_714 ( .ZN(net_687), .A(net_649) );
NAND2_X2 inst_381 ( .ZN(net_468), .A1(net_387), .A2(net_343) );
INV_X2 inst_726 ( .A(net_102), .ZN(net_83) );
NAND2_X2 inst_295 ( .ZN(net_279), .A1(net_224), .A2(net_223) );
NAND2_X2 inst_349 ( .ZN(net_386), .A1(net_385), .A2(net_242) );
NAND2_X2 inst_483 ( .ZN(net_647), .A2(net_642), .A1(net_143) );
INV_X4 inst_576 ( .ZN(net_64), .A(net_45) );
NAND2_X4 inst_209 ( .A2(net_749), .ZN(net_192), .A1(net_118) );
NAND2_X2 inst_259 ( .ZN(net_749), .A1(net_125), .A2(net_94) );
NOR3_X2 inst_40 ( .A1(net_520), .ZN(net_476), .A3(net_388), .A2(net_119) );
NAND2_X2 inst_320 ( .ZN(net_313), .A1(net_224), .A2(net_218) );
NAND3_X2 inst_167 ( .ZN(net_413), .A3(net_412), .A2(net_344), .A1(net_149) );
INV_X4 inst_607 ( .A(net_210), .ZN(net_103) );
NAND2_X2 inst_246 ( .A2(net_761), .ZN(net_61), .A1(net_27) );
INV_X16 inst_756 ( .ZN(net_526), .A(net_152) );
INV_X4 inst_635 ( .ZN(net_535), .A(net_363) );
NOR2_X2 inst_95 ( .ZN(net_395), .A1(net_364), .A2(net_107) );
INV_X4 inst_705 ( .ZN(net_611), .A(net_456) );
OR3_X2 inst_1 ( .ZN(net_704), .A2(net_137), .A1(net_31), .A3(net_17) );
NOR2_X2 inst_72 ( .ZN(net_145), .A2(net_87), .A1(net_71) );
INV_X8 inst_519 ( .A(net_255), .ZN(net_211) );
NAND2_X2 inst_439 ( .ZN(net_583), .A1(net_564), .A2(net_521) );
NAND2_X2 inst_331 ( .ZN(net_342), .A1(net_341), .A2(net_340) );
INV_X4 inst_582 ( .ZN(net_117), .A(net_52) );
INV_X2 inst_735 ( .ZN(net_153), .A(net_120) );
INV_X4 inst_683 ( .A(net_314), .ZN(net_296) );
NOR2_X2 inst_115 ( .ZN(net_615), .A2(net_587), .A1(net_239) );
NAND2_X2 inst_235 ( .A2(net_760), .A1(net_42), .ZN(net_19) );
INV_X2 inst_750 ( .A(net_404), .ZN(net_318) );
NAND2_X4 inst_210 ( .ZN(net_739), .A1(net_686), .A2(net_193) );
NAND2_X2 inst_317 ( .ZN(net_298), .A2(net_297), .A1(net_214) );
INV_X4 inst_667 ( .ZN(net_236), .A(net_139) );
NAND2_X2 inst_278 ( .ZN(net_188), .A2(net_187), .A1(net_116) );
NAND2_X2 inst_467 ( .ZN(net_628), .A2(net_607), .A1(net_453) );
DFFR_X2 inst_761 ( .QN(net_759), .RN(net_657), .D(net_652), .CK(net_776) );
NAND2_X2 inst_239 ( .ZN(net_41), .A2(net_24), .A1(v0) );
NOR2_X2 inst_105 ( .ZN(net_524), .A2(net_463), .A1(net_402) );
NAND2_X1 inst_488 ( .ZN(net_220), .A2(net_47), .A1(net_29) );
NAND2_X2 inst_387 ( .ZN(net_484), .A1(net_385), .A2(net_370) );
INV_X2 inst_725 ( .ZN(net_67), .A(net_66) );
INV_X4 inst_593 ( .ZN(net_443), .A(net_72) );
NAND3_X2 inst_175 ( .ZN(net_477), .A1(net_409), .A3(net_329), .A2(net_177) );
INV_X2 inst_747 ( .ZN(net_264), .A(net_263) );
NAND2_X2 inst_254 ( .ZN(net_698), .A2(net_322), .A1(net_36) );
INV_X4 inst_654 ( .ZN(net_344), .A(net_175) );
INV_X4 inst_625 ( .ZN(net_260), .A(net_168) );
NAND2_X4 inst_225 ( .A2(net_742), .A1(net_741), .ZN(net_715) );
INV_X4 inst_601 ( .ZN(net_330), .A(net_189) );
NAND4_X2 inst_133 ( .A1(net_578), .ZN(net_500), .A2(net_499), .A4(net_346), .A3(net_318) );
INV_X8 inst_508 ( .ZN(net_161), .A(net_19) );
INV_X4 inst_568 ( .ZN(net_59), .A(net_10) );
NOR2_X2 inst_112 ( .A2(net_530), .A1(net_489), .ZN(v13_D_16) );
INV_X4 inst_523 ( .A(net_718), .ZN(net_717) );
NAND2_X2 inst_365 ( .ZN(net_734), .A2(net_361), .A1(net_194) );
DFFR_X2 inst_764 ( .QN(net_760), .RN(net_657), .D(net_656), .CK(net_774) );
NOR2_X2 inst_67 ( .ZN(net_189), .A1(net_57), .A2(net_17) );
NAND3_X2 inst_181 ( .ZN(net_565), .A2(net_564), .A3(net_461), .A1(net_74) );
NAND2_X2 inst_305 ( .A2(net_322), .ZN(net_258), .A1(net_233) );
NAND2_X2 inst_479 ( .ZN(net_646), .A2(net_628), .A1(net_430) );
NOR3_X4 inst_29 ( .ZN(net_295), .A2(net_294), .A1(net_180), .A3(net_85) );
AND2_X4 inst_771 ( .A2(net_760), .ZN(net_142), .A1(net_57) );
NAND2_X2 inst_391 ( .ZN(net_487), .A2(net_365), .A1(net_261) );
INV_X4 inst_661 ( .ZN(net_338), .A(net_265) );
INV_X4 inst_590 ( .A(net_545), .ZN(net_501) );
INV_X4 inst_713 ( .ZN(net_598), .A(net_581) );
NAND2_X4 inst_202 ( .ZN(net_187), .A1(net_135), .A2(net_31) );
NAND4_X4 inst_126 ( .ZN(net_672), .A2(net_598), .A1(net_560), .A4(net_232), .A3(net_228) );
NAND2_X2 inst_480 ( .ZN(net_712), .A1(net_684), .A2(CLR) );
INV_X4 inst_634 ( .ZN(net_334), .A(net_121) );
NAND2_X2 inst_419 ( .ZN(net_548), .A2(net_498), .A1(net_139) );
NAND2_X2 inst_477 ( .ZN(net_644), .A1(net_643), .A2(net_633) );
INV_X4 inst_646 ( .A(net_297), .ZN(net_209) );
INV_X4 inst_564 ( .ZN(net_87), .A(net_27) );
INV_X4 inst_538 ( .A(net_5), .ZN(net_4) );
NAND2_X2 inst_423 ( .A1(net_757), .ZN(net_741), .A2(net_535) );
INV_X2 inst_739 ( .A(net_762), .ZN(net_147) );
NOR3_X2 inst_35 ( .ZN(net_675), .A3(net_46), .A2(net_32), .A1(net_25) );
NAND2_X2 inst_382 ( .ZN(net_470), .A1(net_449), .A2(net_403) );
NOR2_X4 inst_48 ( .A2(net_760), .A1(net_31), .ZN(net_26) );
NAND2_X2 inst_358 ( .ZN(net_415), .A2(net_337), .A1(net_308) );
NOR2_X4 inst_46 ( .A1(net_762), .A2(net_761), .ZN(net_36) );
NAND4_X2 inst_136 ( .ZN(net_573), .A1(net_572), .A2(net_497), .A4(net_496), .A3(net_208) );
NOR3_X4 inst_30 ( .ZN(net_699), .A3(net_541), .A2(net_522), .A1(net_421) );
NAND2_X2 inst_330 ( .ZN(net_397), .A1(net_211), .A2(net_168) );
INV_X4 inst_610 ( .A(net_284), .ZN(net_89) );
NAND2_X4 inst_233 ( .ZN(net_743), .A2(net_673), .A1(net_672) );
INV_X4 inst_710 ( .ZN(net_478), .A(net_428) );
NAND3_X2 inst_165 ( .ZN(net_383), .A2(net_340), .A3(net_245), .A1(net_244) );
CLKBUF_X2 inst_796 ( .A(net_775), .Z(net_777) );
NAND2_X2 inst_271 ( .A1(net_542), .A2(net_176), .ZN(net_165) );
NAND2_X2 inst_443 ( .ZN(net_589), .A2(net_559), .A1(net_108) );
INV_X4 inst_633 ( .ZN(net_160), .A(net_70) );
NOR3_X2 inst_34 ( .A2(net_190), .ZN(net_63), .A1(net_62), .A3(net_8) );
OR2_X4 inst_12 ( .ZN(net_678), .A1(net_363), .A2(net_362) );
INV_X4 inst_529 ( .ZN(net_654), .A(CLR) );
INV_X4 inst_524 ( .ZN(net_32), .A(v3) );
NOR2_X4 inst_56 ( .ZN(net_166), .A2(net_117), .A1(net_97) );
NOR2_X2 inst_71 ( .ZN(net_248), .A2(net_117), .A1(net_106) );
INV_X4 inst_655 ( .ZN(net_320), .A(net_196) );
NAND2_X2 inst_308 ( .ZN(net_266), .A2(net_265), .A1(net_139) );
NOR2_X2 inst_104 ( .ZN(net_517), .A1(net_437), .A2(net_267) );
NAND2_X2 inst_448 ( .ZN(net_604), .A1(net_603), .A2(net_557) );
NOR2_X4 inst_60 ( .ZN(net_528), .A2(net_458), .A1(net_256) );
NAND2_X2 inst_455 ( .ZN(net_616), .A2(net_567), .A1(net_270) );
NAND3_X2 inst_168 ( .ZN(net_424), .A3(net_264), .A1(net_230), .A2(net_183) );
INV_X4 inst_695 ( .ZN(net_603), .A(net_564) );
INV_X2 inst_730 ( .ZN(net_96), .A(net_95) );
INV_X2 inst_727 ( .ZN(net_184), .A(net_136) );
INV_X4 inst_675 ( .A(net_263), .ZN(net_262) );
NAND2_X2 inst_384 ( .ZN(net_474), .A2(net_473), .A1(net_65) );
INV_X1 inst_758 ( .A(net_135), .ZN(net_51) );
NAND2_X2 inst_321 ( .ZN(net_315), .A1(net_314), .A2(net_279) );
NAND2_X1 inst_496 ( .ZN(net_483), .A1(net_454), .A2(net_372) );
INV_X4 inst_653 ( .A(net_334), .ZN(net_324) );
INV_X4 inst_608 ( .ZN(net_499), .A(net_86) );
NAND2_X2 inst_336 ( .A1(net_702), .ZN(net_348), .A2(net_137) );
INV_X4 inst_563 ( .ZN(net_406), .A(net_56) );
INV_X4 inst_583 ( .ZN(net_125), .A(net_87) );
INV_X4 inst_580 ( .ZN(net_322), .A(net_49) );
NAND3_X2 inst_170 ( .ZN(net_428), .A3(net_243), .A1(net_195), .A2(net_163) );
NAND2_X2 inst_258 ( .ZN(net_381), .A1(net_246), .A2(net_121) );
NAND2_X2 inst_376 ( .ZN(net_461), .A1(net_460), .A2(net_331) );
NAND2_X4 inst_199 ( .A1(net_762), .ZN(net_95), .A2(net_48) );
NOR3_X2 inst_41 ( .ZN(net_543), .A1(net_542), .A2(net_435), .A3(net_433) );
INV_X8 inst_511 ( .ZN(net_135), .A(net_40) );
NAND3_X4 inst_143 ( .A2(net_740), .A1(net_739), .ZN(net_708), .A3(net_182) );
INV_X4 inst_708 ( .ZN(net_464), .A(net_402) );
NAND3_X2 inst_152 ( .ZN(net_191), .A2(net_190), .A3(net_189), .A1(net_31) );
NAND2_X2 inst_265 ( .ZN(net_144), .A1(net_132), .A2(net_20) );
NAND2_X2 inst_482 ( .A2(net_644), .A1(net_576), .ZN(v13_D_6) );
NAND2_X2 inst_468 ( .A1(net_643), .ZN(net_629), .A2(net_619) );
INV_X4 inst_682 ( .ZN(net_552), .A(net_347) );
INV_X2 inst_736 ( .ZN(net_223), .A(net_162) );
INV_X4 inst_544 ( .A(net_134), .ZN(net_18) );
NAND2_X2 inst_238 ( .A2(net_761), .ZN(net_30), .A1(net_9) );
INV_X4 inst_540 ( .ZN(net_22), .A(net_6) );
INV_X4 inst_539 ( .ZN(net_42), .A(net_5) );
NAND2_X2 inst_429 ( .ZN(net_562), .A2(net_503), .A1(net_427) );
INV_X2 inst_724 ( .A(net_161), .ZN(net_72) );
NAND2_X2 inst_404 ( .ZN(net_518), .A2(net_447), .A1(net_64) );
NAND3_X2 inst_178 ( .ZN(net_660), .A3(net_596), .A2(net_544), .A1(net_507) );
NOR2_X2 inst_89 ( .A2(net_362), .ZN(net_311), .A1(net_39) );
NOR2_X2 inst_111 ( .ZN(net_584), .A1(net_514), .A2(net_422) );
NOR2_X2 inst_66 ( .A1(net_761), .ZN(net_718), .A2(net_5) );
NAND2_X2 inst_388 ( .A1(net_603), .ZN(net_485), .A2(net_321) );
INV_X2 inst_734 ( .A(net_326), .ZN(net_112) );
OR2_X4 inst_7 ( .A1(net_760), .A2(net_287), .ZN(net_16) );
NAND3_X2 inst_182 ( .ZN(net_713), .A1(net_499), .A3(net_417), .A2(CLR) );
NAND2_X2 inst_392 ( .ZN(net_488), .A2(net_413), .A1(net_289) );
NOR2_X2 inst_120 ( .A1(net_701), .A2(net_654), .ZN(net_652) );
NAND2_X2 inst_273 ( .A1(net_287), .ZN(net_172), .A2(net_100) );
CLKBUF_X2 inst_788 ( .A(net_768), .Z(net_769) );
NAND2_X2 inst_294 ( .ZN(net_222), .A2(net_220), .A1(net_141) );
NAND2_X4 inst_222 ( .A2(net_762), .A1(net_676), .ZN(net_479) );
NAND2_X2 inst_284 ( .A1(net_762), .ZN(net_201), .A2(net_131) );
NAND2_X1 inst_489 ( .A1(net_762), .ZN(net_122), .A2(net_121) );
NAND3_X2 inst_192 ( .A1(net_641), .A2(net_640), .A3(net_620), .ZN(v13_D_13) );
NAND2_X2 inst_280 ( .ZN(net_194), .A2(net_136), .A1(net_132) );
DFFR_X2 inst_763 ( .QN(net_761), .RN(net_657), .D(net_655), .CK(net_771) );
NAND2_X2 inst_366 ( .A1(net_578), .ZN(net_438), .A2(net_353) );
NAND2_X2 inst_346 ( .ZN(net_373), .A1(net_334), .A2(net_277) );
NAND2_X1 inst_491 ( .ZN(net_205), .A2(net_132), .A1(net_123) );
INV_X4 inst_567 ( .A(net_56), .ZN(net_35) );
NAND3_X1 inst_193 ( .A3(net_643), .ZN(net_592), .A2(net_546), .A1(net_540) );
NAND3_X4 inst_149 ( .A3(net_744), .A1(net_743), .ZN(net_649), .A2(net_539) );
NAND2_X2 inst_318 ( .A1(net_344), .ZN(net_301), .A2(net_215) );
NOR3_X2 inst_39 ( .ZN(net_389), .A3(net_388), .A2(net_355), .A1(net_283) );
NAND2_X4 inst_230 ( .A2(net_700), .A1(net_699), .ZN(net_694) );

endmodule
