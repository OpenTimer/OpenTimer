module c2670 (
n2678,
n8,
n651,
n2,
n123,
n34,
n1971,
n94,
n4,
n543,
n61,
n53,
n120,
n1341,
n16,
n55,
n63,
n95,
n452,
n136,
n65,
n1961,
n27,
n113,
n92,
n2443,
n74,
n2427,
n1,
n14,
n1384,
n128,
n101,
n80,
n1348,
n2106,
n116,
n43,
n49,
n78,
n567,
n142,
n119,
n89,
n114,
n11,
n1956,
n141,
n21,
n105,
n36,
n124,
n103,
n69,
n81,
n40,
n32,
n25,
n1976,
n76,
n131,
n2430,
n661,
n57,
n2104,
n111,
n1991,
n67,
n20,
n29,
n126,
n47,
n107,
n50,
n2066,
n1981,
n73,
n62,
n52,
n91,
n87,
n129,
n139,
n23,
n130,
n127,
n137,
n22,
n72,
n118,
n2096,
n88,
n54,
n19,
n2100,
n75,
n28,
n60,
n64,
n82,
n7,
n2067,
n1966,
n2078,
n2084,
n51,
n140,
n112,
n48,
n2438,
n35,
n135,
n104,
n2454,
n85,
n132,
n117,
n2105,
n93,
n2435,
n37,
n108,
n100,
n3,
n483,
n115,
n102,
n2446,
n99,
n26,
n2451,
n868,
n86,
n5,
n1996,
n68,
n1986,
n1083,
n2090,
n15,
n79,
n96,
n138,
n2474,
n56,
n66,
n77,
n106,
n24,
n125,
n559,
n44,
n2072,
n33,
n6,
n860,
n90,
n227,
n259,
n286,
n223,
n350,
n329,
n319,
n295,
n238,
n217,
n168,
n261,
n237,
n188,
n218,
n311,
n158,
n171,
n288,
n221,
n220,
n321,
n308,
n284,
n297,
n229,
n325,
n282,
n234,
n369,
n145,
n162,
n335,
n367,
n148,
n166,
n409,
n391,
n323,
n290,
n384,
n301,
n164,
n397,
n160,
n401,
n235,
n280,
n411,
n305,
n173,
n156,
n150,
n225,
n176,
n236,
n337,
n331,
n153,
n303,
n219,
n395,
n299);

// Start PIs
input n2678;
input n8;
input n651;
input n2;
input n123;
input n34;
input n1971;
input n94;
input n4;
input n543;
input n61;
input n53;
input n120;
input n1341;
input n16;
input n55;
input n63;
input n95;
input n452;
input n136;
input n65;
input n1961;
input n27;
input n113;
input n92;
input n2443;
input n74;
input n2427;
input n1;
input n14;
input n1384;
input n128;
input n101;
input n80;
input n1348;
input n2106;
input n116;
input n43;
input n49;
input n78;
input n567;
input n142;
input n119;
input n89;
input n114;
input n11;
input n1956;
input n141;
input n21;
input n105;
input n36;
input n124;
input n103;
input n69;
input n81;
input n40;
input n32;
input n25;
input n1976;
input n76;
input n131;
input n2430;
input n661;
input n57;
input n2104;
input n111;
input n1991;
input n67;
input n20;
input n29;
input n126;
input n47;
input n107;
input n50;
input n2066;
input n1981;
input n73;
input n62;
input n52;
input n91;
input n87;
input n129;
input n139;
input n23;
input n130;
input n127;
input n137;
input n22;
input n72;
input n118;
input n2096;
input n88;
input n54;
input n19;
input n2100;
input n75;
input n28;
input n60;
input n64;
input n82;
input n7;
input n2067;
input n1966;
input n2078;
input n2084;
input n51;
input n140;
input n112;
input n48;
input n2438;
input n35;
input n135;
input n104;
input n2454;
input n85;
input n132;
input n117;
input n2105;
input n93;
input n2435;
input n37;
input n108;
input n100;
input n3;
input n483;
input n115;
input n102;
input n2446;
input n99;
input n26;
input n2451;
input n868;
input n86;
input n5;
input n1996;
input n68;
input n1986;
input n1083;
input n2090;
input n15;
input n79;
input n96;
input n138;
input n2474;
input n56;
input n66;
input n77;
input n106;
input n24;
input n125;
input n559;
input n44;
input n2072;
input n33;
input n6;
input n860;
input n90;

// Start POs
output n227;
output n259;
output n286;
output n223;
output n350;
output n329;
output n319;
output n295;
output n238;
output n217;
output n168;
output n261;
output n237;
output n188;
output n218;
output n311;
output n158;
output n171;
output n288;
output n221;
output n220;
output n321;
output n308;
output n284;
output n297;
output n229;
output n325;
output n282;
output n234;
output n369;
output n145;
output n162;
output n335;
output n367;
output n148;
output n166;
output n409;
output n391;
output n323;
output n290;
output n384;
output n301;
output n164;
output n397;
output n160;
output n401;
output n235;
output n280;
output n411;
output n305;
output n173;
output n156;
output n150;
output n225;
output n176;
output n236;
output n337;
output n331;
output n153;
output n303;
output n219;
output n395;
output n299;

// Start wires
wire n2678;
wire net_47;
wire n2;
wire net_176;
wire n319;
wire net_215;
wire net_137;
wire n1971;
wire net_132;
wire net_54;
wire net_237;
wire n94;
wire net_105;
wire n543;
wire n61;
wire n53;
wire net_129;
wire net_119;
wire net_98;
wire n1341;
wire net_12;
wire net_151;
wire net_53;
wire net_93;
wire net_210;
wire n63;
wire n220;
wire net_168;
wire n136;
wire n1961;
wire n27;
wire n113;
wire net_259;
wire net_269;
wire net_127;
wire n74;
wire n391;
wire n1;
wire n14;
wire net_76;
wire n128;
wire n101;
wire net_101;
wire n160;
wire net_187;
wire n1348;
wire net_111;
wire net_264;
wire net_90;
wire net_225;
wire n116;
wire net_100;
wire n150;
wire n43;
wire net_85;
wire n78;
wire n567;
wire net_263;
wire net_252;
wire net_124;
wire n142;
wire n119;
wire n176;
wire net_240;
wire net_160;
wire n1956;
wire n141;
wire net_221;
wire n21;
wire net_115;
wire n153;
wire n105;
wire net_4;
wire n36;
wire n124;
wire net_17;
wire n286;
wire n223;
wire net_164;
wire n81;
wire net_87;
wire net_0;
wire n32;
wire net_35;
wire n25;
wire n1976;
wire net_16;
wire n131;
wire net_239;
wire net_193;
wire net_157;
wire net_257;
wire n57;
wire net_233;
wire net_42;
wire net_120;
wire n308;
wire net_201;
wire net_109;
wire n67;
wire net_80;
wire net_65;
wire net_50;
wire n297;
wire n234;
wire net_234;
wire net_96;
wire net_66;
wire net_38;
wire net_167;
wire n409;
wire n47;
wire net_207;
wire net_136;
wire net_280;
wire net_19;
wire net_126;
wire net_278;
wire n173;
wire n73;
wire net_34;
wire net_108;
wire net_270;
wire n87;
wire n129;
wire n139;
wire net_183;
wire n130;
wire n303;
wire net_150;
wire net_63;
wire net_274;
wire n22;
wire n72;
wire n118;
wire n350;
wire n238;
wire net_30;
wire n2096;
wire net_189;
wire n19;
wire net_99;
wire net_24;
wire net_186;
wire net_46;
wire n60;
wire n64;
wire net_118;
wire n82;
wire n7;
wire net_216;
wire n2067;
wire net_146;
wire n171;
wire n2078;
wire net_122;
wire net_7;
wire n51;
wire net_224;
wire n2438;
wire n35;
wire net_172;
wire net_52;
wire net_165;
wire n166;
wire n290;
wire n384;
wire n2454;
wire net_13;
wire net_246;
wire net_94;
wire n85;
wire n132;
wire n2105;
wire n93;
wire net_219;
wire n2435;
wire net_18;
wire net_131;
wire net_114;
wire net_196;
wire net_29;
wire n331;
wire n108;
wire net_149;
wire net_142;
wire net_248;
wire net_31;
wire n3;
wire n483;
wire net_36;
wire net_158;
wire n115;
wire n102;
wire net_41;
wire net_198;
wire net_253;
wire net_276;
wire n26;
wire net_209;
wire n261;
wire net_3;
wire net_154;
wire n868;
wire n86;
wire net_213;
wire n1996;
wire n158;
wire net_238;
wire net_260;
wire net_28;
wire n321;
wire n1986;
wire n1083;
wire n284;
wire n15;
wire n79;
wire n96;
wire net_97;
wire n229;
wire n325;
wire n2474;
wire n66;
wire n335;
wire net_182;
wire net_192;
wire net_60;
wire net_267;
wire net_273;
wire net_256;
wire n397;
wire net_58;
wire net_82;
wire n280;
wire n235;
wire net_64;
wire net_121;
wire net_73;
wire n44;
wire net_200;
wire n236;
wire net_177;
wire net_86;
wire net_75;
wire net_206;
wire net_195;
wire net_125;
wire n860;
wire net_166;
wire net_107;
wire net_223;
wire n651;
wire n8;
wire net_179;
wire net_235;
wire net_159;
wire n123;
wire net_61;
wire n34;
wire n4;
wire net_62;
wire n188;
wire net_6;
wire n120;
wire net_217;
wire n311;
wire net_271;
wire net_23;
wire net_117;
wire n16;
wire net_74;
wire n55;
wire net_250;
wire net_205;
wire net_135;
wire n95;
wire n452;
wire net_265;
wire net_242;
wire n65;
wire net_130;
wire n92;
wire net_147;
wire n2443;
wire n162;
wire n367;
wire net_220;
wire n323;
wire net_14;
wire n2427;
wire net_113;
wire net_26;
wire n1384;
wire net_32;
wire n80;
wire n2106;
wire net_40;
wire n411;
wire n49;
wire net_69;
wire net_161;
wire n114;
wire n89;
wire net_141;
wire n11;
wire net_83;
wire net_95;
wire net_173;
wire n103;
wire net_78;
wire net_27;
wire n69;
wire n295;
wire net_56;
wire n40;
wire net_155;
wire net_261;
wire net_191;
wire net_22;
wire net_181;
wire n76;
wire n2430;
wire net_39;
wire net_245;
wire net_227;
wire net_144;
wire net_102;
wire net_2;
wire net_59;
wire n661;
wire net_9;
wire n111;
wire n2104;
wire n288;
wire n1991;
wire net_162;
wire n20;
wire n29;
wire n145;
wire net_230;
wire net_44;
wire n126;
wire net_277;
wire n301;
wire net_199;
wire net_134;
wire n107;
wire n50;
wire n2066;
wire net_89;
wire net_45;
wire n1981;
wire n305;
wire net_185;
wire n52;
wire n62;
wire n91;
wire net_272;
wire n23;
wire net_178;
wire n337;
wire n127;
wire n219;
wire net_236;
wire net_208;
wire n137;
wire net_212;
wire net_243;
wire n299;
wire n227;
wire net_222;
wire net_152;
wire n329;
wire net_116;
wire n54;
wire n88;
wire net_175;
wire net_91;
wire n2100;
wire n237;
wire n75;
wire net_106;
wire net_55;
wire n28;
wire net_258;
wire net_255;
wire net_140;
wire net_266;
wire net_247;
wire net_279;
wire net_148;
wire net_104;
wire n1966;
wire net_72;
wire n221;
wire net_25;
wire net_229;
wire n2084;
wire net_70;
wire n140;
wire net_251;
wire n48;
wire n112;
wire net_194;
wire net_241;
wire n369;
wire net_5;
wire net_244;
wire net_128;
wire n135;
wire n104;
wire n164;
wire net_138;
wire net_184;
wire n117;
wire net_11;
wire net_123;
wire n37;
wire net_262;
wire net_170;
wire net_68;
wire net_214;
wire net_77;
wire net_249;
wire net_20;
wire n100;
wire net_49;
wire n259;
wire net_15;
wire net_275;
wire net_57;
wire n2446;
wire n217;
wire n168;
wire net_71;
wire n99;
wire net_153;
wire net_156;
wire net_218;
wire net_84;
wire net_174;
wire net_231;
wire n2451;
wire n218;
wire net_112;
wire net_92;
wire net_1;
wire net_103;
wire net_226;
wire net_139;
wire n5;
wire net_43;
wire net_228;
wire net_10;
wire net_180;
wire n68;
wire net_169;
wire net_21;
wire net_51;
wire n2090;
wire net_171;
wire net_79;
wire net_143;
wire n138;
wire n282;
wire net_190;
wire n56;
wire net_88;
wire n148;
wire net_145;
wire net_197;
wire n77;
wire net_204;
wire net_81;
wire n24;
wire n106;
wire net_232;
wire net_163;
wire n401;
wire n559;
wire n125;
wire net_254;
wire net_67;
wire net_202;
wire net_37;
wire n156;
wire net_268;
wire net_188;
wire net_110;
wire n225;
wire net_48;
wire net_33;
wire n2072;
wire net_8;
wire net_211;
wire net_133;
wire n6;
wire n33;
wire net_203;
wire n395;
wire n90;

// Start cells
MUX2_X2 inst_257 ( .A(n299), .Z(n297), .B(n286), .S(n868) );
INV_X1 inst_290 ( .ZN(net_61), .A(n2104) );
NAND3_X1 inst_145 ( .ZN(net_17), .A3(n76), .A2(n651), .A1(n543) );
MUX2_X2 inst_272 ( .B(net_212), .Z(net_150), .A(n4), .S(n16) );
NOR2_X1 inst_103 ( .ZN(net_168), .A2(net_157), .A1(n1996) );
MUX2_X2 inst_248 ( .Z(net_29), .S(n2104), .A(n123), .B(n111) );
NAND2_X1 inst_228 ( .ZN(net_241), .A2(n286), .A1(n8) );
NAND4_X1 inst_125 ( .ZN(net_131), .A3(net_88), .A2(net_71), .A4(net_63), .A1(net_35) );
NAND2_X1 inst_207 ( .ZN(net_81), .A2(net_80), .A1(n62) );
NAND4_X1 inst_138 ( .ZN(net_215), .A4(net_197), .A2(net_179), .A3(net_166), .A1(net_161) );
NAND3_X1 inst_159 ( .A3(net_60), .ZN(net_50), .A1(n2104), .A2(n105) );
NAND4_X1 inst_134 ( .ZN(net_246), .A2(net_102), .A3(net_98), .A4(net_44), .A1(net_20) );
NAND2_X1 inst_244 ( .ZN(net_272), .A1(net_257), .A2(net_254) );
AND3_X4 inst_333 ( .ZN(net_234), .A1(net_187), .A3(net_186), .A2(n290) );
NAND4_X1 inst_131 ( .A3(net_73), .A4(net_72), .A2(net_41), .A1(net_1), .ZN(n305) );
NAND2_X1 inst_214 ( .ZN(net_90), .A2(net_27), .A1(n543) );
NAND3_X1 inst_180 ( .ZN(net_270), .A1(net_269), .A3(net_262), .A2(net_250) );
NAND3_X1 inst_160 ( .A3(net_53), .ZN(net_51), .A1(n543), .A2(n54) );
XNOR2_X1 inst_33 ( .ZN(net_112), .B(net_105), .A(net_4) );
CLKBUF_X1 inst_328 ( .A(n297), .Z(n280) );
INV_X1 inst_312 ( .A(net_266), .ZN(net_259) );
XNOR2_X1 inst_47 ( .ZN(net_192), .B(net_191), .A(net_149) );
XOR2_X1 inst_19 ( .Z(net_179), .B(net_137), .A(n1991) );
INV_X1 inst_309 ( .A(net_186), .ZN(net_182) );
XOR2_X1 inst_8 ( .Z(net_13), .A(n1986), .B(n1981) );
NAND2_X1 inst_232 ( .ZN(net_160), .A2(net_159), .A1(n2072) );
INV_X1 inst_301 ( .A(net_125), .ZN(n162) );
INV_X1 inst_297 ( .A(net_109), .ZN(n164) );
MUX2_X2 inst_247 ( .Z(net_28), .S(n2104), .A(n130), .B(n118) );
XNOR2_X1 inst_27 ( .ZN(net_104), .A(net_9), .B(net_2) );
NOR2_X1 inst_100 ( .A2(net_212), .ZN(net_191), .A1(n559) );
INV_X1 inst_302 ( .A(net_126), .ZN(n160) );
CLKBUF_X1 inst_322 ( .Z(n350), .A(n452) );
INV_X1 inst_310 ( .ZN(net_202), .A(net_201) );
MUX2_X2 inst_279 ( .B(net_246), .A(net_206), .Z(n145), .S(n860) );
MUX2_X2 inst_253 ( .Z(net_109), .A(net_31), .B(net_30), .S(n2105) );
NAND2_X1 inst_211 ( .A2(net_87), .ZN(net_86), .A1(n117) );
NAND3_X1 inst_162 ( .ZN(net_54), .A3(net_53), .A1(n543), .A2(n51) );
NOR2_X1 inst_93 ( .ZN(net_83), .A1(net_60), .A2(n2104) );
NOR3_X1 inst_81 ( .ZN(net_209), .A1(net_200), .A3(net_171), .A2(net_146) );
NAND4_X1 inst_139 ( .A2(net_264), .A1(net_219), .A3(net_158), .A4(net_156), .ZN(n150) );
NAND3_X1 inst_155 ( .A1(net_61), .ZN(net_34), .A2(n2105), .A3(n127) );
XNOR2_X1 inst_59 ( .ZN(net_273), .A(net_232), .B(net_231) );
AND2_X4 inst_341 ( .ZN(net_239), .A1(net_238), .A2(net_236) );
NAND4_X1 inst_135 ( .A2(net_0), .A4(n319), .ZN(n188), .A3(n661), .A1(n483) );
NAND2_X1 inst_196 ( .ZN(net_67), .A2(net_42), .A1(n139) );
XNOR2_X1 inst_55 ( .ZN(net_247), .A(net_203), .B(n299) );
XNOR2_X1 inst_37 ( .ZN(net_134), .A(net_133), .B(n303) );
NAND2_X1 inst_237 ( .ZN(net_198), .A2(net_186), .A1(n8) );
NAND3_X1 inst_148 ( .ZN(net_20), .A3(n80), .A2(n651), .A1(n543) );
MUX2_X2 inst_264 ( .Z(net_151), .B(n290), .A(n24), .S(n16) );
NAND2_X1 inst_191 ( .A2(net_64), .ZN(net_45), .A1(n85) );
NOR3_X1 inst_84 ( .A1(net_239), .A3(net_237), .ZN(n397), .A2(n37) );
XNOR2_X1 inst_51 ( .ZN(net_222), .B(net_180), .A(net_124) );
NAND4_X1 inst_142 ( .ZN(net_278), .A2(net_277), .A4(net_276), .A1(net_270), .A3(net_253) );
INV_X1 inst_315 ( .A(n308), .ZN(n225) );
NOR4_X1 inst_80 ( .ZN(net_262), .A4(net_261), .A2(net_259), .A3(net_210), .A1(n301) );
INV_X1 inst_303 ( .A(n301), .ZN(n171) );
INV_X1 inst_298 ( .A(net_189), .ZN(net_110) );
NAND3_X1 inst_173 ( .ZN(net_186), .A1(net_116), .A3(n160), .A2(n40) );
NAND2_X1 inst_224 ( .ZN(net_102), .A2(net_101), .A1(n67) );
NAND2_X1 inst_216 ( .ZN(net_94), .A2(net_93), .A1(n2106) );
NOR4_X1 inst_78 ( .ZN(net_248), .A4(net_247), .A3(net_214), .A1(net_189), .A2(net_185) );
CLKBUF_X1 inst_323 ( .Z(n337), .A(n2066) );
INV_X1 inst_287 ( .ZN(net_5), .A(n543) );
XNOR2_X1 inst_42 ( .B(net_246), .ZN(net_195), .A(net_189) );
NAND2_X1 inst_241 ( .ZN(net_205), .A1(net_187), .A2(net_186) );
NAND3_X1 inst_177 ( .ZN(net_200), .A1(net_170), .A3(net_163), .A2(net_130) );
NAND2_X1 inst_231 ( .ZN(net_158), .A2(net_157), .A1(n1996) );
MUX2_X2 inst_270 ( .Z(net_164), .B(n305), .A(n6), .S(n16) );
NAND2_X1 inst_183 ( .ZN(net_48), .A2(net_5), .A1(n651) );
XNOR2_X1 inst_26 ( .ZN(net_16), .A(n1996), .B(n1991) );
NAND3_X1 inst_151 ( .ZN(net_23), .A3(n79), .A2(n651), .A1(n543) );
OR4_X1 inst_64 ( .ZN(net_274), .A2(net_273), .A4(net_272), .A1(net_234), .A3(net_233) );
NOR2_X1 inst_107 ( .ZN(net_220), .A2(net_198), .A1(net_147) );
OR2_X4 inst_70 ( .ZN(net_231), .A2(net_205), .A1(n1996) );
NAND4_X1 inst_129 ( .A4(net_81), .A3(net_57), .A2(net_46), .A1(net_18), .ZN(n303) );
NOR2_X1 inst_92 ( .ZN(net_78), .A1(net_61), .A2(n2105) );
NAND2_X1 inst_189 ( .ZN(net_43), .A2(net_42), .A1(n131) );
NAND2_X1 inst_223 ( .ZN(net_100), .A2(net_80), .A1(n64) );
XOR2_X1 inst_11 ( .A(net_131), .B(net_128), .Z(net_124) );
NAND2_X1 inst_188 ( .A2(net_64), .ZN(net_41), .A1(n86) );
XOR2_X1 inst_14 ( .A(net_212), .Z(net_193), .B(n299) );
AND2_X4 inst_340 ( .ZN(net_224), .A1(net_223), .A2(net_222) );
XNOR2_X1 inst_31 ( .ZN(net_107), .B(net_16), .A(net_13) );
AND4_X1 inst_329 ( .ZN(net_264), .A1(net_245), .A2(net_209), .A4(net_173), .A3(net_154) );
MUX2_X2 inst_252 ( .Z(net_108), .A(net_32), .B(net_28), .S(n2105) );
NAND3_X1 inst_158 ( .A3(net_53), .ZN(net_49), .A1(n543), .A2(n49) );
NAND4_X1 inst_141 ( .ZN(net_279), .A4(net_274), .A2(net_258), .A3(net_256), .A1(net_218) );
XNOR2_X1 inst_62 ( .ZN(net_240), .A(net_238), .B(net_207) );
NAND2_X1 inst_200 ( .A2(net_78), .ZN(net_71), .A1(n104) );
MUX2_X2 inst_251 ( .Z(net_32), .S(n2104), .A(n142), .B(n106) );
INV_X1 inst_286 ( .ZN(n220), .A(n82) );
XNOR2_X1 inst_57 ( .ZN(net_214), .A(net_213), .B(net_212) );
AND2_X4 inst_338 ( .ZN(net_146), .A2(net_120), .A1(n2078) );
INV_X1 inst_300 ( .ZN(net_133), .A(n288) );
NOR2_X1 inst_102 ( .ZN(net_165), .A2(net_164), .A1(n1981) );
XNOR2_X1 inst_32 ( .ZN(net_142), .A(net_104), .B(net_6) );
NAND3_X1 inst_144 ( .ZN(n259), .A2(n661), .A3(n2), .A1(n15) );
NAND2_X1 inst_195 ( .ZN(net_66), .A2(net_64), .A1(n81) );
XOR2_X1 inst_21 ( .Z(net_266), .A(net_227), .B(net_226) );
MUX2_X2 inst_281 ( .B(net_280), .A(net_279), .S(net_278), .Z(n329) );
NOR2_X1 inst_97 ( .A2(net_93), .A1(net_91), .ZN(n325) );
NAND4_X1 inst_124 ( .ZN(net_126), .A3(net_89), .A2(net_84), .A4(net_62), .A1(net_56) );
XOR2_X1 inst_18 ( .Z(net_178), .B(net_141), .A(n1956) );
NAND2_X1 inst_208 ( .A2(net_83), .ZN(net_82), .A1(n124) );
NOR3_X1 inst_88 ( .A1(net_271), .A3(n401), .ZN(n308), .A2(n227) );
CLKBUF_X1 inst_316 ( .Z(n411), .A(n2066) );
NAND2_X1 inst_220 ( .A2(net_97), .ZN(n234), .A1(n567) );
XOR2_X1 inst_9 ( .Z(net_14), .A(n2090), .B(n2084) );
NOR2_X1 inst_113 ( .ZN(net_221), .A2(net_220), .A1(net_202) );
NAND2_X1 inst_198 ( .A2(net_78), .ZN(net_69), .A1(n103) );
XNOR2_X1 inst_50 ( .ZN(net_238), .B(net_148), .A(net_134) );
NAND4_X1 inst_137 ( .ZN(net_208), .A1(net_190), .A2(net_178), .A3(net_177), .A4(net_176) );
MUX2_X2 inst_245 ( .Z(net_26), .B(n68), .A(n56), .S(n543) );
NAND4_X1 inst_130 ( .A4(net_76), .A3(net_75), .A2(net_39), .A1(net_24), .ZN(n299) );
NAND2_X1 inst_227 ( .A2(net_110), .ZN(n153), .A1(n860) );
NAND2_X1 inst_226 ( .ZN(net_111), .A1(net_94), .A2(net_92) );
MUX2_X2 inst_260 ( .Z(net_159), .B(net_122), .A(n33), .S(n29) );
NAND3_X1 inst_176 ( .ZN(net_199), .A3(net_160), .A2(net_121), .A1(n11) );
XNOR2_X1 inst_58 ( .ZN(net_252), .B(net_220), .A(net_201) );
NAND3_X1 inst_147 ( .ZN(net_19), .A2(n2105), .A1(n2104), .A3(n115) );
INV_X1 inst_313 ( .ZN(net_251), .A(net_250) );
NOR3_X1 inst_87 ( .ZN(net_275), .A2(net_273), .A3(net_272), .A1(net_235) );
INV_X1 inst_293 ( .ZN(n236), .A(n120) );
XNOR2_X1 inst_61 ( .ZN(net_235), .A(net_234), .B(net_233) );
NAND2_X1 inst_203 ( .ZN(net_75), .A2(net_74), .A1(n53) );
NAND2_X1 inst_212 ( .ZN(net_88), .A2(net_87), .A1(n116) );
NAND2_X1 inst_234 ( .ZN(net_166), .A2(net_164), .A1(n1981) );
XOR2_X1 inst_0 ( .Z(net_2), .A(n2446), .B(n2443) );
AND3_X4 inst_335 ( .ZN(net_242), .A3(net_184), .A1(net_174), .A2(n8) );
NAND2_X1 inst_184 ( .A2(net_64), .ZN(net_37), .A1(n90) );
NAND2_X1 inst_236 ( .A2(net_186), .ZN(net_174), .A1(n1966) );
XOR2_X1 inst_10 ( .Z(net_15), .A(n2678), .B(n2067) );
XOR2_X1 inst_4 ( .Z(net_8), .A(n2100), .B(n2096) );
OR3_X4 inst_65 ( .ZN(net_256), .A3(net_255), .A1(net_232), .A2(net_231) );
XNOR2_X1 inst_28 ( .ZN(net_143), .B(net_10), .A(net_7) );
NAND2_X1 inst_242 ( .ZN(net_218), .A1(net_217), .A2(net_216) );
MUX2_X2 inst_275 ( .Z(net_210), .S(net_186), .A(n2078), .B(n1961) );
NOR2_X1 inst_117 ( .A2(net_255), .ZN(net_254), .A1(net_230) );
NOR2_X1 inst_98 ( .ZN(net_116), .A2(n164), .A1(n1384) );
MUX2_X2 inst_263 ( .Z(net_155), .B(net_131), .S(n29), .A(n26) );
NAND2_X1 inst_190 ( .A2(net_64), .ZN(net_44), .A1(n93) );
NAND2_X1 inst_204 ( .A2(net_80), .ZN(net_76), .A1(n65) );
NAND2_X1 inst_185 ( .A2(net_42), .ZN(net_38), .A1(n136) );
XNOR2_X1 inst_49 ( .ZN(net_196), .B(net_195), .A(net_135) );
NAND3_X1 inst_154 ( .A1(net_61), .ZN(net_33), .A2(n2105), .A3(n119) );
XOR2_X1 inst_13 ( .A(net_212), .B(net_189), .Z(net_149) );
OR2_X2 inst_75 ( .ZN(net_173), .A2(net_169), .A1(n2090) );
AND3_X4 inst_332 ( .A3(net_145), .A1(net_144), .ZN(n401), .A2(n14) );
NAND3_X1 inst_166 ( .A1(net_61), .A3(net_60), .ZN(net_58), .A2(n141) );
NOR2_X1 inst_116 ( .A1(net_238), .ZN(net_237), .A2(net_236) );
CLKBUF_X1 inst_324 ( .Z(n335), .A(n452) );
NAND3_X1 inst_163 ( .A3(net_60), .ZN(net_55), .A1(n2104), .A2(n100) );
XNOR2_X1 inst_54 ( .ZN(net_236), .A(net_196), .B(net_193) );
NOR4_X1 inst_79 ( .A4(net_261), .ZN(net_260), .A3(net_259), .A1(net_244), .A2(net_243) );
NOR2_X1 inst_109 ( .ZN(net_226), .A2(net_198), .A1(n1976) );
NOR2_X1 inst_106 ( .ZN(net_197), .A2(net_165), .A1(net_152) );
NAND2_X1 inst_219 ( .A2(net_97), .ZN(n217), .A1(n2106) );
NAND2_X1 inst_201 ( .A2(net_80), .ZN(net_72), .A1(n61) );
XNOR2_X1 inst_43 ( .ZN(net_167), .B(net_119), .A(n1976) );
INV_X1 inst_304 ( .A(n286), .ZN(n168) );
MUX2_X2 inst_255 ( .B(net_189), .Z(net_118), .A(n19), .S(n16) );
NAND4_X1 inst_128 ( .A4(net_70), .A3(net_54), .A2(net_40), .A1(net_17), .ZN(n286) );
OR2_X2 inst_73 ( .ZN(net_121), .A2(net_120), .A1(n2078) );
MUX2_X2 inst_256 ( .Z(net_119), .B(n288), .A(n23), .S(n16) );
XOR2_X1 inst_23 ( .Z(net_269), .A(net_244), .B(net_243) );
AND2_X4 inst_339 ( .ZN(net_162), .A2(net_155), .A1(n2067) );
NOR2_X1 inst_94 ( .ZN(net_74), .A1(net_5), .A2(n651) );
MUX2_X2 inst_262 ( .Z(net_153), .B(net_126), .A(n34), .S(n29) );
CLKBUF_X1 inst_325 ( .A(n331), .Z(n295) );
NAND2_X1 inst_243 ( .ZN(net_257), .A1(net_229), .A2(net_228) );
INV_X1 inst_285 ( .ZN(net_60), .A(n2105) );
XOR2_X1 inst_15 ( .Z(net_163), .B(net_118), .A(n1341) );
NAND2_X1 inst_218 ( .ZN(net_96), .A2(net_26), .A1(n651) );
NAND2_X1 inst_197 ( .A2(net_74), .ZN(net_68), .A1(n52) );
MUX2_X2 inst_250 ( .Z(net_31), .S(n2104), .A(n138), .B(n102) );
NAND3_X1 inst_179 ( .ZN(net_253), .A3(net_252), .A1(net_227), .A2(net_226) );
AND2_X2 inst_343 ( .ZN(n173), .A1(n94), .A2(n452) );
XNOR2_X1 inst_24 ( .ZN(net_3), .A(n1976), .B(n1971) );
XOR2_X1 inst_6 ( .Z(net_10), .A(n1348), .B(n1341) );
NOR2_X1 inst_114 ( .ZN(net_225), .A1(net_223), .A2(net_222) );
NAND2_X1 inst_194 ( .ZN(net_65), .A2(net_64), .A1(n87) );
AND2_X4 inst_337 ( .ZN(net_244), .A2(n303), .A1(n8) );
NOR4_X1 inst_76 ( .ZN(net_219), .A4(net_199), .A2(net_172), .A3(net_168), .A1(net_162) );
NAND3_X1 inst_150 ( .ZN(net_22), .A2(n2105), .A1(n2104), .A3(n112) );
NAND3_X1 inst_172 ( .A1(net_90), .A2(net_77), .A3(net_45), .ZN(n290) );
MUX2_X2 inst_277 ( .A(net_189), .B(net_188), .Z(n323), .S(n868) );
NOR3_X1 inst_83 ( .A1(net_225), .A3(net_224), .ZN(n395), .A2(n37) );
NAND4_X1 inst_121 ( .A4(net_65), .A1(net_49), .A2(net_48), .A3(net_36), .ZN(n288) );
NAND4_X1 inst_123 ( .ZN(net_125), .A2(net_82), .A1(net_55), .A4(net_38), .A3(net_22) );
INV_X1 inst_306 ( .ZN(net_147), .A(n305) );
INV_X1 inst_299 ( .A(net_111), .ZN(n319) );
XOR2_X1 inst_2 ( .Z(net_6), .A(n2438), .B(n2435) );
NOR3_X1 inst_86 ( .ZN(net_268), .A1(net_265), .A2(net_261), .A3(net_251) );
NAND4_X1 inst_118 ( .ZN(n158), .A3(n2090), .A4(n2084), .A1(n2078), .A2(n2072) );
XOR2_X1 inst_20 ( .Z(net_190), .B(net_150), .A(n1348) );
NAND3_X1 inst_153 ( .ZN(net_25), .A2(n2105), .A1(n2104), .A3(n107) );
XNOR2_X1 inst_38 ( .ZN(net_135), .A(n301), .B(n286) );
INV_X1 inst_295 ( .ZN(net_101), .A(net_48) );
XNOR2_X1 inst_52 ( .A(net_246), .ZN(net_206), .B(net_192) );
NOR2_X1 inst_90 ( .ZN(net_64), .A2(n651), .A1(n543) );
MUX2_X2 inst_267 ( .Z(net_139), .B(n301), .A(n5), .S(n16) );
NAND4_X1 inst_140 ( .ZN(net_277), .A3(net_269), .A4(net_268), .A1(net_266), .A2(net_211) );
NAND2_X1 inst_209 ( .ZN(net_84), .A2(net_83), .A1(n125) );
MUX2_X2 inst_259 ( .Z(net_130), .B(net_129), .S(n29), .A(n28) );
NAND2_X1 inst_221 ( .ZN(net_98), .A2(net_74), .A1(n55) );
XNOR2_X1 inst_40 ( .B(net_113), .A(net_107), .ZN(n229) );
CLKBUF_X1 inst_320 ( .Z(n369), .A(n1083) );
NAND3_X1 inst_167 ( .A1(net_61), .A3(net_60), .ZN(net_59), .A2(n135) );
MUX2_X2 inst_246 ( .Z(net_27), .B(n72), .S(n651), .A(n47) );
INV_X1 inst_289 ( .ZN(n219), .A(n132) );
NOR2_X1 inst_95 ( .ZN(net_80), .A1(net_53), .A2(n543) );
XOR2_X1 inst_1 ( .Z(net_4), .A(n2078), .B(n2072) );
INV_X1 inst_282 ( .ZN(n218), .A(n44) );
OR2_X4 inst_72 ( .ZN(net_280), .A2(net_279), .A1(net_275) );
AND3_X4 inst_331 ( .ZN(net_187), .A3(net_117), .A1(n160), .A2(n40) );
XNOR2_X1 inst_44 ( .ZN(net_223), .A(net_129), .B(net_127) );
MUX2_X2 inst_274 ( .Z(net_213), .S(net_186), .A(n2067), .B(n1348) );
NAND3_X1 inst_174 ( .ZN(net_228), .A1(net_187), .A3(net_186), .A2(net_136) );
NOR2_X1 inst_115 ( .ZN(net_230), .A1(net_229), .A2(net_228) );
NAND2_X1 inst_235 ( .ZN(net_170), .A2(net_169), .A1(n2090) );
CLKBUF_X1 inst_317 ( .Z(n409), .A(n452) );
NAND2_X1 inst_210 ( .ZN(net_85), .A2(net_83), .A1(n129) );
INV_X1 inst_314 ( .ZN(n311), .A(n150) );
NAND3_X1 inst_164 ( .A3(net_60), .ZN(net_56), .A1(n2104), .A2(n101) );
XOR2_X1 inst_5 ( .Z(net_9), .A(n2430), .B(n2427) );
MUX2_X2 inst_278 ( .B(net_212), .A(net_188), .Z(n148), .S(n860) );
NAND3_X1 inst_157 ( .ZN(net_36), .A3(n74), .A2(n651), .A1(n543) );
NAND2_X1 inst_239 ( .ZN(net_183), .A2(net_182), .A1(n2090) );
NOR2_X1 inst_105 ( .ZN(net_172), .A2(net_159), .A1(n2072) );
OR2_X4 inst_68 ( .ZN(net_144), .A1(net_143), .A2(net_142) );
NAND2_X1 inst_213 ( .ZN(net_89), .A2(net_87), .A1(n113) );
XNOR2_X1 inst_53 ( .ZN(net_207), .B(net_195), .A(net_194) );
NAND3_X1 inst_175 ( .ZN(net_216), .A1(net_187), .A3(net_186), .A2(net_131) );
NAND2_X1 inst_205 ( .A2(net_80), .ZN(net_77), .A1(n60) );
MUX2_X2 inst_254 ( .Z(net_120), .B(net_109), .S(n29), .A(n27) );
NAND2_X1 inst_225 ( .ZN(net_103), .A2(net_101), .A1(n66) );
NAND4_X1 inst_133 ( .ZN(net_212), .A4(net_103), .A1(net_51), .A2(net_47), .A3(net_23) );
INV_X1 inst_292 ( .ZN(n235), .A(n69) );
NOR2_X1 inst_112 ( .ZN(net_229), .A2(net_205), .A1(n1991) );
OR3_X2 inst_67 ( .A1(net_115), .A3(net_114), .ZN(n156), .A2(n2100) );
INV_X1 inst_305 ( .A(n303), .ZN(n166) );
NAND2_X1 inst_181 ( .ZN(n223), .A1(n7), .A2(n661) );
NAND4_X1 inst_127 ( .A4(net_100), .A3(net_68), .A2(net_37), .A1(net_21), .ZN(n301) );
XNOR2_X1 inst_29 ( .ZN(net_105), .A(net_15), .B(net_14) );
NAND2_X1 inst_186 ( .A2(net_64), .ZN(net_39), .A1(n91) );
XOR2_X1 inst_17 ( .Z(net_177), .B(net_140), .A(n1966) );
NAND3_X1 inst_146 ( .ZN(net_18), .A3(n75), .A2(n651), .A1(n543) );
MUX2_X2 inst_249 ( .Z(net_30), .S(n2104), .A(n126), .B(n114) );
AND3_X4 inst_334 ( .ZN(net_232), .A1(net_187), .A3(net_186), .A2(net_128) );
NAND2_X1 inst_202 ( .A2(net_74), .ZN(net_73), .A1(n48) );
NAND2_X1 inst_187 ( .A2(net_64), .ZN(net_40), .A1(n89) );
NAND2_X1 inst_206 ( .ZN(net_79), .A2(net_78), .A1(n95) );
NAND4_X1 inst_122 ( .ZN(net_128), .A3(net_86), .A2(net_85), .A4(net_58), .A1(net_50) );
NAND4_X1 inst_126 ( .ZN(net_122), .A2(net_69), .A4(net_67), .A1(net_34), .A3(net_19) );
XNOR2_X1 inst_25 ( .ZN(net_11), .A(n1966), .B(n1961) );
NAND2_X1 inst_240 ( .ZN(net_184), .A2(net_182), .A1(n2084) );
CLKBUF_X1 inst_326 ( .A(n321), .Z(n284) );
NOR2_X1 inst_110 ( .ZN(net_204), .A2(net_203), .A1(n299) );
OR2_X2 inst_74 ( .ZN(net_156), .A2(net_155), .A1(n2067) );
INV_X1 inst_288 ( .ZN(n237), .A(n57) );
NAND2_X1 inst_229 ( .ZN(net_145), .A1(net_143), .A2(net_142) );
NOR2_X1 inst_99 ( .A2(net_129), .ZN(net_114), .A1(n2096) );
XNOR2_X1 inst_35 ( .ZN(net_123), .A(net_122), .B(n164) );
OR2_X4 inst_69 ( .ZN(net_227), .A2(net_198), .A1(net_133) );
XNOR2_X1 inst_48 ( .ZN(net_194), .A(net_193), .B(net_191) );
NOR3_X1 inst_82 ( .ZN(net_249), .A3(net_247), .A2(net_213), .A1(net_212) );
XNOR2_X1 inst_46 ( .ZN(net_180), .A(net_132), .B(net_123) );
AND4_X1 inst_330 ( .ZN(net_267), .A4(net_266), .A1(net_263), .A2(net_252), .A3(net_241) );
XNOR2_X1 inst_30 ( .ZN(net_106), .A(net_12), .B(net_3) );
NAND4_X1 inst_136 ( .A4(n319), .ZN(n176), .A1(n661), .A2(n483), .A3(n36) );
NOR2_X1 inst_108 ( .ZN(net_201), .A2(net_198), .A1(n1981) );
NAND2_X1 inst_233 ( .ZN(net_161), .A2(net_151), .A1(n1986) );
NAND3_X1 inst_165 ( .ZN(net_57), .A3(net_53), .A1(n543), .A2(n50) );
MUX2_X2 inst_271 ( .A(net_212), .Z(n321), .B(n301), .S(n868) );
INV_X1 inst_283 ( .ZN(n238), .A(n108) );
XOR2_X1 inst_22 ( .Z(net_250), .A(net_242), .B(net_241) );
INV_X1 inst_311 ( .ZN(net_261), .A(net_252) );
XNOR2_X1 inst_34 ( .ZN(net_113), .B(net_106), .A(net_11) );
XOR2_X1 inst_12 ( .B(net_136), .Z(net_132), .A(net_108) );
OR2_X4 inst_71 ( .ZN(net_233), .A2(net_205), .A1(n1986) );
XNOR2_X1 inst_56 ( .ZN(net_211), .A(net_210), .B(n171) );
INV_X1 inst_308 ( .A(net_191), .ZN(net_188) );
NOR2_X1 inst_104 ( .ZN(net_171), .A2(net_153), .A1(n2084) );
XNOR2_X1 inst_60 ( .ZN(net_255), .A(net_217), .B(net_216) );
NAND3_X1 inst_168 ( .ZN(net_62), .A1(net_61), .A3(net_60), .A2(n137) );
NAND3_X1 inst_169 ( .ZN(net_63), .A1(net_61), .A3(net_60), .A2(n140) );
NAND2_X1 inst_215 ( .ZN(net_92), .A2(net_91), .A1(n567) );
INV_X1 inst_307 ( .ZN(net_117), .A(net_116) );
NAND3_X1 inst_161 ( .A3(net_53), .ZN(net_52), .A1(n543), .A2(n43) );
XOR2_X1 inst_16 ( .Z(net_176), .B(net_139), .A(n1961) );
MUX2_X2 inst_276 ( .S(net_186), .Z(net_185), .A(n1996), .B(n1341) );
CLKBUF_X1 inst_321 ( .Z(n367), .A(n1083) );
AND2_X4 inst_336 ( .A2(net_129), .ZN(net_115), .A1(n2096) );
XOR2_X1 inst_3 ( .Z(net_7), .A(n2454), .B(n2451) );
NAND3_X1 inst_156 ( .A1(net_61), .ZN(net_35), .A2(n2105), .A3(n128) );
NAND3_X1 inst_170 ( .ZN(net_189), .A1(net_96), .A3(net_66), .A2(net_52) );
MUX2_X2 inst_258 ( .Z(net_157), .B(net_128), .A(n32), .S(n29) );
XNOR2_X1 inst_41 ( .ZN(net_148), .B(net_147), .A(n290) );
NAND2_X1 inst_199 ( .A2(net_80), .ZN(net_70), .A1(n63) );
INV_X1 inst_296 ( .A(n325), .ZN(n261) );
NOR2_X1 inst_91 ( .ZN(net_42), .A1(n2105), .A2(n2104) );
NAND4_X1 inst_132 ( .ZN(net_136), .A2(net_79), .A4(net_43), .A1(net_33), .A3(net_25) );
NAND3_X1 inst_143 ( .ZN(net_1), .A3(n73), .A2(n651), .A1(n543) );
AND2_X4 inst_342 ( .A2(net_269), .ZN(net_263), .A1(net_242) );
XNOR2_X1 inst_36 ( .ZN(net_127), .A(net_126), .B(net_125) );
NAND3_X1 inst_152 ( .ZN(net_24), .A3(n78), .A2(n651), .A1(n543) );
MUX2_X2 inst_265 ( .Z(net_137), .B(net_136), .S(n29), .A(n25) );
NOR2_X1 inst_96 ( .ZN(net_87), .A2(net_61), .A1(net_60) );
XNOR2_X1 inst_45 ( .ZN(net_175), .A(net_138), .B(n1971) );
NOR2_X1 inst_101 ( .ZN(net_152), .A2(net_151), .A1(n1986) );
CLKBUF_X1 inst_319 ( .Z(n384), .A(n2066) );
MUX2_X2 inst_269 ( .Z(net_141), .B(n299), .A(n20), .S(n16) );
NAND2_X1 inst_238 ( .A2(net_186), .ZN(net_181), .A1(n1971) );
MUX2_X2 inst_261 ( .Z(net_169), .B(net_125), .A(n35), .S(n29) );
NAND3_X1 inst_178 ( .ZN(net_243), .A3(net_183), .A1(net_181), .A2(n8) );
NOR3_X1 inst_89 ( .ZN(net_276), .A3(net_267), .A2(net_260), .A1(net_221) );
NOR2_X1 inst_111 ( .ZN(net_217), .A2(net_205), .A1(n2067) );
OR3_X4 inst_66 ( .A3(net_273), .ZN(net_258), .A1(net_257), .A2(net_255) );
MUX2_X2 inst_268 ( .Z(net_140), .B(n286), .A(n21), .S(n16) );
XOR2_X1 inst_7 ( .Z(net_12), .A(n2474), .B(n1956) );
OR4_X1 inst_63 ( .ZN(net_271), .A1(net_111), .A4(n397), .A3(n395), .A2(n229) );
NAND2_X1 inst_182 ( .ZN(net_0), .A2(n3), .A1(n1) );
MUX2_X2 inst_273 ( .Z(net_203), .S(net_186), .A(n2072), .B(n1956) );
NAND4_X1 inst_120 ( .ZN(net_93), .A1(n96), .A4(n82), .A2(n44), .A3(n132) );
INV_X1 inst_294 ( .ZN(net_97), .A(n223) );
NAND4_X1 inst_119 ( .ZN(net_91), .A2(n69), .A4(n57), .A3(n120), .A1(n108) );
INV_X1 inst_284 ( .ZN(net_53), .A(n651) );
NAND2_X1 inst_222 ( .ZN(net_99), .A2(net_78), .A1(n99) );
CLKBUF_X1 inst_327 ( .A(n323), .Z(n282) );
NAND2_X1 inst_192 ( .A2(net_64), .ZN(net_46), .A1(n88) );
MUX2_X2 inst_280 ( .A(net_246), .B(net_240), .Z(n331), .S(n868) );
NOR3_X1 inst_85 ( .ZN(net_265), .A1(net_249), .A3(net_248), .A2(net_204) );
INV_X1 inst_291 ( .ZN(n221), .A(n96) );
MUX2_X2 inst_266 ( .Z(net_138), .B(n303), .A(n22), .S(n16) );
NAND3_X1 inst_149 ( .ZN(net_21), .A3(n77), .A2(n651), .A1(n543) );
NAND2_X1 inst_193 ( .A2(net_64), .ZN(net_47), .A1(n92) );
CLKBUF_X1 inst_318 ( .Z(n391), .A(n452) );
XNOR2_X1 inst_39 ( .B(net_112), .A(net_8), .ZN(n227) );
NAND2_X1 inst_230 ( .ZN(net_154), .A2(net_153), .A1(n2084) );
NAND2_X1 inst_217 ( .ZN(net_95), .A2(net_29), .A1(n2105) );
NOR4_X1 inst_77 ( .ZN(net_245), .A3(net_215), .A4(net_208), .A2(net_175), .A1(net_167) );
NAND3_X1 inst_171 ( .ZN(net_129), .A2(net_99), .A1(net_95), .A3(net_59) );

endmodule
