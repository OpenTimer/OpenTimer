module s400 (
TEST,
FM,
blif_clk_net,
CLR,
blif_reset_net,
YLW1,
RED2,
GRN1,
RED1,
YLW2,
GRN2);

// Start PIs
input TEST;
input FM;
input blif_clk_net;
input CLR;
input blif_reset_net;

// Start POs
output YLW1;
output RED2;
output GRN1;
output RED1;
output YLW2;
output GRN2;

// Start wires
wire net_166;
wire net_107;
wire net_47;
wire net_179;
wire GRN1;
wire net_176;
wire net_159;
wire net_61;
wire net_137;
wire net_132;
wire net_54;
wire net_105;
wire net_62;
wire net_6;
wire net_129;
wire net_119;
wire net_98;
wire net_23;
wire net_117;
wire net_12;
wire net_151;
wire net_74;
wire net_53;
wire net_93;
wire net_210;
wire net_205;
wire net_168;
wire net_135;
wire net_130;
wire net_147;
wire net_127;
wire net_14;
wire net_113;
wire net_26;
wire net_76;
wire blif_clk_net;
wire net_101;
wire net_32;
wire net_187;
wire net_111;
wire net_90;
wire net_40;
wire net_100;
wire net_85;
wire net_69;
wire net_124;
wire net_161;
wire CLR;
wire net_141;
wire net_160;
wire net_83;
wire net_115;
wire RED1;
wire net_4;
wire net_95;
wire net_17;
wire net_173;
wire net_78;
wire net_27;
wire net_164;
wire net_56;
wire net_87;
wire net_0;
wire net_155;
wire net_35;
wire net_191;
wire net_16;
wire net_22;
wire net_181;
wire net_193;
wire net_39;
wire net_157;
wire net_144;
wire net_102;
wire net_2;
wire net_59;
wire net_9;
wire net_42;
wire net_120;
wire net_201;
wire net_109;
wire net_80;
wire net_65;
wire blif_reset_net;
wire net_50;
wire net_162;
wire YLW1;
wire FM;
wire net_96;
wire net_66;
wire net_38;
wire net_44;
wire net_167;
wire net_207;
wire net_199;
wire net_136;
wire net_134;
wire net_19;
wire net_89;
wire net_45;
wire net_126;
wire net_185;
wire net_34;
wire net_108;
wire net_183;
wire TEST;
wire net_178;
wire net_208;
wire net_150;
wire net_63;
wire net_212;
wire net_152;
wire net_30;
wire net_116;
wire net_189;
wire net_175;
wire net_91;
wire net_24;
wire net_55;
wire net_99;
wire net_106;
wire net_186;
wire net_46;
wire net_140;
wire net_118;
wire net_148;
wire net_104;
wire net_146;
wire net_72;
wire net_122;
wire net_25;
wire net_7;
wire net_70;
wire net_194;
wire net_172;
wire net_5;
wire net_52;
wire net_165;
wire net_128;
wire net_138;
wire net_13;
wire net_184;
wire net_94;
wire net_11;
wire net_18;
wire net_123;
wire net_131;
wire net_114;
wire net_196;
wire net_170;
wire net_29;
wire net_68;
wire net_214;
wire net_149;
wire net_142;
wire net_77;
wire net_20;
wire net_31;
wire net_36;
wire net_49;
wire net_158;
wire net_15;
wire net_41;
wire net_57;
wire net_198;
wire net_71;
wire net_209;
wire net_153;
wire net_156;
wire net_3;
wire net_84;
wire net_174;
wire net_154;
wire net_1;
wire net_92;
wire net_112;
wire net_103;
wire net_213;
wire net_139;
wire net_43;
wire YLW2;
wire net_10;
wire net_180;
wire net_28;
wire net_169;
wire net_21;
wire net_51;
wire net_171;
wire net_79;
wire net_143;
wire net_97;
wire net_190;
wire net_88;
wire net_182;
wire net_192;
wire net_145;
wire net_60;
wire net_197;
wire net_204;
wire net_81;
wire RED2;
wire net_163;
wire net_58;
wire GRN2;
wire net_67;
wire net_82;
wire net_64;
wire net_202;
wire net_37;
wire net_188;
wire net_110;
wire net_121;
wire net_73;
wire net_200;
wire net_48;
wire net_33;
wire net_177;
wire net_8;
wire net_75;
wire net_86;
wire net_211;
wire net_133;
wire net_206;
wire net_203;
wire net_195;
wire net_125;

// Start cells
AND4_X4 inst_145 ( .ZN(net_86), .A1(net_80), .A4(net_73), .A2(net_47), .A3(net_37) );
INV_X2 inst_103 ( .A(net_136), .ZN(net_135) );
DFFR_X2 inst_125 ( .RN(net_118), .D(net_43), .QN(net_6), .CK(net_209) );
CLKBUF_X2 inst_207 ( .A(net_172), .Z(net_201) );
DFFR_X1 inst_138 ( .RN(net_118), .D(net_97), .QN(RED2), .CK(net_177) );
CLKBUF_X2 inst_159 ( .A(net_152), .Z(net_153) );
CLKBUF_X2 inst_218 ( .A(net_211), .Z(net_212) );
NOR3_X2 inst_15 ( .A1(net_132), .A2(net_112), .ZN(net_75), .A3(net_54) );
CLKBUF_X2 inst_197 ( .A(net_190), .Z(net_191) );
DFFR_X1 inst_134 ( .RN(net_118), .D(net_72), .Q(YLW2), .CK(net_200) );
CLKBUF_X2 inst_179 ( .A(net_172), .Z(net_173) );
NOR2_X4 inst_24 ( .A1(net_130), .ZN(net_100), .A2(net_29) );
INV_X2 inst_114 ( .ZN(net_15), .A(net_10) );
XNOR2_X1 inst_6 ( .ZN(net_101), .A(net_100), .B(net_99) );
CLKBUF_X2 inst_194 ( .A(net_187), .Z(net_188) );
DFFR_X2 inst_131 ( .RN(net_118), .D(net_103), .QN(net_12), .CK(net_173) );
NAND2_X2 inst_76 ( .A1(net_141), .ZN(net_110), .A2(net_109) );
CLKBUF_X2 inst_214 ( .A(net_207), .Z(net_208) );
CLKBUF_X2 inst_180 ( .A(net_145), .Z(net_174) );
CLKBUF_X2 inst_160 ( .A(net_153), .Z(net_154) );
CLKBUF_X2 inst_150 ( .A(blif_clk_net), .Z(net_144) );
NOR2_X2 inst_33 ( .A1(net_126), .A2(net_76), .ZN(net_69) );
CLKBUF_X2 inst_172 ( .A(net_165), .Z(net_166) );
INV_X4 inst_83 ( .ZN(net_16), .A(net_0) );
NAND3_X2 inst_47 ( .ZN(net_102), .A1(net_100), .A2(net_99), .A3(net_66) );
NOR3_X2 inst_19 ( .ZN(net_105), .A3(net_104), .A1(net_90), .A2(net_83) );
INV_X1 inst_123 ( .ZN(net_118), .A(blif_reset_net) );
INV_X2 inst_121 ( .A(net_100), .ZN(net_93) );
XNOR2_X2 inst_2 ( .ZN(net_54), .A(net_53), .B(net_40) );
OR3_X2 inst_8 ( .A2(net_66), .ZN(net_50), .A1(net_49), .A3(net_48) );
INV_X2 inst_118 ( .ZN(net_33), .A(net_32) );
INV_X4 inst_86 ( .ZN(net_29), .A(net_16) );
CLKBUF_X2 inst_153 ( .A(net_145), .Z(net_147) );
NOR3_X2 inst_20 ( .ZN(net_106), .A3(net_104), .A1(net_94), .A2(net_89) );
NOR2_X2 inst_27 ( .ZN(net_80), .A1(net_2), .A2(CLR) );
NOR2_X2 inst_38 ( .A2(net_129), .ZN(net_92), .A1(net_56) );
INV_X4 inst_100 ( .ZN(net_112), .A(net_109) );
NAND2_X4 inst_52 ( .ZN(net_136), .A1(net_131), .A2(net_70) );
INV_X4 inst_90 ( .ZN(net_58), .A(net_19) );
DFFR_X1 inst_140 ( .RN(net_118), .D(net_107), .QN(net_9), .CK(net_160) );
CLKBUF_X2 inst_209 ( .A(net_202), .Z(net_203) );
CLKBUF_X2 inst_211 ( .A(net_189), .Z(net_205) );
NOR2_X1 inst_40 ( .A2(net_90), .ZN(net_89), .A1(net_88) );
CLKBUF_X2 inst_162 ( .A(net_155), .Z(net_156) );
CLKBUF_X2 inst_167 ( .A(net_155), .Z(net_161) );
INV_X4 inst_93 ( .ZN(net_99), .A(net_1) );
INV_X4 inst_81 ( .ZN(net_70), .A(net_12) );
INV_X4 inst_95 ( .A(net_57), .ZN(net_45) );
XNOR2_X2 inst_1 ( .A(net_51), .ZN(net_30), .B(FM) );
NAND2_X2 inst_72 ( .A2(net_128), .ZN(net_104), .A1(net_45) );
DFFR_X1 inst_139 ( .RN(net_118), .D(net_96), .QN(YLW1), .CK(net_146) );
CLKBUF_X2 inst_155 ( .A(net_148), .Z(net_149) );
NAND2_X2 inst_59 ( .ZN(net_48), .A1(net_16), .A2(net_1) );
DFFR_X1 inst_135 ( .RN(net_118), .D(net_79), .Q(RED1), .CK(net_193) );
CLKBUF_X2 inst_196 ( .A(net_189), .Z(net_190) );
NAND3_X2 inst_44 ( .A3(net_80), .A2(net_58), .A1(net_51), .ZN(net_41) );
NAND2_X4 inst_55 ( .A1(net_125), .ZN(net_98), .A2(net_28) );
CLKBUF_X2 inst_174 ( .A(net_167), .Z(net_168) );
INV_X2 inst_115 ( .ZN(net_88), .A(net_10) );
NOR2_X2 inst_37 ( .A1(net_130), .ZN(net_125), .A2(net_1) );
CLKBUF_X2 inst_210 ( .A(net_203), .Z(net_204) );
AND2_X2 inst_148 ( .ZN(net_53), .A2(net_34), .A1(net_26) );
CLKBUF_X2 inst_164 ( .A(net_157), .Z(net_158) );
CLKBUF_X2 inst_191 ( .A(net_184), .Z(net_185) );
XNOR2_X2 inst_5 ( .ZN(net_108), .A(net_102), .B(net_58) );
CLKBUF_X2 inst_157 ( .A(net_150), .Z(net_151) );
INV_X4 inst_84 ( .ZN(net_66), .A(net_2) );
NAND2_X4 inst_51 ( .A2(net_140), .ZN(net_137), .A1(net_131) );
DFFR_X1 inst_142 ( .RN(net_118), .D(net_114), .QN(net_0), .CK(net_154) );
INV_X4 inst_80 ( .ZN(net_49), .A(net_5) );
CLKBUF_X2 inst_173 ( .A(net_166), .Z(net_167) );
INV_X2 inst_105 ( .A(net_133), .ZN(net_132) );
CLKBUF_X2 inst_213 ( .A(net_206), .Z(net_207) );
NAND2_X2 inst_68 ( .ZN(net_84), .A1(net_81), .A2(net_67) );
CLKBUF_X2 inst_216 ( .A(net_195), .Z(net_210) );
INV_X4 inst_78 ( .ZN(net_87), .A(net_9) );
NAND4_X2 inst_42 ( .A1(net_66), .ZN(net_63), .A4(net_62), .A2(net_51), .A3(net_17) );
CLKBUF_X2 inst_175 ( .A(net_168), .Z(net_169) );
NAND2_X4 inst_53 ( .A2(net_137), .A1(net_136), .ZN(net_119) );
CLKBUF_X2 inst_205 ( .A(net_156), .Z(net_199) );
CLKBUF_X2 inst_177 ( .A(net_170), .Z(net_171) );
CLKBUF_X2 inst_183 ( .A(net_176), .Z(net_177) );
DFFR_X2 inst_133 ( .RN(net_118), .D(net_106), .QN(net_10), .CK(net_164) );
NOR2_X2 inst_26 ( .ZN(net_81), .A1(net_5), .A2(CLR) );
CLKBUF_X2 inst_151 ( .A(net_144), .Z(net_145) );
INV_X2 inst_112 ( .ZN(net_13), .A(net_11) );
NAND2_X2 inst_64 ( .ZN(net_55), .A2(net_41), .A1(net_39) );
INV_X2 inst_107 ( .A(net_129), .ZN(net_128) );
NAND2_X2 inst_67 ( .ZN(net_73), .A2(net_65), .A1(net_49) );
CLKBUF_X2 inst_181 ( .A(net_165), .Z(net_175) );
DFFR_X2 inst_127 ( .RN(net_118), .D(net_78), .QN(net_8), .CK(net_198) );
NAND2_X2 inst_70 ( .ZN(net_91), .A2(net_84), .A1(net_63) );
CLKBUF_X2 inst_186 ( .A(net_179), .Z(net_180) );
DFFR_X2 inst_129 ( .QN(net_124), .RN(net_118), .D(net_77), .CK(net_196) );
INV_X4 inst_92 ( .A(net_29), .ZN(net_28) );
NOR2_X2 inst_29 ( .A2(net_34), .ZN(net_27), .A1(net_26) );
CLKBUF_X2 inst_189 ( .A(net_182), .Z(net_183) );
NOR3_X2 inst_17 ( .ZN(net_78), .A3(net_76), .A1(net_53), .A2(net_27) );
NOR3_X2 inst_11 ( .ZN(net_64), .A1(net_51), .A3(net_48), .A2(net_19) );
AND3_X2 inst_146 ( .A3(net_122), .ZN(net_114), .A1(net_111), .A2(net_109) );
CLKBUF_X2 inst_188 ( .A(net_167), .Z(net_182) );
NOR3_X2 inst_14 ( .ZN(net_72), .A3(net_60), .A1(net_33), .A2(net_21) );
CLKBUF_X2 inst_202 ( .A(net_195), .Z(net_196) );
CLKBUF_X2 inst_206 ( .A(net_199), .Z(net_200) );
CLKBUF_X2 inst_187 ( .A(net_180), .Z(net_181) );
INV_X1 inst_122 ( .ZN(net_26), .A(net_8) );
NOR2_X2 inst_31 ( .ZN(net_44), .A1(net_42), .A2(net_30) );
NOR2_X2 inst_25 ( .A2(net_127), .A1(net_124), .ZN(net_34) );
DFFR_X2 inst_126 ( .QN(net_127), .RN(net_118), .D(net_69), .CK(net_204) );
CLKBUF_X2 inst_158 ( .A(net_150), .Z(net_152) );
DFFR_X1 inst_141 ( .RN(net_118), .D(net_117), .QN(net_1), .CK(net_156) );
NAND2_X2 inst_62 ( .A2(net_133), .ZN(net_76), .A1(net_45) );
CLKBUF_X2 inst_200 ( .A(net_174), .Z(net_194) );
INV_X2 inst_110 ( .ZN(net_139), .A(net_125) );
NAND2_X2 inst_74 ( .ZN(net_96), .A1(net_95), .A2(net_85) );
NAND2_X2 inst_57 ( .ZN(net_140), .A2(net_11), .A1(net_10) );
NOR2_X2 inst_35 ( .A1(net_136), .ZN(net_90), .A2(net_11) );
INV_X4 inst_99 ( .A(net_66), .ZN(net_31) );
NAND3_X2 inst_48 ( .A2(net_139), .A1(net_138), .ZN(net_121), .A3(net_93) );
NAND2_X2 inst_69 ( .ZN(net_85), .A1(net_84), .A2(net_68) );
NAND3_X2 inst_46 ( .A2(net_109), .ZN(net_79), .A1(net_50), .A3(net_46) );
INV_X4 inst_82 ( .ZN(net_17), .A(CLR) );
DFFR_X1 inst_136 ( .RN(net_118), .D(net_82), .Q(GRN2), .CK(net_191) );
NOR2_X2 inst_30 ( .ZN(net_43), .A1(net_42), .A2(net_22) );
INV_X4 inst_102 ( .ZN(net_115), .A(net_111) );
INV_X2 inst_108 ( .ZN(net_143), .A(net_128) );
CLKBUF_X2 inst_165 ( .A(net_158), .Z(net_159) );
NOR2_X2 inst_32 ( .ZN(net_61), .A2(net_60), .A1(net_57) );
NOR3_X2 inst_22 ( .A1(net_115), .ZN(net_113), .A2(net_112), .A3(net_108) );
DFFR_X1 inst_144 ( .RN(net_118), .D(net_113), .QN(net_3), .CK(net_174) );
NOR2_X2 inst_34 ( .A2(net_131), .ZN(net_71), .A1(net_70) );
NOR3_X2 inst_12 ( .A2(net_58), .ZN(net_52), .A3(net_38), .A1(net_18) );
CLKBUF_X2 inst_195 ( .A(net_188), .Z(net_189) );
NAND2_X4 inst_56 ( .A1(net_121), .ZN(net_111), .A2(net_36) );
NAND2_X2 inst_71 ( .ZN(net_95), .A2(net_91), .A1(net_88) );
NOR3_X2 inst_21 ( .A3(net_143), .A1(net_142), .A2(net_112), .ZN(net_107) );
INV_X2 inst_104 ( .A(net_136), .ZN(net_134) );
NAND2_X2 inst_60 ( .A1(net_51), .ZN(net_37), .A2(net_36) );
CLKBUF_X2 inst_215 ( .A(net_208), .Z(net_209) );
CLKBUF_X2 inst_169 ( .A(net_162), .Z(net_163) );
CLKBUF_X2 inst_168 ( .A(net_161), .Z(net_162) );
INV_X4 inst_97 ( .ZN(net_35), .A(net_28) );
CLKBUF_X2 inst_161 ( .A(net_144), .Z(net_155) );
DFFR_X2 inst_124 ( .RN(net_118), .D(net_44), .QN(net_4), .CK(net_214) );
NOR3_X2 inst_18 ( .A1(net_134), .A3(net_104), .ZN(net_103), .A2(net_71) );
NOR3_X2 inst_16 ( .ZN(net_77), .A3(net_76), .A1(net_34), .A2(net_24) );
CLKBUF_X2 inst_208 ( .A(net_201), .Z(net_202) );
INV_X4 inst_88 ( .ZN(net_18), .A(net_17) );
CLKBUF_X2 inst_220 ( .A(net_213), .Z(net_214) );
XNOR2_X2 inst_3 ( .ZN(net_142), .A(net_94), .B(net_87) );
CLKBUF_X2 inst_156 ( .A(net_149), .Z(net_150) );
OR2_X4 inst_9 ( .ZN(net_60), .A1(net_35), .A2(net_1) );
INV_X2 inst_113 ( .ZN(net_14), .A(CLR) );
CLKBUF_X2 inst_170 ( .A(net_163), .Z(net_164) );
CLKBUF_X2 inst_198 ( .A(net_158), .Z(net_192) );
NAND2_X4 inst_50 ( .A1(net_133), .ZN(net_131), .A2(net_6) );
DFFR_X1 inst_137 ( .RN(net_118), .D(net_86), .Q(GRN1), .CK(net_181) );
CLKBUF_X2 inst_199 ( .A(net_192), .Z(net_193) );
NOR2_X1 inst_41 ( .ZN(net_122), .A2(net_100), .A1(net_92) );
DFFR_X2 inst_130 ( .RN(net_118), .D(net_91), .QN(net_5), .CK(net_186) );
INV_X4 inst_91 ( .A(net_58), .ZN(net_36) );
DFFR_X2 inst_132 ( .RN(net_118), .D(net_105), .QN(net_11), .CK(net_169) );
DFFR_X1 inst_143 ( .RN(net_118), .D(net_116), .QN(net_2), .CK(net_151) );
CLKBUF_X2 inst_176 ( .A(net_146), .Z(net_170) );
CLKBUF_X2 inst_152 ( .A(net_145), .Z(net_146) );
NAND2_X2 inst_58 ( .ZN(net_38), .A1(net_29), .A2(net_1) );
NOR2_X2 inst_36 ( .A2(net_135), .ZN(net_83), .A1(net_13) );
AND2_X4 inst_147 ( .ZN(net_32), .A2(net_14), .A1(net_2) );
INV_X4 inst_87 ( .ZN(net_57), .A(net_17) );
NAND2_X2 inst_61 ( .ZN(net_39), .A2(net_32), .A1(net_23) );
CLKBUF_X2 inst_203 ( .A(net_179), .Z(net_197) );
NAND3_X2 inst_45 ( .ZN(net_46), .A3(net_31), .A1(net_25), .A2(net_20) );
INV_X4 inst_96 ( .A(net_36), .ZN(net_25) );
CLKBUF_X2 inst_212 ( .A(net_205), .Z(net_206) );
INV_X4 inst_101 ( .ZN(net_62), .A(net_38) );
XOR2_X2 inst_0 ( .Z(net_22), .B(net_6), .A(TEST) );
CLKBUF_X2 inst_184 ( .A(net_174), .Z(net_178) );
NOR4_X2 inst_10 ( .ZN(net_82), .A1(net_81), .A3(net_80), .A2(net_61), .A4(net_59) );
XNOR2_X2 inst_4 ( .ZN(net_141), .A(net_98), .B(net_66) );
NAND2_X2 inst_65 ( .ZN(net_67), .A1(net_66), .A2(net_64) );
CLKBUF_X2 inst_178 ( .A(net_171), .Z(net_172) );
INV_X4 inst_89 ( .A(net_49), .ZN(net_20) );
NOR2_X2 inst_28 ( .A2(net_126), .A1(net_123), .ZN(net_24) );
INV_X2 inst_111 ( .A(net_124), .ZN(net_123) );
NAND2_X2 inst_66 ( .ZN(net_68), .A1(net_62), .A2(net_55) );
INV_X2 inst_117 ( .A(net_58), .ZN(net_23) );
INV_X4 inst_98 ( .A(net_109), .ZN(net_42) );
CLKBUF_X2 inst_190 ( .A(net_183), .Z(net_184) );
NAND2_X2 inst_63 ( .A2(net_62), .A1(net_51), .ZN(net_47) );
OR3_X4 inst_7 ( .A2(net_81), .A1(net_80), .ZN(net_74), .A3(net_52) );
CLKBUF_X2 inst_204 ( .A(net_162), .Z(net_198) );
CLKBUF_X2 inst_185 ( .A(net_178), .Z(net_179) );
CLKBUF_X2 inst_182 ( .A(net_175), .Z(net_176) );
NAND2_X4 inst_49 ( .ZN(net_133), .A1(net_120), .A2(net_40) );
INV_X2 inst_120 ( .ZN(net_65), .A(net_64) );
CLKBUF_X2 inst_154 ( .A(net_147), .Z(net_148) );
NOR3_X2 inst_13 ( .ZN(net_59), .A1(net_58), .A2(net_57), .A3(net_56) );
INV_X2 inst_119 ( .ZN(net_56), .A(net_35) );
NAND2_X2 inst_75 ( .ZN(net_97), .A2(net_95), .A1(net_74) );
CLKBUF_X2 inst_192 ( .A(net_185), .Z(net_186) );
CLKBUF_X2 inst_166 ( .A(net_159), .Z(net_160) );
INV_X2 inst_116 ( .ZN(net_21), .A(net_20) );
CLKBUF_X2 inst_163 ( .A(net_155), .Z(net_157) );
INV_X4 inst_85 ( .ZN(net_40), .A(net_7) );
NAND2_X4 inst_54 ( .ZN(net_130), .A1(net_119), .A2(net_87) );
INV_X4 inst_79 ( .ZN(net_19), .A(net_3) );
INV_X2 inst_109 ( .A(net_127), .ZN(net_126) );
INV_X2 inst_106 ( .A(net_130), .ZN(net_129) );
CLKBUF_X2 inst_219 ( .A(net_212), .Z(net_213) );
CLKBUF_X2 inst_201 ( .A(net_194), .Z(net_195) );
CLKBUF_X2 inst_193 ( .A(net_170), .Z(net_187) );
AND2_X2 inst_149 ( .ZN(net_94), .A2(net_90), .A1(net_15) );
NAND3_X2 inst_43 ( .A2(net_127), .A3(net_124), .ZN(net_120), .A1(net_8) );
NOR2_X2 inst_39 ( .ZN(net_116), .A2(net_115), .A1(net_110) );
DFFR_X2 inst_128 ( .RN(net_118), .D(net_75), .QN(net_7), .CK(net_197) );
NAND2_X2 inst_73 ( .ZN(net_138), .A1(net_129), .A2(net_66) );
CLKBUF_X2 inst_217 ( .A(net_210), .Z(net_211) );
NOR3_X2 inst_23 ( .ZN(net_117), .A1(net_115), .A2(net_112), .A3(net_101) );
CLKBUF_X2 inst_171 ( .A(net_163), .Z(net_165) );
INV_X4 inst_77 ( .ZN(net_51), .A(net_4) );
INV_X4 inst_94 ( .ZN(net_109), .A(net_57) );

endmodule
