module wb_dma (
x6157,
x5755,
x5143,
x3227,
x6456,
x5995,
x4866,
x4033,
x4926,
x3684,
x4435,
x4258,
x6706,
x6372,
x4251,
x3465,
x6678,
x54747,
x3314,
x5181,
x7007,
x6326,
x4066,
x4949,
x3954,
x7383,
x3365,
x4303,
x3067,
x3346,
x5078,
x4752,
x6358,
x5413,
x4148,
x6289,
x5846,
x4821,
x3261,
x4096,
x6367,
x6968,
x6430,
x6312,
x5386,
x4843,
x7215,
x7526,
x4118,
x7369,
x5913,
x7314,
x4008,
x3098,
x3884,
x5338,
x4323,
x4336,
x4129,
x4397,
x7345,
x6573,
x6400,
x3758,
x7329,
x4998,
x3865,
x4051,
x6298,
x5118,
x6623,
x3733,
x6334,
x4549,
x5468,
x3501,
x5370,
x5740,
x4502,
x4353,
x7087,
x5934,
x4283,
x7241,
x6650,
x4107,
x6122,
x6063,
x6503,
x4375,
x3986,
x7145,
x6319,
x4604,
x4790,
x3447,
x7404,
x5686,
x3997,
x7264,
x5058,
x5892,
x3527,
x3932,
x3145,
x6264,
x3819,
x5527,
x4658,
x3947,
x5957,
x4629,
x4080,
x4718,
x6880,
x6936,
x3134,
x3245,
x5247,
x3483,
x6039,
x3618,
x3669,
x7442,
x5507,
x3558,
x3338,
x3295,
x5868,
x3396,
x4040,
x4138,
x4206,
x6343,
x6303,
x6439,
x5712,
x3843,
x5269,
x3796,
x5020,
x5556,
x7509,
x3428,
x5628,
x7418,
x3961,
x3595,
x4524,
x6550,
x3976,
x4184,
x3277,
x6773,
x7169,
x3775,
x6727,
x5581,
x4175,
x5796,
x4476,
x7190,
x4022,
x6188,
x6845,
x5224,
x7120,
x5820,
x4578,
x7297,
x6389,
x3900,
x5294,
x4197,
x4089,
x6799,
x5317,
x6236,
x3907,
x7484,
x3190,
x3921,
x4461,
x6470,
x3580,
x6096,
x5448,
x7033,
x3383,
x6380,
x4974,
x6530,
x4164,
x4232,
x4266,
x3411,
x3636,
x5605,
x6908,
x5493,
x7061,
x6207,
x4155,
x7552,
x5429,
x4899,
x6592,
x7466,
x5779,
x6417,
x4690,
x3699,
x3651,
x4416,
x7544,
x5657,
x4219,
x902,
x1167,
x971,
x140,
x2846,
x2273,
x862,
x1105,
x2471,
x1387,
x2690,
x1144,
x950,
x317,
x1535,
x2706,
x962,
x734,
x125,
x1913,
x44,
x2304,
x1897,
x1587,
x835,
x499,
x1113,
x748,
x510,
x2149,
x2119,
x1285,
x1155,
x8,
x15,
x542,
x169,
x2528,
x2661,
x1071,
x2289,
x1701,
x957,
x2435,
x1007,
x2909,
x1266,
x1434,
x2993,
x1241,
x1097,
x1357,
x1663,
x342,
x1507,
x3041,
x2886,
x297,
x1682,
x2791,
x1029,
x255,
x132,
x108,
x2416,
x679,
x2071,
x535,
x1060,
x1578,
x788,
x651,
x1956,
x702,
x996,
x2016,
x421,
x2260,
x1415,
x910,
x2869,
x0,
x2483,
x722,
x627,
x2674,
x2773,
x491,
x2562,
x2175,
x934,
x2451,
x1230,
x234,
x1332,
x1306,
x2134,
x665,
x1218,
x518,
x1768,
x83,
x1086,
x1559,
x691,
x1520,
x760,
x2220,
x1548,
x2950,
x91,
x817,
x2579,
x1337,
x2098,
x1628,
x450,
x2971,
x1442,
x1811,
x381,
x2496,
x439,
x603,
x989,
x1425,
x1937,
x51,
x1322,
x615,
x1981,
x2592,
x1600,
x1451,
x2355,
x1018,
x2333,
x1693,
x1646,
x101,
x781,
x2739,
x398,
x2928,
x210,
x1402,
x878,
x1997,
x1877,
x596,
x925,
x1346,
x2371,
x2200,
x1854,
x768,
x1036,
x1474,
x807,
x1044,
x1195,
x2649,
x2050,
x192,
x2513,
x2233,
x1713,
x564,
x1277,
x1492,
x1462,
x361,
x828,
x1835,
x528,
x1124,
x2318,
x2403,
x550,
x476,
x1371,
x22,
x2611,
x886,
x2819,
x1176,
x638,
x1314,
x272,
x1739,
x2631,
x1794,
x2722,
x75,
x116,
x854,
x1613,
x1253,
x894,
x1294,
x870,
x582,
x1187,
x2543,
x844,
x406,
x711,
x461,
x1207,
x794,
x2752,
x1136,
x981,
x3020,
x1379);

// Start PIs
input x6157;
input x5755;
input x5143;
input x3227;
input x6456;
input x5995;
input x4866;
input x4033;
input x4926;
input x3684;
input x4435;
input x4258;
input x6706;
input x6372;
input x4251;
input x3465;
input x6678;
input x54747;
input x3314;
input x5181;
input x7007;
input x6326;
input x4066;
input x4949;
input x3954;
input x7383;
input x3365;
input x4303;
input x3067;
input x3346;
input x5078;
input x4752;
input x6358;
input x5413;
input x4148;
input x6289;
input x5846;
input x4821;
input x3261;
input x4096;
input x6367;
input x6968;
input x6430;
input x6312;
input x5386;
input x4843;
input x7215;
input x7526;
input x4118;
input x7369;
input x5913;
input x7314;
input x4008;
input x3098;
input x3884;
input x5338;
input x4323;
input x4336;
input x4129;
input x4397;
input x7345;
input x6573;
input x6400;
input x3758;
input x7329;
input x4998;
input x3865;
input x4051;
input x6298;
input x5118;
input x6623;
input x3733;
input x6334;
input x4549;
input x5468;
input x3501;
input x5370;
input x5740;
input x4502;
input x4353;
input x7087;
input x5934;
input x4283;
input x7241;
input x6650;
input x4107;
input x6122;
input x6063;
input x6503;
input x4375;
input x3986;
input x7145;
input x6319;
input x4604;
input x4790;
input x3447;
input x7404;
input x5686;
input x3997;
input x7264;
input x5058;
input x5892;
input x3527;
input x3932;
input x3145;
input x6264;
input x3819;
input x5527;
input x4658;
input x3947;
input x5957;
input x4629;
input x4080;
input x4718;
input x6880;
input x6936;
input x3134;
input x3245;
input x5247;
input x3483;
input x6039;
input x3618;
input x3669;
input x7442;
input x5507;
input x3558;
input x3338;
input x3295;
input x5868;
input x3396;
input x4040;
input x4138;
input x4206;
input x6343;
input x6303;
input x6439;
input x5712;
input x3843;
input x5269;
input x3796;
input x5020;
input x5556;
input x7509;
input x3428;
input x5628;
input x7418;
input x3961;
input x3595;
input x4524;
input x6550;
input x3976;
input x4184;
input x3277;
input x6773;
input x7169;
input x3775;
input x6727;
input x5581;
input x4175;
input x5796;
input x4476;
input x7190;
input x4022;
input x6188;
input x6845;
input x5224;
input x7120;
input x5820;
input x4578;
input x7297;
input x6389;
input x3900;
input x5294;
input x4197;
input x4089;
input x6799;
input x5317;
input x6236;
input x3907;
input x7484;
input x3190;
input x3921;
input x4461;
input x6470;
input x3580;
input x6096;
input x5448;
input x7033;
input x3383;
input x6380;
input x4974;
input x6530;
input x4164;
input x4232;
input x4266;
input x3411;
input x3636;
input x5605;
input x6908;
input x5493;
input x7061;
input x6207;
input x4155;
input x7552;
input x5429;
input x4899;
input x6592;
input x7466;
input x5779;
input x6417;
input x4690;
input x3699;
input x3651;
input x4416;
input x7544;
input x5657;
input x4219;

// Start POs
output x902;
output x1167;
output x971;
output x140;
output x2846;
output x2273;
output x862;
output x1105;
output x2471;
output x1387;
output x2690;
output x1144;
output x950;
output x317;
output x1535;
output x2706;
output x962;
output x734;
output x125;
output x1913;
output x44;
output x2304;
output x1897;
output x1587;
output x835;
output x499;
output x1113;
output x748;
output x510;
output x2149;
output x2119;
output x1285;
output x1155;
output x8;
output x15;
output x542;
output x169;
output x2528;
output x2661;
output x1071;
output x2289;
output x1701;
output x957;
output x2435;
output x1007;
output x2909;
output x1266;
output x1434;
output x2993;
output x1241;
output x1097;
output x1357;
output x1663;
output x342;
output x1507;
output x3041;
output x2886;
output x297;
output x1682;
output x2791;
output x1029;
output x255;
output x132;
output x108;
output x2416;
output x679;
output x2071;
output x535;
output x1060;
output x1578;
output x788;
output x651;
output x1956;
output x702;
output x996;
output x2016;
output x421;
output x2260;
output x1415;
output x910;
output x2869;
output x0;
output x2483;
output x722;
output x627;
output x2674;
output x2773;
output x491;
output x2562;
output x2175;
output x934;
output x2451;
output x1230;
output x234;
output x1332;
output x1306;
output x2134;
output x665;
output x1218;
output x518;
output x1768;
output x83;
output x1086;
output x1559;
output x691;
output x1520;
output x760;
output x2220;
output x1548;
output x2950;
output x91;
output x817;
output x2579;
output x1337;
output x2098;
output x1628;
output x450;
output x2971;
output x1442;
output x1811;
output x381;
output x2496;
output x439;
output x603;
output x989;
output x1425;
output x1937;
output x51;
output x1322;
output x615;
output x1981;
output x2592;
output x1600;
output x1451;
output x2355;
output x1018;
output x2333;
output x1693;
output x1646;
output x101;
output x781;
output x2739;
output x398;
output x2928;
output x210;
output x1402;
output x878;
output x1997;
output x1877;
output x596;
output x925;
output x1346;
output x2371;
output x2200;
output x1854;
output x768;
output x1036;
output x1474;
output x807;
output x1044;
output x1195;
output x2649;
output x2050;
output x192;
output x2513;
output x2233;
output x1713;
output x564;
output x1277;
output x1492;
output x1462;
output x361;
output x828;
output x1835;
output x528;
output x1124;
output x2318;
output x2403;
output x550;
output x476;
output x1371;
output x22;
output x2611;
output x886;
output x2819;
output x1176;
output x638;
output x1314;
output x272;
output x1739;
output x2631;
output x1794;
output x2722;
output x75;
output x116;
output x854;
output x1613;
output x1253;
output x894;
output x1294;
output x870;
output x582;
output x1187;
output x2543;
output x844;
output x406;
output x711;
output x461;
output x1207;
output x794;
output x2752;
output x1136;
output x981;
output x3020;
output x1379;

// Start wires
wire net_2449;
wire net_1317;
wire net_416;
wire net_215;
wire net_2394;
wire x971;
wire net_2418;
wire net_1382;
wire net_943;
wire net_1897;
wire net_980;
wire net_53;
wire net_3498;
wire net_2542;
wire net_1786;
wire net_1377;
wire net_3996;
wire x3346;
wire net_1393;
wire net_2169;
wire net_1324;
wire net_2256;
wire x1701;
wire net_264;
wire net_3904;
wire net_2207;
wire net_263;
wire net_3527;
wire net_1138;
wire net_2769;
wire net_3483;
wire net_3707;
wire net_1064;
wire net_2082;
wire net_3292;
wire net_1439;
wire x2791;
wire net_1778;
wire net_508;
wire net_1090;
wire net_3685;
wire net_703;
wire net_193;
wire net_201;
wire net_2942;
wire net_3817;
wire net_3280;
wire net_3085;
wire net_2896;
wire net_3281;
wire net_3949;
wire net_3134;
wire net_1852;
wire net_1720;
wire net_1555;
wire net_3818;
wire net_3434;
wire x2562;
wire net_2060;
wire net_2051;
wire net_2780;
wire net_789;
wire net_3756;
wire net_3244;
wire net_593;
wire net_2171;
wire net_2765;
wire x817;
wire net_3833;
wire net_742;
wire net_2425;
wire x2496;
wire net_2830;
wire net_1198;
wire net_2509;
wire net_3975;
wire net_2862;
wire net_1860;
wire x1981;
wire net_2457;
wire net_883;
wire net_2156;
wire net_1432;
wire net_1312;
wire x2333;
wire net_2957;
wire net_446;
wire net_1516;
wire net_1712;
wire x596;
wire net_3063;
wire net_1083;
wire net_3546;
wire net_3343;
wire net_3423;
wire net_1499;
wire net_964;
wire net_3326;
wire net_1453;
wire net_2913;
wire net_3295;
wire x564;
wire net_2239;
wire net_3394;
wire net_3542;
wire net_2268;
wire net_634;
wire net_2846;
wire net_2303;
wire net_371;
wire net_3903;
wire net_1735;
wire net_2787;
wire net_2210;
wire net_2176;
wire net_1571;
wire net_2466;
wire net_997;
wire x116;
wire net_256;
wire net_3959;
wire net_850;
wire net_1140;
wire net_2764;
wire net_1464;
wire net_679;
wire net_1168;
wire net_2680;
wire net_3196;
wire net_308;
wire net_515;
wire net_3090;
wire net_3987;
wire net_223;
wire net_1009;
wire net_715;
wire net_2077;
wire net_890;
wire net_2219;
wire net_2745;
wire net_2546;
wire net_3965;
wire net_1876;
wire net_2471;
wire net_312;
wire net_2404;
wire net_130;
wire net_2627;
wire net_572;
wire net_147;
wire net_481;
wire net_369;
wire net_1662;
wire net_1079;
wire net_3935;
wire net_2444;
wire net_2809;
wire net_1188;
wire x2909;
wire net_3235;
wire net_780;
wire net_3586;
wire net_3184;
wire net_1446;
wire net_541;
wire net_1251;
wire net_2391;
wire net_2802;
wire net_2906;
wire net_456;
wire net_155;
wire net_1697;
wire net_3850;
wire net_1753;
wire x6334;
wire net_349;
wire net_2435;
wire net_245;
wire net_3428;
wire net_1409;
wire net_2383;
wire net_2977;
wire x5934;
wire net_493;
wire net_3491;
wire x996;
wire net_1428;
wire net_987;
wire x910;
wire net_277;
wire net_1965;
wire net_3620;
wire x5058;
wire net_89;
wire net_3071;
wire net_2350;
wire net_3271;
wire net_680;
wire x4080;
wire net_338;
wire x1218;
wire net_2998;
wire net_721;
wire net_243;
wire net_3226;
wire net_3143;
wire net_2757;
wire net_1018;
wire net_3629;
wire net_2854;
wire net_2009;
wire net_2369;
wire net_2038;
wire net_4026;
wire net_823;
wire net_106;
wire net_1380;
wire net_1676;
wire x3295;
wire net_698;
wire net_1915;
wire net_1191;
wire net_2255;
wire net_2485;
wire net_3857;
wire net_1997;
wire net_138;
wire net_749;
wire net_1019;
wire net_1948;
wire net_1616;
wire x4476;
wire net_1006;
wire net_2781;
wire net_2969;
wire net_1418;
wire net_3202;
wire net_2985;
wire net_537;
wire net_3056;
wire net_1713;
wire x272;
wire net_3614;
wire net_2668;
wire net_2677;
wire net_3252;
wire x75;
wire net_2775;
wire net_513;
wire net_3916;
wire net_163;
wire net_1576;
wire net_1421;
wire net_3407;
wire net_2736;
wire net_2127;
wire net_1280;
wire net_459;
wire net_3656;
wire net_737;
wire net_2284;
wire net_3412;
wire net_2113;
wire x7544;
wire net_3990;
wire net_2193;
wire net_3856;
wire x1167;
wire net_3915;
wire net_1886;
wire net_1156;
wire net_2604;
wire net_1966;
wire net_3501;
wire net_101;
wire net_1659;
wire net_1272;
wire net_326;
wire net_2381;
wire net_2109;
wire net_1770;
wire net_4001;
wire net_3505;
wire net_589;
wire net_655;
wire x1007;
wire x5913;
wire net_3536;
wire net_1814;
wire net_3175;
wire net_378;
wire net_2829;
wire net_724;
wire net_3309;
wire net_3142;
wire net_3036;
wire net_423;
wire net_1219;
wire x5118;
wire net_328;
wire net_2384;
wire net_3884;
wire net_1958;
wire net_1931;
wire net_3736;
wire net_2877;
wire net_2480;
wire net_3294;
wire net_1549;
wire net_3016;
wire net_874;
wire net_2929;
wire net_1632;
wire net_3796;
wire net_1661;
wire net_1236;
wire net_818;
wire net_3749;
wire net_3674;
wire net_2746;
wire net_2700;
wire net_1211;
wire net_1183;
wire net_2594;
wire net_1488;
wire net_2812;
wire net_1684;
wire net_811;
wire net_352;
wire net_3920;
wire net_1462;
wire net_436;
wire net_2837;
wire net_2017;
wire net_2824;
wire net_1777;
wire net_1926;
wire x4138;
wire net_3115;
wire net_2735;
wire net_1641;
wire net_3518;
wire x5628;
wire net_1621;
wire net_3680;
wire net_3984;
wire net_3615;
wire net_1702;
wire net_1103;
wire net_1035;
wire net_767;
wire net_3055;
wire net_1838;
wire net_131;
wire net_358;
wire net_1973;
wire net_3593;
wire net_3095;
wire net_2845;
wire net_2016;
wire net_2934;
wire net_2641;
wire net_1763;
wire net_3125;
wire net_1285;
wire net_3112;
wire net_1175;
wire x476;
wire net_2882;
wire net_3278;
wire net_2922;
wire net_1513;
wire net_1742;
wire net_3064;
wire net_2276;
wire x3383;
wire x854;
wire x1613;
wire x6380;
wire x4232;
wire x4266;
wire net_468;
wire net_798;
wire net_3135;
wire net_73;
wire x4899;
wire net_2059;
wire net_3370;
wire net_1899;
wire x4219;
wire net_1336;
wire net_3947;
wire net_3441;
wire net_179;
wire net_61;
wire net_4015;
wire net_3662;
wire net_1843;
wire net_62;
wire net_3261;
wire net_534;
wire net_3793;
wire net_3336;
wire net_2289;
wire net_903;
wire x1913;
wire net_1551;
wire net_486;
wire x1587;
wire x835;
wire net_3539;
wire net_2031;
wire net_1868;
wire net_1560;
wire net_406;
wire net_2378;
wire net_3863;
wire net_3640;
wire net_3382;
wire x4008;
wire net_1545;
wire net_748;
wire net_95;
wire net_990;
wire net_3958;
wire net_2327;
wire net_1003;
wire net_514;
wire net_2332;
wire net_3645;
wire net_3774;
wire net_1604;
wire net_2715;
wire net_1803;
wire net_1941;
wire net_524;
wire net_1134;
wire net_3899;
wire net_3742;
wire net_363;
wire net_445;
wire net_1319;
wire net_776;
wire net_3080;
wire net_2508;
wire x4375;
wire net_44;
wire net_1650;
wire net_1582;
wire net_3748;
wire x2483;
wire net_3149;
wire net_1675;
wire net_4016;
wire net_2247;
wire x3145;
wire net_2333;
wire net_2213;
wire net_1368;
wire net_2575;
wire net_1248;
wire net_2291;
wire net_1097;
wire net_2238;
wire net_845;
wire net_762;
wire net_3589;
wire net_695;
wire net_2525;
wire net_1201;
wire net_3713;
wire net_556;
wire net_2671;
wire net_3330;
wire net_893;
wire net_255;
wire net_3826;
wire net_859;
wire net_620;
wire net_619;
wire x989;
wire net_1167;
wire net_3932;
wire net_2198;
wire net_1044;
wire x3277;
wire net_3444;
wire net_3800;
wire net_2940;
wire x5796;
wire net_2043;
wire net_2095;
wire net_3285;
wire net_68;
wire net_2314;
wire net_2613;
wire net_1493;
wire net_3605;
wire net_976;
wire x4197;
wire net_2709;
wire x1713;
wire net_865;
wire net_611;
wire net_231;
wire net_3514;
wire net_2621;
wire net_2579;
wire net_3024;
wire net_1223;
wire net_2750;
wire net_1866;
wire x4461;
wire net_926;
wire net_3692;
wire net_3211;
wire net_2160;
wire net_3477;
wire net_391;
wire net_2297;
wire net_3325;
wire x3411;
wire net_2048;
wire net_582;
wire x461;
wire net_2341;
wire net_661;
wire net_3633;
wire net_3360;
wire net_2516;
wire x6157;
wire net_2807;
wire net_1141;
wire net_3561;
wire net_3243;
wire net_1543;
wire net_1295;
wire x4435;
wire net_2104;
wire x2690;
wire net_1288;
wire net_2071;
wire net_1923;
wire net_1275;
wire net_210;
wire net_2766;
wire net_3771;
wire net_2417;
wire net_2300;
wire net_916;
wire net_3395;
wire net_741;
wire net_940;
wire net_851;
wire net_3719;
wire net_2426;
wire net_3789;
wire x2661;
wire x6367;
wire net_3310;
wire net_1043;
wire net_671;
wire net_2850;
wire net_770;
wire net_1005;
wire net_1059;
wire net_1630;
wire net_3891;
wire net_1454;
wire net_2956;
wire net_307;
wire net_1796;
wire net_1082;
wire net_3342;
wire net_3547;
wire net_1550;
wire net_3543;
wire net_2310;
wire net_1507;
wire x3501;
wire net_3296;
wire net_257;
wire net_233;
wire x5740;
wire net_474;
wire net_3459;
wire net_2656;
wire net_958;
wire x6650;
wire net_1268;
wire net_3922;
wire net_3212;
wire net_3780;
wire net_1115;
wire net_944;
wire net_1734;
wire net_1764;
wire net_961;
wire net_3513;
wire net_2106;
wire net_3335;
wire x491;
wire net_3682;
wire net_3050;
wire net_1728;
wire net_63;
wire net_3327;
wire x1768;
wire net_3956;
wire net_2667;
wire net_3456;
wire x3134;
wire net_425;
wire net_287;
wire net_189;
wire net_1586;
wire net_2205;
wire net_3755;
wire x1628;
wire net_480;
wire net_216;
wire net_2897;
wire net_433;
wire net_2881;
wire net_836;
wire net_2161;
wire net_368;
wire net_224;
wire net_52;
wire net_1898;
wire x2592;
wire net_608;
wire net_1212;
wire net_3604;
wire net_370;
wire net_2000;
wire net_3706;
wire net_2984;
wire net_1120;
wire net_1020;
wire x6845;
wire net_2848;
wire net_3282;
wire net_3122;
wire net_1169;
wire net_973;
wire net_1139;
wire net_3902;
wire net_2206;
wire net_1392;
wire net_1574;
wire net_2094;
wire net_2543;
wire net_311;
wire net_760;
wire net_2479;
wire net_2083;
wire net_3851;
wire net_873;
wire net_2488;
wire net_1811;
wire net_154;
wire net_3699;
wire net_2588;
wire net_1870;
wire x1314;
wire net_704;
wire net_2520;
wire net_1478;
wire net_2179;
wire net_1696;
wire net_587;
wire net_1262;
wire net_2063;
wire net_3997;
wire net_4027;
wire net_192;
wire net_1739;
wire net_1356;
wire net_2912;
wire net_2197;
wire x870;
wire net_3816;
wire net_735;
wire x4155;
wire net_2905;
wire net_1907;
wire net_3809;
wire net_1711;
wire net_200;
wire net_2084;
wire x4690;
wire x4416;
wire net_195;
wire net_1081;
wire net_1853;
wire net_2037;
wire net_2170;
wire net_1237;
wire net_1420;
wire x3465;
wire net_2678;
wire x962;
wire net_3761;
wire net_3144;
wire net_699;
wire net_242;
wire net_359;
wire net_2526;
wire net_2819;
wire net_1644;
wire net_2864;
wire net_2800;
wire net_882;
wire net_1998;
wire net_1827;
wire net_3225;
wire net_1190;
wire net_3858;
wire net_2795;
wire net_1311;
wire net_2283;
wire net_1207;
wire net_1918;
wire x3758;
wire net_2121;
wire net_2191;
wire net_3236;
wire net_3201;
wire net_3558;
wire net_2252;
wire net_555;
wire net_1613;
wire x4502;
wire net_790;
wire net_2126;
wire x6063;
wire net_1577;
wire net_1417;
wire net_1054;
wire x0;
wire net_2386;
wire net_2727;
wire net_2166;
wire net_3650;
wire net_2465;
wire net_2257;
wire net_3418;
wire net_3655;
wire net_2304;
wire net_898;
wire net_2968;
wire net_2643;
wire net_1593;
wire x3618;
wire net_714;
wire net_2999;
wire net_1309;
wire net_3722;
wire net_3380;
wire net_683;
wire net_1771;
wire net_148;
wire net_1376;
wire net_1517;
wire x5269;
wire net_1980;
wire x615;
wire x7418;
wire net_1302;
wire net_2076;
wire net_244;
wire net_2218;
wire net_2395;
wire net_1690;
wire net_1078;
wire x6188;
wire net_4002;
wire net_1989;
wire x2928;
wire net_2997;
wire net_2855;
wire net_2093;
wire net_1795;
wire net_2403;
wire net_1539;
wire x6389;
wire net_3490;
wire net_3035;
wire net_2355;
wire net_3262;
wire net_1548;
wire net_810;
wire net_92;
wire net_394;
wire net_3778;
wire net_2536;
wire net_1189;
wire net_139;
wire net_409;
wire net_2949;
wire net_3429;
wire net_1469;
wire net_3470;
wire net_88;
wire net_1708;
wire net_2436;
wire net_81;
wire net_3974;
wire x711;
wire net_3419;
wire net_2976;
wire net_722;
wire net_988;
wire net_1254;
wire net_3621;
wire net_621;
wire net_435;
wire net_1830;
wire x140;
wire net_132;
wire x2471;
wire x1387;
wire net_105;
wire net_2838;
wire net_1649;
wire net_1837;
wire net_1841;
wire net_1249;
wire net_2427;
wire net_3378;
wire net_1071;
wire net_3985;
wire x3954;
wire net_3163;
wire net_327;
wire net_3877;
wire net_1701;
wire net_999;
wire x3261;
wire net_353;
wire net_822;
wire net_1633;
wire net_3588;
wire net_1974;
wire net_1480;
wire net_319;
wire net_2670;
wire net_1743;
wire net_3046;
wire net_2597;
wire net_164;
wire x1682;
wire net_377;
wire net_87;
wire net_1544;
wire net_288;
wire net_2649;
wire net_3096;
wire net_1629;
wire net_1459;
wire net_3277;
wire net_805;
wire net_3741;
wire net_3590;
wire net_2923;
wire net_2151;
wire net_540;
wire net_512;
wire net_2688;
wire net_2642;
wire net_1174;
wire net_1622;
wire net_891;
wire net_1109;
wire net_3065;
wire net_3102;
wire net_3457;
wire x3932;
wire net_1102;
wire x5527;
wire x4629;
wire net_3371;
wire net_618;
wire net_2244;
wire net_2692;
wire net_3688;
wire net_3777;
wire net_1875;
wire net_3420;
wire net_783;
wire net_3887;
wire net_1487;
wire net_754;
wire net_2759;
wire net_2605;
wire net_921;
wire net_3634;
wire net_550;
wire x3961;
wire net_3308;
wire net_2835;
wire net_3991;
wire net_2192;
wire net_1533;
wire x1018;
wire net_1240;
wire net_461;
wire net_3000;
wire net_3502;
wire net_2564;
wire net_2821;
wire net_1512;
wire net_1658;
wire net_654;
wire net_858;
wire net_330;
wire net_1330;
wire net_3506;
wire net_3007;
wire net_3015;
wire net_1785;
wire net_3174;
wire net_2876;
wire net_570;
wire net_444;
wire net_525;
wire net_844;
wire net_3829;
wire net_3646;
wire net_1496;
wire net_1210;
wire net_1067;
wire net_325;
wire net_3735;
wire net_1820;
wire net_1427;
wire net_3921;
wire net_985;
wire net_3933;
wire x6530;
wire net_424;
wire net_1521;
wire net_1729;
wire net_3353;
wire net_1677;
wire x3651;
wire net_2991;
wire net_564;
wire net_3639;
wire net_2050;
wire x4866;
wire net_2811;
wire net_3086;
wire net_2058;
wire net_813;
wire net_3045;
wire net_1178;
wire net_2612;
wire net_1027;
wire net_2018;
wire net_3825;
wire net_2042;
wire net_340;
wire net_1408;
wire net_2510;
wire net_265;
wire net_2634;
wire net_434;
wire net_3808;
wire net_1797;
wire net_3488;
wire net_3023;
wire net_1202;
wire net_69;
wire x7526;
wire net_1155;
wire net_925;
wire net_339;
wire net_2279;
wire net_3447;
wire net_3468;
wire net_2695;
wire net_864;
wire x6400;
wire net_2710;
wire net_2660;
wire net_2298;
wire net_660;
wire x2071;
wire net_3671;
wire net_102;
wire net_2313;
wire net_59;
wire net_3691;
wire net_1908;
wire net_3217;
wire net_1291;
wire net_230;
wire net_1865;
wire net_3383;
wire net_678;
wire net_3349;
wire net_1222;
wire net_3404;
wire net_928;
wire net_3810;
wire net_3914;
wire net_2578;
wire net_208;
wire net_2744;
wire net_2377;
wire net_1433;
wire net_415;
wire net_116;
wire net_3251;
wire net_2786;
wire net_347;
wire net_3794;
wire x7442;
wire net_3440;
wire net_3358;
wire net_1776;
wire net_2145;
wire x6343;
wire net_3368;
wire net_1335;
wire net_2574;
wire net_4014;
wire net_3311;
wire net_3531;
wire net_3747;
wire net_2212;
wire net_2132;
wire net_2292;
wire net_1880;
wire net_3862;
wire net_184;
wire net_3571;
wire net_610;
wire net_1844;
wire net_389;
wire net_3538;
wire net_902;
wire net_1867;
wire net_2344;
wire net_1323;
wire net_2650;
wire net_1949;
wire net_1506;
wire x1474;
wire net_1583;
wire net_736;
wire net_1804;
wire net_539;
wire net_2331;
wire net_692;
wire net_1563;
wire net_3898;
wire x528;
wire net_3361;
wire net_1365;
wire net_1135;
wire x3190;
wire net_1346;
wire net_43;
wire x2819;
wire net_1942;
wire net_1801;
wire net_1400;
wire net_885;
wire x1739;
wire net_1267;
wire net_3944;
wire net_3661;
wire x894;
wire net_869;
wire net_3714;
wire net_669;
wire net_937;
wire net_2441;
wire net_3517;
wire net_2349;
wire net_761;
wire net_496;
wire x5429;
wire net_1554;
wire x1207;
wire net_479;
wire net_1294;
wire x981;
wire net_2459;
wire net_2030;
wire net_3520;
wire net_1587;
wire x5755;
wire net_1354;
wire net_2904;
wire net_796;
wire net_1308;
wire net_2249;
wire net_648;
wire net_1389;
wire net_739;
wire net_3250;
wire net_2548;
wire net_2075;
wire net_826;
wire net_1738;
wire net_3658;
wire net_548;
wire net_3359;
wire net_2402;
wire net_2624;
wire net_636;
wire net_343;
wire net_511;
wire net_3967;
wire net_1961;
wire net_1260;
wire net_2654;
wire net_2487;
wire net_2911;
wire net_1819;
wire net_1185;
wire x6298;
wire net_239;
wire net_310;
wire net_2975;
wire x788;
wire net_2437;
wire net_2779;
wire net_1912;
wire net_1490;
wire net_682;
wire net_989;
wire net_1963;
wire x3527;
wire net_1538;
wire net_108;
wire net_458;
wire x2175;
wire net_685;
wire x4718;
wire net_3560;
wire x1520;
wire net_1007;
wire x1548;
wire net_1579;
wire net_1292;
wire net_1999;
wire net_1014;
wire net_2796;
wire net_1444;
wire net_2679;
wire net_4024;
wire net_3410;
wire net_2111;
wire net_1946;
wire net_2733;
wire net_538;
wire net_3612;
wire net_1605;
wire net_1937;
wire net_2535;
wire net_3191;
wire x3775;
wire x7169;
wire net_366;
wire net_1956;
wire net_1854;
wire net_1917;
wire x1693;
wire net_1614;
wire net_1755;
wire net_747;
wire net_1359;
wire net_2305;
wire net_1653;
wire net_2460;
wire net_2983;
wire net_3209;
wire net_2258;
wire net_1647;
wire net_198;
wire x2233;
wire x2513;
wire x4089;
wire net_209;
wire net_1282;
wire net_294;
wire net_2367;
wire net_2892;
wire net_2810;
wire net_2429;
wire net_3204;
wire net_1265;
wire net_1053;
wire net_1004;
wire net_3471;
wire net_848;
wire net_1080;
wire net_1619;
wire net_3232;
wire net_2124;
wire net_1890;
wire net_3512;
wire net_1161;
wire net_82;
wire net_3228;
wire net_2282;
wire net_2430;
wire net_2357;
wire x406;
wire net_1395;
wire net_1546;
wire net_3481;
wire net_1589;
wire net_1046;
wire x4926;
wire x2273;
wire net_606;
wire net_3906;
wire net_623;
wire net_2396;
wire net_663;
wire net_1213;
wire net_1891;
wire net_2265;
wire net_3998;
wire net_579;
wire net_2445;
wire net_769;
wire net_3396;
wire net_1780;
wire net_2062;
wire net_2856;
wire x8;
wire net_787;
wire net_3603;
wire net_2894;
wire net_1025;
wire net_3758;
wire net_1988;
wire net_3718;
wire net_1518;
wire net_1089;
wire net_1194;
wire net_1437;
wire net_3579;
wire net_3525;
wire net_1664;
wire net_705;
wire net_2139;
wire net_1608;
wire net_506;
wire net_3769;
wire net_2948;
wire net_1910;
wire net_3775;
wire net_1036;
wire net_3544;
wire net_3034;
wire net_1196;
wire net_3973;
wire net_2493;
wire net_919;
wire net_3626;
wire net_290;
wire net_4008;
wire net_3313;
wire net_3136;
wire net_2209;
wire net_1372;
wire net_1757;
wire net_3834;
wire net_3591;
wire net_3152;
wire net_2682;
wire x2098;
wire net_3648;
wire net_140;
wire net_740;
wire net_1722;
wire net_2329;
wire x5868;
wire net_3790;
wire net_2150;
wire net_2008;
wire net_2065;
wire net_3183;
wire net_2927;
wire net_2808;
wire x5020;
wire net_3908;
wire net_194;
wire net_2178;
wire net_730;
wire net_1128;
wire net_3073;
wire net_2713;
wire net_2105;
wire net_1127;
wire net_804;
wire net_1119;
wire net_3548;
wire net_1314;
wire net_957;
wire net_1287;
wire x210;
wire net_2726;
wire net_531;
wire x1346;
wire net_77;
wire net_499;
wire net_3345;
wire net_2752;
wire net_49;
wire net_1340;
wire net_3123;
wire net_2955;
wire net_71;
wire net_3328;
wire x828;
wire net_771;
wire net_3534;
wire net_1765;
wire net_2844;
wire net_2301;
wire net_2978;
wire x7484;
wire x22;
wire net_2107;
wire net_180;
wire net_3950;
wire net_51;
wire net_2774;
wire net_2420;
wire net_4028;
wire net_2860;
wire net_432;
wire net_1979;
wire x7033;
wire net_1062;
wire net_3731;
wire net_3290;
wire net_3293;
wire net_1142;
wire net_1460;
wire net_1475;
wire net_1451;
wire net_3159;
wire x6908;
wire net_67;
wire net_2240;
wire net_2416;
wire x2752;
wire x6417;
wire net_203;
wire net_1411;
wire net_2173;
wire net_505;
wire net_3723;
wire x6456;
wire net_1602;
wire net_4013;
wire net_992;
wire net_237;
wire net_613;
wire net_782;
wire net_2144;
wire net_2236;
wire net_3744;
wire x3314;
wire net_1095;
wire net_3443;
wire net_578;
wire net_3314;
wire net_3945;
wire net_2971;
wire x510;
wire net_1558;
wire net_2743;
wire net_2836;
wire net_1505;
wire net_1805;
wire net_2159;
wire net_388;
wire net_3952;
wire net_3669;
wire net_1861;
wire net_3647;
wire net_3635;
wire net_536;
wire net_455;
wire net_1332;
wire x1663;
wire net_221;
wire net_1594;
wire net_115;
wire net_3339;
wire net_3276;
wire net_1110;
wire net_393;
wire net_442;
wire net_542;
wire net_1832;
wire net_408;
wire net_1026;
wire net_3246;
wire net_2215;
wire net_1845;
wire net_2573;
wire net_3087;
wire net_2376;
wire net_1520;
wire net_1821;
wire net_3993;
wire net_3390;
wire net_1401;
wire net_3865;
wire net_2372;
wire net_1588;
wire net_3909;
wire net_66;
wire net_3937;
wire net_868;
wire net_1495;
wire net_2992;
wire net_3664;
wire net_3233;
wire x627;
wire net_443;
wire net_3522;
wire net_270;
wire net_522;
wire net_922;
wire net_2638;
wire net_668;
wire net_3079;
wire net_1584;
wire net_1990;
wire net_2330;
wire net_2264;
wire x6039;
wire net_977;
wire net_643;
wire net_3397;
wire net_1070;
wire net_1225;
wire net_622;
wire net_812;
wire x3558;
wire net_3587;
wire net_3762;
wire x6439;
wire x5712;
wire net_3687;
wire net_2857;
wire net_1107;
wire net_2767;
wire net_1338;
wire net_3874;
wire net_2045;
wire net_2053;
wire net_3384;
wire net_2180;
wire net_1203;
wire net_2869;
wire net_3332;
wire net_825;
wire net_3446;
wire net_1892;
wire net_1798;
wire net_3220;
wire net_2119;
wire net_309;
wire x1997;
wire net_1366;
wire net_837;
wire net_3469;
wire net_2615;
wire x7297;
wire x1036;
wire net_927;
wire net_2007;
wire net_1151;
wire net_713;
wire net_693;
wire net_1519;
wire x6236;
wire net_729;
wire net_3964;
wire net_3213;
wire net_2818;
wire net_863;
wire net_3164;
wire net_580;
wire net_2136;
wire net_904;
wire net_2339;
wire net_341;
wire net_58;
wire net_1879;
wire net_970;
wire net_488;
wire net_2319;
wire net_3044;
wire net_1532;
wire net_1160;
wire net_159;
wire net_3268;
wire net_2163;
wire net_3417;
wire net_3307;
wire net_553;
wire net_1093;
wire net_2592;
wire net_2875;
wire net_763;
wire net_3580;
wire net_3259;
wire x2149;
wire net_1740;
wire net_324;
wire x4148;
wire x6289;
wire net_710;
wire net_418;
wire net_462;
wire net_872;
wire net_3097;
wire net_161;
wire net_3066;
wire net_3970;
wire x2886;
wire net_3018;
wire net_2606;
wire net_173;
wire net_1486;
wire net_3880;
wire net_78;
wire net_2320;
wire net_1839;
wire net_1665;
wire net_3006;
wire net_376;
wire net_2133;
wire net_1681;
wire x535;
wire x1060;
wire net_3550;
wire net_2515;
wire net_1812;
wire net_3173;
wire net_3738;
wire net_2224;
wire net_3203;
wire net_422;
wire net_1345;
wire net_1450;
wire net_561;
wire net_2659;
wire net_2589;
wire net_1700;
wire net_591;
wire net_746;
wire net_2290;
wire net_1274;
wire net_2458;
wire net_1682;
wire net_2851;
wire net_178;
wire net_3435;
wire net_2843;
wire net_3466;
wire net_2635;
wire net_3374;
wire net_3772;
wire net_3807;
wire net_2698;
wire net_809;
wire net_1663;
wire net_629;
wire net_3450;
wire net_635;
wire net_266;
wire net_1235;
wire net_2691;
wire net_1037;
wire net_3528;
wire net_2019;
wire net_350;
wire net_3019;
wire net_3460;
wire net_2351;
wire x4524;
wire net_3117;
wire x2355;
wire net_1350;
wire net_3482;
wire net_3198;
wire net_1648;
wire net_1626;
wire net_2822;
wire net_1258;
wire net_2982;
wire net_1623;
wire net_631;
wire net_3369;
wire net_1101;
wire net_994;
wire net_318;
wire net_3927;
wire net_4007;
wire net_1971;
wire net_2409;
wire net_3192;
wire net_1900;
wire net_1779;
wire net_2647;
wire net_670;
wire net_3340;
wire net_103;
wire net_3844;
wire net_2687;
wire net_1849;
wire net_228;
wire net_3554;
wire net_2640;
wire net_966;
wire net_3372;
wire net_1920;
wire net_2201;
wire net_3928;
wire net_1108;
wire net_2827;
wire net_2025;
wire net_2010;
wire net_3854;
wire net_2936;
wire net_1878;
wire x6207;
wire net_755;
wire net_1723;
wire net_3890;
wire net_2900;
wire x5779;
wire net_133;
wire net_4025;
wire net_3151;
wire x3684;
wire net_3628;
wire net_2306;
wire net_3882;
wire net_3272;
wire net_2873;
wire net_557;
wire net_3043;
wire x1535;
wire net_2254;
wire net_2861;
wire net_1652;
wire net_3652;
wire net_2669;
wire net_1429;
wire net_1991;
wire net_1611;
wire net_1173;
wire x15;
wire net_1209;
wire net_1754;
wire net_1431;
wire net_2725;
wire x542;
wire net_3613;
wire net_2328;
wire net_1714;
wire x4096;
wire net_727;
wire net_847;
wire net_283;
wire x5386;
wire net_3190;
wire net_240;
wire x1241;
wire net_3757;
wire x342;
wire net_295;
wire net_344;
wire net_3951;
wire net_2269;
wire x679;
wire net_884;
wire net_712;
wire net_2281;
wire net_1422;
wire net_2259;
wire net_1106;
wire x7241;
wire net_1394;
wire net_2963;
wire net_2972;
wire net_2739;
wire net_1281;
wire net_2110;
wire net_2463;
wire net_2919;
wire x5686;
wire net_2893;
wire net_2241;
wire net_3227;
wire net_2358;
wire x722;
wire net_278;
wire x2773;
wire net_3057;
wire net_1547;
wire net_571;
wire x1332;
wire net_3509;
wire net_1162;
wire net_3934;
wire net_2443;
wire net_2472;
wire net_1307;
wire net_2790;
wire net_2742;
wire net_1877;
wire net_720;
wire net_2199;
wire x51;
wire net_3320;
wire net_2625;
wire net_684;
wire net_2648;
wire x3976;
wire net_3657;
wire net_3720;
wire net_510;
wire net_1353;
wire net_1595;
wire net_114;
wire net_3581;
wire net_3776;
wire net_2653;
wire net_1300;
wire net_3432;
wire x2371;
wire net_2974;
wire net_2960;
wire net_1252;
wire net_3895;
wire net_2734;
wire x1277;
wire net_2782;
wire net_494;
wire net_547;
wire x1835;
wire net_1098;
wire net_3146;
wire net_507;
wire net_1902;
wire net_238;
wire net_3074;
wire net_2438;
wire net_2600;
wire net_1911;
wire net_3022;
wire net_3563;
wire net_3461;
wire net_649;
wire net_1374;
wire net_1962;
wire net_457;
wire net_291;
wire net_2246;
wire net_1964;
wire net_772;
wire net_2494;
wire net_857;
wire net_867;
wire net_396;
wire net_3700;
wire x902;
wire net_107;
wire net_1277;
wire net_2661;
wire net_530;
wire x4258;
wire net_1541;
wire net_3893;
wire x4251;
wire net_594;
wire net_271;
wire net_3329;
wire net_673;
wire x5181;
wire net_3611;
wire net_2064;
wire net_2797;
wire net_2852;
wire net_1721;
wire net_3846;
wire net_1925;
wire net_3549;
wire net_1445;
wire net_2074;
wire net_1909;
wire net_2577;
wire net_1410;
wire net_2954;
wire net_1073;
wire net_365;
wire net_3274;
wire net_1947;
wire net_3913;
wire x4118;
wire net_3344;
wire x7369;
wire net_2953;
wire net_141;
wire net_3787;
wire net_467;
wire net_1810;
wire net_879;
wire net_1118;
wire net_2910;
wire net_2415;
wire net_372;
wire net_2990;
wire net_2081;
wire net_803;
wire net_3165;
wire x2416;
wire net_3595;
wire net_3197;
wire net_2788;
wire net_1348;
wire net_1476;
wire net_3489;
wire net_1293;
wire net_2883;
wire net_2302;
wire net_563;
wire net_1147;
wire net_3422;
wire net_199;
wire net_2789;
wire net_2681;
wire net_3835;
wire net_431;
wire net_2158;
wire net_1266;
wire net_3684;
wire net_2368;
wire net_1452;
wire net_2773;
wire net_2428;
wire net_909;
wire net_222;
wire net_152;
wire net_3105;
wire net_3999;
wire net_3966;
wire net_2895;
wire net_1788;
wire net_2138;
wire x5507;
wire net_258;
wire net_607;
wire net_2477;
wire x3338;
wire x381;
wire net_2935;
wire x1425;
wire net_1045;
wire net_2446;
wire net_3497;
wire net_3905;
wire x1600;
wire net_585;
wire net_3516;
wire net_3601;
wire net_1438;
wire net_3759;
wire net_3511;
wire net_374;
wire net_1143;
wire net_1987;
wire net_788;
wire net_214;
wire net_3602;
wire net_249;
wire net_3578;
wire net_1088;
wire x2050;
wire net_3885;
wire net_2079;
wire net_1731;
wire net_706;
wire net_2052;
wire net_4009;
wire net_2768;
wire net_2565;
wire net_2632;
wire net_551;
wire x2611;
wire net_2547;
wire net_3636;
wire net_2118;
wire net_463;
wire net_2295;
wire net_1536;
wire net_1817;
wire net_197;
wire net_2560;
wire net_3478;
wire net_1498;
wire net_1381;
wire net_3709;
wire net_202;
wire net_1199;
wire net_3312;
wire net_1756;
wire net_2208;
wire net_3627;
wire net_2595;
wire net_1383;
wire net_2751;
wire net_918;
wire net_949;
wire net_450;
wire net_289;
wire net_2614;
wire net_1642;
wire net_1683;
wire net_978;
wire net_2524;
wire x125;
wire net_1313;
wire net_1129;
wire net_3331;
wire x7007;
wire net_1056;
wire x4949;
wire net_1224;
wire net_2296;
wire net_768;
wire x1155;
wire net_3385;
wire net_357;
wire net_2044;
wire net_2181;
wire net_908;
wire net_1789;
wire net_3451;
wire net_519;
wire net_838;
wire net_3219;
wire x7314;
wire net_2694;
wire net_3118;
wire net_2096;
wire net_2697;
wire net_2576;
wire net_3827;
wire net_2352;
wire net_1829;
wire net_1038;
wire net_1204;
wire net_2342;
wire net_3763;
wire net_3515;
wire net_662;
wire net_3214;
wire net_1986;
wire net_862;
wire net_50;
wire net_3398;
wire net_2277;
wire net_2307;
wire net_342;
wire net_975;
wire net_612;
wire net_738;
wire net_892;
wire net_1150;
wire net_504;
wire net_2006;
wire net_3406;
wire net_1331;
wire net_1537;
wire x5247;
wire net_2130;
wire net_4000;
wire net_3362;
wire net_1148;
wire x1337;
wire net_3120;
wire net_2214;
wire net_3338;
wire net_2382;
wire x3396;
wire net_1561;
wire net_3442;
wire net_3864;
wire net_2728;
wire net_417;
wire net_122;
wire net_3269;
wire x1322;
wire x3595;
wire x1451;
wire net_1940;
wire net_3337;
wire net_2662;
wire net_94;
wire net_3752;
wire net_482;
wire net_991;
wire net_3258;
wire net_3912;
wire net_149;
wire net_3088;
wire net_387;
wire net_1473;
wire net_3275;
wire net_2979;
wire net_2772;
wire x1195;
wire net_1893;
wire net_1932;
wire net_1674;
wire net_1651;
wire net_3836;
wire net_577;
wire net_3401;
wire net_2375;
wire net_1806;
wire net_3234;
wire net_2550;
wire net_797;
wire net_2347;
wire net_3545;
wire net_1957;
wire net_1799;
wire net_1363;
wire net_1869;
wire net_3806;
wire net_2684;
wire net_2572;
wire net_3972;
wire net_521;
wire net_60;
wire net_2414;
wire net_2754;
wire net_337;
wire net_267;
wire net_1585;
wire net_1846;
wire net_690;
wire net_4012;
wire net_3743;
wire net_3663;
wire net_523;
wire net_3260;
wire net_3681;
wire net_3815;
wire net_3555;
wire net_2716;
wire net_2371;
wire net_3375;
wire net_3467;
wire net_351;
wire x950;
wire x734;
wire net_3982;
wire net_1388;
wire net_2842;
wire net_3158;
wire net_2828;
wire net_1257;
wire net_939;
wire net_824;
wire net_3458;
wire net_3391;
wire net_1822;
wire net_2730;
wire net_1631;
wire x6430;
wire net_1337;
wire net_1182;
wire net_1624;
wire net_2791;
wire net_1972;
wire net_1638;
wire x1097;
wire net_1950;
wire net_3126;
wire net_993;
wire net_3875;
wire x4336;
wire net_2421;
wire net_317;
wire net_856;
wire net_880;
wire net_1100;
wire net_1402;
wire net_2153;
wire net_3845;
wire net_1939;
wire net_2817;
wire net_3098;
wire net_2026;
wire x651;
wire net_2901;
wire net_162;
wire net_653;
wire net_1326;
wire net_3033;
wire x6319;
wire net_134;
wire net_546;
wire x3997;
wire net_3373;
wire net_3052;
wire net_2672;
wire net_3145;
wire net_588;
wire net_3694;
wire net_2200;
wire net_1157;
wire net_3701;
wire net_3855;
wire net_236;
wire x518;
wire net_487;
wire net_3883;
wire net_552;
wire net_1787;
wire net_1542;
wire net_1172;
wire net_3551;
wire x2950;
wire net_756;
wire net_104;
wire net_1065;
wire net_2237;
wire x6303;
wire net_3416;
wire x603;
wire net_72;
wire net_2566;
wire net_3953;
wire net_3795;
wire x5556;
wire net_3100;
wire net_241;
wire net_917;
wire net_3730;
wire net_3537;
wire net_2874;
wire x4175;
wire net_599;
wire net_711;
wire net_2225;
wire net_2993;
wire net_3067;
wire net_3111;
wire net_323;
wire net_963;
wire net_846;
wire x3900;
wire net_3017;
wire net_3737;
wire net_153;
wire net_2389;
wire net_174;
wire net_2607;
wire net_562;
wire net_375;
wire x3907;
wire net_364;
wire net_3172;
wire net_1831;
wire net_1482;
wire x6470;
wire net_79;
wire net_3291;
wire net_2168;
wire net_3306;
wire net_2928;
wire net_2849;
wire net_1885;
wire net_1030;
wire net_1485;
wire net_3245;
wire x582;
wire net_3171;
wire net_1247;
wire net_3673;
wire net_1969;
wire net_745;
wire net_2388;
wire net_933;
wire net_1244;
wire net_1215;
wire net_3496;
wire net_429;
wire net_129;
wire net_3377;
wire net_98;
wire net_373;
wire net_151;
wire net_356;
wire net_452;
wire net_1625;
wire net_545;
wire net_3683;
wire net_284;
wire net_1483;
wire net_2147;
wire x3365;
wire net_560;
wire net_439;
wire net_3031;
wire net_259;
wire net_2513;
wire net_3351;
wire net_3582;
wire x6358;
wire net_2645;
wire net_3119;
wire net_187;
wire net_1231;
wire net_3305;
wire x957;
wire net_2674;
wire net_160;
wire net_2872;
wire net_2432;
wire net_832;
wire net_322;
wire net_815;
wire net_1671;
wire net_420;
wire net_665;
wire net_1746;
wire net_2222;
wire x4998;
wire net_2322;
wire net_2825;
wire net_586;
wire net_3670;
wire net_1347;
wire net_1091;
wire net_3341;
wire net_3838;
wire net_1072;
wire net_3745;
wire net_120;
wire net_292;
wire net_109;
wire net_1706;
wire net_3708;
wire net_3574;
wire net_96;
wire net_1730;
wire net_2921;
wire net_167;
wire net_3289;
wire net_651;
wire net_2931;
wire net_3114;
wire net_3415;
wire net_744;
wire net_598;
wire net_2556;
wire x934;
wire x4658;
wire net_3519;
wire net_2740;
wire net_2806;
wire net_2011;
wire net_3455;
wire net_672;
wire net_777;
wire net_3157;
wire net_2820;
wire net_490;
wire net_2027;
wire x2971;
wire net_3068;
wire net_3892;
wire net_2456;
wire net_2753;
wire net_3610;
wire net_1232;
wire net_3462;
wire x3796;
wire net_1953;
wire net_3059;
wire x6550;
wire net_632;
wire net_3860;
wire net_843;
wire net_3925;
wire net_464;
wire net_3847;
wire net_2841;
wire x781;
wire net_1977;
wire net_2100;
wire net_2938;
wire net_2122;
wire x1402;
wire x4578;
wire net_1171;
wire net_1540;
wire net_248;
wire net_3594;
wire net_1725;
wire x1492;
wire net_3541;
wire net_1256;
wire net_802;
wire net_1413;
wire net_3532;
wire net_1767;
wire net_3556;
wire net_4010;
wire net_1840;
wire net_3041;
wire net_1640;
wire net_2724;
wire net_3427;
wire x4974;
wire net_1031;
wire x1294;
wire net_503;
wire net_1741;
wire x5493;
wire net_1636;
wire net_1672;
wire net_2103;
wire net_996;
wire net_3091;
wire net_3257;
wire net_2994;
wire net_75;
wire net_959;
wire net_1334;
wire net_206;
wire net_757;
wire net_1688;
wire net_2020;
wire net_3051;
wire net_4004;
wire net_2345;
wire net_235;
wire net_2973;
wire net_3106;
wire net_2961;
wire net_2374;
wire net_2503;
wire net_2164;
wire net_3644;
wire net_250;
wire net_3600;
wire net_3751;
wire net_3081;
wire net_2055;
wire net_2630;
wire net_2338;
wire net_3721;
wire net_403;
wire net_1985;
wire net_2340;
wire net_3524;
wire net_2616;
wire x6312;
wire net_282;
wire net_1596;
wire net_2275;
wire net_3976;
wire net_841;
wire net_1750;
wire net_794;
wire net_2370;
wire net_2397;
wire net_2047;
wire net_3346;
wire net_2469;
wire net_2693;
wire net_528;
wire x7329;
wire net_1012;
wire net_1404;
wire x3865;
wire net_335;
wire net_3433;
wire net_907;
wire net_1468;
wire net_3464;
wire net_181;
wire net_3333;
wire x5468;
wire net_3076;
wire net_395;
wire net_2036;
wire net_2539;
wire net_3649;
wire net_1130;
wire net_2719;
wire net_386;
wire net_2323;
wire net_3867;
wire x1415;
wire net_3677;
wire net_641;
wire net_1790;
wire net_2798;
wire net_3869;
wire net_1152;
wire net_1226;
wire net_2318;
wire net_3449;
wire net_1901;
wire net_3021;
wire net_3711;
wire net_1039;
wire net_1709;
wire net_3805;
wire x6936;
wire net_400;
wire net_3942;
wire net_1935;
wire net_602;
wire net_2379;
wire net_175;
wire net_1818;
wire net_2918;
wire net_1850;
wire net_2925;
wire net_1497;
wire net_1800;
wire x450;
wire net_1855;
wire net_279;
wire x4040;
wire net_1163;
wire net_1177;
wire net_1523;
wire net_1992;
wire net_3347;
wire net_897;
wire net_1656;
wire x7509;
wire net_2853;
wire net_691;
wire net_2705;
wire net_615;
wire net_3273;
wire net_441;
wire net_1559;
wire net_3178;
wire net_2701;
wire net_1620;
wire net_1863;
wire net_2833;
wire net_2608;
wire net_2561;
wire net_2663;
wire net_2813;
wire net_728;
wire net_1276;
wire net_719;
wire net_170;
wire net_2519;
wire net_471;
wire net_3813;
wire net_1055;
wire net_2571;
wire net_3894;
wire net_878;
wire net_1531;
wire net_1159;
wire net_518;
wire net_861;
wire net_57;
wire net_3479;
wire net_3222;
wire net_929;
wire net_3321;
wire net_708;
wire net_2523;
wire net_3552;
wire net_696;
wire net_3954;
wire net_3216;
wire net_1565;
wire net_169;
wire net_171;
wire net_2234;
wire x4164;
wire net_3821;
wire net_604;
wire net_967;
wire net_1527;
wire net_268;
wire net_3486;
wire net_48;
wire net_483;
wire net_3386;
wire net_1149;
wire net_1645;
wire net_2962;
wire x4033;
wire net_176;
wire net_3638;
wire net_1298;
wire net_2570;
wire net_296;
wire net_2131;
wire net_3354;
wire net_614;
wire net_2712;
wire net_2005;
wire net_1123;
wire net_2771;
wire net_3194;
wire net_3572;
wire x7383;
wire net_2228;
wire net_3020;
wire net_786;
wire net_1192;
wire net_127;
wire net_984;
wire net_1339;
wire net_3363;
wire x2528;
wire net_3781;
wire net_1105;
wire net_906;
wire net_2172;
wire net_2422;
wire net_3156;
wire net_2482;
wire net_707;
wire net_3577;
wire net_652;
wire net_3840;
wire net_1815;
wire net_3782;
wire net_1856;
wire net_830;
wire net_575;
wire net_2505;
wire net_877;
wire net_1279;
wire net_1047;
wire net_2799;
wire net_3697;
wire net_3734;
wire net_2683;
wire net_2631;
wire net_2165;
wire net_3618;
wire net_3284;
wire net_1467;
wire net_1474;
wire net_1061;
wire net_2784;
wire net_3181;
wire net_765;
wire net_675;
wire net_1342;
wire net_2562;
wire net_2633;
wire net_2867;
wire net_1666;
wire net_3837;
wire x7264;
wire net_3472;
wire net_2288;
wire net_2099;
wire net_1768;
wire net_2182;
wire net_150;
wire net_304;
wire net_2021;
wire net_1068;
wire net_1703;
wire net_186;
wire net_3983;
wire net_2495;
wire net_3814;
wire net_3693;
wire net_1050;
wire net_2072;
wire net_2760;
wire net_1316;
wire net_1872;
wire net_792;
wire net_2271;
wire net_3070;
wire net_3409;
wire net_2203;
wire x6773;
wire net_1716;
wire net_1904;
wire net_3907;
wire net_1607;
wire net_219;
wire net_3609;
wire net_1263;
wire net_2187;
wire net_196;
wire net_2476;
wire net_3452;
wire net_913;
wire net_2067;
wire net_3130;
wire net_3387;
wire net_1479;
wire net_4019;
wire net_1639;
wire net_3094;
wire net_360;
wire net_1927;
wire net_3625;
wire net_213;
wire net_2324;
wire net_260;
wire net_947;
wire net_2947;
wire net_3137;
wire net_732;
wire net_1126;
wire net_2152;
wire net_2004;
wire net_1325;
wire net_3316;
wire net_3032;
wire net_1597;
wire net_1352;
wire net_1373;
wire net_2567;
wire net_2885;
wire net_2088;
wire net_1187;
wire net_2689;
wire net_3988;
wire net_2761;
wire net_3206;
wire net_1303;
wire net_3788;
wire net_2858;
wire x3020;
wire net_1503;
wire net_3961;
wire net_2102;
wire net_1442;
wire net_449;
wire net_1807;
wire net_1930;
wire net_1943;
wire net_1087;
wire net_3995;
wire net_733;
wire net_887;
wire net_1894;
wire x5078;
wire net_2431;
wire net_2308;
wire net_633;
wire net_113;
wire net_2989;
wire net_497;
wire net_1914;
wire net_2770;
wire net_2408;
wire net_3889;
wire net_1424;
wire net_2636;
wire net_1414;
wire net_300;
wire net_3567;
wire net_2652;
wire x3884;
wire net_1233;
wire net_1457;
wire net_2720;
wire net_2741;
wire net_1834;
wire net_950;
wire net_4011;
wire net_1436;
wire net_2448;
wire net_3400;
wire net_3392;
wire net_2551;
wire net_2816;
wire net_646;
wire net_2731;
wire net_1214;
wire net_2601;
wire net_3641;
wire x6503;
wire net_866;
wire net_2891;
wire net_520;
wire net_3150;
wire x3447;
wire net_1032;
wire net_567;
wire net_3726;
wire net_3979;
wire net_3231;
wire net_981;
wire net_272;
wire x234;
wire net_2401;
wire net_3939;
wire x2134;
wire net_1024;
wire x1086;
wire net_1566;
wire net_1590;
wire net_1305;
wire net_1612;
wire net_2354;
wire net_839;
wire net_1387;
wire net_814;
wire net_1581;
wire net_2413;
wire net_559;
wire net_345;
wire net_2792;
wire net_3042;
wire net_2128;
wire net_2965;
wire net_3930;
wire net_1717;
wire net_2586;
wire net_3299;
wire net_398;
wire net_1655;
wire net_3399;
wire net_954;
wire net_2365;
wire net_2117;
wire net_2461;
wire net_1766;
wire x7190;
wire net_2582;
wire net_2361;
wire net_2598;
wire net_3872;
wire net_2879;
wire net_1572;
wire net_1680;
wire x925;
wire net_3302;
wire net_3187;
wire net_2134;
wire net_2622;
wire net_316;
wire net_84;
wire x1371;
wire net_1759;
wire net_3764;
wire x6096;
wire net_2262;
wire net_4022;
wire net_3011;
wire net_2087;
wire net_2541;
wire net_3689;
wire net_533;
wire net_1002;
wire net_1695;
wire x3636;
wire net_911;
wire net_1617;
wire net_3188;
wire net_1993;
wire net_3010;
wire net_881;
wire net_2805;
wire net_1397;
wire net_2903;
wire net_568;
wire x3227;
wire net_47;
wire net_1227;
wire net_1008;
wire net_1443;
wire net_1954;
wire net_3873;
wire net_3069;
wire net_3170;
wire net_2840;
wire x6326;
wire net_3463;
wire net_2155;
wire net_4005;
wire net_168;
wire net_2041;
wire net_3199;
wire net_3597;
wire net_385;
wire net_269;
wire net_2609;
wire net_3193;
wire net_469;
wire net_3131;
wire net_1945;
wire net_1978;
wire net_3179;
wire x4821;
wire net_3167;
wire net_1170;
wire net_1833;
wire net_2423;
wire net_2280;
wire net_2831;
wire net_3029;
wire net_778;
wire net_2366;
wire net_2380;
wire net_3393;
wire net_1455;
wire net_2930;
wire net_895;
wire net_1412;
wire x6623;
wire net_1255;
wire net_3980;
wire net_1250;
wire net_1481;
wire net_995;
wire net_207;
wire net_3040;
wire net_3557;
wire x7404;
wire net_3643;
wire net_700;
wire net_1246;
wire net_3004;
wire x6264;
wire net_1689;
wire net_1774;
wire net_1673;
wire net_3830;
wire net_3060;
wire net_274;
wire net_2568;
wire net_3480;
wire net_321;
wire net_1075;
wire x3669;
wire net_833;
wire net_930;
wire net_2387;
wire net_2995;
wire net_99;
wire net_3526;
wire net_2945;
wire net_2267;
wire net_934;
wire x1811;
wire net_3103;
wire net_544;
wire net_717;
wire net_3665;
wire net_1399;
wire net_3630;
wire net_1824;
wire net_3350;
wire net_3402;
wire net_2223;
wire net_3553;
wire x1646;
wire net_2673;
wire net_3500;
wire net_3166;
wire net_3304;
wire net_1245;
wire net_2549;
wire net_860;
wire net_1781;
wire net_3660;
wire net_3465;
wire net_870;
wire net_2046;
wire net_3049;
wire net_637;
wire net_2878;
wire net_2514;
wire net_2871;
wire x1124;
wire x5317;
wire net_2390;
wire net_3267;
wire net_2321;
wire net_2686;
wire net_3474;
wire net_2013;
wire net_817;
wire net_1509;
wire net_529;
wire net_3414;
wire net_3495;
wire net_97;
wire net_2028;
wire net_2553;
wire net_3766;
wire net_1889;
wire net_1591;
wire net_2920;
wire net_2981;
wire net_1747;
wire net_650;
wire net_1164;
wire net_2012;
wire x844;
wire net_121;
wire net_597;
wire net_743;
wire net_3770;
wire net_1922;
wire net_2583;
wire net_3820;
wire net_3799;
wire net_2664;
wire x862;
wire x6706;
wire net_2706;
wire net_849;
wire net_603;
wire net_2451;
wire net_2602;
wire net_401;
wire net_642;
wire net_1522;
wire net_2699;
wire net_3798;
wire net_1158;
wire net_2714;
wire net_2926;
wire net_2183;
wire net_2557;
wire net_440;
wire x1113;
wire net_470;
wire net_758;
wire x5846;
wire net_2702;
wire net_430;
wire net_2834;
wire net_718;
wire x4843;
wire net_3943;
wire net_83;
wire x4323;
wire net_3129;
wire net_56;
wire net_3255;
wire x132;
wire net_1063;
wire net_968;
wire x108;
wire net_336;
wire net_1578;
wire net_2534;
wire net_2917;
wire x1956;
wire net_3221;
wire net_1504;
wire net_697;
wire net_475;
wire net_2003;
wire net_3732;
wire net_605;
wire net_3411;
wire net_2309;
wire net_502;
wire net_2470;
wire net_1564;
wire net_3426;
wire net_1568;
wire net_3804;
wire net_924;
wire net_1526;
wire net_1884;
wire net_1333;
wire net_3919;
wire net_2348;
wire net_489;
wire x91;
wire net_2646;
wire net_3868;
wire net_3082;
wire net_3936;
wire net_3676;
wire net_2628;
wire net_2748;
wire net_251;
wire net_1360;
wire net_2054;
wire net_3364;
wire net_664;
wire net_128;
wire net_840;
wire net_1364;
wire net_549;
wire net_827;
wire net_2793;
wire net_411;
wire net_2137;
wire net_1836;
wire net_2337;
wire net_1369;
wire x768;
wire net_3430;
wire net_1862;
wire x2649;
wire net_2317;
wire x1462;
wire net_1013;
wire net_1530;
wire net_3075;
wire net_3583;
wire net_112;
wire net_842;
wire net_2952;
wire net_1705;
wire net_2336;
wire net_2035;
wire x886;
wire net_2373;
wire net_2826;
wire net_3739;
wire net_2398;
wire net_492;
wire net_3678;
wire net_2141;
wire net_2639;
wire net_3315;
wire net_2455;
wire net_1609;
wire net_402;
wire x2543;
wire net_3453;
wire net_3695;
wire net_1327;
wire net_3448;
wire net_110;
wire net_1403;
wire net_3248;
wire net_2248;
wire net_2270;
wire net_2274;
wire net_1667;
wire net_3866;
wire x5143;
wire net_1386;
wire net_1606;
wire net_3710;
wire net_2359;
wire net_3054;
wire net_3978;
wire net_2186;
wire x2304;
wire net_3696;
wire net_3473;
wire x499;
wire net_1430;
wire net_2029;
wire net_2868;
wire net_569;
wire net_2478;
wire net_3698;
wire x2119;
wire net_2563;
wire net_2946;
wire net_2587;
wire net_1284;
wire net_3408;
wire net_630;
wire net_76;
wire net_2959;
wire net_2202;
wire net_1888;
wire net_2490;
wire net_4018;
wire net_3929;
wire net_1791;
wire net_1471;
wire net_1792;
wire x2993;
wire net_2496;
wire x1357;
wire net_3109;
wire net_2066;
wire net_3608;
wire x3041;
wire net_1598;
wire net_3124;
wire net_1903;
wire net_2407;
wire net_731;
wire net_1146;
wire net_912;
wire net_1733;
wire net_2078;
wire x5370;
wire net_779;
wire net_3841;
wire net_1928;
wire x2016;
wire net_1328;
wire net_234;
wire net_2859;
wire net_3848;
wire net_2884;
wire net_2762;
wire net_3205;
wire net_1094;
wire net_3487;
wire net_2749;
wire net_855;
wire net_1724;
wire net_674;
wire net_3703;
wire x83;
wire net_303;
wire net_2089;
wire net_491;
wire net_2475;
wire net_965;
wire net_3797;
wire net_1299;
wire net_948;
wire net_2937;
wire net_3535;
wire net_1195;
wire net_2916;
wire net_421;
wire net_1396;
wire net_2502;
wire net_1104;
wire net_764;
wire net_876;
wire net_2593;
wire net_2162;
wire net_2737;
wire net_2439;
wire net_172;
wire net_2481;
wire net_1117;
wire net_1458;
wire x101;
wire net_3955;
wire net_905;
wire net_1060;
wire net_2617;
wire net_142;
wire x2200;
wire net_2229;
wire net_2235;
wire net_158;
wire x1854;
wire net_1715;
wire net_3200;
wire net_3733;
wire net_3881;
wire net_2080;
wire net_3675;
wire net_2711;
wire net_2097;
wire net_2504;
wire net_3619;
wire net_3784;
wire net_1216;
wire net_2175;
wire net_2815;
wire net_3785;
wire net_1086;
wire net_1271;
wire net_2116;
wire net_1758;
wire net_1782;
wire net_1769;
wire net_1197;
wire net_1967;
wire net_273;
wire net_1278;
wire net_1567;
wire net_576;
wire net_3182;
wire net_1654;
wire net_2098;
wire net_465;
wire x794;
wire net_177;
wire net_3355;
wire net_3005;
wire net_1883;
wire net_476;
wire net_2783;
wire net_2803;
wire net_382;
wire net_3058;
wire net_3301;
wire x5995;
wire net_725;
wire net_3931;
wire net_583;
wire net_1315;
wire net_953;
wire net_894;
wire net_1074;
wire net_1058;
wire x44;
wire net_1423;
wire net_1871;
wire net_2902;
wire net_517;
wire net_628;
wire net_2489;
wire net_3494;
wire net_220;
wire net_1465;
wire net_293;
wire net_3666;
wire net_1938;
wire net_543;
wire net_3160;
wire net_625;
wire net_2125;
wire net_3760;
wire net_1823;
wire x4397;
wire net_1289;
wire x7345;
wire net_3138;
wire net_2623;
wire net_261;
wire net_191;
wire net_3576;
wire net_2909;
wire net_558;
wire net_2069;
wire x3733;
wire net_2362;
wire net_1618;
wire net_2497;
wire net_1955;
wire net_2723;
wire net_2552;
wire net_3562;
wire net_1001;
wire net_3229;
wire net_3765;
wire net_781;
wire net_1694;
wire net_910;
wire x4790;
wire net_3012;
wire net_3754;
wire net_2412;
wire net_185;
wire net_4023;
wire net_3989;
wire x6880;
wire net_1984;
wire net_1994;
wire net_315;
wire net_1015;
wire net_1375;
wire net_2980;
wire x1559;
wire net_1944;
wire net_4006;
wire net_3897;
wire net_1351;
wire net_1775;
wire net_3960;
wire net_346;
wire net_297;
wire net_91;
wire net_1535;
wire net_3992;
wire net_2400;
wire x1442;
wire net_2287;
wire x4206;
wire net_448;
wire net_2034;
wire x1937;
wire net_886;
wire net_229;
wire net_3189;
wire net_1808;
wire net_2146;
wire net_2988;
wire net_3256;
wire net_687;
wire net_405;
wire net_3266;
wire net_1111;
wire net_2651;
wire net_3888;
wire net_3651;
wire net_3971;
wire x4022;
wire net_3155;
wire net_3322;
wire net_2533;
wire net_1470;
wire net_3566;
wire x878;
wire net_1913;
wire x1877;
wire x5820;
wire net_831;
wire net_3596;
wire net_451;
wire net_750;
wire net_1234;
wire x807;
wire x192;
wire net_1760;
wire net_1184;
wire x361;
wire net_2778;
wire net_3926;
wire net_2756;
wire x550;
wire net_3403;
wire net_1085;
wire net_1960;
wire net_592;
wire net_3093;
wire net_647;
wire net_3247;
wire net_773;
wire net_2266;
wire net_2464;
wire net_281;
wire net_828;
wire net_3839;
wire net_1603;
wire net_2732;
wire x7552;
wire net_3521;
wire net_1096;
wire net_3727;
wire x1136;
wire net_795;
wire net_982;
wire net_1580;
wire net_1406;
wire net_54;
wire x2846;
wire net_3896;
wire net_526;
wire net_2718;
wire net_834;
wire net_694;
wire net_1434;
wire net_2747;
wire net_3668;
wire net_1570;
wire net_974;
wire net_774;
wire net_923;
wire x1285;
wire net_1707;
wire net_2190;
wire net_1881;
wire net_501;
wire net_111;
wire x6968;
wire net_3679;
wire net_225;
wire net_252;
wire net_124;
wire net_3128;
wire net_3323;
wire x3098;
wire net_2399;
wire x1507;
wire x4129;
wire net_901;
wire net_447;
wire net_871;
wire net_2611;
wire net_3425;
wire net_410;
wire net_1492;
wire net_390;
wire net_1154;
wire net_2537;
wire net_3767;
wire net_80;
wire net_2951;
wire net_2603;
wire net_3631;
wire net_1132;
wire net_2442;
wire net_2293;
wire net_280;
wire net_3026;
wire net_495;
wire net_1802;
wire x1230;
wire net_2140;
wire net_2356;
wire x1306;
wire net_971;
wire net_3288;
wire net_2049;
wire net_2273;
wire net_617;
wire net_2517;
wire net_2316;
wire net_2184;
wire net_554;
wire x760;
wire net_2755;
wire net_3740;
wire net_1678;
wire net_2703;
wire net_46;
wire net_3366;
wire net_584;
wire net_1441;
wire net_969;
wire net_1525;
wire net_3870;
wire net_2411;
wire net_165;
wire net_4003;
wire net_821;
wire net_3438;
wire net_3824;
wire x398;
wire net_3436;
wire net_2335;
wire net_3940;
wire net_384;
wire net_3911;
wire net_3823;
wire net_2618;
wire net_3503;
wire net_3365;
wire net_3859;
wire net_2599;
wire net_2665;
wire net_3642;
wire net_3803;
wire net_1114;
wire net_2707;
wire net_3388;
wire net_485;
wire net_1748;
wire net_3078;
wire net_3218;
wire x1253;
wire net_2964;
wire x1187;
wire net_3334;
wire net_3224;
wire net_64;
wire net_1719;
wire net_2232;
wire net_2343;
wire net_726;
wire net_3811;
wire net_1028;
wire net_1529;
wire net_600;
wire net_3237;
wire net_701;
wire net_125;
wire net_397;
wire net_808;
wire net_1685;
wire net_1704;
wire net_2440;
wire net_1384;
wire net_2738;
wire net_3918;
wire net_1379;
wire net_320;
wire x317;
wire x6678;
wire net_1322;
wire net_2644;
wire net_2944;
wire net_1301;
wire net_986;
wire net_1242;
wire net_286;
wire x4752;
wire net_1241;
wire net_3690;
wire net_3584;
wire net_935;
wire net_3001;
wire net_1511;
wire net_3116;
wire net_645;
wire net_426;
wire net_3121;
wire net_1634;
wire net_609;
wire net_414;
wire x5338;
wire net_1048;
wire net_3048;
wire net_799;
wire net_3083;
wire net_3475;
wire net_1816;
wire net_2014;
wire net_1221;
wire net_1951;
wire net_331;
wire x7087;
wire x702;
wire net_816;
wire net_3264;
wire net_2092;
wire net_2558;
wire net_2454;
wire net_2040;
wire net_2220;
wire net_2823;
wire net_1217;
wire net_1508;
wire net_3379;
wire net_2933;
wire net_3728;
wire net_931;
wire net_3381;
wire net_2242;
wire net_759;
wire x3245;
wire net_1575;
wire net_3279;
wire net_657;
wire net_1727;
wire net_247;
wire net_329;
wire net_1259;
wire net_1924;
wire net_2143;
wire net_2839;
wire net_1825;
wire net_3791;
wire net_2196;
wire net_70;
wire net_3168;
wire net_3413;
wire net_1341;
wire net_962;
wire net_478;
wire net_1934;
wire net_3242;
wire net_1835;
wire net_596;
wire net_1848;
wire net_1261;
wire net_333;
wire net_639;
wire net_2120;
wire net_1975;
wire net_1238;
wire net_565;
wire net_2569;
wire net_2832;
wire net_1033;
wire net_3923;
wire net_2149;
wire net_3028;
wire net_2554;
wire net_1692;
wire net_2528;
wire net_2655;
wire net_3107;
wire net_1686;
wire net_1361;
wire net_367;
wire net_3303;
wire net_2450;
wire net_1842;
wire net_1208;
wire net_204;
wire net_232;
wire net_3957;
wire net_1180;
wire net_1627;
wire net_2002;
wire net_1069;
wire x6592;
wire net_2022;
wire net_2167;
wire net_2880;
wire net_2385;
wire net_2996;
wire net_2889;
wire net_3431;
wire net_3565;
wire net_1416;
wire net_137;
wire x6372;
wire net_3154;
wire net_2433;
wire net_532;
wire net_2501;
wire net_3530;
wire net_3622;
wire net_4029;
wire net_1601;
wire net_93;
wire x4066;
wire net_1916;
wire net_2729;
wire net_2468;
wire net_302;
wire net_1131;
wire net_889;
wire net_1116;
wire net_348;
wire net_753;
wire net_626;
wire x2289;
wire net_100;
wire net_1809;
wire net_686;
wire net_2195;
wire net_1615;
wire net_3421;
wire net_2814;
wire net_1691;
wire net_689;
wire net_751;
wire net_2112;
wire net_595;
wire net_2363;
wire net_1320;
wire net_1828;
wire net_1466;
wire net_3659;
wire net_3724;
wire net_157;
wire net_1710;
wire net_1228;
wire net_1205;
wire x6122;
wire net_466;
wire net_1179;
wire x2869;
wire net_2722;
wire net_1426;
wire net_3039;
wire net_2217;
wire net_1407;
wire net_938;
wire net_3147;
wire net_1610;
wire net_1761;
wire net_3569;
wire net_183;
wire net_3263;
wire net_1440;
wire net_4020;
wire net_1057;
wire net_2915;
wire net_1011;
wire net_1355;
wire net_800;
wire net_644;
wire x2579;
wire net_852;
wire net_2987;
wire net_2253;
wire net_2580;
wire net_1699;
wire net_1042;
wire net_1385;
wire net_1643;
wire net_1534;
wire net_1919;
wire net_1000;
wire net_1995;
wire net_2521;
wire x6727;
wire net_2545;
wire net_1016;
wire x2739;
wire x5224;
wire net_659;
wire net_3977;
wire net_899;
wire net_1744;
wire net_1010;
wire net_516;
wire net_1693;
wire net_2870;
wire net_3176;
wire net_3654;
wire net_3585;
wire net_3779;
wire x1044;
wire net_956;
wire net_2908;
wire net_3963;
wire net_2068;
wire net_2596;
wire net_3705;
wire net_2970;
wire x638;
wire net_438;
wire net_2675;
wire net_2794;
wire net_2584;
wire x2631;
wire net_314;
wire net_1752;
wire net_2250;
wire net_2527;
wire net_3013;
wire net_952;
wire net_3110;
wire net_2091;
wire net_2967;
wire net_2406;
wire net_3185;
wire net_807;
wire net_3300;
wire net_3405;
wire net_86;
wire net_3270;
wire net_2245;
wire x5657;
wire net_3484;
wire net_2474;
wire net_945;
wire net_2530;
wire net_2101;
wire net_383;
wire net_3570;
wire net_217;
wire net_3140;
wire net_427;
wire net_135;
wire x1897;
wire net_2785;
wire net_915;
wire net_1121;
wire net_2226;
wire net_3849;
wire x3067;
wire net_473;
wire net_3599;
wire x169;
wire net_2777;
wire net_1049;
wire net_3901;
wire net_454;
wire net_1784;
wire net_1296;
wire net_709;
wire net_2484;
wire net_2863;
wire net_3507;
wire net_1165;
wire net_1066;
wire net_677;
wire net_1472;
wire net_2939;
wire net_1113;
wire net_2424;
wire net_1968;
wire net_2591;
wire net_1344;
wire x4051;
wire net_3968;
wire net_1283;
wire net_1084;
wire net_1500;
wire net_354;
wire net_2507;
wire net_1136;
wire net_3008;
wire net_2685;
wire net_2763;
wire net_573;
wire net_2658;
wire net_2898;
wire net_1391;
wire net_2174;
wire net_784;
wire net_3356;
wire x4604;
wire net_1772;
wire net_3529;
wire net_45;
wire net_3616;
wire net_381;
wire x2674;
wire net_2498;
wire net_3886;
wire net_2326;
wire net_1592;
wire net_3540;
wire net_3783;
wire net_2085;
wire net_3672;
wire net_1857;
wire net_1637;
wire net_3702;
wire net_1318;
wire net_3238;
wire net_941;
wire net_55;
wire net_1557;
wire net_3852;
wire net_1514;
wire x439;
wire net_3092;
wire net_2070;
wire net_2311;
wire net_3575;
wire net_1599;
wire net_306;
wire net_3981;
wire net_3828;
wire net_3132;
wire net_3161;
wire net_1290;
wire net_500;
wire net_1906;
wire net_3053;
wire net_2610;
wire net_3297;
wire net_2023;
wire net_1329;
wire net_123;
wire net_527;
wire net_362;
wire net_262;
wire net_1668;
wire net_3424;
wire net_3127;
wire net_1052;
wire net_3139;
wire net_3831;
wire net_1793;
wire net_3786;
wire net_3104;
wire x2318;
wire net_2189;
wire net_3632;
wire net_2057;
wire net_2278;
wire net_3072;
wire net_1124;
wire net_226;
wire net_1021;
wire x1176;
wire net_1737;
wire net_143;
wire x1794;
wire net_1859;
wire net_190;
wire net_2887;
wire net_1447;
wire net_145;
wire net_1929;
wire net_3607;
wire net_1983;
wire net_1145;
wire net_2061;
wire net_3030;
wire net_3493;
wire net_2804;
wire x7061;
wire net_2261;
wire net_3842;
wire net_188;
wire net_1553;
wire net_3753;
wire net_1895;
wire net_3061;
wire net_509;
wire net_3319;
wire net_211;
wire net_2491;
wire net_2958;
wire net_1077;
wire net_3208;
wire net_2704;
wire net_2924;
wire x1105;
wire net_3910;
wire net_2410;
wire net_1851;
wire net_3941;
wire net_119;
wire net_3108;
wire x2706;
wire net_2185;
wire net_1321;
wire net_2233;
wire net_3445;
wire net_2941;
wire net_2033;
wire net_477;
wire net_3348;
wire net_2123;
wire net_1099;
wire x5413;
wire net_2943;
wire net_3861;
wire net_2532;
wire net_90;
wire net_2315;
wire net_85;
wire net_2231;
wire net_1864;
wire x1266;
wire net_404;
wire net_3812;
wire net_1200;
wire net_2518;
wire net_2666;
wire net_1239;
wire x255;
wire net_1463;
wire net_1646;
wire net_2056;
wire net_2776;
wire net_3389;
wire net_3437;
wire x4353;
wire net_1562;
wire net_3822;
wire x4283;
wire net_472;
wire net_2522;
wire net_1510;
wire net_65;
wire net_1628;
wire net_3476;
wire net_3077;
wire x421;
wire net_896;
wire net_484;
wire net_2512;
wire x7145;
wire net_3223;
wire net_136;
wire net_1524;
wire net_1936;
wire net_3802;
wire net_1528;
wire net_126;
wire net_2708;
wire net_1749;
wire net_3367;
wire x2451;
wire net_2211;
wire net_601;
wire net_1362;
wire x691;
wire net_1896;
wire net_2346;
wire net_1732;
wire net_1982;
wire net_829;
wire net_2511;
wire net_2626;
wire net_2115;
wire net_2294;
wire net_2299;
wire net_2393;
wire net_3917;
wire x3843;
wire net_3376;
wire net_900;
wire net_1405;
wire net_3253;
wire net_1882;
wire x5581;
wire net_413;
wire net_2001;
wire net_1491;
wire net_716;
wire x7120;
wire net_1269;
wire net_3750;
wire net_2419;
wire net_1034;
wire net_3715;
wire net_3533;
wire net_2696;
wire net_253;
wire net_276;
wire net_1449;
wire net_3439;
wire net_666;
wire net_1959;
wire net_616;
wire net_1220;
wire net_4017;
wire net_3946;
wire net_1847;
wire net_2717;
wire net_793;
wire net_460;
wire net_1657;
wire net_3084;
wire net_2353;
wire net_2272;
wire net_2334;
wire net_3994;
wire net_1367;
wire net_1133;
wire net_3287;
wire net_166;
wire net_1976;
wire net_2866;
wire net_3169;
wire net_3025;
wire net_3871;
wire net_3792;
wire net_1371;
wire net_2758;
wire net_3352;
wire net_117;
wire net_74;
wire net_3832;
wire net_1826;
wire net_205;
wire net_1286;
wire x748;
wire net_2142;
wire net_920;
wire net_334;
wire net_1952;
wire net_1461;
wire net_2453;
wire net_3009;
wire net_3062;
wire x7215;
wire net_820;
wire net_3177;
wire net_380;
wire x1434;
wire net_2847;
wire net_1556;
wire net_3768;
wire net_437;
wire net_1270;
wire net_3573;
wire net_2286;
wire net_566;
wire net_1552;
wire x1029;
wire net_3878;
wire x4549;
wire net_624;
wire net_2148;
wire net_3215;
wire net_3717;
wire net_298;
wire net_1933;
wire net_2108;
wire net_2529;
wire net_688;
wire x4107;
wire net_3241;
wire net_998;
wire net_2157;
wire net_2555;
wire net_3504;
wire net_3027;
wire net_2405;
wire net_835;
wire net_1687;
wire net_1762;
wire x3947;
wire net_1181;
wire x665;
wire net_1357;
wire net_638;
wire net_3986;
wire net_3637;
wire net_932;
wire x2220;
wire net_313;
wire net_1243;
wire net_1660;
wire net_1484;
wire net_1783;
wire net_3667;
wire net_419;
wire net_1874;
wire x3428;
wire net_1635;
wire net_972;
wire net_936;
wire net_819;
wire net_3499;
wire net_785;
wire net_3002;
wire net_1489;
wire net_854;
wire net_2619;
wire net_3141;
wire net_1670;
wire net_3746;
wire net_2221;
wire net_1349;
wire net_2801;
wire net_3265;
wire net_979;
wire net_2392;
wire net_2932;
wire net_156;
wire net_2015;
wire net_1264;
wire x3921;
wire net_1040;
wire net_332;
wire net_1745;
wire net_1679;
wire net_3089;
wire net_3101;
wire net_3037;
wire net_3148;
wire net_1229;
wire net_656;
wire net_3876;
wire net_766;
wire x5605;
wire net_2907;
wire net_3686;
wire net_1153;
wire net_1887;
wire net_3014;
wire net_379;
wire net_2243;
wire net_1569;
wire x7466;
wire net_3113;
wire net_3454;
wire net_3133;
wire net_3047;
wire net_2559;
wire net_3969;
wire net_2657;
wire net_1358;
wire net_3729;
wire net_2629;
wire net_2486;
wire net_2251;
wire net_1698;
wire net_1017;
wire net_955;
wire net_1206;
wire net_2585;
wire net_3653;
wire net_960;
wire net_1996;
wire net_3704;
wire net_1166;
wire net_1029;
wire net_801;
wire net_412;
wire net_2620;
wire net_1718;
wire net_2581;
wire x2435;
wire net_2986;
wire net_3162;
wire net_1873;
wire net_2129;
wire net_3801;
wire x297;
wire net_453;
wire net_581;
wire net_2899;
wire net_3510;
wire net_3180;
wire net_658;
wire net_3249;
wire net_2263;
wire net_734;
wire net_3624;
wire net_2544;
wire net_2090;
wire net_2325;
wire x1578;
wire net_951;
wire net_2086;
wire net_806;
wire net_3186;
wire x2260;
wire x3986;
wire net_4021;
wire x5892;
wire net_946;
wire net_1176;
wire net_2676;
wire net_2966;
wire net_1253;
wire net_2194;
wire net_2500;
wire net_1076;
wire net_3900;
wire net_1751;
wire net_3559;
wire x3483;
wire net_681;
wire net_3153;
wire net_3508;
wire net_2434;
wire net_3564;
wire net_1448;
wire net_2032;
wire net_392;
wire net_118;
wire net_3598;
wire net_2467;
wire net_146;
wire net_2452;
wire net_3938;
wire net_3523;
wire net_3712;
wire net_1502;
wire net_428;
wire net_246;
wire net_1186;
wire net_640;
wire net_2216;
wire net_2888;
wire net_775;
wire net_1378;
wire net_752;
wire net_3773;
wire net_1773;
wire net_1600;
wire net_2531;
wire net_3716;
wire net_888;
wire net_498;
wire net_535;
wire net_676;
wire net_2721;
wire net_2637;
wire net_1023;
wire net_2538;
wire net_2447;
wire net_3623;
wire net_301;
wire net_2360;
wire net_3617;
wire net_299;
wire net_1343;
wire net_2285;
wire x5448;
wire net_3492;
wire x2722;
wire net_182;
wire net_2462;
wire net_590;
wire net_3879;
wire net_2024;
wire net_3240;
wire net_3324;
wire net_3254;
wire net_3725;
wire net_1435;
wire net_1370;
wire x3699;
wire net_407;
wire x1379;
wire net_3568;
wire net_1736;
wire net_3207;
wire net_2204;
wire net_2492;
wire net_2312;
wire x1144;
wire net_1970;
wire net_1306;
wire net_3843;
wire net_1669;
wire net_1858;
wire net_1041;
wire net_2073;
wire net_3038;
wire net_2690;
wire net_2950;
wire net_3924;
wire x4303;
wire net_791;
wire net_1419;
wire net_3239;
wire net_2188;
wire net_1051;
wire net_2364;
wire x1071;
wire net_942;
wire net_1981;
wire net_1515;
wire net_1218;
wire net_1573;
wire net_1494;
wire net_361;
wire net_3286;
wire net_2890;
wire net_2154;
wire net_1726;
wire x6573;
wire net_305;
wire net_1905;
wire net_1398;
wire net_2540;
wire net_3099;
wire net_3298;
wire net_1125;
wire net_2230;
wire net_144;
wire net_227;
wire net_1144;
wire net_1794;
wire net_3592;
wire net_1022;
wire net_1415;
wire net_3485;
wire net_2260;
wire net_2865;
wire net_3606;
wire net_2886;
wire net_3317;
wire net_702;
wire net_1921;
wire x3819;
wire net_1477;
wire net_3195;
wire net_3853;
wire net_3210;
wire x5957;
wire net_3318;
wire net_1230;
wire net_2135;
wire net_667;
wire net_853;
wire net_212;
wire net_914;
wire net_1193;
wire net_1425;
wire net_1122;
wire net_875;
wire net_1813;
wire net_1092;
wire net_627;
wire x4184;
wire net_2039;
wire net_983;
wire net_355;
wire net_1456;
wire net_723;
wire net_2227;
wire net_2483;
wire net_3962;
wire net_2473;
wire x5294;
wire net_275;
wire net_399;
wire x6799;
wire net_2914;
wire net_1390;
wire net_218;
wire net_2590;
wire net_1112;
wire x2403;
wire net_1273;
wire net_3283;
wire net_1137;
wire net_3948;
wire net_2114;
wire net_2506;
wire x3580;
wire net_3230;
wire net_285;
wire net_3819;
wire net_1310;
wire net_254;
wire net_2499;
wire net_1501;
wire net_1297;
wire net_3003;
wire net_1304;
wire net_574;
wire net_2177;
wire net_3357;

// Start cells
DFF_X2 inst_1783 ( .QN(net_2423), .D(net_757), .CK(net_3451) );
CLKBUF_X2 inst_2685 ( .A(net_2476), .Z(net_2477) );
OAI211_X2 inst_481 ( .C2(net_2314), .C1(net_1052), .ZN(net_1027), .A(net_890), .B(net_860) );
CLKBUF_X2 inst_4123 ( .A(net_3914), .Z(net_3915) );
DFF_X2 inst_1751 ( .QN(net_2345), .D(net_1446), .CK(net_4012) );
AOI22_X2 inst_2235 ( .B2(net_2162), .A1(net_1967), .B1(net_1474), .ZN(net_1395), .A2(net_1199) );
NAND2_X2 inst_779 ( .ZN(net_1348), .A2(net_1292), .A1(net_1278) );
AOI22_X2 inst_2205 ( .A2(net_2178), .B2(net_2145), .A1(net_1916), .ZN(net_1476), .B1(net_1474) );
CLKBUF_X2 inst_2858 ( .A(net_2649), .Z(net_2650) );
CLKBUF_X2 inst_4131 ( .A(net_3464), .Z(net_3923) );
OAI211_X2 inst_452 ( .C1(net_1639), .ZN(net_1103), .A(net_827), .B(net_669), .C2(net_395) );
OAI22_X2 inst_214 ( .A2(net_2235), .A1(net_2013), .B1(net_1404), .B2(net_207), .ZN(x1897) );
CLKBUF_X2 inst_3061 ( .A(net_2852), .Z(net_2853) );
CLKBUF_X2 inst_4228 ( .A(net_2861), .Z(net_4020) );
NOR2_X2 inst_548 ( .A2(net_2413), .ZN(net_608), .A1(net_603) );
CLKBUF_X2 inst_4144 ( .A(net_3935), .Z(net_3936) );
NAND2_X4 inst_728 ( .A2(net_1982), .ZN(net_1780), .A1(net_1779) );
CLKBUF_X2 inst_3121 ( .A(net_2912), .Z(net_2913) );
CLKBUF_X2 inst_2780 ( .A(net_2571), .Z(net_2572) );
AOI222_X1 inst_2485 ( .B1(net_1995), .A1(net_1749), .B2(net_1565), .ZN(net_1015), .C1(net_782), .A2(net_167), .C2(x3383) );
CLKBUF_X2 inst_4152 ( .A(net_3943), .Z(net_3944) );
AOI22_X2 inst_2217 ( .A2(net_2386), .B2(net_2109), .A1(net_1960), .B1(net_1915), .ZN(net_1463) );
NAND2_X2 inst_850 ( .A2(net_1908), .A1(net_1840), .ZN(net_1256) );
CLKBUF_X2 inst_3347 ( .A(net_3138), .Z(net_3139) );
CLKBUF_X2 inst_3130 ( .A(net_2921), .Z(net_2922) );
CLKBUF_X2 inst_2844 ( .A(net_2635), .Z(net_2636) );
AOI222_X1 inst_2492 ( .B1(net_1995), .A1(net_1751), .B2(net_1559), .C1(net_1020), .ZN(net_1008), .A2(net_161), .C2(x3483) );
CLKBUF_X2 inst_4136 ( .A(net_3927), .Z(net_3928) );
CLKBUF_X2 inst_3582 ( .A(net_2772), .Z(net_3374) );
INV_X4 inst_1228 ( .ZN(net_410), .A(net_397) );
CLKBUF_X2 inst_3480 ( .A(net_3271), .Z(net_3272) );
CLKBUF_X2 inst_4221 ( .A(net_2452), .Z(net_4013) );
NOR2_X4 inst_521 ( .ZN(net_416), .A1(net_380), .A2(net_378) );
INV_X16 inst_1685 ( .ZN(net_961), .A(net_633) );
AOI221_X2 inst_2511 ( .B2(net_2248), .A(net_2056), .B1(net_1893), .ZN(net_1770), .C1(net_910), .C2(net_815) );
AOI22_X2 inst_2438 ( .B1(net_2096), .ZN(net_1856), .A2(net_1855), .A1(net_1769), .B2(net_1539) );
INV_X2 inst_1655 ( .A(net_2290), .ZN(net_344) );
CLKBUF_X2 inst_3578 ( .A(net_2581), .Z(net_3370) );
CLKBUF_X2 inst_2772 ( .A(net_2488), .Z(net_2564) );
AOI21_X2 inst_2543 ( .A(net_1971), .ZN(net_595), .B1(net_514), .B2(net_356) );
OAI22_X2 inst_237 ( .B2(net_2259), .ZN(net_748), .A2(net_747), .A1(net_745), .B1(net_534) );
NAND2_X2 inst_813 ( .ZN(net_1300), .A1(net_1267), .A2(net_1224) );
SDFF_X2 inst_51 ( .SE(net_1768), .SI(net_1528), .Q(net_78), .D(net_78), .CK(net_3201) );
DFF_X2 inst_1837 ( .Q(net_1526), .CK(net_3096), .D(x5370) );
NAND2_X2 inst_1066 ( .A1(net_2027), .ZN(net_1732), .A2(net_1156) );
NAND2_X2 inst_974 ( .A2(net_1566), .A1(net_961), .ZN(net_865) );
CLKBUF_X2 inst_3392 ( .A(net_2830), .Z(net_3184) );
AOI22_X2 inst_2342 ( .B1(net_2197), .A1(net_2038), .A2(net_1572), .B2(net_1522), .ZN(net_822) );
CLKBUF_X2 inst_3291 ( .A(net_2518), .Z(net_3083) );
AOI22_X2 inst_2294 ( .B2(net_1573), .A2(net_1284), .ZN(net_963), .A1(net_962), .B1(net_961) );
INV_X2 inst_1617 ( .ZN(net_200), .A(x4752) );
OR2_X1 inst_151 ( .A1(net_2168), .A2(x3921), .ZN(x1322) );
SDFF_X2 inst_64 ( .Q(net_1574), .D(net_1574), .SE(net_498), .CK(net_3122), .SI(x6727) );
AOI22_X2 inst_2256 ( .B2(net_2120), .A1(net_1967), .B1(net_1474), .ZN(net_1374), .A2(net_1240) );
NAND2_X2 inst_1001 ( .A2(net_2123), .A1(net_979), .ZN(net_672) );
CLKBUF_X2 inst_4051 ( .A(net_3842), .Z(net_3843) );
DFFR_X1 inst_2106 ( .QN(net_2296), .RN(net_1347), .D(net_954), .CK(net_3082) );
NAND2_X4 inst_743 ( .ZN(net_2198), .A1(net_1962), .A2(net_1593) );
CLKBUF_X2 inst_2723 ( .A(net_2503), .Z(net_2515) );
CLKBUF_X2 inst_3931 ( .A(net_2657), .Z(net_3723) );
CLKBUF_X2 inst_3033 ( .A(net_2447), .Z(net_2825) );
CLKBUF_X2 inst_2925 ( .A(net_2716), .Z(net_2717) );
CLKBUF_X2 inst_3867 ( .A(net_3658), .Z(net_3659) );
DFF_X2 inst_1828 ( .QN(net_2206), .CK(net_2866), .D(x6550) );
DFFR_X2 inst_2072 ( .QN(net_1754), .RN(net_1347), .D(net_1247), .CK(net_3988) );
INV_X2 inst_1603 ( .ZN(net_208), .A(x6334) );
DFF_X2 inst_1809 ( .Q(net_1524), .CK(net_2456), .D(x5317) );
OAI21_X2 inst_340 ( .B1(net_1507), .ZN(net_1490), .A(net_1466), .B2(net_1048) );
CLKBUF_X2 inst_3388 ( .A(net_3179), .Z(net_3180) );
CLKBUF_X2 inst_3735 ( .A(net_2749), .Z(net_3527) );
CLKBUF_X2 inst_2675 ( .A(net_2466), .Z(net_2467) );
OAI22_X2 inst_158 ( .B1(net_1427), .A1(net_1426), .B2(net_235), .A2(net_96), .ZN(x1548) );
OR2_X2 inst_141 ( .ZN(net_407), .A2(x6207), .A1(x6188) );
AOI21_X2 inst_2520 ( .B1(net_1669), .A(net_1139), .ZN(net_1138), .B2(net_302) );
INV_X2 inst_1490 ( .A(net_2352), .ZN(net_1213) );
NOR2_X4 inst_507 ( .A2(net_2329), .ZN(net_1161), .A1(net_1146) );
NOR2_X2 inst_571 ( .A2(net_2331), .A1(net_2329), .ZN(net_321) );
CLKBUF_X2 inst_4011 ( .A(net_2562), .Z(net_3803) );
CLKBUF_X2 inst_3709 ( .A(net_3500), .Z(net_3501) );
DFF_X1 inst_1974 ( .Q(net_2140), .D(net_1042), .CK(net_3111) );
DFF_X1 inst_2017 ( .QN(net_2224), .D(net_1847), .CK(net_3099) );
NAND2_X2 inst_884 ( .ZN(net_1164), .A1(net_761), .A2(net_84) );
INV_X8 inst_1154 ( .A(net_1741), .ZN(net_1740) );
NAND2_X4 inst_711 ( .ZN(net_1171), .A1(net_1161), .A2(net_285) );
NAND2_X2 inst_827 ( .A1(net_1840), .ZN(net_1288), .A2(net_327) );
OAI211_X2 inst_469 ( .C2(net_2322), .C1(net_1054), .ZN(net_1042), .A(net_905), .B(net_877) );
CLKBUF_X2 inst_3040 ( .A(net_2831), .Z(net_2832) );
CLKBUF_X2 inst_2980 ( .A(net_2771), .Z(net_2772) );
CLKBUF_X2 inst_4191 ( .A(net_3123), .Z(net_3983) );
CLKBUF_X2 inst_3870 ( .A(net_2805), .Z(net_3662) );
XNOR2_X2 inst_18 ( .B(net_2337), .ZN(net_1179), .A(net_1166) );
NAND2_X2 inst_915 ( .A1(net_975), .A2(net_778), .ZN(x2971) );
CLKBUF_X2 inst_4128 ( .A(net_3919), .Z(net_3920) );
AOI22_X2 inst_2263 ( .ZN(net_1691), .A2(net_1543), .A1(net_1000), .B1(net_999), .B2(net_318) );
AOI22_X2 inst_2339 ( .B1(net_2197), .A1(net_2038), .A2(net_1565), .B2(net_1529), .ZN(net_825) );
CLKBUF_X2 inst_3549 ( .A(net_3293), .Z(net_3341) );
CLKBUF_X2 inst_3501 ( .A(net_3292), .Z(net_3293) );
INV_X4 inst_1216 ( .ZN(net_515), .A(net_499) );
CLKBUF_X2 inst_3936 ( .A(net_3727), .Z(net_3728) );
NAND2_X2 inst_952 ( .A1(net_1830), .A2(net_1747), .ZN(net_985) );
CLKBUF_X2 inst_4175 ( .A(net_3966), .Z(net_3967) );
INV_X2 inst_1668 ( .A(net_2335), .ZN(net_1812) );
NAND2_X4 inst_721 ( .A1(net_1873), .ZN(net_1595), .A2(net_442) );
OAI22_X2 inst_293 ( .A1(net_1615), .B1(net_1406), .B2(net_262), .A2(net_137), .ZN(x210) );
CLKBUF_X2 inst_3744 ( .A(net_3535), .Z(net_3536) );
CLKBUF_X2 inst_3009 ( .A(net_2800), .Z(net_2801) );
INV_X2 inst_1366 ( .A(net_1018), .ZN(x2543) );
CLKBUF_X2 inst_3102 ( .A(net_2893), .Z(net_2894) );
CLKBUF_X2 inst_2695 ( .A(net_2483), .Z(net_2487) );
CLKBUF_X2 inst_3860 ( .A(net_3651), .Z(net_3652) );
DFF_X1 inst_1915 ( .D(net_1318), .QN(net_128), .CK(net_3794) );
CLKBUF_X2 inst_2794 ( .A(net_2525), .Z(net_2586) );
DFF_X1 inst_2063 ( .QN(net_2375), .D(net_415), .CK(net_3961) );
INV_X4 inst_1254 ( .A(net_1580), .ZN(net_958) );
CLKBUF_X2 inst_2953 ( .A(net_2744), .Z(net_2745) );
CLKBUF_X2 inst_3553 ( .A(net_3344), .Z(net_3345) );
CLKBUF_X2 inst_3723 ( .A(net_3148), .Z(net_3515) );
CLKBUF_X2 inst_3521 ( .A(net_3312), .Z(net_3313) );
DFF_X2 inst_1811 ( .Q(net_1519), .CK(net_2599), .D(x5868) );
SDFF_X2 inst_98 ( .SE(net_488), .Q(net_168), .D(net_168), .CK(net_2708), .SI(x4461) );
CLKBUF_X2 inst_3440 ( .A(net_3231), .Z(net_3232) );
CLKBUF_X2 inst_3985 ( .A(net_3776), .Z(net_3777) );
CLKBUF_X2 inst_3087 ( .A(net_2878), .Z(net_2879) );
DFF_X1 inst_2036 ( .Q(net_2397), .D(net_847), .CK(net_3032) );
NAND2_X2 inst_959 ( .A2(net_2165), .A1(net_1829), .ZN(net_926) );
CLKBUF_X2 inst_4001 ( .A(net_3792), .Z(net_3793) );
DFF_X1 inst_2049 ( .QN(net_2405), .D(net_540), .CK(net_3750) );
NAND2_X2 inst_868 ( .A1(net_1838), .ZN(net_1214), .A2(net_1213) );
OAI22_X2 inst_163 ( .A1(net_1408), .B1(net_1406), .B2(net_227), .A2(net_133), .ZN(x297) );
OAI21_X2 inst_394 ( .B1(net_1829), .ZN(net_1113), .B2(net_953), .A(net_930) );
OAI22_X2 inst_201 ( .A2(net_2230), .B1(net_1406), .A1(net_1405), .B2(net_196), .ZN(x1997) );
NOR2_X2 inst_605 ( .A2(net_2258), .ZN(net_1926), .A1(net_520) );
CLKBUF_X2 inst_3627 ( .A(net_3418), .Z(net_3419) );
NAND2_X2 inst_1084 ( .A1(net_1840), .ZN(net_1839), .A2(net_331) );
OAI22_X2 inst_304 ( .A2(net_2215), .B1(net_1895), .A1(net_1405), .B2(net_230), .ZN(x2304) );
DFF_X2 inst_1814 ( .Q(net_1533), .CK(net_2500), .D(x5493) );
CLKBUF_X2 inst_2799 ( .A(net_2529), .Z(net_2591) );
CLKBUF_X2 inst_4157 ( .A(net_3948), .Z(net_3949) );
NAND2_X2 inst_1027 ( .ZN(net_519), .A2(net_507), .A1(net_501) );
INV_X8 inst_1143 ( .A(net_2018), .ZN(net_589) );
INV_X4 inst_1345 ( .A(net_2339), .ZN(net_2076) );
CLKBUF_X2 inst_2947 ( .A(net_2738), .Z(net_2739) );
DFF_X1 inst_2048 ( .Q(net_2391), .D(net_546), .CK(net_3280) );
CLKBUF_X2 inst_2948 ( .A(net_2739), .Z(net_2740) );
OAI21_X2 inst_361 ( .B2(net_2405), .B1(net_1441), .ZN(net_1433), .A(net_1371) );
CLKBUF_X2 inst_3608 ( .A(net_2883), .Z(net_3400) );
CLKBUF_X2 inst_3400 ( .A(net_2664), .Z(net_3192) );
NAND2_X2 inst_1016 ( .ZN(net_766), .A1(net_611), .A2(net_513) );
CLKBUF_X2 inst_4147 ( .A(net_3938), .Z(net_3939) );
INV_X2 inst_1538 ( .ZN(net_257), .A(x6417) );
NAND2_X2 inst_848 ( .A2(net_1913), .A1(net_1840), .ZN(net_1258) );
DFF_X1 inst_1931 ( .D(net_1119), .QN(net_60), .CK(net_3502) );
CLKBUF_X2 inst_3002 ( .A(net_2793), .Z(net_2794) );
AOI222_X1 inst_2479 ( .B1(net_1995), .A1(net_1751), .B2(net_1573), .ZN(net_1022), .C1(net_1020), .A2(net_175), .C2(x3245) );
AND2_X4 inst_2578 ( .A1(net_1668), .ZN(net_513), .A2(net_512) );
NAND2_X2 inst_786 ( .A1(net_1822), .ZN(net_1327), .A2(net_1212) );
CLKBUF_X2 inst_2940 ( .A(net_2731), .Z(net_2732) );
DFF_X1 inst_1996 ( .Q(net_2160), .D(net_1085), .CK(net_3519) );
INV_X2 inst_1554 ( .ZN(net_246), .A(x4926) );
INV_X2 inst_1542 ( .ZN(net_254), .A(x4658) );
XOR2_X2 inst_2 ( .A(net_1199), .Z(net_415), .B(net_414) );
CLKBUF_X2 inst_3340 ( .A(net_3131), .Z(net_3132) );
NAND4_X2 inst_644 ( .ZN(net_2084), .A4(net_2076), .A3(net_1284), .A2(net_1186), .A1(net_1184) );
CLKBUF_X2 inst_3474 ( .A(net_2673), .Z(net_3266) );
INV_X2 inst_1380 ( .A(net_1004), .ZN(x2773) );
CLKBUF_X2 inst_2806 ( .A(net_2572), .Z(net_2598) );
NOR2_X2 inst_578 ( .A1(net_1896), .ZN(net_1724), .A2(net_46) );
NAND2_X2 inst_888 ( .ZN(net_1135), .A1(net_998), .A2(net_850) );
DFF_X2 inst_1769 ( .QN(net_2432), .D(net_1646), .CK(net_3031) );
CLKBUF_X2 inst_3891 ( .A(net_3550), .Z(net_3683) );
CLKBUF_X2 inst_3625 ( .A(net_3416), .Z(net_3417) );
CLKBUF_X2 inst_4008 ( .A(net_3012), .Z(net_3800) );
CLKBUF_X2 inst_3472 ( .A(net_3263), .Z(net_3264) );
AND2_X4 inst_2581 ( .A2(net_2379), .A1(net_2200), .ZN(net_422) );
CLKBUF_X2 inst_4110 ( .A(net_3901), .Z(net_3902) );
INV_X2 inst_1498 ( .A(net_2423), .ZN(net_646) );
OAI21_X2 inst_432 ( .ZN(net_1844), .B2(net_1843), .B1(net_1842), .A(net_1839) );
OAI22_X2 inst_282 ( .A2(net_2237), .A1(net_2017), .B1(net_1406), .B2(net_228), .ZN(x1854) );
INV_X2 inst_1358 ( .ZN(net_1163), .A(net_1162) );
AOI22_X2 inst_2322 ( .A2(net_2159), .B1(net_2096), .A1(net_1769), .B2(net_1541), .ZN(net_887) );
NOR2_X4 inst_513 ( .ZN(net_511), .A2(net_492), .A1(net_464) );
CLKBUF_X2 inst_3266 ( .A(net_3057), .Z(net_3058) );
CLKBUF_X2 inst_3171 ( .A(net_2962), .Z(net_2963) );
INV_X2 inst_1630 ( .A(net_1590), .ZN(net_191) );
INV_X2 inst_1586 ( .A(net_1587), .ZN(net_222) );
CLKBUF_X2 inst_3385 ( .A(net_3176), .Z(net_3177) );
CLKBUF_X2 inst_3182 ( .A(net_2973), .Z(net_2974) );
INV_X2 inst_1572 ( .ZN(net_231), .A(x4578) );
CLKBUF_X2 inst_2866 ( .A(net_2657), .Z(net_2658) );
NAND2_X2 inst_774 ( .A2(net_1758), .A1(net_1714), .ZN(net_1397) );
AOI22_X2 inst_2292 ( .B2(net_1574), .ZN(net_967), .A1(net_962), .B1(net_961), .A2(net_309) );
NAND2_X2 inst_838 ( .A1(net_1745), .ZN(net_1275), .A2(net_1265) );
CLKBUF_X2 inst_2766 ( .A(net_2557), .Z(net_2558) );
INV_X2 inst_1508 ( .A(net_2421), .ZN(net_357) );
INV_X4 inst_1222 ( .ZN(net_450), .A(net_449) );
INV_X2 inst_1405 ( .A(net_571), .ZN(x1029) );
CLKBUF_X2 inst_3407 ( .A(net_2459), .Z(net_3199) );
CLKBUF_X2 inst_4058 ( .A(net_3849), .Z(net_3850) );
NAND2_X2 inst_1073 ( .A1(net_2104), .ZN(net_1814), .A2(net_327) );
AOI22_X2 inst_2323 ( .A2(net_2158), .B1(net_2096), .A1(net_1769), .B2(net_1542), .ZN(net_886) );
CLKBUF_X2 inst_3741 ( .A(net_3532), .Z(net_3533) );
CLKBUF_X2 inst_2749 ( .A(net_2455), .Z(net_2541) );
INV_X2 inst_1449 ( .ZN(net_378), .A(net_321) );
OR3_X4 inst_127 ( .ZN(net_2174), .A1(net_2026), .A2(net_2023), .A3(net_1575) );
DFF_X1 inst_2013 ( .QN(net_2215), .D(net_1072), .CK(net_3330) );
OAI22_X2 inst_187 ( .B1(net_1427), .A1(net_529), .B2(net_212), .A2(net_87), .ZN(x1682) );
OAI22_X2 inst_206 ( .A2(net_2224), .B1(net_1406), .A1(net_1405), .B2(net_241), .ZN(x2134) );
CLKBUF_X2 inst_3739 ( .A(net_3517), .Z(net_3531) );
CLKBUF_X2 inst_3029 ( .A(net_2777), .Z(net_2821) );
INV_X4 inst_1268 ( .A(net_2334), .ZN(net_1276) );
SDFFR_X1 inst_122 ( .SE(net_1829), .D(net_1537), .RN(net_1347), .SI(net_50), .Q(net_50), .CK(net_3054) );
CLKBUF_X2 inst_2756 ( .A(net_2547), .Z(net_2548) );
OAI21_X2 inst_405 ( .B2(net_2422), .ZN(net_881), .B1(net_880), .A(net_631) );
DFF_X2 inst_1731 ( .QN(net_2319), .D(net_1498), .CK(net_3055) );
NOR3_X4 inst_492 ( .ZN(net_2024), .A2(net_2023), .A1(net_2022), .A3(net_1575) );
CLKBUF_X2 inst_2960 ( .A(net_2632), .Z(net_2752) );
DFF_X1 inst_1909 ( .D(net_1314), .QN(net_132), .CK(net_3441) );
CLKBUF_X2 inst_3912 ( .A(net_3062), .Z(net_3704) );
AOI22_X2 inst_2306 ( .A2(net_2141), .B1(net_2096), .A1(net_1769), .B2(net_1537), .ZN(net_903) );
SDFF_X2 inst_82 ( .SE(net_487), .Q(net_164), .D(net_164), .CK(net_2742), .SI(x4549) );
CLKBUF_X2 inst_4187 ( .A(net_3978), .Z(net_3979) );
INV_X2 inst_1646 ( .A(net_2298), .ZN(net_306) );
CLKBUF_X2 inst_2892 ( .A(net_2683), .Z(net_2684) );
NAND2_X2 inst_1121 ( .ZN(net_2106), .A2(net_2105), .A1(net_2104) );
NAND2_X2 inst_1102 ( .ZN(net_1989), .A1(net_1988), .A2(net_507) );
CLKBUF_X2 inst_3161 ( .A(net_2952), .Z(net_2953) );
CLKBUF_X2 inst_3187 ( .A(net_2978), .Z(net_2979) );
OAI22_X2 inst_307 ( .B1(net_1895), .A1(net_1408), .B2(net_198), .A2(net_116), .ZN(x535) );
CLKBUF_X2 inst_2816 ( .A(net_2562), .Z(net_2608) );
NAND3_X2 inst_702 ( .ZN(net_2057), .A1(net_1810), .A3(net_799), .A2(net_653) );
DFF_X1 inst_2034 ( .QN(net_2403), .D(net_916), .CK(net_4029) );
INV_X2 inst_1505 ( .A(net_2066), .ZN(net_287) );
NAND2_X4 inst_717 ( .ZN(net_522), .A1(net_485), .A2(net_480) );
OAI22_X2 inst_276 ( .B2(net_2306), .B1(net_1865), .ZN(net_1608), .A1(net_1597), .A2(net_713) );
AOI222_X1 inst_2482 ( .B1(net_1995), .A1(net_1751), .B2(net_1569), .C1(net_1020), .ZN(net_1018), .A2(net_171), .C2(x3314) );
CLKBUF_X2 inst_2957 ( .A(net_2748), .Z(net_2749) );
CLKBUF_X2 inst_3339 ( .A(net_3130), .Z(net_3131) );
CLKBUF_X2 inst_3791 ( .A(net_3582), .Z(net_3583) );
CLKBUF_X2 inst_2711 ( .A(net_2502), .Z(net_2503) );
CLKBUF_X2 inst_3531 ( .A(net_2800), .Z(net_3323) );
CLKBUF_X2 inst_2753 ( .A(net_2544), .Z(net_2545) );
CLKBUF_X2 inst_3672 ( .A(net_3320), .Z(net_3464) );
SDFF_X2 inst_91 ( .SE(net_488), .Q(net_152), .D(net_152), .CK(net_2572), .SI(x4899) );
DFF_X2 inst_1762 ( .QN(net_1591), .D(net_1149), .CK(net_3960) );
OR2_X4 inst_132 ( .ZN(net_1976), .A1(net_1754), .A2(net_1581) );
DFF_X1 inst_2023 ( .QN(net_2236), .D(net_2057), .CK(net_3222) );
CLKBUF_X2 inst_2779 ( .A(net_2470), .Z(net_2571) );
CLKBUF_X2 inst_3686 ( .A(net_3477), .Z(net_3478) );
CLKBUF_X2 inst_3842 ( .A(net_3633), .Z(net_3634) );
INV_X1 inst_1703 ( .A(net_2028), .ZN(net_1296) );
CLKBUF_X2 inst_3545 ( .A(net_3336), .Z(net_3337) );
CLKBUF_X2 inst_3611 ( .A(net_3402), .Z(net_3403) );
CLKBUF_X2 inst_2928 ( .A(net_2719), .Z(net_2720) );
CLKBUF_X2 inst_3813 ( .A(net_3457), .Z(net_3605) );
OAI21_X2 inst_400 ( .ZN(net_991), .A(net_845), .B1(net_843), .B2(net_593) );
CLKBUF_X2 inst_2991 ( .A(net_2782), .Z(net_2783) );
NOR2_X2 inst_614 ( .ZN(net_2005), .A2(net_1945), .A1(net_1155) );
CLKBUF_X2 inst_3513 ( .A(net_3118), .Z(net_3305) );
DFF_X1 inst_1896 ( .D(net_1319), .QN(net_125), .CK(net_3802) );
OAI22_X2 inst_261 ( .B2(net_2254), .A2(net_939), .A1(net_714), .ZN(net_701), .B1(net_534) );
NAND2_X2 inst_1031 ( .ZN(net_464), .A1(net_447), .A2(net_349) );
NAND2_X2 inst_945 ( .ZN(net_997), .A1(net_842), .A2(net_764) );
OAI22_X2 inst_268 ( .B2(net_2307), .B1(net_1865), .ZN(net_1599), .A1(net_951), .A2(net_711) );
INV_X2 inst_1518 ( .ZN(net_265), .A(x3986) );
OAI21_X2 inst_369 ( .B1(net_1443), .ZN(net_1420), .A(net_1386), .B2(net_1157) );
DFF_X1 inst_1900 ( .D(net_1311), .QN(net_137), .CK(net_3648) );
CLKBUF_X2 inst_3975 ( .A(net_3766), .Z(net_3767) );
OAI21_X2 inst_327 ( .B1(net_2041), .ZN(net_1503), .A(net_1469), .B2(net_352) );
CLKBUF_X2 inst_3509 ( .A(net_2874), .Z(net_3301) );
CLKBUF_X2 inst_2916 ( .A(net_2707), .Z(net_2708) );
INV_X4 inst_1286 ( .ZN(net_323), .A(net_47) );
OAI22_X2 inst_266 ( .B2(net_2202), .A2(net_958), .ZN(net_652), .B1(net_554), .A1(net_553) );
DFF_X1 inst_2051 ( .QN(net_2404), .D(net_2183), .CK(net_3746) );
CLKBUF_X2 inst_3853 ( .A(net_2885), .Z(net_3645) );
INV_X4 inst_1198 ( .A(net_1970), .ZN(net_680) );
SDFF_X2 inst_77 ( .Q(net_1545), .D(net_1545), .SE(net_491), .CK(net_2670), .SI(x7484) );
OAI22_X2 inst_171 ( .B1(net_2168), .A1(net_775), .B2(net_390), .A2(net_112), .ZN(x1357) );
CLKBUF_X2 inst_3097 ( .A(net_2888), .Z(net_2889) );
CLKBUF_X2 inst_3661 ( .A(net_2469), .Z(net_3453) );
OAI21_X2 inst_374 ( .B2(net_2402), .B1(net_1443), .ZN(net_1415), .A(net_1374) );
NOR2_X4 inst_502 ( .ZN(net_1250), .A1(net_1192), .A2(net_411) );
SDFF_X2 inst_103 ( .SE(net_487), .Q(net_150), .D(net_150), .CK(net_2570), .SI(x4949) );
CLKBUF_X2 inst_3690 ( .A(net_3481), .Z(net_3482) );
CLKBUF_X2 inst_3221 ( .A(net_3012), .Z(net_3013) );
CLKBUF_X2 inst_3645 ( .A(net_3436), .Z(net_3437) );
INV_X2 inst_1598 ( .ZN(net_212), .A(x4232) );
CLKBUF_X2 inst_3738 ( .A(net_3529), .Z(net_3530) );
OAI21_X2 inst_357 ( .B2(net_2400), .B1(net_1441), .ZN(net_1437), .A(net_1376) );
CLKBUF_X2 inst_2855 ( .A(net_2646), .Z(net_2647) );
CLKBUF_X2 inst_4092 ( .A(net_3883), .Z(net_3884) );
DFF_X1 inst_2058 ( .Q(net_2386), .D(net_474), .CK(net_3365) );
NAND2_X2 inst_809 ( .A2(net_1681), .ZN(net_1304), .A1(net_1269) );
CLKBUF_X2 inst_3980 ( .A(net_3771), .Z(net_3772) );
CLKBUF_X2 inst_3675 ( .A(net_3466), .Z(net_3467) );
CLKBUF_X2 inst_3152 ( .A(net_2943), .Z(net_2944) );
CLKBUF_X2 inst_4161 ( .A(net_3599), .Z(net_3953) );
CLKBUF_X2 inst_3758 ( .A(net_2542), .Z(net_3550) );
AOI211_X2 inst_2562 ( .C2(net_2136), .C1(net_1929), .A(net_1882), .B(net_1785), .ZN(net_676) );
INV_X4 inst_1234 ( .A(net_2329), .ZN(net_1262) );
NAND2_X2 inst_912 ( .A1(net_978), .A2(net_781), .ZN(x2886) );
AOI22_X2 inst_2398 ( .B1(net_2197), .ZN(net_1626), .A1(net_1621), .B2(net_1515), .A2(net_1201) );
AND2_X4 inst_2595 ( .A2(net_2202), .ZN(net_2169), .A1(net_277) );
NAND2_X2 inst_1022 ( .A1(net_1915), .A2(net_786), .ZN(net_548) );
CLKBUF_X2 inst_3196 ( .A(net_2506), .Z(net_2988) );
AOI22_X2 inst_2371 ( .B2(net_2163), .A1(net_2038), .A2(net_1562), .B1(net_979), .ZN(net_685) );
CLKBUF_X2 inst_2939 ( .A(net_2730), .Z(net_2731) );
CLKBUF_X2 inst_4025 ( .A(net_2987), .Z(net_3817) );
OAI21_X2 inst_322 ( .ZN(net_1509), .B1(net_1507), .A(net_1473), .B2(net_1036) );
INV_X4 inst_1223 ( .A(net_492), .ZN(net_446) );
CLKBUF_X2 inst_3516 ( .A(net_3307), .Z(net_3308) );
CLKBUF_X2 inst_2785 ( .A(net_2576), .Z(net_2577) );
CLKBUF_X2 inst_3906 ( .A(net_3697), .Z(net_3698) );
CLKBUF_X2 inst_4200 ( .A(net_3991), .Z(net_3992) );
CLKBUF_X2 inst_4188 ( .A(net_3979), .Z(net_3980) );
NAND3_X2 inst_681 ( .A3(net_2423), .A2(net_2176), .ZN(net_449), .A1(net_351) );
CLKBUF_X2 inst_4169 ( .A(net_2921), .Z(net_3961) );
CLKBUF_X2 inst_3902 ( .A(net_3693), .Z(net_3694) );
DFF_X1 inst_2010 ( .QN(net_2218), .D(net_1069), .CK(net_3332) );
CLKBUF_X2 inst_2915 ( .A(net_2706), .Z(net_2707) );
CLKBUF_X2 inst_3296 ( .A(net_3087), .Z(net_3088) );
CLKBUF_X2 inst_4181 ( .A(net_3582), .Z(net_3973) );
NAND2_X2 inst_871 ( .A1(net_1838), .ZN(net_1210), .A2(net_322) );
AOI22_X2 inst_2315 ( .A2(net_2147), .B1(net_2096), .A1(net_1769), .B2(net_1529), .ZN(net_894) );
CLKBUF_X2 inst_2684 ( .A(net_2475), .Z(net_2476) );
NAND2_X2 inst_962 ( .A2(net_1545), .A1(net_961), .ZN(net_878) );
NOR2_X4 inst_532 ( .A2(net_2204), .ZN(net_2064), .A1(net_1659) );
CLKBUF_X2 inst_3164 ( .A(net_2655), .Z(net_2956) );
CLKBUF_X2 inst_2965 ( .A(net_2496), .Z(net_2757) );
AOI22_X2 inst_2382 ( .A1(net_1718), .B1(net_1450), .B2(net_788), .ZN(net_643), .A2(net_356) );
DFF_X1 inst_2008 ( .QN(net_2225), .D(net_1081), .CK(net_3294) );
INV_X8 inst_1171 ( .A(net_2075), .ZN(net_2001) );
NAND4_X2 inst_641 ( .ZN(net_1940), .A3(net_1914), .A4(net_1845), .A2(net_1835), .A1(net_1760) );
CLKBUF_X2 inst_2969 ( .A(net_2725), .Z(net_2761) );
NOR3_X2 inst_498 ( .A2(net_2352), .A1(net_2351), .A3(net_2348), .ZN(net_385) );
CLKBUF_X2 inst_3314 ( .A(net_3105), .Z(net_3106) );
DFF_X1 inst_1988 ( .Q(net_2152), .D(net_1044), .CK(net_2968) );
AND2_X4 inst_2594 ( .A1(net_2418), .ZN(net_2167), .A2(net_1582) );
CLKBUF_X2 inst_4037 ( .A(net_3520), .Z(net_3829) );
DFF_X1 inst_1912 ( .D(net_1316), .QN(net_130), .CK(net_3506) );
CLKBUF_X2 inst_3976 ( .A(net_3767), .Z(net_3768) );
DFF_X2 inst_1831 ( .QN(net_2208), .CK(net_2695), .D(x6503) );
INV_X4 inst_1327 ( .A(net_2011), .ZN(net_1961) );
CLKBUF_X2 inst_3468 ( .A(net_3259), .Z(net_3260) );
OAI21_X2 inst_350 ( .B2(net_2374), .ZN(net_1446), .B1(net_1443), .A(net_1395) );
AOI22_X2 inst_2395 ( .B1(net_2197), .ZN(net_1623), .A1(net_1621), .B2(net_1537), .A2(net_1238) );
OAI22_X2 inst_231 ( .B2(net_2281), .B1(net_1865), .A1(net_1603), .ZN(net_943), .A2(net_707) );
NAND2_X2 inst_1119 ( .ZN(net_2097), .A1(net_2095), .A2(net_2035) );
CLKBUF_X2 inst_3309 ( .A(net_3100), .Z(net_3101) );
CLKBUF_X2 inst_3699 ( .A(net_3490), .Z(net_3491) );
INV_X4 inst_1255 ( .A(net_2364), .ZN(net_1196) );
AOI22_X2 inst_2317 ( .A2(net_2151), .B1(net_2096), .A1(net_1769), .B2(net_1523), .ZN(net_892) );
DFF_X2 inst_1791 ( .QN(net_2431), .D(net_1786), .CK(net_3888) );
INV_X2 inst_1452 ( .A(net_2429), .ZN(net_377) );
CLKBUF_X2 inst_3420 ( .A(net_3211), .Z(net_3212) );
CLKBUF_X2 inst_4077 ( .A(net_3868), .Z(net_3869) );
CLKBUF_X2 inst_3139 ( .A(net_2930), .Z(net_2931) );
NOR2_X4 inst_528 ( .ZN(net_1997), .A1(net_1983), .A2(net_372) );
AOI21_X2 inst_2558 ( .ZN(net_2187), .B2(net_1936), .A(net_1935), .B1(net_1339) );
NAND2_X2 inst_903 ( .ZN(net_1116), .A1(net_982), .A2(net_915) );
DFF_X2 inst_1725 ( .QN(net_2312), .D(net_1505), .CK(net_3134) );
INV_X2 inst_1396 ( .A(net_579), .ZN(x1018) );
OAI21_X2 inst_352 ( .B1(net_1736), .ZN(net_1444), .B2(net_1443), .A(net_1379) );
NAND2_X2 inst_846 ( .A1(net_1745), .ZN(net_1267), .A2(net_371) );
OAI22_X2 inst_286 ( .A1(net_1615), .B1(net_1407), .B2(net_247), .A2(net_118), .ZN(x518) );
CLKBUF_X2 inst_3504 ( .A(net_2493), .Z(net_3296) );
CLKBUF_X2 inst_3924 ( .A(net_3715), .Z(net_3716) );
DFF_X2 inst_1734 ( .QN(net_2318), .D(net_1497), .CK(net_3552) );
CLKBUF_X2 inst_3003 ( .A(net_2680), .Z(net_2795) );
CLKBUF_X2 inst_3841 ( .A(net_2656), .Z(net_3633) );
CLKBUF_X2 inst_3464 ( .A(net_3255), .Z(net_3256) );
CLKBUF_X2 inst_4050 ( .A(net_3841), .Z(net_3842) );
NAND2_X2 inst_1044 ( .A1(net_1743), .ZN(net_1671), .A2(net_1227) );
CLKBUF_X2 inst_3354 ( .A(net_3145), .Z(net_3146) );
AOI22_X2 inst_2370 ( .B2(net_2128), .A1(net_2038), .A2(net_1558), .B1(net_979), .ZN(net_686) );
CLKBUF_X2 inst_3882 ( .A(net_3673), .Z(net_3674) );
CLKBUF_X2 inst_2811 ( .A(net_2602), .Z(net_2603) );
CLKBUF_X2 inst_3014 ( .A(net_2805), .Z(net_2806) );
OR2_X2 inst_137 ( .A2(net_2202), .A1(net_1582), .ZN(net_512) );
OAI21_X2 inst_425 ( .ZN(net_427), .B1(net_426), .B2(x6207), .A(x5995) );
AOI211_X2 inst_2567 ( .C2(net_2140), .C1(net_1974), .ZN(net_1862), .A(net_1861), .B(net_557) );
CLKBUF_X2 inst_3206 ( .A(net_2460), .Z(net_2998) );
INV_X2 inst_1532 ( .ZN(net_261), .A(x4718) );
OAI22_X2 inst_227 ( .B2(net_2302), .B1(net_1865), .A1(net_951), .ZN(net_947), .A2(net_722) );
DFFR_X1 inst_2136 ( .QN(net_2268), .RN(net_1347), .D(net_729), .CK(net_2514) );
CLKBUF_X2 inst_3927 ( .A(net_2915), .Z(net_3719) );
CLKBUF_X2 inst_2891 ( .A(net_2682), .Z(net_2683) );
CLKBUF_X2 inst_2718 ( .A(net_2459), .Z(net_2510) );
AND4_X2 inst_2572 ( .A2(net_2050), .ZN(net_1908), .A3(net_1905), .A1(net_522), .A4(net_346) );
SDFF_X2 inst_58 ( .Q(net_1563), .D(net_1563), .SE(net_396), .CK(net_2936), .SI(x7087) );
CLKBUF_X2 inst_3633 ( .A(net_3424), .Z(net_3425) );
CLKBUF_X2 inst_4046 ( .A(net_3837), .Z(net_3838) );
CLKBUF_X2 inst_3365 ( .A(net_3156), .Z(net_3157) );
INV_X2 inst_1469 ( .A(net_1513), .ZN(net_848) );
CLKBUF_X2 inst_3254 ( .A(net_2657), .Z(net_3046) );
NAND2_X2 inst_983 ( .A2(net_1551), .A1(net_961), .ZN(net_856) );
DFF_X1 inst_1897 ( .D(net_1320), .QN(net_124), .CK(net_3801) );
CLKBUF_X2 inst_3159 ( .A(net_2809), .Z(net_2951) );
AOI21_X2 inst_2551 ( .ZN(net_441), .B2(net_370), .A(net_351), .B1(net_318) );
NOR2_X2 inst_581 ( .A2(net_2044), .ZN(net_1738), .A1(net_1737) );
XNOR2_X2 inst_28 ( .B(net_1213), .ZN(net_916), .A(net_642) );
AOI22_X2 inst_2424 ( .B2(net_2150), .B1(net_1974), .ZN(net_1798), .A1(net_1791), .A2(net_312) );
INV_X2 inst_1569 ( .A(net_2288), .ZN(net_284) );
CLKBUF_X2 inst_3144 ( .A(net_2935), .Z(net_2936) );
AND2_X2 inst_2633 ( .A1(net_594), .A2(x7215), .ZN(x768) );
DFF_X2 inst_1772 ( .QN(net_2379), .D(net_988), .CK(net_3861) );
NOR2_X2 inst_592 ( .A2(net_2253), .ZN(net_1881), .A1(net_520) );
CLKBUF_X2 inst_3666 ( .A(net_2562), .Z(net_3458) );
NAND2_X2 inst_993 ( .ZN(net_844), .A1(net_843), .A2(net_772) );
DFFR_X1 inst_2143 ( .QN(net_2277), .RN(net_1347), .D(net_710), .CK(net_2721) );
INV_X4 inst_1291 ( .ZN(net_811), .A(net_69) );
DFFR_X1 inst_2130 ( .QN(net_2261), .RN(net_1347), .D(net_743), .CK(net_2644) );
OAI21_X2 inst_359 ( .B2(net_2401), .B1(net_1443), .ZN(net_1435), .A(net_1375) );
NAND2_X2 inst_1055 ( .A1(net_1741), .ZN(net_1683), .A2(net_932) );
DFFR_X1 inst_2100 ( .QN(net_2289), .D(net_1612), .RN(net_1347), .CK(net_2850) );
CLKBUF_X2 inst_3948 ( .A(net_3739), .Z(net_3740) );
AOI22_X2 inst_2284 ( .A1(net_1996), .B1(net_1749), .A2(net_1550), .ZN(net_978), .B2(net_152) );
DFF_X1 inst_1962 ( .Q(net_2128), .D(net_1061), .CK(net_3491) );
NAND4_X2 inst_630 ( .A2(net_1918), .A1(net_1739), .ZN(net_1363), .A3(net_1296), .A4(net_421) );
INV_X4 inst_1273 ( .ZN(net_307), .A(net_55) );
NAND2_X2 inst_923 ( .A2(net_1635), .ZN(net_1091), .A1(net_690) );
NOR2_X4 inst_512 ( .A2(net_2354), .ZN(net_541), .A1(net_526) );
INV_X4 inst_1301 ( .ZN(net_1615), .A(net_1614) );
DFFR_X1 inst_2151 ( .QN(net_2254), .RN(net_1347), .D(net_701), .CK(net_2828) );
CLKBUF_X2 inst_2830 ( .A(net_2621), .Z(net_2622) );
NAND3_X4 inst_647 ( .ZN(net_2095), .A3(net_2064), .A1(net_1961), .A2(net_1831) );
CLKBUF_X2 inst_3054 ( .A(net_2845), .Z(net_2846) );
OAI22_X2 inst_194 ( .A2(net_2438), .B1(net_1427), .A1(net_529), .B2(net_458), .ZN(x1294) );
CLKBUF_X2 inst_3453 ( .A(net_2813), .Z(net_3245) );
CLKBUF_X2 inst_2985 ( .A(net_2776), .Z(net_2777) );
CLKBUF_X2 inst_3766 ( .A(net_2963), .Z(net_3558) );
NAND2_X2 inst_833 ( .A1(net_1745), .ZN(net_1281), .A2(net_1242) );
CLKBUF_X2 inst_3772 ( .A(net_3563), .Z(net_3564) );
CLKBUF_X2 inst_4210 ( .A(net_2721), .Z(net_4002) );
AOI21_X2 inst_2536 ( .A(net_1785), .B1(net_910), .ZN(net_795), .B2(net_794) );
DFF_X1 inst_2043 ( .QN(net_2406), .D(net_2182), .CK(net_3753) );
NAND2_X2 inst_960 ( .A1(net_1829), .ZN(net_925), .A2(net_324) );
SDFF_X2 inst_118 ( .Q(net_1550), .D(net_1550), .SE(net_491), .CK(net_2658), .SI(x7383) );
AOI22_X2 inst_2411 ( .B1(net_2197), .ZN(net_1640), .A1(net_1619), .B2(net_1540), .A2(net_1239) );
OAI21_X1 inst_442 ( .B2(net_2417), .ZN(net_1251), .B1(net_1250), .A(net_468) );
AOI221_X2 inst_2507 ( .B2(net_2123), .B1(net_1929), .A(net_1884), .C1(net_1863), .ZN(net_1761), .C2(net_323) );
AOI22_X2 inst_2245 ( .B2(net_2131), .A1(net_1967), .B1(net_1915), .ZN(net_1385), .A2(net_1190) );
XNOR2_X2 inst_38 ( .A(net_1205), .ZN(net_465), .B(net_457) );
AND2_X4 inst_2601 ( .A1(net_2422), .A2(net_2421), .ZN(net_2176) );
DFF_X1 inst_2037 ( .QN(net_2402), .D(net_692), .CK(net_3790) );
OAI21_X2 inst_381 ( .A(net_1939), .B2(net_1356), .ZN(net_1355), .B1(net_1335) );
CLKBUF_X2 inst_3837 ( .A(net_3628), .Z(net_3629) );
DFF_X1 inst_1925 ( .D(net_1120), .QN(net_63), .CK(net_3503) );
NAND2_X2 inst_883 ( .ZN(net_1165), .A1(net_762), .A2(net_84) );
XNOR2_X2 inst_40 ( .A(net_2172), .ZN(net_1736), .B(net_1735) );
INV_X4 inst_1249 ( .ZN(net_1036), .A(net_846) );
NAND2_X4 inst_756 ( .ZN(net_2012), .A1(net_451), .A2(x5995) );
CLKBUF_X2 inst_4099 ( .A(net_3514), .Z(net_3891) );
INV_X2 inst_1416 ( .A(net_560), .ZN(x1144) );
INV_X4 inst_1318 ( .ZN(net_1851), .A(net_1850) );
OAI21_X2 inst_439 ( .ZN(net_2082), .B1(net_2081), .A(net_2078), .B2(net_2076) );
INV_X4 inst_1188 ( .ZN(net_1146), .A(net_1145) );
INV_X8 inst_1165 ( .ZN(net_1960), .A(net_1959) );
AND2_X2 inst_2644 ( .ZN(net_394), .A2(net_393), .A1(net_286) );
NAND2_X2 inst_1070 ( .ZN(net_1777), .A2(net_82), .A1(x5181) );
AND2_X2 inst_2626 ( .A1(net_594), .A2(x7526), .ZN(x902) );
AOI222_X2 inst_2454 ( .C1(net_2014), .A2(net_1569), .A1(net_590), .B1(net_589), .ZN(net_582), .B2(net_171), .C2(x5338) );
CLKBUF_X2 inst_3601 ( .A(net_2964), .Z(net_3393) );
CLKBUF_X2 inst_3873 ( .A(net_2817), .Z(net_3665) );
NAND2_X2 inst_992 ( .A1(net_1717), .ZN(net_845), .A2(net_377) );
NOR4_X2 inst_488 ( .A4(net_2363), .A3(net_2362), .A2(net_2361), .A1(net_2360), .ZN(net_2189) );
OAI21_X2 inst_387 ( .B1(net_1842), .ZN(net_1342), .A(net_1341), .B2(net_336) );
OAI22_X2 inst_254 ( .B2(net_2275), .ZN(net_715), .A1(net_714), .A2(net_713), .B1(net_534) );
NAND3_X2 inst_654 ( .A3(net_2167), .A1(net_2003), .A2(net_1667), .ZN(net_1180) );
INV_X2 inst_1673 ( .ZN(net_1864), .A(net_49) );
DFFR_X1 inst_2129 ( .QN(net_2259), .RN(net_1347), .D(net_748), .CK(net_2880) );
INV_X2 inst_1412 ( .A(net_564), .ZN(x1176) );
INV_X1 inst_1708 ( .A(net_2090), .ZN(net_1786) );
INV_X4 inst_1181 ( .A(net_2040), .ZN(net_1507) );
INV_X8 inst_1153 ( .ZN(net_1639), .A(net_1619) );
CLKBUF_X2 inst_3823 ( .A(net_3037), .Z(net_3615) );
OAI21_X2 inst_391 ( .B2(net_2372), .B1(net_1740), .ZN(net_1334), .A(net_1333) );
NAND3_X2 inst_661 ( .A1(net_1763), .A2(net_1662), .ZN(net_1081), .A3(net_810) );
CLKBUF_X2 inst_4107 ( .A(net_3898), .Z(net_3899) );
INV_X2 inst_1548 ( .ZN(net_813), .A(net_68) );
DFFR_X2 inst_2073 ( .QN(net_2418), .D(net_2052), .RN(net_1347), .CK(net_3949) );
CLKBUF_X2 inst_2738 ( .A(net_2529), .Z(net_2530) );
CLKBUF_X2 inst_3984 ( .A(net_3775), .Z(net_3776) );
NAND4_X2 inst_634 ( .A2(net_2050), .ZN(net_1906), .A3(net_1905), .A4(net_1276), .A1(net_522) );
OAI21_X2 inst_419 ( .ZN(net_662), .B2(net_661), .B1(net_606), .A(net_333) );
CLKBUF_X2 inst_3122 ( .A(net_2518), .Z(net_2914) );
INV_X2 inst_1477 ( .A(net_1520), .ZN(net_705) );
CLKBUF_X2 inst_3717 ( .A(net_3508), .Z(net_3509) );
XNOR2_X2 inst_34 ( .B(net_1242), .ZN(net_649), .A(net_597) );
DFF_X2 inst_1799 ( .QN(net_2310), .D(net_278), .CK(net_3956) );
XOR2_X1 inst_12 ( .Z(net_2185), .B(net_1291), .A(net_365) );
NOR2_X4 inst_529 ( .ZN(net_2003), .A1(net_2001), .A2(net_1158) );
INV_X2 inst_1528 ( .ZN(net_262), .A(x6312) );
CLKBUF_X2 inst_3458 ( .A(net_3102), .Z(net_3250) );
INV_X2 inst_1424 ( .A(net_1780), .ZN(net_501) );
INV_X4 inst_1313 ( .ZN(net_1825), .A(net_372) );
INV_X2 inst_1425 ( .ZN(net_497), .A(net_479) );
NAND3_X2 inst_675 ( .A2(net_1792), .ZN(net_919), .A1(net_787), .A3(net_658) );
CLKBUF_X2 inst_4068 ( .A(net_3859), .Z(net_3860) );
CLKBUF_X2 inst_4116 ( .A(net_3135), .Z(net_3908) );
CLKBUF_X2 inst_2886 ( .A(net_2677), .Z(net_2678) );
CLKBUF_X2 inst_2705 ( .A(net_2475), .Z(net_2497) );
AOI22_X2 inst_2307 ( .A2(net_2142), .B1(net_2096), .A1(net_1769), .B2(net_1536), .ZN(net_902) );
OAI22_X2 inst_258 ( .B2(net_2278), .A1(net_740), .ZN(net_706), .A2(net_705), .B1(net_534) );
AND2_X2 inst_2611 ( .A1(net_609), .A2(x6799), .ZN(x603) );
CLKBUF_X2 inst_2773 ( .A(net_2564), .Z(net_2565) );
DFFR_X2 inst_2081 ( .RN(net_1347), .D(net_1144), .QN(net_57), .CK(net_3518) );
CLKBUF_X2 inst_3261 ( .A(net_2899), .Z(net_3053) );
AOI22_X2 inst_2405 ( .B1(net_2197), .ZN(net_1633), .A1(net_1621), .B2(net_1519), .A2(net_934) );
CLKBUF_X2 inst_2994 ( .A(net_2785), .Z(net_2786) );
CLKBUF_X2 inst_3023 ( .A(net_2814), .Z(net_2815) );
INV_X4 inst_1243 ( .A(net_2319), .ZN(net_371) );
CLKBUF_X2 inst_3076 ( .A(net_2621), .Z(net_2868) );
INV_X4 inst_1211 ( .A(net_1614), .ZN(net_1403) );
OAI211_X2 inst_482 ( .C2(net_2315), .C1(net_1052), .ZN(net_1026), .A(net_884), .B(net_859) );
CLKBUF_X2 inst_3751 ( .A(net_2589), .Z(net_3543) );
INV_X4 inst_1192 ( .A(net_913), .ZN(net_759) );
NAND3_X2 inst_682 ( .ZN(net_433), .A2(net_393), .A1(net_360), .A3(net_279) );
CLKBUF_X2 inst_3534 ( .A(net_3325), .Z(net_3326) );
OAI22_X2 inst_238 ( .B2(net_2260), .ZN(net_746), .A1(net_745), .A2(net_744), .B1(net_534) );
CLKBUF_X2 inst_3276 ( .A(net_3047), .Z(net_3068) );
CLKBUF_X2 inst_3996 ( .A(net_2476), .Z(net_3788) );
NAND2_X2 inst_1093 ( .A1(net_2418), .ZN(net_1903), .A2(net_1754) );
NOR2_X2 inst_539 ( .A2(net_2361), .ZN(net_1153), .A1(net_1147) );
AOI22_X2 inst_2222 ( .A2(net_2391), .B2(net_2158), .A1(net_1916), .B1(net_1915), .ZN(net_1458) );
CLKBUF_X2 inst_3333 ( .A(net_3124), .Z(net_3125) );
NAND2_X2 inst_895 ( .A2(net_1709), .A1(net_1708), .ZN(net_1125) );
CLKBUF_X2 inst_4059 ( .A(net_3225), .Z(net_3851) );
CLKBUF_X2 inst_3109 ( .A(net_2900), .Z(net_2901) );
CLKBUF_X2 inst_3271 ( .A(net_2912), .Z(net_3063) );
INV_X2 inst_1430 ( .ZN(net_412), .A(net_402) );
DFF_X2 inst_1755 ( .QN(net_2348), .D(net_1438), .CK(net_3773) );
CLKBUF_X2 inst_3257 ( .A(net_3048), .Z(net_3049) );
AOI22_X2 inst_2240 ( .B2(net_2161), .A1(net_1967), .B1(net_1450), .ZN(net_1390), .A2(net_366) );
INV_X4 inst_1210 ( .ZN(net_1427), .A(net_529) );
AOI22_X2 inst_2341 ( .B1(net_2197), .A1(net_2038), .A2(net_1570), .B2(net_1524), .ZN(net_823) );
AOI22_X2 inst_2437 ( .B2(net_2109), .B1(net_1974), .ZN(net_1811), .A1(net_1789), .A2(net_316) );
NAND2_X2 inst_806 ( .A2(net_1675), .ZN(net_1307), .A1(net_1271) );
CLKBUF_X2 inst_4122 ( .A(net_3380), .Z(net_3914) );
DFF_X1 inst_1981 ( .Q(net_2146), .D(net_1053), .CK(net_3232) );
NAND2_X4 inst_763 ( .ZN(net_2094), .A2(net_2093), .A1(net_2092) );
AOI22_X2 inst_2330 ( .A2(net_2108), .B1(net_2096), .A1(net_1769), .B2(net_1522), .ZN(net_838) );
NOR3_X4 inst_491 ( .A2(net_2020), .ZN(net_2006), .A3(net_2005), .A1(net_2004) );
CLKBUF_X2 inst_3636 ( .A(net_3316), .Z(net_3428) );
CLKBUF_X2 inst_3775 ( .A(net_2523), .Z(net_3567) );
NOR2_X2 inst_537 ( .A2(net_2363), .ZN(net_1172), .A1(net_1162) );
AOI222_X2 inst_2472 ( .C1(net_2016), .A2(net_1551), .A1(net_590), .B1(net_589), .ZN(net_564), .B2(net_153), .C2(x5755) );
NAND2_X2 inst_826 ( .A2(net_2105), .A1(net_1840), .ZN(net_1289) );
CLKBUF_X2 inst_3086 ( .A(net_2877), .Z(net_2878) );
CLKBUF_X2 inst_4002 ( .A(net_3793), .Z(net_3794) );
CLKBUF_X2 inst_2791 ( .A(net_2582), .Z(net_2583) );
OAI22_X2 inst_159 ( .B1(net_1428), .A1(net_1426), .B2(net_184), .A2(net_93), .ZN(x1587) );
NAND2_X2 inst_872 ( .A1(net_1838), .ZN(net_1209), .A2(net_932) );
INV_X2 inst_1667 ( .A(net_1873), .ZN(net_1783) );
INV_X4 inst_1349 ( .A(net_2321), .ZN(net_2105) );
CLKBUF_X2 inst_3950 ( .A(net_3666), .Z(net_3742) );
OAI211_X2 inst_462 ( .C2(net_2331), .ZN(net_1053), .C1(net_1052), .A(net_896), .B(net_851) );
NAND2_X2 inst_869 ( .A1(net_1838), .A2(net_1239), .ZN(net_1212) );
AND2_X2 inst_2646 ( .ZN(net_278), .A1(x3098), .A2(x3067) );
XNOR2_X2 inst_19 ( .B(net_1235), .ZN(net_1177), .A(net_1163) );
CLKBUF_X2 inst_3745 ( .A(net_2757), .Z(net_3537) );
AOI22_X2 inst_2224 ( .B2(net_2151), .A1(net_1960), .ZN(net_1456), .B1(net_1450), .A2(net_1187) );
CLKBUF_X2 inst_3830 ( .A(net_2683), .Z(net_3622) );
CLKBUF_X2 inst_3267 ( .A(net_3058), .Z(net_3059) );
CLKBUF_X2 inst_3205 ( .A(net_2538), .Z(net_2997) );
INV_X16 inst_1686 ( .ZN(net_979), .A(net_556) );
DFF_X1 inst_1914 ( .D(net_1309), .QN(net_140), .CK(net_3644) );
DFF_X1 inst_1975 ( .D(net_1058), .QN(net_43), .CK(net_3107) );
DFF_X1 inst_1890 ( .D(net_1334), .Q(net_144), .CK(net_3009) );
AOI22_X2 inst_2308 ( .A2(net_2143), .B1(net_2096), .A1(net_1769), .B2(net_1535), .ZN(net_901) );
CLKBUF_X2 inst_4093 ( .A(net_2589), .Z(net_3885) );
NOR2_X2 inst_612 ( .A2(net_2255), .ZN(net_1992), .A1(net_520) );
CLKBUF_X2 inst_2879 ( .A(net_2613), .Z(net_2671) );
DFF_X2 inst_1789 ( .QN(net_1588), .D(net_511), .CK(net_3889) );
INV_X16 inst_1692 ( .A(net_1990), .ZN(net_1785) );
CLKBUF_X2 inst_3986 ( .A(net_3430), .Z(net_3778) );
AOI22_X2 inst_2338 ( .B1(net_2197), .A1(net_2038), .A2(net_1571), .B2(net_1523), .ZN(net_826) );
CLKBUF_X2 inst_3475 ( .A(net_3266), .Z(net_3267) );
CLKBUF_X2 inst_3017 ( .A(net_2808), .Z(net_2809) );
CLKBUF_X2 inst_3441 ( .A(net_2765), .Z(net_3233) );
NAND2_X2 inst_845 ( .A1(net_1840), .ZN(net_1268), .A2(net_1259) );
CLKBUF_X2 inst_3554 ( .A(net_3345), .Z(net_3346) );
AOI222_X2 inst_2455 ( .C1(net_2017), .A2(net_1568), .A1(net_590), .B1(net_589), .ZN(net_581), .B2(net_170), .C2(x5370) );
INV_X2 inst_1367 ( .A(net_1017), .ZN(x2562) );
DFF_X1 inst_2016 ( .QN(net_2228), .D(net_1078), .CK(net_3244) );
CLKBUF_X2 inst_3687 ( .A(net_3478), .Z(net_3479) );
AOI22_X2 inst_2287 ( .A1(net_1996), .B1(net_1749), .A2(net_1546), .ZN(net_975), .B2(net_148) );
INV_X2 inst_1460 ( .A(net_2362), .ZN(net_1190) );
INV_X4 inst_1344 ( .ZN(net_2079), .A(net_2078) );
NAND2_X2 inst_885 ( .A2(net_1190), .ZN(net_1162), .A1(net_1153) );
AND2_X2 inst_2630 ( .A1(net_594), .A2(x4266), .ZN(x1713) );
CLKBUF_X2 inst_4012 ( .A(net_2540), .Z(net_3804) );
CLKBUF_X2 inst_3053 ( .A(net_2814), .Z(net_2845) );
INV_X2 inst_1443 ( .A(net_1518), .ZN(net_696) );
NAND2_X2 inst_1028 ( .A2(net_1198), .ZN(net_526), .A1(net_486) );
OAI21_X2 inst_393 ( .A(net_2047), .B1(net_1829), .ZN(net_1134), .B2(net_958) );
CLKBUF_X2 inst_3935 ( .A(net_3726), .Z(net_3727) );
CLKBUF_X2 inst_3610 ( .A(net_3401), .Z(net_3402) );
CLKBUF_X2 inst_2999 ( .A(net_2790), .Z(net_2791) );
DFF_X2 inst_1813 ( .Q(net_1542), .CK(net_2780), .D(x5712) );
SDFF_X2 inst_92 ( .SE(net_487), .Q(net_157), .D(net_157), .CK(net_2546), .SI(x4752) );
OAI21_X2 inst_345 ( .A(net_2083), .B1(net_2082), .B2(net_1484), .ZN(net_1483) );
INV_X4 inst_1271 ( .A(net_2377), .ZN(net_313) );
CLKBUF_X2 inst_3103 ( .A(net_2894), .Z(net_2895) );
AOI22_X2 inst_2321 ( .A2(net_2107), .B1(net_2096), .A1(net_1769), .B2(net_1513), .ZN(net_888) );
CLKBUF_X2 inst_3304 ( .A(net_3095), .Z(net_3096) );
CLKBUF_X2 inst_4156 ( .A(net_3602), .Z(net_3948) );
OAI22_X2 inst_200 ( .A2(net_2231), .A1(net_2013), .B1(net_1407), .B2(net_245), .ZN(x1981) );
SDFF_X2 inst_57 ( .Q(net_1572), .D(net_1572), .SE(net_396), .CK(net_2855), .SI(x6799) );
CLKBUF_X2 inst_3655 ( .A(net_2830), .Z(net_3447) );
DFF_X2 inst_1750 ( .QN(net_2351), .D(net_1415), .CK(net_3777) );
AOI22_X2 inst_2236 ( .B2(net_2125), .A1(net_1967), .B1(net_1450), .ZN(net_1394), .A2(net_1239) );
CLKBUF_X2 inst_3368 ( .A(net_3159), .Z(net_3160) );
INV_X2 inst_1553 ( .ZN(net_247), .A(x6573) );
CLKBUF_X2 inst_2843 ( .A(net_2634), .Z(net_2635) );
DFF_X1 inst_1888 ( .D(net_1844), .QN(net_126), .CK(net_3709) );
CLKBUF_X2 inst_4130 ( .A(net_3921), .Z(net_3922) );
CLKBUF_X2 inst_3379 ( .A(net_3019), .Z(net_3171) );
DFF_X2 inst_1763 ( .D(net_1140), .QN(net_83), .CK(net_4001) );
INV_X2 inst_1635 ( .ZN(net_187), .A(x6503) );
INV_X4 inst_1307 ( .A(net_1743), .ZN(net_1742) );
INV_X2 inst_1500 ( .A(net_2383), .ZN(net_376) );
CLKBUF_X2 inst_2805 ( .A(net_2546), .Z(net_2597) );
NAND2_X2 inst_1094 ( .ZN(net_1909), .A2(net_1904), .A1(net_1903) );
CLKBUF_X2 inst_3499 ( .A(net_3290), .Z(net_3291) );
CLKBUF_X2 inst_4145 ( .A(net_2576), .Z(net_3937) );
CLKBUF_X2 inst_2932 ( .A(net_2660), .Z(net_2724) );
NAND2_X2 inst_893 ( .A2(net_1701), .A1(net_1700), .ZN(net_1127) );
CLKBUF_X2 inst_3680 ( .A(net_2733), .Z(net_3472) );
CLKBUF_X2 inst_3048 ( .A(net_2839), .Z(net_2840) );
INV_X16 inst_1699 ( .ZN(net_1974), .A(net_1973) );
NAND2_X2 inst_851 ( .ZN(net_1249), .A1(net_1193), .A2(net_440) );
NAND2_X2 inst_831 ( .A1(net_1840), .ZN(net_1283), .A2(net_846) );
SDFF_X2 inst_50 ( .SE(net_1768), .SI(net_1529), .Q(net_77), .D(net_77), .CK(net_3204) );
CLKBUF_X2 inst_3346 ( .A(net_3137), .Z(net_3138) );
NOR2_X2 inst_569 ( .A2(net_2333), .A1(net_2330), .ZN(net_342) );
CLKBUF_X2 inst_2992 ( .A(net_2783), .Z(net_2784) );
AND2_X4 inst_2589 ( .A1(net_1953), .ZN(net_1830), .A2(net_552) );
NAND2_X2 inst_1080 ( .A1(net_2104), .ZN(net_1821), .A2(net_1263) );
AOI22_X2 inst_2374 ( .B2(net_2164), .B1(net_1929), .ZN(net_658), .A1(net_655), .A2(net_338) );
NAND2_X2 inst_1103 ( .ZN(net_1987), .A2(net_1982), .A1(net_443) );
INV_X2 inst_1650 ( .ZN(net_295), .A(net_54) );
NOR2_X2 inst_549 ( .A2(net_2378), .A1(net_2196), .ZN(net_607) );
CLKBUF_X2 inst_4220 ( .A(net_3229), .Z(net_4012) );
INV_X2 inst_1497 ( .A(net_2313), .ZN(net_328) );
NOR2_X4 inst_522 ( .A2(net_2416), .A1(net_1872), .ZN(net_431) );
CLKBUF_X2 inst_2872 ( .A(net_2663), .Z(net_2664) );
NAND2_X2 inst_1002 ( .A2(net_2129), .A1(net_979), .ZN(net_671) );
CLKBUF_X2 inst_2809 ( .A(net_2600), .Z(net_2601) );
OAI211_X2 inst_478 ( .C2(net_2312), .C1(net_1052), .ZN(net_1030), .A(net_906), .B(net_878) );
CLKBUF_X2 inst_3380 ( .A(net_3171), .Z(net_3172) );
CLKBUF_X2 inst_2673 ( .A(net_2454), .Z(net_2465) );
INV_X2 inst_1618 ( .ZN(net_199), .A(x6380) );
DFFR_X1 inst_2126 ( .QN(net_2300), .D(net_1610), .RN(net_1347), .CK(net_2802) );
NAND2_X2 inst_804 ( .ZN(net_1309), .A1(net_1290), .A2(net_1226) );
CLKBUF_X2 inst_3290 ( .A(net_2669), .Z(net_3082) );
XOR2_X1 inst_13 ( .Z(net_2188), .B(net_1238), .A(net_659) );
AND2_X4 inst_2584 ( .A1(net_1592), .A2(net_1591), .ZN(net_417) );
CLKBUF_X2 inst_3600 ( .A(net_3391), .Z(net_3392) );
CLKBUF_X2 inst_2765 ( .A(net_2478), .Z(net_2557) );
NAND2_X2 inst_799 ( .A2(net_1679), .ZN(net_1314), .A1(net_1274) );
CLKBUF_X2 inst_3481 ( .A(net_3208), .Z(net_3273) );
OAI22_X2 inst_219 ( .A1(net_1829), .B1(net_1596), .B2(net_1583), .ZN(net_995), .A2(net_938) );
NAND2_X4 inst_738 ( .ZN(net_2194), .A2(net_1933), .A1(net_525) );
NAND2_X4 inst_719 ( .A2(net_2426), .ZN(net_514), .A1(net_479) );
CLKBUF_X2 inst_4166 ( .A(net_3957), .Z(net_3958) );
CLKBUF_X2 inst_2755 ( .A(net_2529), .Z(net_2547) );
DFF_X2 inst_1819 ( .Q(net_1528), .CK(net_2451), .D(x5413) );
CLKBUF_X2 inst_3868 ( .A(net_3659), .Z(net_3660) );
OAI22_X2 inst_255 ( .B2(net_2276), .A1(net_714), .ZN(net_712), .A2(net_711), .B1(net_534) );
CLKBUF_X2 inst_2726 ( .A(net_2517), .Z(net_2518) );
OAI211_X2 inst_453 ( .C1(net_1639), .ZN(net_1101), .A(net_826), .B(net_668), .C2(net_359) );
INV_X8 inst_1134 ( .ZN(net_1054), .A(net_962) );
NOR3_X2 inst_493 ( .A1(net_2432), .A2(net_2335), .A3(net_2332), .ZN(net_1142) );
CLKBUF_X2 inst_2674 ( .A(net_2465), .Z(net_2466) );
AOI22_X2 inst_2204 ( .A2(net_2398), .B2(net_2143), .A1(net_1960), .ZN(net_1477), .B1(net_1450) );
XNOR2_X2 inst_23 ( .B(net_2329), .ZN(net_1160), .A(net_1145) );
NAND2_X2 inst_1113 ( .ZN(net_2050), .A1(net_2049), .A2(net_383) );
DFF_X2 inst_1822 ( .Q(net_1536), .CK(net_2497), .D(x5556) );
INV_X2 inst_1609 ( .ZN(net_205), .A(x6456) );
CLKBUF_X2 inst_4105 ( .A(net_3896), .Z(net_3897) );
CLKBUF_X2 inst_3790 ( .A(net_3581), .Z(net_3582) );
CLKBUF_X2 inst_4206 ( .A(net_3997), .Z(net_3998) );
CLKBUF_X2 inst_3546 ( .A(net_3337), .Z(net_3338) );
OAI21_X2 inst_408 ( .B2(net_2029), .ZN(net_767), .B1(net_766), .A(net_531) );
INV_X8 inst_1144 ( .A(net_2019), .ZN(net_590) );
NAND2_X2 inst_812 ( .A2(net_1676), .ZN(net_1301), .A1(net_1279) );
AOI211_X2 inst_2568 ( .C2(net_2125), .ZN(net_2098), .C1(net_1929), .A(net_1894), .B(net_1785) );
AOI22_X2 inst_2295 ( .B2(net_1567), .A2(net_1276), .A1(net_962), .B1(net_961), .ZN(net_960) );
OAI22_X2 inst_179 ( .B1(net_1428), .A1(net_529), .B2(net_209), .A2(net_98), .ZN(x1520) );
DFF_X2 inst_1730 ( .QN(net_2314), .D(net_1501), .CK(net_3353) );
CLKBUF_X2 inst_3799 ( .A(net_3590), .Z(net_3591) );
CLKBUF_X2 inst_3814 ( .A(net_3127), .Z(net_3606) );
CLKBUF_X2 inst_3734 ( .A(net_3525), .Z(net_3526) );
CLKBUF_X2 inst_3532 ( .A(net_3323), .Z(net_3324) );
CLKBUF_X2 inst_3028 ( .A(net_2819), .Z(net_2820) );
SDFF_X2 inst_76 ( .Q(net_1566), .D(net_1566), .SE(net_491), .CK(net_2623), .SI(x7007) );
CLKBUF_X2 inst_3854 ( .A(net_3069), .Z(net_3646) );
NAND2_X1 inst_1127 ( .A2(net_2440), .A1(net_1404), .ZN(x44) );
CLKBUF_X2 inst_3514 ( .A(net_3305), .Z(net_3306) );
OAI22_X2 inst_172 ( .B1(net_1427), .A1(net_529), .B2(net_265), .A2(net_110), .ZN(x1379) );
OAI21_X2 inst_362 ( .B2(net_2410), .B1(net_1441), .ZN(net_1432), .A(net_1390) );
INV_X2 inst_1530 ( .ZN(net_301), .A(net_70) );
OAI22_X2 inst_277 ( .B2(net_2301), .B1(net_1865), .ZN(net_1609), .A1(net_951), .A2(net_724) );
INV_X2 inst_1510 ( .A(net_2418), .ZN(net_358) );
SDFF_X2 inst_83 ( .SE(net_487), .Q(net_154), .D(net_154), .CK(net_2550), .SI(x4843) );
SDFFR_X1 inst_121 ( .SE(net_1829), .D(net_1538), .RN(net_1347), .SI(net_49), .Q(net_49), .CK(net_2863) );
OAI22_X2 inst_306 ( .A2(net_2225), .B1(net_1895), .A1(net_1408), .B2(net_254), .ZN(x2119) );
CLKBUF_X2 inst_4186 ( .A(net_3629), .Z(net_3978) );
NAND2_X2 inst_1065 ( .A2(net_2073), .ZN(net_1731), .A1(net_931) );
CLKBUF_X2 inst_4119 ( .A(net_3910), .Z(net_3911) );
CLKBUF_X2 inst_3386 ( .A(net_2606), .Z(net_3178) );
CLKBUF_X2 inst_3095 ( .A(net_2886), .Z(net_2887) );
HA_X1 inst_1715 ( .B(net_1260), .S(net_474), .CO(net_473), .A(net_394) );
OR2_X2 inst_140 ( .ZN(net_426), .A2(x6264), .A1(x6236) );
OAI22_X2 inst_267 ( .B2(net_2283), .B1(net_1865), .ZN(net_1598), .A1(net_951), .A2(net_696) );
CLKBUF_X2 inst_2824 ( .A(net_2615), .Z(net_2616) );
NAND2_X4 inst_716 ( .A1(net_1918), .ZN(net_621), .A2(net_413) );
CLKBUF_X2 inst_3594 ( .A(net_3385), .Z(net_3386) );
CLKBUF_X2 inst_4174 ( .A(net_3684), .Z(net_3966) );
DFF_X1 inst_1906 ( .D(net_1305), .QN(net_116), .CK(net_3566) );
NOR2_X4 inst_530 ( .ZN(net_2035), .A1(net_2033), .A2(net_1977) );
NAND2_X2 inst_792 ( .A1(net_1823), .ZN(net_1321), .A2(net_1202) );
DFF_X1 inst_2024 ( .QN(net_2235), .D(net_2058), .CK(net_3218) );
CLKBUF_X2 inst_3124 ( .A(net_2915), .Z(net_2916) );
CLKBUF_X2 inst_2952 ( .A(net_2509), .Z(net_2744) );
INV_X32 inst_1353 ( .A(net_1840), .ZN(net_1741) );
AOI221_X2 inst_2502 ( .B2(net_2130), .B1(net_1929), .A(net_1890), .C1(net_1863), .ZN(net_969), .C2(net_307) );
AOI22_X2 inst_2216 ( .A2(net_2387), .B2(net_2155), .A1(net_1960), .B1(net_1915), .ZN(net_1464) );
NAND2_X2 inst_769 ( .ZN(net_1486), .A2(net_1447), .A1(net_1370) );
OAI22_X2 inst_174 ( .B1(net_1428), .A1(net_1426), .B2(net_236), .A2(net_103), .ZN(x1451) );
INV_X4 inst_1200 ( .ZN(net_554), .A(net_553) );
CLKBUF_X2 inst_2988 ( .A(net_2779), .Z(net_2780) );
DFFR_X1 inst_2105 ( .QN(net_2295), .RN(net_1347), .D(net_955), .CK(net_2566) );
INV_X4 inst_1199 ( .ZN(net_768), .A(net_630) );
XOR2_X1 inst_5 ( .Z(net_2178), .A(net_1161), .B(net_285) );
CLKBUF_X2 inst_3974 ( .A(net_3214), .Z(net_3766) );
CLKBUF_X2 inst_3021 ( .A(net_2812), .Z(net_2813) );
NAND2_X4 inst_729 ( .A2(net_1984), .ZN(net_1827), .A1(net_1826) );
DFFR_X1 inst_2157 ( .QN(net_2260), .RN(net_1347), .D(net_746), .CK(net_2872) );
INV_X2 inst_1662 ( .A(net_1753), .ZN(net_1752) );
CLKBUF_X2 inst_2783 ( .A(net_2574), .Z(net_2575) );
OAI22_X2 inst_213 ( .A2(net_2210), .B1(net_1407), .A1(net_1405), .B2(net_202), .ZN(x2403) );
NOR2_X2 inst_604 ( .A2(net_2260), .ZN(net_1894), .A1(net_520) );
OAI22_X2 inst_205 ( .A2(net_2226), .B1(net_1614), .A1(net_1405), .B2(net_215), .ZN(x2098) );
INV_X2 inst_1645 ( .A(net_2248), .ZN(net_182) );
INV_X4 inst_1285 ( .A(net_2347), .ZN(net_1291) );
OAI21_X2 inst_380 ( .A(net_1942), .ZN(net_1357), .B2(net_1356), .B1(net_1341) );
CLKBUF_X2 inst_4057 ( .A(net_3848), .Z(net_3849) );
INV_X4 inst_1179 ( .A(net_1916), .ZN(net_1484) );
CLKBUF_X2 inst_3722 ( .A(net_3513), .Z(net_3514) );
OAI22_X2 inst_292 ( .A1(net_1615), .B1(net_1407), .B2(net_199), .A2(net_129), .ZN(x381) );
CLKBUF_X2 inst_3650 ( .A(net_2456), .Z(net_3442) );
DFF_X1 inst_2012 ( .QN(net_2216), .D(net_1071), .CK(net_3291) );
CLKBUF_X2 inst_3911 ( .A(net_3702), .Z(net_3703) );
INV_X2 inst_1515 ( .A(net_2299), .ZN(net_320) );
NAND3_X2 inst_706 ( .A2(net_2206), .A3(net_2203), .ZN(net_2086), .A1(net_2085) );
DFF_X2 inst_1782 ( .QN(net_2425), .D(net_752), .CK(net_3664) );
CLKBUF_X2 inst_2951 ( .A(net_2670), .Z(net_2743) );
CLKBUF_X2 inst_3890 ( .A(net_3681), .Z(net_3682) );
NAND2_X2 inst_839 ( .A1(net_1840), .ZN(net_1274), .A2(net_1262) );
NAND2_X2 inst_1015 ( .A2(net_2114), .ZN(net_616), .A1(net_536) );
OAI22_X2 inst_240 ( .B2(net_2262), .ZN(net_741), .A1(net_740), .A2(net_739), .B1(net_534) );
CLKBUF_X2 inst_3966 ( .A(net_2486), .Z(net_3758) );
SDFF_X2 inst_110 ( .SE(net_487), .Q(net_145), .D(net_145), .CK(net_3018), .SI(x5078) );
CLKBUF_X2 inst_3899 ( .A(net_3495), .Z(net_3691) );
DFF_X1 inst_2047 ( .QN(net_2401), .D(net_551), .CK(net_3787) );
CLKBUF_X2 inst_3213 ( .A(net_2718), .Z(net_3005) );
CLKBUF_X2 inst_3825 ( .A(net_3438), .Z(net_3617) );
AOI21_X2 inst_2535 ( .A(net_1785), .B1(net_910), .ZN(net_797), .B2(net_796) );
SDFF_X2 inst_99 ( .SE(net_488), .Q(net_176), .D(net_176), .CK(net_2950), .SI(x4303) );
INV_X2 inst_1661 ( .A(net_1748), .ZN(net_1747) );
DFF_X1 inst_2059 ( .QN(net_2399), .D(net_465), .CK(net_3782) );
CLKBUF_X2 inst_2949 ( .A(net_2740), .Z(net_2741) );
AOI22_X2 inst_2414 ( .A2(net_2153), .B2(net_2115), .A1(net_1974), .B1(net_1929), .ZN(net_1660) );
OAI22_X2 inst_283 ( .A2(net_2236), .A1(net_1615), .B1(net_1407), .B2(net_224), .ZN(x1877) );
OAI22_X2 inst_311 ( .B1(net_1895), .A1(net_1405), .B2(net_186), .A2(net_115), .ZN(x542) );
CLKBUF_X2 inst_3406 ( .A(net_3197), .Z(net_3198) );
AOI21_X2 inst_2519 ( .A(net_2044), .B1(net_1739), .ZN(net_1362), .B2(net_282) );
INV_X2 inst_1597 ( .ZN(net_213), .A(x4033) );
CLKBUF_X2 inst_3502 ( .A(net_3293), .Z(net_3294) );
AOI22_X2 inst_2203 ( .A2(net_2177), .B2(net_2147), .A1(net_1960), .B1(net_1915), .ZN(net_1478) );
CLKBUF_X2 inst_3473 ( .A(net_3264), .Z(net_3265) );
OAI21_X2 inst_431 ( .B1(net_2416), .ZN(net_1719), .B2(net_1581), .A(net_1579) );
OAI21_X2 inst_348 ( .B1(net_2080), .B2(net_1484), .ZN(net_1480), .A(net_1449) );
DFF_X1 inst_1930 ( .D(net_1124), .QN(net_69), .CK(net_3475) );
NAND2_X2 inst_889 ( .ZN(net_1131), .A1(net_1002), .A2(net_911) );
NOR2_X2 inst_577 ( .A2(net_2412), .A1(net_1746), .ZN(net_1682) );
CLKBUF_X2 inst_2686 ( .A(net_2456), .Z(net_2478) );
CLKBUF_X2 inst_3740 ( .A(net_3531), .Z(net_3532) );
AOI22_X2 inst_2293 ( .A1(net_1996), .B1(net_1749), .A2(net_1549), .ZN(net_964), .B2(net_151) );
AOI22_X2 inst_2379 ( .A1(net_1718), .B1(net_1474), .B2(net_796), .ZN(net_647), .A2(net_646) );
INV_X2 inst_1364 ( .A(net_1021), .ZN(x2513) );
CLKBUF_X2 inst_3938 ( .A(net_3729), .Z(net_3730) );
CLKBUF_X2 inst_2865 ( .A(net_2656), .Z(net_2657) );
NAND3_X4 inst_645 ( .ZN(net_1159), .A2(net_1142), .A1(net_416), .A3(net_342) );
CLKBUF_X2 inst_3571 ( .A(net_3362), .Z(net_3363) );
CLKBUF_X2 inst_3041 ( .A(net_2755), .Z(net_2833) );
CLKBUF_X2 inst_2719 ( .A(net_2510), .Z(net_2511) );
AOI22_X2 inst_2352 ( .A1(net_783), .B1(net_782), .ZN(net_780), .A2(net_355), .B2(x3684) );
OAI22_X2 inst_269 ( .B2(net_2298), .B1(net_1865), .ZN(net_1600), .A1(net_951), .A2(net_949) );
INV_X4 inst_1190 ( .ZN(net_1168), .A(net_931) );
OAI21_X1 inst_444 ( .B2(net_1752), .B1(net_1250), .ZN(net_1247), .A(net_437) );
AOI21_X2 inst_2544 ( .B2(net_1933), .A(net_839), .ZN(net_661), .B1(net_550) );
NOR2_X4 inst_514 ( .A2(net_1595), .A1(net_1594), .ZN(net_507) );
INV_X2 inst_1541 ( .ZN(net_255), .A(x4148) );
CLKBUF_X2 inst_4236 ( .A(net_4027), .Z(net_4028) );
NAND3_X2 inst_685 ( .A1(net_2443), .ZN(net_462), .A3(x3865), .A2(x3843) );
SDFF_X2 inst_63 ( .Q(net_1552), .D(net_1552), .SE(net_396), .CK(net_2688), .SI(x7345) );
SDFF_X2 inst_119 ( .Q(net_1560), .D(net_1560), .SE(net_491), .CK(net_2892), .SI(x7169) );
CLKBUF_X2 inst_3181 ( .A(net_2972), .Z(net_2973) );
NAND2_X2 inst_939 ( .A2(net_1623), .ZN(net_1061), .A1(net_686) );
INV_X4 inst_1233 ( .ZN(net_400), .A(net_285) );
CLKBUF_X2 inst_2924 ( .A(x7552), .Z(net_2716) );
CLKBUF_X2 inst_3432 ( .A(net_3223), .Z(net_3224) );
NAND2_X2 inst_1019 ( .A2(net_2415), .ZN(net_612), .A1(net_552) );
DFF_X1 inst_2006 ( .QN(net_2227), .D(net_1079), .CK(net_3295) );
DFF_X2 inst_1827 ( .Q(net_1540), .CK(net_2590), .D(x5657) );
NAND2_X4 inst_742 ( .A1(net_2192), .ZN(net_1957), .A2(net_1945) );
OAI21_X2 inst_427 ( .ZN(net_408), .B1(net_407), .B2(x6264), .A(x5995) );
CLKBUF_X2 inst_3840 ( .A(net_3631), .Z(net_3632) );
AND2_X2 inst_2619 ( .A1(net_594), .A2(x7190), .ZN(x760) );
CLKBUF_X2 inst_3465 ( .A(net_3256), .Z(net_3257) );
DFF_X1 inst_2033 ( .QN(net_2237), .D(net_837), .CK(net_2984) );
DFFR_X1 inst_2144 ( .QN(net_2250), .RN(net_1347), .D(net_708), .CK(net_2876) );
AOI21_X1 inst_2559 ( .ZN(net_518), .A(net_502), .B1(net_492), .B2(net_374) );
OR2_X2 inst_138 ( .A2(net_2371), .A1(net_2370), .ZN(net_420) );
DFF_X1 inst_1955 ( .Q(net_2121), .D(net_1089), .CK(net_3467) );
CLKBUF_X2 inst_2810 ( .A(net_2601), .Z(net_2602) );
CLKBUF_X2 inst_3618 ( .A(net_3409), .Z(net_3410) );
INV_X4 inst_1269 ( .A(net_2419), .ZN(net_318) );
NAND2_X2 inst_899 ( .A2(net_1689), .A1(net_1688), .ZN(net_1120) );
OAI22_X2 inst_312 ( .B2(net_2293), .ZN(net_1972), .A1(net_1864), .A2(net_1851), .B1(net_1848) );
CLKBUF_X2 inst_3241 ( .A(net_2691), .Z(net_3033) );
CLKBUF_X2 inst_2704 ( .A(net_2495), .Z(net_2496) );
INV_X2 inst_1620 ( .ZN(net_388), .A(x3947) );
OAI22_X2 inst_309 ( .B1(net_1895), .A1(net_1408), .B2(net_240), .A2(net_138), .ZN(x192) );
CLKBUF_X2 inst_3416 ( .A(net_3207), .Z(net_3208) );
OAI21_X2 inst_347 ( .ZN(net_1481), .B1(net_1424), .A(net_1396), .B2(net_395) );
DFFR_X1 inst_2149 ( .QN(net_2256), .RN(net_1347), .D(net_699), .CK(net_3384) );
NAND2_X4 inst_755 ( .A2(net_2209), .ZN(net_2011), .A1(net_2008) );
DFF_X2 inst_1724 ( .QN(net_2328), .D(net_1488), .CK(net_2959) );
AND2_X2 inst_2610 ( .A1(net_594), .A2(x6727), .ZN(x582) );
CLKBUF_X2 inst_2694 ( .A(net_2485), .Z(net_2486) );
NAND2_X2 inst_1043 ( .A1(net_1841), .ZN(net_1670), .A2(net_934) );
CLKBUF_X2 inst_4030 ( .A(net_3130), .Z(net_3822) );
DFF_X1 inst_1968 ( .Q(net_2134), .D(net_1090), .CK(net_3190) );
CLKBUF_X2 inst_4078 ( .A(net_3869), .Z(net_3870) );
CLKBUF_X2 inst_4067 ( .A(net_3858), .Z(net_3859) );
DFF_X2 inst_1792 ( .QN(net_2439), .D(net_490), .CK(net_2784) );
INV_X4 inst_1330 ( .ZN(net_1996), .A(net_1994) );
CLKBUF_X2 inst_3928 ( .A(net_2573), .Z(net_3720) );
CLKBUF_X2 inst_3353 ( .A(net_3144), .Z(net_3145) );
DFF_X1 inst_1898 ( .D(net_1310), .QN(net_138), .CK(net_3447) );
CLKBUF_X2 inst_3634 ( .A(net_3425), .Z(net_3426) );
CLKBUF_X2 inst_3883 ( .A(net_3674), .Z(net_3675) );
CLKBUF_X2 inst_4017 ( .A(net_3808), .Z(net_3809) );
HA_X1 inst_1714 ( .B(net_1203), .S(net_504), .CO(net_503), .A(net_435) );
INV_X2 inst_1496 ( .A(net_2336), .ZN(net_363) );
INV_X2 inst_1565 ( .ZN(net_235), .A(x4138) );
NAND2_X2 inst_924 ( .A2(net_1629), .ZN(net_1090), .A1(net_828) );
OAI22_X2 inst_287 ( .A1(net_1615), .B1(net_1406), .B2(net_214), .A2(net_119), .ZN(x510) );
OAI21_X2 inst_426 ( .ZN(net_425), .B1(net_407), .B2(x6236), .A(x5995) );
CLKBUF_X2 inst_3145 ( .A(net_2550), .Z(net_2937) );
AND2_X4 inst_2577 ( .A2(net_2415), .A1(net_1976), .ZN(net_543) );
NAND3_X2 inst_648 ( .ZN(net_1455), .A1(net_1401), .A2(net_1369), .A3(net_616) );
CLKBUF_X2 inst_3094 ( .A(net_2885), .Z(net_2886) );
CLKBUF_X2 inst_2903 ( .A(net_2694), .Z(net_2695) );
OAI22_X2 inst_270 ( .B2(net_2293), .B1(net_1865), .ZN(net_1601), .A1(net_1597), .A2(net_739) );
CLKBUF_X2 inst_4045 ( .A(net_3836), .Z(net_3837) );
DFF_X1 inst_1901 ( .D(net_1302), .QN(net_121), .CK(net_3578) );
NAND2_X2 inst_984 ( .A2(net_1553), .A1(net_961), .ZN(net_855) );
CLKBUF_X2 inst_3804 ( .A(net_3595), .Z(net_3596) );
DFF_X1 inst_2064 ( .Q(net_2344), .D(net_392), .CK(net_3141) );
CLKBUF_X2 inst_4104 ( .A(net_3737), .Z(net_3896) );
AOI22_X2 inst_2266 ( .B1(net_1768), .ZN(net_1692), .B2(net_1532), .A1(net_1001), .A2(net_660) );
INV_X4 inst_1292 ( .ZN(net_796), .A(net_62) );
AOI21_X2 inst_2552 ( .B1(net_1924), .ZN(net_1727), .A(net_1726), .B2(net_303) );
DFF_X1 inst_1963 ( .Q(net_2129), .D(net_1093), .CK(net_3639) );
NAND4_X2 inst_631 ( .A3(net_2167), .A1(net_1978), .ZN(net_521), .A2(net_489), .A4(net_448) );
NAND2_X2 inst_1056 ( .ZN(net_1686), .A1(net_1685), .A2(net_399) );
CLKBUF_X2 inst_3648 ( .A(net_3439), .Z(net_3440) );
CLKBUF_X2 inst_3674 ( .A(net_3465), .Z(net_3466) );
AOI221_X2 inst_2514 ( .B2(net_2161), .ZN(net_1986), .A(net_1985), .B1(net_1929), .C1(net_1863), .C2(net_51) );
CLKBUF_X2 inst_3995 ( .A(net_3786), .Z(net_3787) );
NAND2_X1 inst_1128 ( .ZN(net_2048), .A2(net_2045), .A1(net_760) );
CLKBUF_X2 inst_4211 ( .A(net_4002), .Z(net_4003) );
CLKBUF_X2 inst_3759 ( .A(net_3550), .Z(net_3551) );
CLKBUF_X2 inst_3222 ( .A(net_2843), .Z(net_3014) );
DFF_X2 inst_1745 ( .QN(net_2361), .D(net_1420), .CK(net_3588) );
CLKBUF_X2 inst_3831 ( .A(net_3622), .Z(net_3623) );
DFFR_X2 inst_2079 ( .QN(net_1577), .RN(net_1347), .D(net_1165), .CK(net_3730) );
SDFF_X2 inst_102 ( .SE(net_487), .Q(net_169), .D(net_169), .CK(net_2736), .SI(x4435) );
AOI21_X2 inst_2527 ( .A(net_1785), .B1(net_910), .ZN(net_806), .B2(net_74) );
CLKBUF_X2 inst_3277 ( .A(net_3068), .Z(net_3069) );
CLKBUF_X2 inst_4070 ( .A(net_3383), .Z(net_3862) );
CLKBUF_X2 inst_2786 ( .A(net_2548), .Z(net_2578) );
INV_X4 inst_1224 ( .ZN(net_1656), .A(net_443) );
CLKBUF_X2 inst_3905 ( .A(net_2702), .Z(net_3697) );
DFF_X1 inst_1924 ( .Q(net_2435), .D(net_1726), .CK(net_3924) );
INV_X8 inst_1170 ( .ZN(net_1995), .A(net_1994) );
AND2_X4 inst_2596 ( .A1(net_2413), .ZN(net_2170), .A2(net_1582) );
CLKBUF_X2 inst_3022 ( .A(net_2491), .Z(net_2814) );
NAND3_X2 inst_680 ( .A2(net_2170), .ZN(net_484), .A3(net_448), .A1(net_384) );
NAND2_X2 inst_785 ( .A1(net_1813), .ZN(net_1328), .A2(net_1200) );
AOI22_X2 inst_2362 ( .B2(net_2115), .A1(net_2038), .A2(net_1574), .B1(net_979), .ZN(net_695) );
CLKBUF_X2 inst_3299 ( .A(net_3090), .Z(net_3091) );
CLKBUF_X2 inst_4160 ( .A(net_3951), .Z(net_3952) );
CLKBUF_X2 inst_3255 ( .A(net_3046), .Z(net_3047) );
CLKBUF_X2 inst_2856 ( .A(net_2518), .Z(net_2648) );
NAND2_X2 inst_961 ( .A2(net_933), .ZN(net_915), .A1(net_913) );
INV_X2 inst_1590 ( .ZN(net_219), .A(x3997) );
AOI22_X2 inst_2318 ( .B2(net_2242), .A2(net_2153), .B1(net_2096), .A1(net_1769), .ZN(net_891) );
OAI21_X2 inst_399 ( .B1(net_1829), .ZN(net_1108), .B2(net_936), .A(net_925) );
NOR2_X4 inst_527 ( .ZN(net_1865), .A1(net_1848), .A2(net_372) );
CLKBUF_X2 inst_3957 ( .A(net_3748), .Z(net_3749) );
CLKBUF_X2 inst_3567 ( .A(net_2700), .Z(net_3359) );
OAI22_X2 inst_226 ( .B2(net_2299), .B1(net_1865), .A1(net_1597), .ZN(net_948), .A2(net_728) );
INV_X4 inst_1180 ( .ZN(net_1424), .A(net_1423) );
CLKBUF_X2 inst_4020 ( .A(net_3286), .Z(net_3812) );
OAI21_X2 inst_414 ( .B1(net_2196), .ZN(net_755), .A(net_624), .B2(net_518) );
NOR2_X4 inst_531 ( .A2(net_2415), .ZN(net_2049), .A1(net_500) );
CLKBUF_X2 inst_2737 ( .A(net_2528), .Z(net_2529) );
AOI22_X2 inst_2316 ( .A2(net_2148), .B1(net_2096), .A1(net_1769), .B2(net_1527), .ZN(net_893) );
OAI22_X2 inst_212 ( .A2(net_2214), .B1(net_1407), .A1(net_1405), .B2(net_223), .ZN(x2318) );
CLKBUF_X2 inst_2732 ( .A(net_2464), .Z(net_2524) );
INV_X4 inst_1299 ( .ZN(net_788), .A(net_66) );
NOR3_X2 inst_499 ( .A2(net_2318), .A1(net_2317), .A3(net_2314), .ZN(net_360) );
DFF_X1 inst_1952 ( .Q(net_2118), .D(net_1096), .CK(net_3565) );
NAND3_X2 inst_674 ( .ZN(net_923), .A2(net_682), .A1(net_641), .A3(net_548) );
AOI22_X2 inst_2400 ( .B1(net_2197), .ZN(net_1628), .A1(net_1621), .B2(net_1525), .A2(net_1227) );
INV_X2 inst_1451 ( .A(net_2349), .ZN(net_1203) );
CLKBUF_X2 inst_4082 ( .A(net_3873), .Z(net_3874) );
CLKBUF_X2 inst_3698 ( .A(net_3489), .Z(net_3490) );
AOI22_X2 inst_2253 ( .B2(net_2117), .A1(net_1967), .B1(net_1474), .ZN(net_1377), .A2(net_1205) );
CLKBUF_X2 inst_4155 ( .A(net_3946), .Z(net_3947) );
CLKBUF_X2 inst_2966 ( .A(net_2757), .Z(net_2758) );
DFF_X1 inst_2009 ( .QN(net_2221), .D(net_1082), .CK(net_3486) );
CLKBUF_X2 inst_3246 ( .A(net_3037), .Z(net_3038) );
CLKBUF_X2 inst_2868 ( .A(net_2659), .Z(net_2660) );
NOR3_X1 inst_501 ( .ZN(net_456), .A1(net_455), .A3(net_454), .A2(net_451) );
DFFR_X2 inst_2093 ( .QN(net_2202), .RN(net_1347), .D(net_652), .CK(net_3543) );
NAND2_X2 inst_1081 ( .A1(net_2104), .ZN(net_1822), .A2(net_1265) );
CLKBUF_X2 inst_3195 ( .A(net_2986), .Z(net_2987) );
AOI22_X2 inst_2381 ( .A1(net_1718), .B1(net_1450), .B2(net_792), .ZN(net_644), .A2(net_355) );
CLKBUF_X2 inst_2905 ( .A(net_2696), .Z(net_2697) );
DFF_X2 inst_1832 ( .Q(net_2242), .CK(net_2955), .D(x5224) );
NOR2_X2 inst_570 ( .A2(net_2313), .A1(net_2312), .ZN(net_393) );
CLKBUF_X2 inst_2819 ( .A(net_2610), .Z(net_2611) );
INV_X2 inst_1570 ( .ZN(net_232), .A(x4323) );
NAND4_X2 inst_640 ( .ZN(net_1939), .A3(net_1914), .A2(net_1835), .A1(net_1760), .A4(net_1735) );
INV_X2 inst_1612 ( .A(net_2307), .ZN(net_299) );
INV_X2 inst_1478 ( .A(net_1540), .ZN(net_744) );
NAND2_X2 inst_1114 ( .ZN(net_2054), .A2(net_1948), .A1(net_517) );
OAI211_X2 inst_454 ( .C2(net_2370), .C1(net_1639), .ZN(net_1100), .A(net_822), .B(net_663) );
CLKBUF_X2 inst_4163 ( .A(net_2920), .Z(net_3955) );
DFF_X1 inst_1982 ( .Q(net_2147), .D(net_1040), .CK(net_2996) );
DFFR_X2 inst_2089 ( .QN(net_1585), .RN(net_1347), .D(net_1110), .CK(net_3546) );
CLKBUF_X2 inst_3718 ( .A(net_3509), .Z(net_3510) );
DFF_X1 inst_1849 ( .QN(net_2372), .D(net_1453), .CK(net_3404) );
INV_X2 inst_1679 ( .ZN(net_1968), .A(net_514) );
DFF_X1 inst_1976 ( .Q(net_2141), .D(net_1055), .CK(net_3067) );
CLKBUF_X2 inst_3681 ( .A(net_3472), .Z(net_3473) );
CLKBUF_X2 inst_2744 ( .A(net_2535), .Z(net_2536) );
AOI22_X2 inst_2215 ( .A2(net_2342), .B2(net_2154), .A1(net_1960), .B1(net_1915), .ZN(net_1465) );
CLKBUF_X2 inst_3077 ( .A(net_2868), .Z(net_2869) );
DFF_X1 inst_1855 ( .QN(net_2357), .D(net_1429), .CK(net_3722) );
OAI21_X2 inst_337 ( .B2(net_2331), .B1(net_2041), .ZN(net_1493), .A(net_1459) );
AOI22_X2 inst_2384 ( .A1(net_2195), .B1(net_839), .ZN(net_637), .A2(net_422), .B2(net_73) );
INV_X4 inst_1212 ( .ZN(net_1428), .A(net_609) );
NAND3_X2 inst_670 ( .A2(net_1811), .ZN(net_1072), .A1(net_965), .A3(net_795) );
INV_X2 inst_1423 ( .A(net_510), .ZN(net_502) );
CLKBUF_X2 inst_4180 ( .A(net_3971), .Z(net_3972) );
AOI22_X2 inst_2419 ( .B2(net_2157), .B1(net_1974), .ZN(net_1793), .A1(net_1791), .A2(net_319) );
NAND2_X2 inst_1034 ( .A1(net_2208), .A2(net_2207), .ZN(net_418) );
INV_X4 inst_1207 ( .A(net_1614), .ZN(net_1405) );
CLKBUF_X2 inst_3901 ( .A(net_3692), .Z(net_3693) );
NOR2_X2 inst_613 ( .ZN(net_2004), .A2(net_484), .A1(net_481) );
AOI22_X2 inst_2396 ( .B1(net_2197), .ZN(net_1624), .A1(net_1621), .B2(net_1521), .A2(net_1199) );
INV_X2 inst_1428 ( .A(net_2310), .ZN(net_423) );
OAI211_X2 inst_483 ( .C2(net_2317), .C1(net_1052), .ZN(net_1025), .A(net_875), .B(net_854) );
CLKBUF_X2 inst_2739 ( .A(net_2530), .Z(net_2531) );
OAI22_X2 inst_259 ( .B2(net_2251), .A1(net_740), .ZN(net_704), .A2(net_703), .B1(net_534) );
NAND2_X2 inst_1046 ( .A1(net_1743), .ZN(net_1673), .A2(net_1218) );
OAI22_X2 inst_246 ( .B2(net_2249), .ZN(net_731), .A2(net_730), .A1(net_714), .B1(net_534) );
NAND4_X2 inst_635 ( .A2(net_2050), .ZN(net_1907), .A3(net_1905), .A1(net_522), .A4(net_330) );
NAND2_X2 inst_807 ( .A2(net_1674), .ZN(net_1306), .A1(net_1285) );
NAND3_X2 inst_705 ( .ZN(net_2061), .A1(net_2060), .A3(net_1920), .A2(net_802) );
NAND2_X2 inst_911 ( .A1(net_980), .A2(net_785), .ZN(x2869) );
NOR2_X4 inst_519 ( .ZN(net_447), .A1(net_402), .A2(net_333) );
CLKBUF_X2 inst_3796 ( .A(net_3587), .Z(net_3588) );
NAND2_X2 inst_909 ( .A1(net_922), .A2(net_773), .ZN(x2791) );
NAND2_X2 inst_1003 ( .A2(net_2133), .A1(net_979), .ZN(net_669) );
AOI222_X1 inst_2484 ( .B1(net_1995), .A1(net_1751), .B2(net_1566), .C1(net_1020), .ZN(net_1016), .A2(net_168), .C2(x3365) );
NAND2_X2 inst_1053 ( .A1(net_1746), .ZN(net_1680), .A2(net_1239) );
CLKBUF_X2 inst_2919 ( .A(net_2710), .Z(net_2711) );
NAND2_X2 inst_894 ( .A2(net_1705), .A1(net_1704), .ZN(net_1126) );
AOI22_X2 inst_2425 ( .B2(net_2110), .B1(net_1974), .ZN(net_1799), .A1(net_1791), .A2(net_283) );
DFF_X1 inst_1872 ( .D(net_2069), .QN(net_100), .CK(net_3878) );
CLKBUF_X2 inst_3469 ( .A(net_3260), .Z(net_3261) );
NAND2_X2 inst_994 ( .A1(net_1798), .ZN(net_837), .A2(net_677) );
CLKBUF_X2 inst_2774 ( .A(net_2565), .Z(net_2566) );
OAI22_X2 inst_239 ( .B2(net_2261), .ZN(net_743), .A2(net_742), .A1(net_740), .B1(net_534) );
CLKBUF_X2 inst_4028 ( .A(net_3819), .Z(net_3820) );
DFFR_X2 inst_2080 ( .RN(net_1347), .D(net_1164), .QN(net_55), .CK(net_3078) );
DFF_X1 inst_1879 ( .D(net_1325), .QN(net_103), .CK(net_3828) );
INV_X4 inst_1193 ( .A(net_1766), .ZN(net_1000) );
INV_X2 inst_1625 ( .A(net_2295), .ZN(net_290) );
DFF_X1 inst_1863 ( .D(net_1353), .QN(net_106), .CK(net_3839) );
NOR2_X2 inst_593 ( .A2(net_2276), .ZN(net_1882), .A1(net_520) );
AOI22_X2 inst_2223 ( .A2(net_2392), .B2(net_2159), .A1(net_1960), .ZN(net_1457), .B1(net_1450) );
DFFR_X1 inst_2135 ( .QN(net_2267), .RN(net_1347), .D(net_732), .CK(net_2516) );
NOR2_X2 inst_601 ( .A2(net_2268), .ZN(net_1890), .A1(net_520) );
CLKBUF_X2 inst_3119 ( .A(net_2826), .Z(net_2911) );
CLKBUF_X2 inst_3777 ( .A(net_3568), .Z(net_3569) );
NAND2_X4 inst_764 ( .ZN(net_2092), .A1(net_2091), .A2(net_83) );
DFF_X2 inst_1773 ( .QN(net_2428), .D(net_923), .CK(net_3463) );
OAI211_X2 inst_479 ( .C2(net_2328), .C1(net_1054), .ZN(net_1029), .A(net_899), .B(net_870) );
AOI22_X2 inst_2344 ( .B1(net_2197), .A1(net_2038), .A2(net_1548), .B2(net_1517), .ZN(net_820) );
INV_X2 inst_1547 ( .ZN(net_252), .A(x6319) );
XNOR2_X2 inst_29 ( .A(net_1643), .ZN(net_847), .B(net_846) );
CLKBUF_X2 inst_3326 ( .A(net_3014), .Z(net_3118) );
INV_X2 inst_1583 ( .ZN(net_917), .A(net_61) );
NAND2_X2 inst_771 ( .ZN(net_1447), .A1(net_1423), .A2(net_1228) );
AOI22_X2 inst_2369 ( .B2(net_2161), .A1(net_2038), .A2(net_1559), .B1(net_979), .ZN(net_687) );
DFFR_X1 inst_2152 ( .QN(net_2278), .RN(net_1347), .D(net_706), .CK(net_2720) );
CLKBUF_X2 inst_3947 ( .A(net_2462), .Z(net_3739) );
INV_X4 inst_1274 ( .A(net_2345), .ZN(net_1199) );
CLKBUF_X2 inst_3838 ( .A(net_3629), .Z(net_3630) );
NOR2_X2 inst_538 ( .A2(net_2201), .ZN(net_1149), .A1(net_482) );
CLKBUF_X2 inst_2831 ( .A(net_2528), .Z(net_2623) );
AND2_X2 inst_2651 ( .ZN(net_2077), .A2(net_2076), .A1(net_1186) );
INV_X4 inst_1319 ( .A(net_2203), .ZN(net_1873) );
INV_X4 inst_1300 ( .A(net_1829), .ZN(net_1596) );
CLKBUF_X2 inst_4201 ( .A(net_2948), .Z(net_3993) );
XNOR2_X2 inst_35 ( .B(net_2317), .ZN(net_617), .A(net_596) );
OAI21_X2 inst_358 ( .B1(net_1441), .ZN(net_1436), .A(net_1388), .B2(net_1141) );
SDFF_X2 inst_48 ( .SE(net_1768), .SI(net_1533), .Q(net_74), .D(net_74), .CK(net_3419) );
AOI22_X2 inst_2246 ( .B2(net_2160), .A1(net_1967), .B1(net_1450), .ZN(net_1384), .A2(net_934) );
DFF_X2 inst_1756 ( .QN(net_2350), .D(net_1435), .CK(net_3769) );
AOI22_X2 inst_2279 ( .ZN(net_1709), .A2(net_1551), .A1(net_1000), .B1(net_999), .B2(net_356) );
OAI21_X1 inst_443 ( .B2(net_2416), .B1(net_1250), .ZN(net_1248), .A(net_439) );
AND2_X4 inst_2600 ( .ZN(net_2175), .A2(net_1904), .A1(net_1748) );
DFF_X1 inst_2038 ( .Q(net_2396), .D(net_2181), .CK(net_3092) );
DFF_X1 inst_2044 ( .Q(net_2395), .D(net_1654), .CK(net_3088) );
NAND3_X2 inst_655 ( .A1(net_2189), .ZN(net_1151), .A2(net_1143), .A3(net_386) );
AOI22_X2 inst_2274 ( .B1(net_1768), .ZN(net_1708), .B2(net_1514), .A1(net_1001), .A2(net_788) );
INV_X16 inst_1700 ( .ZN(net_2041), .A(net_2040) );
AND4_X4 inst_2571 ( .A4(net_2430), .A3(net_2429), .A2(net_2420), .A1(net_2419), .ZN(net_2088) );
NAND3_X2 inst_695 ( .ZN(net_1900), .A3(net_1899), .A2(net_1898), .A1(net_1897) );
NAND2_X4 inst_730 ( .ZN(net_1829), .A1(net_1828), .A2(net_1825) );
CLKBUF_X2 inst_4038 ( .A(net_3829), .Z(net_3830) );
OAI21_X2 inst_321 ( .B2(net_2441), .B1(net_2015), .A(net_545), .ZN(x22) );
AOI222_X1 inst_2493 ( .B1(net_1995), .A1(net_1749), .B2(net_1558), .C1(net_1020), .ZN(net_1007), .A2(net_160), .C2(x3501) );
NOR2_X4 inst_511 ( .ZN(net_534), .A1(net_520), .A2(net_372) );
XNOR2_X2 inst_41 ( .ZN(net_2080), .A(net_2079), .B(net_1284) );
CLKBUF_X2 inst_3131 ( .A(net_2922), .Z(net_2923) );
CLKBUF_X2 inst_3559 ( .A(net_3350), .Z(net_3351) );
AND2_X2 inst_2645 ( .A1(net_2430), .A2(net_2429), .ZN(net_379) );
DFF_X1 inst_1989 ( .Q(net_2153), .D(net_1059), .CK(net_3389) );
INV_X8 inst_1164 ( .A(net_1964), .ZN(net_1918) );
CLKBUF_X2 inst_3112 ( .A(net_2903), .Z(net_2904) );
OAI22_X2 inst_152 ( .A1(net_1408), .B1(net_1406), .B2(net_203), .A2(net_117), .ZN(x528) );
INV_X8 inst_1152 ( .ZN(net_1621), .A(net_1618) );
INV_X4 inst_1242 ( .A(net_2381), .ZN(net_374) );
INV_X2 inst_1400 ( .A(net_575), .ZN(x1060) );
SDFF_X2 inst_89 ( .Q(net_1555), .D(net_1555), .SE(net_491), .CK(net_2665), .SI(x7297) );
INV_X2 inst_1520 ( .ZN(net_458), .A(x3884) );
OAI21_X2 inst_388 ( .B1(net_1742), .ZN(net_1340), .A(net_1339), .B2(net_1105) );
CLKBUF_X2 inst_3872 ( .A(net_3663), .Z(net_3664) );
INV_X2 inst_1535 ( .ZN(net_259), .A(x4790) );
OAI22_X2 inst_182 ( .B1(net_1427), .A1(net_529), .B2(net_190), .A2(net_92), .ZN(x1600) );
NAND2_X2 inst_788 ( .A1(net_1819), .ZN(net_1325), .A2(net_1209) );
NOR4_X1 inst_489 ( .A1(net_455), .ZN(net_452), .A3(net_451), .A2(net_275), .A4(x6039) );
NAND2_X2 inst_931 ( .A2(net_1632), .ZN(net_1083), .A1(net_695) );
CLKBUF_X2 inst_3174 ( .A(net_2965), .Z(net_2966) );
CLKBUF_X2 inst_3824 ( .A(net_3156), .Z(net_3616) );
INV_X2 inst_1674 ( .ZN(net_1870), .A(net_1866) );
CLKBUF_X2 inst_3622 ( .A(net_3413), .Z(net_3414) );
INV_X2 inst_1579 ( .ZN(net_227), .A(x6343) );
INV_X2 inst_1411 ( .A(net_565), .ZN(x1167) );
OR2_X1 inst_149 ( .A1(net_2168), .A2(x3932), .ZN(x1332) );
OAI22_X2 inst_193 ( .B1(net_1428), .A1(net_1426), .B2(net_250), .A2(net_105), .ZN(x1434) );
XNOR2_X2 inst_39 ( .A(net_2314), .ZN(net_432), .B(net_393) );
CLKBUF_X2 inst_4089 ( .A(net_2707), .Z(net_3881) );
INV_X2 inst_1415 ( .A(net_561), .ZN(x1218) );
AND2_X2 inst_2627 ( .A1(net_594), .A2(x7404), .ZN(x854) );
INV_X1 inst_1709 ( .ZN(net_1924), .A(net_1923) );
CLKBUF_X2 inst_3301 ( .A(net_2647), .Z(net_3093) );
AOI22_X2 inst_2320 ( .A2(net_2157), .B1(net_2096), .A1(net_1769), .B2(net_1514), .ZN(net_889) );
CLKBUF_X2 inst_3173 ( .A(net_2455), .Z(net_2965) );
SDFFR_X1 inst_125 ( .Q(net_2248), .D(net_2248), .SI(net_1580), .RN(net_1347), .SE(net_534), .CK(net_3313) );
AOI21_X2 inst_2534 ( .A(net_1785), .B1(net_910), .ZN(net_799), .B2(net_81) );
AOI22_X2 inst_2202 ( .B2(net_2112), .A1(net_1916), .B1(net_1915), .ZN(net_1479), .A2(net_1150) );
CLKBUF_X2 inst_3180 ( .A(net_2886), .Z(net_2972) );
CLKBUF_X2 inst_2987 ( .A(net_2778), .Z(net_2779) );
CLKBUF_X2 inst_3737 ( .A(net_3528), .Z(net_3529) );
INV_X2 inst_1636 ( .ZN(net_186), .A(x6650) );
OAI21_X2 inst_430 ( .A(net_1917), .ZN(net_1717), .B1(net_680), .B2(net_621) );
NOR2_X4 inst_515 ( .ZN(net_485), .A1(net_484), .A2(net_431) );
INV_X2 inst_1501 ( .A(net_2365), .ZN(net_364) );
AOI222_X2 inst_2473 ( .C1(net_2016), .A2(net_1548), .A1(net_590), .B1(net_589), .ZN(net_563), .B2(net_150), .C2(x5820) );
CLKBUF_X2 inst_3212 ( .A(net_3003), .Z(net_3004) );
INV_X16 inst_1698 ( .ZN(net_1967), .A(net_1966) );
AOI211_X2 inst_2565 ( .C2(net_2127), .C1(net_1929), .A(net_1886), .ZN(net_1846), .B(net_1785) );
NAND2_X2 inst_944 ( .A1(net_2046), .A2(net_1829), .ZN(net_998) );
CLKBUF_X2 inst_2945 ( .A(net_2532), .Z(net_2737) );
INV_X2 inst_1584 ( .ZN(net_224), .A(x4397) );
NAND4_X2 inst_642 ( .ZN(net_1941), .A3(net_1914), .A2(net_1835), .A1(net_1760), .A4(net_1196) );
OAI211_X2 inst_459 ( .C2(net_2323), .A(net_1856), .ZN(net_1058), .C1(net_1054), .B(net_876) );
CLKBUF_X2 inst_2993 ( .A(net_2658), .Z(net_2785) );
CLKBUF_X2 inst_2864 ( .A(net_2446), .Z(net_2656) );
CLKBUF_X2 inst_3476 ( .A(net_2884), .Z(net_3268) );
NAND2_X2 inst_1018 ( .A2(net_1264), .ZN(net_597), .A1(net_596) );
CLKBUF_X2 inst_3789 ( .A(net_3516), .Z(net_3581) );
CLKBUF_X2 inst_2933 ( .A(net_2724), .Z(net_2725) );
NAND3_X2 inst_700 ( .A2(net_1984), .ZN(net_1953), .A1(net_1826), .A3(net_1825) );
CLKBUF_X2 inst_3393 ( .A(net_3184), .Z(net_3185) );
OAI21_X2 inst_367 ( .B1(net_1443), .ZN(net_1422), .A(net_1380), .B2(net_1170) );
NAND2_X2 inst_957 ( .A1(net_1829), .ZN(net_928), .A2(net_295) );
NAND2_X2 inst_979 ( .A2(net_1547), .A1(net_961), .ZN(net_860) );
CLKBUF_X2 inst_2713 ( .A(net_2504), .Z(net_2505) );
NAND2_X2 inst_1008 ( .A2(net_2138), .A1(net_979), .ZN(net_664) );
CLKBUF_X2 inst_3409 ( .A(net_3200), .Z(net_3201) );
NOR2_X2 inst_559 ( .ZN(net_508), .A1(net_466), .A2(net_182) );
DFF_X1 inst_1871 ( .D(net_1824), .QN(net_108), .CK(net_3830) );
AOI22_X2 inst_2296 ( .B1(net_1768), .ZN(net_1696), .B2(net_1541), .A1(net_999), .A2(net_772) );
CLKBUF_X2 inst_3591 ( .A(net_3382), .Z(net_3383) );
AOI22_X2 inst_2300 ( .A1(net_1996), .B1(net_1749), .A2(net_1554), .ZN(net_922), .B2(net_156) );
OAI211_X2 inst_450 ( .C1(net_1639), .ZN(net_1106), .C2(net_1105), .A(net_824), .B(net_665) );
NOR2_X4 inst_520 ( .A1(net_1779), .A2(net_1757), .ZN(net_443) );
NAND2_X4 inst_745 ( .A2(net_2028), .ZN(net_1966), .A1(net_1965) );
CLKBUF_X2 inst_3658 ( .A(net_2992), .Z(net_3450) );
CLKBUF_X2 inst_3405 ( .A(net_3196), .Z(net_3197) );
CLKBUF_X2 inst_3888 ( .A(net_2769), .Z(net_3680) );
DFF_X1 inst_2032 ( .QN(net_2238), .D(net_836), .CK(net_2987) );
CLKBUF_X2 inst_4113 ( .A(net_2762), .Z(net_3905) );
CLKBUF_X2 inst_3623 ( .A(net_3414), .Z(net_3415) );
SDFF_X2 inst_80 ( .Q(net_1543), .D(net_1543), .SE(net_491), .CK(net_3120), .SI(x7526) );
DFF_X1 inst_2026 ( .QN(net_2233), .D(net_2061), .CK(net_3213) );
NAND2_X2 inst_836 ( .A1(net_1840), .ZN(net_1278), .A2(net_1261) );
INV_X2 inst_1556 ( .ZN(net_244), .A(x6430) );
CLKBUF_X2 inst_4040 ( .A(net_3831), .Z(net_3832) );
OAI22_X2 inst_241 ( .B2(net_2263), .A1(net_745), .ZN(net_738), .A2(net_737), .B1(net_534) );
NAND2_X2 inst_1059 ( .ZN(net_1715), .A1(net_1713), .A2(net_1361) );
NAND2_X2 inst_1075 ( .A1(net_2104), .ZN(net_1816), .A2(net_1260) );
NAND2_X2 inst_862 ( .A1(net_1838), .ZN(net_1221), .A2(net_366) );
CLKBUF_X2 inst_3918 ( .A(net_2936), .Z(net_3710) );
CLKBUF_X2 inst_2758 ( .A(net_2549), .Z(net_2550) );
NAND2_X2 inst_1116 ( .A1(net_2100), .ZN(net_2068), .A2(net_2067) );
AOI22_X2 inst_2257 ( .B2(net_2164), .A1(net_1967), .B1(net_1450), .ZN(net_1373), .A2(net_1213) );
CLKBUF_X2 inst_4173 ( .A(net_3964), .Z(net_3965) );
CLKBUF_X2 inst_3753 ( .A(net_3544), .Z(net_3545) );
DFF_X2 inst_1764 ( .D(net_1121), .QN(net_84), .CK(net_3238) );
NAND2_X2 inst_1104 ( .ZN(net_1998), .A2(net_1997), .A1(net_1782) );
INV_X8 inst_1159 ( .A(net_1848), .ZN(net_1791) );
AOI22_X2 inst_2355 ( .A1(net_783), .B1(net_782), .ZN(net_777), .A2(net_357), .B2(x3775) );
CLKBUF_X2 inst_3136 ( .A(net_2927), .Z(net_2928) );
OAI21_X2 inst_402 ( .B2(net_2380), .ZN(net_921), .B1(net_920), .A(net_629) );
OAI21_X2 inst_329 ( .B2(net_2314), .B1(net_2041), .ZN(net_1501), .A(net_1465) );
NOR3_X2 inst_494 ( .A3(net_2413), .A1(net_531), .ZN(net_489), .A2(net_271) );
NOR2_X2 inst_574 ( .A2(net_2346), .A1(net_2345), .ZN(net_365) );
NAND2_X2 inst_938 ( .A2(net_1640), .ZN(net_1062), .A1(net_832) );
AOI22_X2 inst_2347 ( .B1(net_2197), .A1(net_2038), .A2(net_1554), .B2(net_1541), .ZN(net_817) );
CLKBUF_X2 inst_4102 ( .A(net_3893), .Z(net_3894) );
INV_X4 inst_1229 ( .ZN(net_498), .A(net_411) );
INV_X4 inst_1288 ( .A(net_2325), .ZN(net_327) );
CLKBUF_X2 inst_3844 ( .A(net_3635), .Z(net_3636) );
CLKBUF_X2 inst_2894 ( .A(net_2685), .Z(net_2686) );
AOI22_X2 inst_2358 ( .A1(net_783), .B1(net_782), .ZN(net_773), .A2(net_772), .B2(x3595) );
DFFR_X1 inst_2125 ( .QN(net_2308), .D(net_1607), .RN(net_1347), .CK(net_2723) );
CLKBUF_X2 inst_3638 ( .A(net_3028), .Z(net_3430) );
CLKBUF_X2 inst_2959 ( .A(net_2750), .Z(net_2751) );
NOR2_X2 inst_599 ( .A2(net_2252), .ZN(net_1888), .A1(net_520) );
NAND2_X2 inst_1033 ( .ZN(net_424), .A1(net_385), .A2(net_273) );
INV_X2 inst_1683 ( .ZN(net_2193), .A(net_1584) );
CLKBUF_X2 inst_3865 ( .A(net_3656), .Z(net_3657) );
INV_X4 inst_1348 ( .ZN(net_2093), .A(net_1585) );
DFFR_X1 inst_2102 ( .QN(net_2291), .D(net_1613), .RN(net_1347), .CK(net_2651) );
DFF_X2 inst_1748 ( .QN(net_2352), .D(net_1425), .CK(net_4016) );
NOR2_X2 inst_541 ( .A2(net_2433), .A1(net_2359), .ZN(net_1143) );
CLKBUF_X2 inst_4047 ( .A(net_3838), .Z(net_3839) );
NOR2_X4 inst_505 ( .A2(net_2331), .ZN(net_1175), .A1(net_1171) );
INV_X2 inst_1365 ( .A(net_1019), .ZN(x2528) );
OAI22_X2 inst_198 ( .B2(net_2366), .ZN(net_1189), .A1(net_1188), .A2(net_404), .B1(net_364) );
CLKBUF_X2 inst_4125 ( .A(net_3916), .Z(net_3917) );
INV_X2 inst_1371 ( .A(net_1013), .ZN(x2649) );
INV_X2 inst_1644 ( .A(net_2283), .ZN(net_340) );
CLKBUF_X2 inst_3543 ( .A(net_3334), .Z(net_3335) );
NAND2_X2 inst_784 ( .A1(net_1817), .ZN(net_1329), .A2(net_1215) );
CLKBUF_X2 inst_3237 ( .A(net_3028), .Z(net_3029) );
INV_X4 inst_1264 ( .A(net_2355), .ZN(net_1239) );
CLKBUF_X2 inst_3461 ( .A(net_2773), .Z(net_3253) );
NAND3_X2 inst_690 ( .ZN(net_1737), .A1(net_1735), .A2(net_1734), .A3(net_1225) );
CLKBUF_X2 inst_3511 ( .A(net_3243), .Z(net_3303) );
DFF_X1 inst_2025 ( .QN(net_2234), .D(net_2059), .CK(net_3215) );
AOI222_X2 inst_2461 ( .C1(net_2016), .A2(net_1562), .A1(net_590), .B1(net_589), .ZN(net_575), .B2(net_164), .C2(x5493) );
NAND2_X4 inst_732 ( .A2(net_2073), .ZN(net_1835), .A1(net_931) );
OAI22_X2 inst_263 ( .B2(net_2256), .A2(net_936), .A1(net_745), .ZN(net_699), .B1(net_534) );
OAI22_X2 inst_185 ( .B1(net_1427), .A1(net_1426), .B2(net_201), .A2(net_89), .ZN(x1646) );
SDFF_X2 inst_75 ( .Q(net_1571), .D(net_1571), .SE(net_491), .CK(net_2628), .SI(x6845) );
OAI22_X2 inst_166 ( .A1(net_1408), .B1(net_1404), .B2(net_210), .A2(net_127), .ZN(x406) );
CLKBUF_X2 inst_3815 ( .A(net_3606), .Z(net_3607) );
SDFF_X2 inst_79 ( .SE(net_487), .Q(net_155), .D(net_155), .CK(net_2553), .SI(x4821) );
DFF_X2 inst_1757 ( .QN(net_2349), .D(net_1437), .CK(net_3765) );
CLKBUF_X2 inst_3851 ( .A(net_3642), .Z(net_3643) );
CLKBUF_X2 inst_2654 ( .A(net_2445), .Z(net_2446) );
CLKBUF_X2 inst_4118 ( .A(net_3909), .Z(net_3910) );
INV_X2 inst_1605 ( .ZN(net_207), .A(x4416) );
CLKBUF_X2 inst_2975 ( .A(net_2506), .Z(net_2767) );
DFF_X2 inst_1741 ( .QN(net_2335), .D(net_1482), .CK(net_3168) );
NAND2_X2 inst_1024 ( .A1(net_2015), .ZN(net_545), .A2(x5957) );
AOI22_X2 inst_2232 ( .ZN(net_1410), .A2(net_425), .A1(net_141), .B2(x6264), .B1(x5995) );
INV_X2 inst_1658 ( .ZN(net_177), .A(x4022) );
INV_X16 inst_1689 ( .A(net_1935), .ZN(net_1760) );
CLKBUF_X2 inst_3965 ( .A(net_3756), .Z(net_3757) );
CLKBUF_X2 inst_2846 ( .A(net_2480), .Z(net_2638) );
CLKBUF_X2 inst_3584 ( .A(net_3375), .Z(net_3376) );
INV_X2 inst_1448 ( .A(net_1519), .ZN(net_703) );
OAI21_X1 inst_440 ( .B2(net_2437), .B1(net_775), .A(net_530), .ZN(x1277) );
DFF_X2 inst_1816 ( .Q(net_1525), .CK(net_2454), .D(x5338) );
CLKBUF_X2 inst_3898 ( .A(net_3689), .Z(net_3690) );
AOI22_X2 inst_2373 ( .B2(net_2124), .A1(net_2038), .A2(net_1569), .B1(net_979), .ZN(net_683) );
CLKBUF_X2 inst_3381 ( .A(net_2819), .Z(net_3173) );
CLKBUF_X2 inst_3503 ( .A(net_3040), .Z(net_3295) );
NAND2_X2 inst_1091 ( .ZN(net_1898), .A1(net_910), .A2(net_660) );
DFF_X1 inst_1887 ( .D(net_1299), .QN(net_99), .CK(net_3874) );
INV_X4 inst_1331 ( .ZN(net_2002), .A(net_2001) );
CLKBUF_X2 inst_4138 ( .A(net_3929), .Z(net_3930) );
SDFF_X2 inst_52 ( .SE(net_1768), .SI(net_1527), .Q(net_79), .D(net_79), .CK(net_3387) );
NAND3_X2 inst_668 ( .A1(net_1947), .A2(net_1801), .ZN(net_1074), .A3(net_803) );
CLKBUF_X2 inst_3223 ( .A(net_3014), .Z(net_3015) );
CLKBUF_X2 inst_3579 ( .A(net_3370), .Z(net_3371) );
CLKBUF_X2 inst_3049 ( .A(net_2797), .Z(net_2841) );
CLKBUF_X2 inst_4154 ( .A(net_2534), .Z(net_3946) );
CLKBUF_X2 inst_3560 ( .A(net_3258), .Z(net_3352) );
CLKBUF_X2 inst_4159 ( .A(net_3950), .Z(net_3951) );
CLKBUF_X2 inst_2683 ( .A(net_2449), .Z(net_2475) );
INV_X2 inst_1672 ( .ZN(net_1855), .A(net_43) );
CLKBUF_X2 inst_4223 ( .A(net_4014), .Z(net_4015) );
CLKBUF_X2 inst_3349 ( .A(net_3140), .Z(net_3141) );
DFF_X1 inst_2015 ( .QN(net_2411), .D(net_1116), .CK(net_3922) );
CLKBUF_X2 inst_3179 ( .A(net_2667), .Z(net_2971) );
AOI21_X2 inst_2545 ( .A(net_1968), .ZN(net_544), .B1(net_497), .B2(net_398) );
CLKBUF_X2 inst_3059 ( .A(net_2676), .Z(net_2851) );
CLKBUF_X2 inst_3937 ( .A(net_3728), .Z(net_3729) );
CLKBUF_X2 inst_2970 ( .A(net_2761), .Z(net_2762) );
CLKBUF_X2 inst_2768 ( .A(net_2559), .Z(net_2560) );
DFF_X2 inst_1835 ( .QN(net_2204), .CK(net_2938), .D(x6623) );
CLKBUF_X2 inst_4085 ( .A(net_3876), .Z(net_3877) );
DFF_X1 inst_1910 ( .D(net_1315), .QN(net_131), .CK(net_3645) );
AND2_X4 inst_2587 ( .A1(net_2416), .A2(net_1754), .ZN(net_1666) );
NOR2_X1 inst_621 ( .ZN(net_341), .A2(net_56), .A1(net_53) );
CLKBUF_X2 inst_3115 ( .A(net_2906), .Z(net_2907) );
AOI211_X2 inst_2560 ( .C2(net_2126), .C1(net_1929), .A(net_1892), .B(net_1785), .ZN(net_678) );
CLKBUF_X2 inst_3219 ( .A(net_3010), .Z(net_3011) );
NAND2_X2 inst_815 ( .ZN(net_1298), .A2(net_1257), .A1(net_1216) );
CLKBUF_X2 inst_3031 ( .A(net_2822), .Z(net_2823) );
NAND2_X2 inst_875 ( .A1(net_1838), .ZN(net_1204), .A2(net_1203) );
INV_X4 inst_1257 ( .A(net_2425), .ZN(net_355) );
CLKBUF_X2 inst_3298 ( .A(net_3089), .Z(net_3090) );
CLKBUF_X2 inst_3482 ( .A(net_3273), .Z(net_3274) );
CLKBUF_X2 inst_3081 ( .A(net_2514), .Z(net_2873) );
INV_X2 inst_1387 ( .A(net_588), .ZN(x1266) );
DFF_X1 inst_1991 ( .Q(net_2155), .D(net_1023), .CK(net_3376) );
DFFR_X2 inst_2069 ( .QN(net_1575), .RN(net_1347), .D(net_1345), .CK(net_3954) );
AOI22_X2 inst_2365 ( .B2(net_2120), .A1(net_2038), .A2(net_1551), .B1(net_979), .ZN(net_691) );
DFFR_X1 inst_2108 ( .QN(net_2280), .D(net_1611), .RN(net_1347), .CK(net_2523) );
CLKBUF_X2 inst_3572 ( .A(net_3363), .Z(net_3364) );
CLKBUF_X2 inst_3066 ( .A(net_2857), .Z(net_2858) );
CLKBUF_X2 inst_4098 ( .A(net_2776), .Z(net_3890) );
AOI22_X2 inst_2250 ( .B2(net_2135), .A1(net_1967), .B1(net_1474), .ZN(net_1380), .A2(net_1225) );
CLKBUF_X2 inst_2978 ( .A(net_2769), .Z(net_2770) );
OAI21_X2 inst_413 ( .B1(net_2196), .ZN(net_756), .A(net_626), .B2(net_313) );
NAND2_X2 inst_859 ( .A1(net_1741), .ZN(net_1226), .A2(net_1225) );
CLKBUF_X2 inst_2672 ( .A(net_2463), .Z(net_2464) );
XNOR2_X2 inst_25 ( .ZN(net_1152), .B(net_1143), .A(net_322) );
CLKBUF_X2 inst_3323 ( .A(net_2836), .Z(net_3115) );
DFF_X1 inst_2019 ( .QN(net_2222), .D(net_2099), .CK(net_2446) );
CLKBUF_X2 inst_3527 ( .A(net_3254), .Z(net_3319) );
AOI221_X2 inst_2500 ( .B2(net_2121), .B1(net_1929), .A(net_1885), .C1(net_1863), .ZN(net_971), .C2(net_298) );
SDFF_X2 inst_69 ( .Q(net_1547), .D(net_1547), .SE(net_498), .CK(net_2914), .SI(x7442) );
CLKBUF_X2 inst_3434 ( .A(net_3225), .Z(net_3226) );
CLKBUF_X2 inst_3764 ( .A(net_2579), .Z(net_3556) );
CLKBUF_X2 inst_2669 ( .A(x7552), .Z(net_2461) );
INV_X16 inst_1691 ( .A(net_2034), .ZN(net_1769) );
NAND2_X2 inst_844 ( .A1(net_1840), .ZN(net_1269), .A2(net_1260) );
AOI222_X1 inst_2489 ( .B1(net_1995), .A1(net_1751), .B2(net_1562), .ZN(net_1011), .C1(net_782), .A2(net_164), .C2(x3428) );
CLKBUF_X2 inst_3688 ( .A(net_2921), .Z(net_3480) );
CLKBUF_X2 inst_3619 ( .A(net_2731), .Z(net_3411) );
AOI22_X2 inst_2340 ( .B1(net_2197), .A1(net_2038), .A2(net_1564), .B2(net_1530), .ZN(net_824) );
OAI211_X2 inst_460 ( .ZN(net_1057), .C2(net_1056), .C1(net_1052), .A(net_904), .B(net_874) );
INV_X2 inst_1455 ( .A(net_1529), .ZN(net_724) );
CLKBUF_X2 inst_3204 ( .A(net_2995), .Z(net_2996) );
AOI222_X1 inst_2497 ( .B1(net_1995), .A1(net_1751), .B2(net_1567), .ZN(net_1003), .C1(net_782), .A2(net_169), .C2(x3346) );
CLKBUF_X2 inst_3660 ( .A(net_2986), .Z(net_3452) );
CLKBUF_X2 inst_3421 ( .A(net_3212), .Z(net_3213) );
NOR2_X2 inst_560 ( .ZN(net_490), .A1(net_455), .A2(net_438) );
CLKBUF_X2 inst_2679 ( .A(net_2470), .Z(net_2471) );
XNOR2_X2 inst_16 ( .ZN(net_1187), .B(net_1186), .A(net_1173) );
CLKBUF_X2 inst_4230 ( .A(net_4021), .Z(net_4022) );
CLKBUF_X2 inst_3949 ( .A(net_3740), .Z(net_3741) );
CLKBUF_X2 inst_2808 ( .A(net_2521), .Z(net_2600) );
OAI22_X2 inst_156 ( .B1(net_1428), .A1(net_529), .B2(net_248), .A2(net_104), .ZN(x1442) );
DFF_X2 inst_1777 ( .QN(net_2433), .D(net_914), .CK(net_3621) );
DFF_X2 inst_1802 ( .Q(net_1517), .CK(net_2604), .D(x5820) );
NAND2_X2 inst_950 ( .A1(net_1830), .ZN(net_987), .A2(net_291) );
NAND2_X2 inst_1068 ( .A1(net_1999), .ZN(net_1767), .A2(net_613) );
NAND2_X2 inst_886 ( .ZN(net_1155), .A1(net_303), .A2(net_84) );
CLKBUF_X2 inst_3442 ( .A(net_2907), .Z(net_3234) );
CLKBUF_X2 inst_3955 ( .A(net_2930), .Z(net_3747) );
CLKBUF_X2 inst_2982 ( .A(net_2773), .Z(net_2774) );
CLKBUF_X2 inst_2693 ( .A(net_2484), .Z(net_2485) );
CLKBUF_X2 inst_3359 ( .A(net_3101), .Z(net_3151) );
INV_X4 inst_1218 ( .A(net_2168), .ZN(net_775) );
SDFF_X2 inst_96 ( .SE(net_488), .Q(net_147), .D(net_147), .CK(net_2540), .SI(x5020) );
CLKBUF_X2 inst_3020 ( .A(net_2444), .Z(net_2812) );
SDFF_X2 inst_101 ( .SE(net_488), .Q(net_146), .D(net_146), .CK(net_2537), .SI(x5058) );
INV_X2 inst_1549 ( .ZN(net_251), .A(x4604) );
CLKBUF_X2 inst_3555 ( .A(net_3083), .Z(net_3347) );
DFF_X1 inst_1969 ( .Q(net_2135), .D(net_1102), .CK(net_3397) );
CLKBUF_X2 inst_2881 ( .A(net_2672), .Z(net_2673) );
NAND2_X2 inst_821 ( .A1(net_1840), .ZN(net_1341), .A2(net_369) );
NAND2_X2 inst_980 ( .A2(net_1548), .A1(net_961), .ZN(net_859) );
NOR2_X4 inst_510 ( .A1(net_1781), .ZN(net_542), .A2(net_516) );
AOI22_X2 inst_2436 ( .B2(net_2149), .B1(net_1974), .ZN(net_1810), .A1(net_1789), .A2(net_329) );
CLKBUF_X2 inst_2832 ( .A(net_2472), .Z(net_2624) );
INV_X2 inst_1677 ( .A(net_2414), .ZN(net_1922) );
NOR2_X2 inst_603 ( .A2(net_2261), .ZN(net_1892), .A1(net_520) );
NAND2_X2 inst_830 ( .A1(net_1840), .ZN(net_1285), .A2(net_1284) );
DFF_X2 inst_1785 ( .QN(net_2381), .D(net_755), .CK(net_3856) );
OAI22_X2 inst_291 ( .A1(net_1615), .B1(net_1404), .B2(net_211), .A2(net_128), .ZN(x398) );
CLKBUF_X2 inst_2878 ( .A(net_2611), .Z(net_2670) );
CLKBUF_X2 inst_4213 ( .A(net_4004), .Z(net_4005) );
CLKBUF_X2 inst_3150 ( .A(net_2941), .Z(net_2942) );
AOI222_X1 inst_2494 ( .B1(net_1995), .A1(net_1749), .B2(net_1557), .ZN(net_1006), .C1(net_782), .A2(net_159), .C2(x3527) );
NAND2_X2 inst_776 ( .ZN(net_1365), .A1(net_1350), .A2(net_538) );
AOI21_X2 inst_2526 ( .A(net_1785), .B1(net_910), .ZN(net_807), .B2(net_73) );
AOI22_X2 inst_2286 ( .A1(net_1996), .B1(net_1749), .A2(net_1547), .ZN(net_976), .B2(net_149) );
NAND2_X2 inst_866 ( .A1(net_1838), .A2(net_1225), .ZN(net_1216) );
DFFR_X1 inst_2137 ( .QN(net_2269), .RN(net_1347), .D(net_727), .CK(net_2794) );
INV_X2 inst_1439 ( .A(net_1537), .ZN(net_737) );
DFF_X1 inst_1972 ( .Q(net_2138), .D(net_1104), .CK(net_3427) );
NOR2_X2 inst_558 ( .ZN(net_550), .A1(net_510), .A2(net_281) );
CLKBUF_X2 inst_3640 ( .A(net_3431), .Z(net_3432) );
OAI22_X2 inst_248 ( .B2(net_2269), .A1(net_745), .ZN(net_727), .A2(net_726), .B1(net_534) );
INV_X2 inst_1613 ( .ZN(net_203), .A(x6592) );
CLKBUF_X2 inst_3107 ( .A(net_2898), .Z(net_2899) );
OAI21_X2 inst_389 ( .B2(net_2364), .B1(net_1842), .ZN(net_1338), .A(net_1337) );
DFF_X1 inst_1919 ( .D(net_1245), .QN(net_109), .CK(net_3816) );
CLKBUF_X2 inst_2712 ( .A(net_2503), .Z(net_2504) );
INV_X2 inst_1382 ( .ZN(net_641), .A(net_640) );
CLKBUF_X2 inst_2795 ( .A(net_2586), .Z(net_2587) );
INV_X8 inst_1141 ( .A(net_1918), .ZN(net_1474) );
DFF_X2 inst_1807 ( .QN(net_2205), .CK(net_2637), .D(x6573) );
CLKBUF_X2 inst_3589 ( .A(net_3380), .Z(net_3381) );
AOI222_X1 inst_2488 ( .B1(net_1995), .A1(net_1751), .B2(net_1574), .ZN(net_1012), .C1(net_782), .A2(net_176), .C2(x3227) );
NAND2_X2 inst_932 ( .A2(net_1626), .ZN(net_1068), .A1(net_693) );
OAI22_X2 inst_180 ( .B1(net_1428), .A1(net_529), .B2(net_255), .A2(net_95), .ZN(x1559) );
NAND2_X2 inst_913 ( .A1(net_964), .A2(net_780), .ZN(x2909) );
DFF_X1 inst_1960 ( .Q(net_2126), .D(net_1087), .CK(net_3526) );
OAI22_X2 inst_302 ( .A2(net_2234), .A1(net_2013), .B1(net_1895), .B2(net_237), .ZN(x1913) );
NAND3_X2 inst_673 ( .A2(net_1793), .ZN(net_1069), .A1(net_983), .A3(net_789) );
CLKBUF_X2 inst_3585 ( .A(net_2987), .Z(net_3377) );
CLKBUF_X2 inst_3287 ( .A(net_2539), .Z(net_3079) );
OAI22_X2 inst_211 ( .A2(net_2217), .A1(net_1408), .B1(net_1406), .B2(net_204), .ZN(x2273) );
AOI222_X1 inst_2483 ( .B1(net_1995), .A1(net_1751), .B2(net_1568), .C1(net_1020), .ZN(net_1017), .A2(net_170), .C2(x3338) );
INV_X8 inst_1151 ( .A(net_2017), .ZN(net_1614) );
CLKBUF_X2 inst_3120 ( .A(net_2911), .Z(net_2912) );
INV_X2 inst_1414 ( .A(net_562), .ZN(x1113) );
NOR2_X2 inst_561 ( .A2(net_2279), .ZN(net_493), .A1(net_466) );
CLKBUF_X2 inst_3994 ( .A(net_2675), .Z(net_3786) );
OAI211_X4 inst_449 ( .A(net_1944), .C1(net_1741), .B(net_1617), .ZN(net_1293), .C2(net_1114) );
CLKBUF_X2 inst_4212 ( .A(net_4003), .Z(net_4004) );
AOI221_X2 inst_2505 ( .B2(net_2160), .B1(net_1929), .A(net_1887), .ZN(net_918), .C2(net_917), .C1(net_910) );
CLKBUF_X2 inst_2790 ( .A(net_2447), .Z(net_2582) );
DFFR_X1 inst_2138 ( .QN(net_2270), .RN(net_1347), .D(net_725), .CK(net_2509) );
INV_X2 inst_1641 ( .A(net_2285), .ZN(net_292) );
CLKBUF_X2 inst_2736 ( .A(x7552), .Z(net_2528) );
CLKBUF_X2 inst_3249 ( .A(net_3040), .Z(net_3041) );
OAI22_X2 inst_196 ( .A2(net_2363), .B2(net_1907), .B1(net_1841), .A1(net_1836), .ZN(net_1244) );
INV_X2 inst_1567 ( .ZN(net_233), .A(x4155) );
CLKBUF_X2 inst_3451 ( .A(net_3242), .Z(net_3243) );
AOI22_X2 inst_2417 ( .B2(net_2152), .B1(net_1974), .ZN(net_1790), .A1(net_1789), .A2(net_296) );
AOI22_X2 inst_2309 ( .A2(net_2110), .B1(net_2096), .A1(net_1769), .B2(net_1526), .ZN(net_900) );
INV_X2 inst_1403 ( .A(net_610), .ZN(x1086) );
OAI22_X2 inst_298 ( .A2(net_2211), .B1(net_1895), .A1(net_1615), .B2(net_193), .ZN(x2371) );
DFF_X1 inst_1856 ( .QN(net_2355), .D(net_1445), .CK(net_3759) );
CLKBUF_X2 inst_3614 ( .A(net_3405), .Z(net_3406) );
AND2_X2 inst_2603 ( .A2(net_2093), .ZN(net_1140), .A1(net_1139) );
XNOR2_X2 inst_42 ( .B(net_2333), .ZN(net_2186), .A(net_1182) );
DFFR_X1 inst_2153 ( .QN(net_2275), .RN(net_1347), .D(net_715), .CK(net_2460) );
CLKBUF_X2 inst_4084 ( .A(net_3588), .Z(net_3876) );
NOR2_X2 inst_588 ( .A2(net_2263), .ZN(net_1877), .A1(net_520) );
INV_X2 inst_1479 ( .A(net_2314), .ZN(net_1261) );
CLKBUF_X2 inst_3529 ( .A(net_3320), .Z(net_3321) );
DFF_X1 inst_2040 ( .QN(net_2407), .D(net_657), .CK(net_3755) );
OAI21_X2 inst_437 ( .B1(net_2417), .A(net_2415), .ZN(net_2032), .B2(net_1581) );
INV_X2 inst_1356 ( .A(net_1411), .ZN(x125) );
INV_X1 inst_1706 ( .ZN(net_1347), .A(x7544) );
AND2_X2 inst_2628 ( .A1(net_594), .A2(x7418), .ZN(x862) );
CLKBUF_X2 inst_3485 ( .A(net_3067), .Z(net_3277) );
AOI22_X2 inst_2220 ( .A2(net_2390), .B2(net_2107), .A1(net_1916), .ZN(net_1460), .B1(net_1450) );
NAND2_X2 inst_1045 ( .A1(net_1746), .ZN(net_1672), .A2(net_1228) );
CLKBUF_X2 inst_2743 ( .A(net_2534), .Z(net_2535) );
OAI22_X2 inst_252 ( .B2(net_2273), .A1(net_740), .ZN(net_719), .A2(net_718), .B1(net_534) );
NAND2_X2 inst_865 ( .A1(net_1838), .A2(net_1228), .ZN(net_1217) );
DFFR_X2 inst_2083 ( .QN(net_1578), .RN(net_1347), .D(net_1134), .CK(net_3763) );
NAND2_X2 inst_956 ( .A1(net_1829), .ZN(net_929), .A2(net_276) );
INV_X2 inst_1470 ( .A(net_1528), .ZN(net_722) );
AOI22_X2 inst_2247 ( .B2(net_2138), .A1(net_1967), .B1(net_1450), .ZN(net_1383), .A2(net_1235) );
INV_X4 inst_1213 ( .A(net_1402), .ZN(net_609) );
CLKBUF_X2 inst_3072 ( .A(net_2836), .Z(net_2864) );
OAI211_X2 inst_484 ( .C2(net_2319), .C1(net_1052), .ZN(net_1024), .A(net_888), .B(net_857) );
AOI222_X2 inst_2452 ( .C1(net_2017), .A2(net_1571), .A1(net_590), .B1(net_589), .ZN(net_584), .B2(net_173), .C2(x5294) );
XNOR2_X2 inst_32 ( .B(net_2323), .A(net_1650), .ZN(net_673) );
OAI21_X2 inst_428 ( .B2(net_2281), .B1(net_1848), .ZN(net_1664), .A(net_1663) );
DFF_X2 inst_1821 ( .Q(net_1530), .CK(net_2498), .D(x5448) );
CLKBUF_X2 inst_3418 ( .A(net_3209), .Z(net_3210) );
CLKBUF_X2 inst_3334 ( .A(net_3125), .Z(net_3126) );
OAI21_X2 inst_407 ( .ZN(net_769), .B1(net_768), .A(net_627), .B2(net_544) );
CLKBUF_X2 inst_3558 ( .A(net_3349), .Z(net_3350) );
INV_X4 inst_1208 ( .A(net_1614), .ZN(net_1408) );
SDFF_X2 inst_97 ( .SE(net_488), .Q(net_165), .D(net_165), .CK(net_2737), .SI(x4524) );
NOR2_X2 inst_616 ( .ZN(net_2036), .A2(net_2033), .A1(net_1978) );
NAND2_X2 inst_775 ( .A1(net_2166), .ZN(net_1366), .A2(net_1351) );
NOR2_X1 inst_620 ( .A1(net_1918), .A2(net_813), .ZN(net_593) );
NAND3_X2 inst_652 ( .A2(net_1918), .ZN(net_1195), .A1(net_1194), .A3(net_537) );
DFF_X2 inst_1784 ( .QN(net_2377), .D(net_756), .CK(net_3890) );
CLKBUF_X2 inst_3118 ( .A(net_2909), .Z(net_2910) );
DFFR_X2 inst_2071 ( .QN(net_2416), .RN(net_1347), .D(net_1248), .CK(net_3989) );
NAND3_X2 inst_677 ( .A2(net_2169), .A1(net_603), .ZN(net_602), .A3(net_601) );
OR2_X4 inst_130 ( .A2(net_1904), .A1(net_1752), .ZN(net_440) );
INV_X2 inst_1427 ( .ZN(net_434), .A(net_433) );
INV_X2 inst_1566 ( .ZN(net_234), .A(x4219) );
INV_X2 inst_1409 ( .A(net_567), .ZN(x1136) );
AOI22_X2 inst_2242 ( .B2(net_2129), .A1(net_1967), .B1(net_1474), .ZN(net_1388), .A2(net_1218) );
SDFF_X2 inst_87 ( .Q(net_1568), .D(net_1568), .SE(net_491), .CK(net_2613), .SI(x6936) );
CLKBUF_X2 inst_2996 ( .A(net_2787), .Z(net_2788) );
NAND2_X2 inst_1054 ( .A1(net_1741), .ZN(net_1681), .A2(net_1205) );
CLKBUF_X2 inst_2918 ( .A(net_2709), .Z(net_2710) );
NAND2_X2 inst_972 ( .A2(net_1546), .A1(net_961), .ZN(net_867) );
CLKBUF_X2 inst_2721 ( .A(net_2512), .Z(net_2513) );
INV_X2 inst_1671 ( .ZN(net_1852), .A(net_1851) );
CLKBUF_X2 inst_3074 ( .A(net_2865), .Z(net_2866) );
NAND2_X2 inst_800 ( .A2(net_1683), .ZN(net_1313), .A1(net_1273) );
DFF_X1 inst_1843 ( .QN(net_2325), .D(net_1503), .CK(net_3072) );
XOR2_X1 inst_10 ( .Z(net_2183), .B(net_1198), .A(net_486) );
CLKBUF_X2 inst_3795 ( .A(net_2805), .Z(net_3587) );
XOR2_X1 inst_4 ( .Z(net_2177), .A(net_1175), .B(net_330) );
CLKBUF_X2 inst_2884 ( .A(net_2504), .Z(net_2676) );
NOR2_X2 inst_600 ( .A2(net_2250), .ZN(net_1889), .A1(net_520) );
CLKBUF_X2 inst_3272 ( .A(net_3063), .Z(net_3064) );
INV_X4 inst_1194 ( .ZN(net_840), .A(net_650) );
OAI22_X2 inst_204 ( .A2(net_2227), .B1(net_1614), .A1(net_1405), .B2(net_251), .ZN(x2071) );
SDFF_X2 inst_49 ( .SE(net_1768), .SI(net_1531), .Q(net_75), .D(net_75), .CK(net_3208) );
DFF_X1 inst_1866 ( .D(net_1358), .QN(net_96), .CK(net_3655) );
INV_X2 inst_1550 ( .ZN(net_250), .A(x4040) );
DFF_X1 inst_1878 ( .D(net_1324), .QN(net_112), .CK(net_3607) );
NAND2_X2 inst_910 ( .A1(net_968), .A2(net_771), .ZN(x2819) );
CLKBUF_X2 inst_4097 ( .A(net_3263), .Z(net_3889) );
NAND3_X2 inst_693 ( .A2(net_2090), .A1(net_2073), .ZN(net_1788), .A3(net_1776) );
NAND2_X4 inst_765 ( .ZN(net_2103), .A2(net_2102), .A1(net_2100) );
INV_X4 inst_1276 ( .A(net_2359), .ZN(net_1218) );
OAI22_X2 inst_256 ( .B2(net_2277), .A1(net_714), .ZN(net_710), .A2(net_709), .B1(net_534) );
DFF_X1 inst_1902 ( .D(net_1301), .QN(net_120), .CK(net_3574) );
NAND2_X2 inst_937 ( .A2(net_1642), .ZN(net_1063), .A1(net_829) );
NAND2_X2 inst_908 ( .A1(net_981), .A2(net_784), .ZN(x2846) );
OAI21_X2 inst_355 ( .B2(net_2373), .B1(net_1443), .ZN(net_1439), .A(net_1378) );
OAI22_X2 inst_218 ( .A2(net_2238), .A1(net_2013), .B1(net_1404), .B2(net_242), .ZN(x1835) );
CLKBUF_X2 inst_3647 ( .A(net_2872), .Z(net_3439) );
CLKBUF_X2 inst_3498 ( .A(net_3289), .Z(net_3290) );
CLKBUF_X2 inst_3422 ( .A(net_2869), .Z(net_3214) );
CLKBUF_X2 inst_3978 ( .A(net_3447), .Z(net_3770) );
CLKBUF_X2 inst_3832 ( .A(net_2978), .Z(net_3624) );
CLKBUF_X2 inst_4039 ( .A(net_2936), .Z(net_3831) );
CLKBUF_X2 inst_3693 ( .A(net_2593), .Z(net_3485) );
CLKBUF_X2 inst_2967 ( .A(net_2758), .Z(net_2759) );
CLKBUF_X2 inst_3769 ( .A(net_3560), .Z(net_3561) );
CLKBUF_X2 inst_4053 ( .A(net_3843), .Z(net_3845) );
DFFR_X2 inst_2078 ( .QN(net_2415), .RN(net_1347), .D(net_1176), .CK(net_3945) );
DFF_X2 inst_1747 ( .QN(net_2359), .D(net_1436), .CK(net_3632) );
NAND3_X2 inst_699 ( .A1(net_2006), .ZN(net_1944), .A2(net_1835), .A3(net_1199) );
CLKBUF_X2 inst_3917 ( .A(net_3708), .Z(net_3709) );
INV_X2 inst_1462 ( .A(net_2333), .ZN(net_368) );
AOI22_X2 inst_2273 ( .ZN(net_1707), .B1(net_1001), .A1(net_999), .B2(net_790), .A2(net_398) );
CLKBUF_X2 inst_2682 ( .A(net_2448), .Z(net_2474) );
AND4_X2 inst_2574 ( .A2(net_2050), .ZN(net_1913), .A4(net_1909), .A3(net_846), .A1(net_522) );
AOI22_X2 inst_2229 ( .ZN(net_1413), .A2(net_427), .A1(net_144), .B2(x6188), .B1(x5995) );
DFF_X1 inst_2003 ( .QN(net_2231), .D(net_1075), .CK(net_3252) );
NAND2_X2 inst_964 ( .A2(net_1556), .A1(net_961), .ZN(net_876) );
CLKBUF_X2 inst_2787 ( .A(net_2578), .Z(net_2579) );
CLKBUF_X2 inst_3372 ( .A(net_3163), .Z(net_3164) );
AND2_X4 inst_2599 ( .A2(net_2380), .A1(net_2379), .ZN(net_2173) );
AOI22_X2 inst_2426 ( .B2(net_2148), .B1(net_1974), .ZN(net_1800), .A1(net_1791), .A2(net_274) );
INV_X4 inst_1245 ( .ZN(net_1098), .A(net_367) );
AOI22_X2 inst_2313 ( .A2(net_2146), .B1(net_2096), .A1(net_1769), .B2(net_1530), .ZN(net_896) );
CLKBUF_X2 inst_3971 ( .A(net_3762), .Z(net_3763) );
CLKBUF_X2 inst_3788 ( .A(net_3579), .Z(net_3580) );
INV_X2 inst_1485 ( .A(net_1539), .ZN(net_742) );
CLKBUF_X2 inst_3663 ( .A(net_3454), .Z(net_3455) );
CLKBUF_X2 inst_3001 ( .A(net_2792), .Z(net_2793) );
CLKBUF_X2 inst_2818 ( .A(net_2520), .Z(net_2610) );
CLKBUF_X2 inst_3008 ( .A(net_2799), .Z(net_2800) );
CLKBUF_X2 inst_3198 ( .A(net_2484), .Z(net_2990) );
OAI21_X4 inst_317 ( .ZN(net_1990), .B2(net_1988), .A(net_1782), .B1(net_1665) );
NAND2_X4 inst_750 ( .ZN(net_1983), .A2(net_1982), .A1(net_1980) );
NAND2_X1 inst_1123 ( .A2(net_1238), .ZN(net_670), .A1(net_659) );
CLKBUF_X2 inst_2904 ( .A(net_2660), .Z(net_2696) );
OAI22_X2 inst_278 ( .B2(net_2300), .B1(net_1865), .ZN(net_1610), .A1(net_1603), .A2(net_726) );
AOI22_X2 inst_2383 ( .B1(net_839), .A1(net_661), .ZN(net_639), .A2(net_376), .B2(net_77) );
INV_X16 inst_1701 ( .ZN(net_2096), .A(net_2095) );
OAI211_X2 inst_467 ( .C1(net_1052), .ZN(net_1046), .C2(net_1045), .A(net_892), .B(net_852) );
CLKBUF_X2 inst_3677 ( .A(net_3468), .Z(net_3469) );
CLKBUF_X2 inst_4071 ( .A(net_3862), .Z(net_3863) );
CLKBUF_X2 inst_3456 ( .A(net_3247), .Z(net_3248) );
CLKBUF_X2 inst_2963 ( .A(net_2754), .Z(net_2755) );
INV_X2 inst_1628 ( .ZN(net_193), .A(x5058) );
INV_X4 inst_1329 ( .ZN(net_1988), .A(net_1987) );
AOI222_X2 inst_2469 ( .C1(net_2014), .A2(net_1555), .A1(net_590), .B1(net_589), .ZN(net_567), .B2(net_157), .C2(x5657) );
INV_X4 inst_1204 ( .A(net_1402), .ZN(net_594) );
CLKBUF_X2 inst_4066 ( .A(net_3857), .Z(net_3858) );
OAI22_X2 inst_225 ( .B2(net_2297), .B1(net_1865), .ZN(net_952), .A1(net_951), .A2(net_950) );
NOR2_X4 inst_508 ( .A2(net_2356), .ZN(net_659), .A1(net_598) );
AND2_X2 inst_2618 ( .A1(net_609), .A2(x7145), .ZN(x734) );
INV_X8 inst_1135 ( .A(net_1765), .ZN(net_999) );
CLKBUF_X2 inst_3715 ( .A(net_2976), .Z(net_3507) );
NOR2_X2 inst_590 ( .A2(net_2254), .ZN(net_1879), .A1(net_520) );
AOI21_X2 inst_2553 ( .A(net_1935), .ZN(net_1759), .B2(net_1352), .B1(net_1246) );
CLKBUF_X2 inst_3127 ( .A(net_2918), .Z(net_2919) );
CLKBUF_X2 inst_3042 ( .A(net_2833), .Z(net_2834) );
CLKBUF_X2 inst_3243 ( .A(net_3034), .Z(net_3035) );
DFF_X2 inst_1729 ( .QN(net_2313), .D(net_1502), .CK(net_3358) );
NAND2_X2 inst_1105 ( .ZN(net_2009), .A1(net_2008), .A2(net_1873) );
CLKBUF_X2 inst_2746 ( .A(net_2483), .Z(net_2538) );
NAND2_X2 inst_981 ( .A2(net_1549), .A1(net_961), .ZN(net_858) );
INV_X4 inst_1266 ( .ZN(net_324), .A(net_45) );
DFFR_X1 inst_2094 ( .QN(net_1584), .RN(net_1347), .D(net_1136), .CK(net_3733) );
OAI21_X2 inst_330 ( .B2(net_2316), .B1(net_1507), .ZN(net_1500), .A(net_1464) );
CLKBUF_X2 inst_3417 ( .A(net_2670), .Z(net_3209) );
CLKBUF_X2 inst_3733 ( .A(net_3524), .Z(net_3525) );
OAI22_X2 inst_165 ( .A1(net_1408), .B1(net_1407), .B2(net_225), .A2(net_131), .ZN(x342) );
CLKBUF_X2 inst_3491 ( .A(net_2771), .Z(net_3283) );
CLKBUF_X2 inst_3566 ( .A(net_3357), .Z(net_3358) );
AOI22_X2 inst_2393 ( .B1(net_2197), .ZN(net_1620), .A1(net_1619), .B2(net_1531), .A2(net_932) );
INV_X8 inst_1176 ( .ZN(net_2040), .A(net_2039) );
DFF_X2 inst_1838 ( .Q(net_1521), .CK(net_2585), .D(x5892) );
SDFF_X2 inst_71 ( .Q(net_1548), .D(net_1548), .SE(net_396), .CK(net_2913), .SI(x7418) );
INV_X2 inst_1454 ( .A(net_2416), .ZN(net_375) );
CLKBUF_X2 inst_4079 ( .A(net_3870), .Z(net_3871) );
INV_X4 inst_1232 ( .A(net_1778), .ZN(net_487) );
CLKBUF_X2 inst_3231 ( .A(net_3022), .Z(net_3023) );
CLKBUF_X2 inst_3147 ( .A(net_2880), .Z(net_2939) );
DFF_X1 inst_1945 ( .Q(net_2111), .D(net_1034), .CK(net_3161) );
CLKBUF_X2 inst_4172 ( .A(net_3963), .Z(net_3964) );
CLKBUF_X2 inst_2657 ( .A(net_2448), .Z(net_2449) );
AND2_X2 inst_2605 ( .A1(net_609), .A2(x6936), .ZN(x651) );
NAND2_X4 inst_758 ( .ZN(net_2034), .A2(net_2033), .A1(net_1963) );
OAI21_X2 inst_336 ( .B1(net_2041), .ZN(net_1494), .A(net_1457), .B2(net_1031) );
DFFR_X1 inst_2146 ( .QN(net_2252), .RN(net_1347), .D(net_697), .CK(net_2832) );
CLKBUF_X2 inst_3437 ( .A(net_3228), .Z(net_3229) );
CLKBUF_X2 inst_2703 ( .A(net_2494), .Z(net_2495) );
OAI21_X2 inst_376 ( .B1(net_1746), .ZN(net_1409), .A(net_1366), .B2(net_82) );
DFF_X1 inst_1939 ( .QN(net_2220), .D(net_1133), .CK(net_3304) );
CLKBUF_X2 inst_3268 ( .A(net_2993), .Z(net_3060) );
CLKBUF_X2 inst_2902 ( .A(net_2693), .Z(net_2694) );
OR2_X2 inst_143 ( .ZN(net_2199), .A1(net_763), .A2(net_651) );
DFF_X1 inst_1953 ( .Q(net_2119), .D(net_1068), .CK(net_3562) );
CLKBUF_X2 inst_3016 ( .A(net_2807), .Z(net_2808) );
DFF_X1 inst_1958 ( .Q(net_2124), .D(net_1084), .CK(net_3438) );
AOI22_X2 inst_2337 ( .B1(net_2197), .A1(net_2038), .A2(net_1567), .B2(net_1527), .ZN(net_827) );
CLKBUF_X2 inst_3250 ( .A(net_2465), .Z(net_3042) );
CLKBUF_X2 inst_3240 ( .A(net_3031), .Z(net_3032) );
DFF_X2 inst_1778 ( .QN(net_2427), .D(net_798), .CK(net_3671) );
DFF_X2 inst_1736 ( .QN(net_2316), .D(net_1500), .CK(net_3346) );
NAND2_X2 inst_1040 ( .A2(net_2066), .ZN(net_1645), .A1(net_1644) );
CLKBUF_X2 inst_4027 ( .A(net_3818), .Z(net_3819) );
CLKBUF_X2 inst_3880 ( .A(net_3605), .Z(net_3672) );
CLKBUF_X2 inst_3100 ( .A(net_2891), .Z(net_2892) );
CLKBUF_X2 inst_4052 ( .A(net_3843), .Z(net_3844) );
SDFF_X2 inst_111 ( .SE(net_487), .Q(net_175), .D(net_175), .CK(net_2704), .SI(x4323) );
INV_X2 inst_1596 ( .ZN(net_214), .A(x6550) );
CLKBUF_X2 inst_3146 ( .A(net_2937), .Z(net_2938) );
DFF_X2 inst_1723 ( .QN(net_2336), .D(net_1490), .CK(net_2981) );
CLKBUF_X2 inst_3278 ( .A(net_3069), .Z(net_3070) );
DFF_X1 inst_2056 ( .Q(net_2390), .D(net_506), .CK(net_3277) );
CLKBUF_X2 inst_3752 ( .A(net_2885), .Z(net_3544) );
DFFR_X1 inst_2116 ( .QN(net_2307), .D(net_1599), .RN(net_1347), .CK(net_2474) );
AOI22_X2 inst_2265 ( .ZN(net_1697), .A2(net_1554), .B1(net_1001), .A1(net_1000), .B2(net_811) );
OAI22_X2 inst_284 ( .A2(net_2212), .A1(net_1615), .B1(net_1404), .B2(net_263), .ZN(x2355) );
CLKBUF_X2 inst_2825 ( .A(net_2616), .Z(net_2617) );
INV_X2 inst_1555 ( .ZN(net_245), .A(x4502) );
CLKBUF_X2 inst_4031 ( .A(net_3822), .Z(net_3823) );
INV_X4 inst_1293 ( .ZN(net_792), .A(net_64) );
CLKBUF_X2 inst_3805 ( .A(net_3453), .Z(net_3597) );
AND2_X4 inst_2579 ( .ZN(net_466), .A1(net_387), .A2(net_381) );
OAI22_X2 inst_280 ( .B2(net_2289), .B1(net_1865), .ZN(net_1612), .A1(net_1603), .A2(net_749) );
OAI21_X2 inst_346 ( .B2(net_1484), .ZN(net_1482), .A(net_1451), .B1(net_1346) );
CLKBUF_X2 inst_3157 ( .A(net_2948), .Z(net_2949) );
NAND2_X2 inst_978 ( .A2(net_1572), .A1(net_961), .ZN(net_861) );
HA_X1 inst_1713 ( .S(net_506), .CO(net_505), .A(net_434), .B(net_346) );
CLKBUF_X2 inst_2955 ( .A(net_2746), .Z(net_2747) );
CLKBUF_X2 inst_3926 ( .A(net_2629), .Z(net_3718) );
CLKBUF_X2 inst_3929 ( .A(net_3720), .Z(net_3721) );
CLKBUF_X2 inst_3137 ( .A(net_2928), .Z(net_2929) );
CLKBUF_X2 inst_3852 ( .A(net_3643), .Z(net_3644) );
AOI211_X2 inst_2566 ( .C2(net_2111), .C1(net_1974), .ZN(net_1860), .A(net_1859), .B(net_558) );
NOR3_X2 inst_495 ( .A3(net_2310), .A2(net_1583), .ZN(net_470), .A1(net_45) );
NAND2_X2 inst_1051 ( .A1(net_1746), .ZN(net_1678), .A2(net_1238) );
NAND2_X2 inst_951 ( .A2(net_2193), .A1(net_1830), .ZN(net_986) );
DFF_X1 inst_1864 ( .D(net_2187), .QN(net_104), .CK(net_3835) );
CLKBUF_X2 inst_3603 ( .A(net_3394), .Z(net_3395) );
CLKBUF_X2 inst_3224 ( .A(net_3015), .Z(net_3016) );
CLKBUF_X2 inst_3043 ( .A(net_2834), .Z(net_2835) );
INV_X2 inst_1359 ( .ZN(net_1156), .A(net_1155) );
CLKBUF_X2 inst_3188 ( .A(net_2627), .Z(net_2980) );
CLKBUF_X2 inst_3129 ( .A(net_2920), .Z(net_2921) );
CLKBUF_X2 inst_2893 ( .A(net_2612), .Z(net_2685) );
NOR2_X2 inst_573 ( .A2(net_2350), .A1(net_2349), .ZN(net_273) );
CLKBUF_X2 inst_3797 ( .A(net_3189), .Z(net_3589) );
SDFF_X2 inst_100 ( .SE(net_487), .Q(net_174), .D(net_174), .CK(net_2947), .SI(x4336) );
NAND2_X2 inst_921 ( .A1(net_1637), .ZN(net_1096), .A2(net_819) );
INV_X2 inst_1453 ( .A(net_2105), .ZN(net_1031) );
OAI22_X2 inst_279 ( .B2(net_2280), .B1(net_1865), .ZN(net_1611), .A1(net_951), .A2(net_730) );
CLKBUF_X2 inst_3970 ( .A(net_3761), .Z(net_3762) );
CLKBUF_X2 inst_3387 ( .A(net_2768), .Z(net_3179) );
CLKBUF_X2 inst_3007 ( .A(net_2798), .Z(net_2799) );
SDFF_X2 inst_81 ( .SE(net_488), .Q(net_153), .D(net_153), .CK(net_2577), .SI(x4866) );
CLKBUF_X2 inst_4185 ( .A(net_3976), .Z(net_3977) );
CLKBUF_X2 inst_3544 ( .A(net_2750), .Z(net_3336) );
CLKBUF_X2 inst_3512 ( .A(net_3303), .Z(net_3304) );
NAND2_X2 inst_790 ( .A1(net_1816), .ZN(net_1323), .A2(net_1206) );
NAND2_X2 inst_1009 ( .A2(net_2137), .A1(net_979), .ZN(net_663) );
INV_X4 inst_1206 ( .A(net_2015), .ZN(net_1406) );
CLKBUF_X2 inst_2954 ( .A(net_2677), .Z(net_2746) );
NAND2_X4 inst_733 ( .A2(net_1989), .ZN(net_1850), .A1(net_1827) );
CLKBUF_X2 inst_3466 ( .A(net_2645), .Z(net_3258) );
DFF_X1 inst_1959 ( .Q(net_2125), .D(net_1062), .CK(net_3530) );
AND2_X4 inst_2582 ( .ZN(net_382), .A1(net_83), .A2(x3098) );
OR2_X2 inst_142 ( .A2(net_2326), .ZN(net_1644), .A1(net_1643) );
SDFF_X2 inst_78 ( .Q(net_1573), .D(net_1573), .SE(net_491), .CK(net_2622), .SI(x6773) );
INV_X2 inst_1487 ( .A(net_2319), .ZN(net_346) );
CLKBUF_X2 inst_2813 ( .A(net_2571), .Z(net_2605) );
OAI22_X2 inst_177 ( .B1(net_1427), .A1(net_529), .B2(net_195), .A2(net_102), .ZN(x1462) );
NAND2_X2 inst_783 ( .A1(net_1821), .ZN(net_1330), .A2(net_1219) );
CLKBUF_X2 inst_3522 ( .A(net_3118), .Z(net_3314) );
DFF_X1 inst_1933 ( .D(net_1118), .QN(net_62), .CK(net_3471) );
DFF_X1 inst_2014 ( .QN(net_2214), .D(net_1073), .CK(net_3286) );
INV_X8 inst_1142 ( .A(net_1931), .ZN(net_525) );
DFF_X2 inst_1758 ( .QN(net_2353), .D(net_1434), .CK(net_3738) );
NOR2_X2 inst_615 ( .A2(net_2414), .ZN(net_2031), .A1(net_2030) );
CLKBUF_X2 inst_3816 ( .A(net_3560), .Z(net_3608) );
CLKBUF_X2 inst_2822 ( .A(net_2599), .Z(net_2614) );
AOI222_X2 inst_2467 ( .C1(net_2016), .A2(net_1556), .A1(net_590), .B1(net_589), .ZN(net_569), .B2(net_158), .C2(x5628) );
CLKBUF_X2 inst_3843 ( .A(net_3634), .Z(net_3635) );
INV_X2 inst_1381 ( .A(net_1003), .ZN(x2579) );
DFF_X1 inst_2031 ( .QN(net_2239), .D(net_835), .CK(net_2989) );
NAND4_X2 inst_643 ( .ZN(net_1942), .A3(net_1914), .A2(net_1835), .A1(net_1760), .A4(net_1197) );
OAI21_X2 inst_338 ( .B2(net_2329), .B1(net_2041), .ZN(net_1492), .A(net_1467) );
AOI22_X2 inst_2412 ( .B2(net_2117), .ZN(net_1641), .A1(net_1619), .A2(net_1205), .B1(net_979) );
CLKBUF_X2 inst_4005 ( .A(net_3796), .Z(net_3797) );
AOI22_X2 inst_2214 ( .A2(net_2179), .B2(net_2149), .A1(net_1960), .B1(net_1915), .ZN(net_1466) );
CLKBUF_X2 inst_4146 ( .A(net_3937), .Z(net_3938) );
DFF_X1 inst_1997 ( .Q(net_2161), .D(net_1086), .CK(net_3257) );
AOI222_X2 inst_2474 ( .C1(net_2017), .A2(net_1557), .A1(net_590), .B1(net_589), .ZN(net_562), .B2(net_159), .C2(x5605) );
NAND2_X2 inst_1017 ( .A2(net_1239), .ZN(net_599), .A1(net_541) );
NOR2_X2 inst_579 ( .A1(net_1896), .ZN(net_1725), .A2(net_82) );
CLKBUF_X2 inst_3736 ( .A(net_3527), .Z(net_3528) );
AOI222_X1 inst_2495 ( .B1(net_1995), .A1(net_1751), .B2(net_1556), .ZN(net_1005), .C1(net_782), .A2(net_158), .C2(x3558) );
AOI22_X2 inst_2297 ( .B1(net_1768), .ZN(net_1688), .B2(net_1517), .A1(net_999), .A2(net_373) );
CLKBUF_X2 inst_4019 ( .A(net_3810), .Z(net_3811) );
CLKBUF_X2 inst_3341 ( .A(net_3132), .Z(net_3133) );
OAI22_X2 inst_281 ( .B2(net_2291), .B1(net_1865), .ZN(net_1613), .A1(net_1597), .A2(net_744) );
CLKBUF_X2 inst_3236 ( .A(net_2610), .Z(net_3028) );
NAND3_X2 inst_698 ( .A1(net_2006), .ZN(net_1943), .A2(net_1835), .A3(net_414) );
DFF_X2 inst_1836 ( .Q(net_1529), .CK(net_2743), .D(x5429) );
CLKBUF_X2 inst_3964 ( .A(net_3379), .Z(net_3756) );
CLKBUF_X2 inst_3944 ( .A(net_3735), .Z(net_3736) );
CLKBUF_X2 inst_3394 ( .A(net_2895), .Z(net_3186) );
CLKBUF_X2 inst_3408 ( .A(net_3199), .Z(net_3200) );
SDFF_X2 inst_88 ( .Q(net_1549), .D(net_1549), .SE(net_491), .CK(net_2896), .SI(x7404) );
CLKBUF_X2 inst_2863 ( .A(net_2654), .Z(net_2655) );
AOI221_X2 inst_2508 ( .B2(net_2131), .B1(net_1929), .A(net_1891), .C1(net_1863), .ZN(net_1762), .C2(net_317) );
OAI21_X2 inst_360 ( .B2(net_2404), .B1(net_1441), .ZN(net_1434), .A(net_1372) );
CLKBUF_X2 inst_3897 ( .A(net_3688), .Z(net_3689) );
NAND2_X2 inst_773 ( .A1(net_1715), .A2(net_1686), .ZN(net_1398) );
CLKBUF_X2 inst_2946 ( .A(net_2669), .Z(net_2738) );
CLKBUF_X2 inst_3908 ( .A(net_3308), .Z(net_3700) );
CLKBUF_X2 inst_3620 ( .A(net_3411), .Z(net_3412) );
CLKBUF_X2 inst_3754 ( .A(net_3545), .Z(net_3546) );
OAI22_X2 inst_260 ( .B2(net_2253), .A2(net_941), .A1(net_745), .ZN(net_702), .B1(net_534) );
NAND2_X1 inst_1129 ( .ZN(net_2055), .A2(net_1988), .A1(net_493) );
NAND2_X2 inst_837 ( .A1(net_1742), .ZN(net_1277), .A2(net_1276) );
NAND2_X4 inst_744 ( .ZN(net_1963), .A2(net_1961), .A1(net_1832) );
CLKBUF_X2 inst_3211 ( .A(net_3002), .Z(net_3003) );
CLKBUF_X2 inst_3827 ( .A(net_3618), .Z(net_3619) );
CLKBUF_X2 inst_4139 ( .A(net_3930), .Z(net_3931) );
CLKBUF_X2 inst_4112 ( .A(net_2721), .Z(net_3904) );
CLKBUF_X2 inst_3889 ( .A(net_3680), .Z(net_3681) );
SDFF_X2 inst_65 ( .Q(net_1569), .D(net_1569), .SE(net_498), .CK(net_2919), .SI(x6908) );
NOR2_X2 inst_536 ( .A1(net_1188), .ZN(net_1183), .A2(net_364) );
CLKBUF_X2 inst_3592 ( .A(net_3383), .Z(net_3384) );
AOI22_X2 inst_2386 ( .B1(net_1450), .B2(net_917), .ZN(net_631), .A1(net_630), .A2(net_476) );
NOR2_X4 inst_516 ( .A2(net_2086), .A1(net_1656), .ZN(net_1593) );
CLKBUF_X2 inst_3732 ( .A(net_2500), .Z(net_3524) );
AOI22_X2 inst_2258 ( .B2(net_2122), .A1(net_1967), .B1(net_1450), .ZN(net_1372), .A2(net_1198) );
OAI22_X2 inst_190 ( .B1(net_1402), .A1(net_775), .B2(net_389), .A2(net_113), .ZN(x1346) );
CLKBUF_X2 inst_4103 ( .A(net_3894), .Z(net_3895) );
INV_X4 inst_1267 ( .A(net_2371), .ZN(net_367) );
INV_X2 inst_1507 ( .A(net_2370), .ZN(net_282) );
DFF_X1 inst_2027 ( .QN(net_2219), .D(net_919), .CK(net_3282) );
CLKBUF_X2 inst_2926 ( .A(net_2641), .Z(net_2718) );
OAI21_X2 inst_416 ( .B1(net_768), .ZN(net_753), .A(net_628), .B2(net_441) );
INV_X8 inst_1158 ( .A(net_1848), .ZN(net_1789) );
DFF_X1 inst_1870 ( .D(net_1682), .QN(net_1587), .CK(net_3907) );
DFF_X1 inst_2062 ( .Q(net_2342), .D(net_432), .CK(net_3360) );
CLKBUF_X2 inst_3786 ( .A(net_3577), .Z(net_3578) );
AOI22_X2 inst_2350 ( .ZN(net_784), .A1(net_783), .B1(net_782), .A2(net_681), .B2(x3636) );
INV_X2 inst_1406 ( .A(net_570), .ZN(x1105) );
CLKBUF_X2 inst_3404 ( .A(net_3195), .Z(net_3196) );
NOR2_X2 inst_542 ( .A1(net_1725), .A2(net_1664), .ZN(net_1002) );
OR3_X2 inst_128 ( .A1(net_2247), .ZN(net_1121), .A2(x5143), .A3(x3145) );
AOI22_X2 inst_2445 ( .B2(net_2108), .ZN(net_2083), .A2(net_2076), .A1(net_2040), .B1(net_1450) );
CLKBUF_X2 inst_3039 ( .A(net_2830), .Z(net_2831) );
NAND2_X2 inst_973 ( .A2(net_1565), .A1(net_961), .ZN(net_866) );
CLKBUF_X2 inst_4000 ( .A(net_3791), .Z(net_3792) );
CLKBUF_X2 inst_3435 ( .A(net_3226), .Z(net_3227) );
CLKBUF_X2 inst_3058 ( .A(net_2849), .Z(net_2850) );
OAI211_X2 inst_461 ( .ZN(net_1055), .C1(net_1054), .A(net_903), .B(net_873), .C2(net_352) );
CLKBUF_X2 inst_3218 ( .A(net_2450), .Z(net_3010) );
NAND2_X2 inst_829 ( .A1(net_1745), .ZN(net_1286), .A2(net_363) );
OAI22_X2 inst_197 ( .B2(net_1906), .B1(net_1841), .A1(net_1836), .ZN(net_1243), .A2(net_395) );
CLKBUF_X2 inst_2958 ( .A(net_2749), .Z(net_2750) );
DFF_X1 inst_1973 ( .Q(net_2139), .D(net_1030), .CK(net_3157) );
CLKBUF_X2 inst_3089 ( .A(net_2663), .Z(net_2881) );
XNOR2_X2 inst_24 ( .ZN(net_1157), .B(net_1148), .A(net_932) );
CLKBUF_X2 inst_3051 ( .A(net_2842), .Z(net_2843) );
CLKBUF_X2 inst_2668 ( .A(net_2459), .Z(net_2460) );
NAND2_X1 inst_1122 ( .A2(net_1784), .A1(net_1660), .ZN(net_912) );
CLKBUF_X2 inst_3324 ( .A(net_3115), .Z(net_3116) );
INV_X4 inst_1209 ( .ZN(net_527), .A(net_515) );
OR2_X1 inst_150 ( .A1(net_2168), .A2(x3907), .ZN(x1314) );
INV_X2 inst_1611 ( .ZN(net_204), .A(x4899) );
NAND2_X2 inst_887 ( .ZN(net_1147), .A2(net_1143), .A1(net_322) );
CLKBUF_X2 inst_2981 ( .A(net_2772), .Z(net_2773) );
INV_X2 inst_1669 ( .ZN(net_1833), .A(x3190) );
INV_X2 inst_1663 ( .A(net_1754), .ZN(net_1753) );
CLKBUF_X2 inst_2714 ( .A(net_2505), .Z(net_2506) );
CLKBUF_X2 inst_3162 ( .A(net_2953), .Z(net_2954) );
CLKBUF_X2 inst_3956 ( .A(net_3747), .Z(net_3748) );
SDFF_X2 inst_90 ( .SE(net_487), .Q(net_159), .D(net_159), .CK(net_2813), .SI(x4690) );
AOI22_X2 inst_2357 ( .A1(net_783), .B1(net_775), .ZN(net_774), .A2(net_318), .B2(x3819) );
DFF_X2 inst_1801 ( .Q(net_1580), .CK(net_3027), .D(x5934) );
CLKBUF_X2 inst_3833 ( .A(net_3624), .Z(net_3625) );
NAND2_X4 inst_720 ( .A1(net_1687), .ZN(net_481), .A2(net_480) );
NAND2_X2 inst_958 ( .A2(net_2093), .A1(net_1829), .ZN(net_927) );
DFF_X1 inst_1961 ( .Q(net_2127), .D(net_1088), .CK(net_3523) );
AOI222_X2 inst_2460 ( .C1(net_2017), .A2(net_1563), .A1(net_590), .B1(net_589), .ZN(net_576), .B2(net_165), .C2(x5468) );
INV_X4 inst_1217 ( .A(net_2168), .ZN(net_782) );
OAI21_X2 inst_368 ( .B2(net_1443), .ZN(net_1421), .A(net_1383), .B1(net_1177) );
NAND2_X2 inst_1010 ( .ZN(net_913), .A1(net_659), .A2(net_268) );
INV_X16 inst_1697 ( .A(net_2102), .ZN(net_1935) );
NAND2_X2 inst_867 ( .A1(net_1838), .A2(net_1291), .ZN(net_1215) );
CLKBUF_X2 inst_3027 ( .A(net_2818), .Z(net_2819) );
NAND2_X2 inst_820 ( .A1(net_1840), .ZN(net_1343), .A2(net_345) );
CLKBUF_X2 inst_3689 ( .A(net_3480), .Z(net_3481) );
CLKBUF_X2 inst_3556 ( .A(net_3347), .Z(net_3348) );
OAI22_X2 inst_157 ( .B1(net_1427), .A1(net_529), .B2(net_221), .A2(net_97), .ZN(x1535) );
INV_X2 inst_1441 ( .A(net_1530), .ZN(net_726) );
CLKBUF_X2 inst_2929 ( .A(net_2520), .Z(net_2721) );
CLKBUF_X2 inst_3443 ( .A(net_3234), .Z(net_3235) );
CLKBUF_X2 inst_3568 ( .A(net_3359), .Z(net_3360) );
SDFF_X2 inst_68 ( .Q(net_1551), .D(net_1551), .SE(net_498), .CK(net_2680), .SI(x7369) );
DFF_X1 inst_1966 ( .Q(net_2132), .D(net_1063), .CK(net_3429) );
CLKBUF_X2 inst_3914 ( .A(net_3705), .Z(net_3706) );
INV_X4 inst_1253 ( .ZN(net_399), .A(net_82) );
CLKBUF_X2 inst_2793 ( .A(net_2584), .Z(net_2585) );
DFF_X1 inst_1884 ( .D(net_1323), .QN(net_88), .CK(net_3712) );
DFF_X1 inst_2018 ( .QN(net_2223), .D(net_1854), .CK(net_3062) );
AOI22_X2 inst_2435 ( .B2(net_2146), .B1(net_1974), .ZN(net_1809), .A1(net_1789), .A2(net_335) );
CLKBUF_X2 inst_4158 ( .A(net_2629), .Z(net_3950) );
INV_X2 inst_1643 ( .A(net_2353), .ZN(net_1198) );
CLKBUF_X2 inst_3410 ( .A(net_2729), .Z(net_3202) );
INV_X16 inst_1690 ( .A(net_1998), .ZN(net_1768) );
CLKBUF_X2 inst_2678 ( .A(net_2451), .Z(net_2470) );
DFFR_X1 inst_2120 ( .QN(net_2284), .D(net_1605), .RN(net_1347), .CK(net_3118) );
INV_X2 inst_1678 ( .A(net_1991), .ZN(net_1928) );
AND2_X2 inst_2613 ( .A1(net_609), .A2(x6908), .ZN(x638) );
XNOR2_X2 inst_17 ( .B(net_1196), .ZN(net_1185), .A(net_1172) );
OAI22_X2 inst_249 ( .B2(net_2270), .A1(net_745), .ZN(net_725), .A2(net_724), .B1(net_534) );
INV_X4 inst_1287 ( .A(net_2338), .ZN(net_1186) );
AOI22_X2 inst_2233 ( .A2(net_2370), .B2(net_2137), .A1(net_1738), .B1(net_1474), .ZN(net_1400) );
CLKBUF_X2 inst_4231 ( .A(net_4022), .Z(net_4023) );
CLKBUF_X2 inst_3866 ( .A(net_3220), .Z(net_3658) );
AOI22_X2 inst_2234 ( .B2(net_2133), .B1(net_1915), .ZN(net_1396), .A2(net_1367), .A1(net_1183) );
INV_X8 inst_1169 ( .ZN(net_1982), .A(net_1981) );
INV_X2 inst_1649 ( .A(net_2431), .ZN(net_267) );
CLKBUF_X2 inst_3483 ( .A(net_3274), .Z(net_3275) );
INV_X2 inst_1480 ( .A(net_2427), .ZN(net_356) );
OAI21_X2 inst_396 ( .B1(net_1829), .ZN(net_1111), .B2(net_949), .A(net_928) );
CLKBUF_X2 inst_3382 ( .A(net_3173), .Z(net_3174) );
CLKBUF_X2 inst_3377 ( .A(net_2980), .Z(net_3169) );
CLKBUF_X2 inst_2877 ( .A(net_2668), .Z(net_2669) );
NAND3_X2 inst_669 ( .A2(net_1795), .A1(net_1764), .ZN(net_1073), .A3(net_797) );
NAND3_X2 inst_664 ( .A2(net_1804), .ZN(net_1078), .A1(net_970), .A3(net_807) );
DFF_X1 inst_1918 ( .D(net_1837), .QN(net_113), .CK(net_3821) );
CLKBUF_X2 inst_2845 ( .A(net_2636), .Z(net_2637) );
INV_X2 inst_1418 ( .ZN(net_613), .A(net_612) );
DFF_X2 inst_1740 ( .QN(net_2365), .D(net_1481), .CK(net_3596) );
CLKBUF_X2 inst_2977 ( .A(net_2768), .Z(net_2769) );
NAND2_X2 inst_1092 ( .ZN(net_1899), .A1(net_1863), .A2(net_1747) );
CLKBUF_X2 inst_4064 ( .A(net_3855), .Z(net_3856) );
DFF_X1 inst_2001 ( .QN(net_2210), .D(net_1771), .CK(net_3333) );
INV_X2 inst_1657 ( .A(net_2274), .ZN(net_304) );
CLKBUF_X2 inst_3839 ( .A(net_3630), .Z(net_3631) );
DFF_X1 inst_1844 ( .QN(net_2340), .D(net_1480), .CK(net_3193) );
DFF_X1 inst_1913 ( .D(net_1317), .QN(net_129), .CK(net_3707) );
DFFR_X2 inst_2077 ( .QN(net_2414), .D(net_1925), .RN(net_1347), .CK(net_3947) );
AOI22_X2 inst_2368 ( .B2(net_2121), .A1(net_2038), .A2(net_1560), .B1(net_979), .ZN(net_688) );
DFF_X1 inst_1990 ( .Q(net_2154), .D(net_1027), .CK(net_3378) );
CLKBUF_X2 inst_2735 ( .A(net_2526), .Z(net_2527) );
XNOR2_X2 inst_36 ( .B(net_2320), .ZN(net_546), .A(net_505) );
CLKBUF_X2 inst_2934 ( .A(net_2559), .Z(net_2726) );
CLKBUF_X2 inst_2767 ( .A(net_2541), .Z(net_2559) );
INV_X2 inst_1370 ( .A(net_1014), .ZN(x2631) );
AOI221_X2 inst_2512 ( .B2(net_2138), .ZN(net_1947), .A(net_1946), .B1(net_1929), .C1(net_1863), .C2(net_302) );
OAI211_X2 inst_451 ( .C2(net_2363), .C1(net_1639), .ZN(net_1104), .A(net_825), .B(net_664) );
NAND2_X2 inst_797 ( .ZN(net_1316), .A1(net_1287), .A2(net_1229) );
INV_X2 inst_1495 ( .A(net_2332), .ZN(net_330) );
CLKBUF_X2 inst_4124 ( .A(net_3348), .Z(net_3916) );
CLKBUF_X2 inst_3067 ( .A(net_2858), .Z(net_2859) );
CLKBUF_X2 inst_3032 ( .A(net_2823), .Z(net_2824) );
CLKBUF_X2 inst_3657 ( .A(net_2625), .Z(net_3449) );
DFF_X1 inst_1998 ( .Q(net_2162), .D(net_1066), .CK(net_3488) );
CLKBUF_X2 inst_3302 ( .A(net_3093), .Z(net_3094) );
CLKBUF_X2 inst_2870 ( .A(net_2661), .Z(net_2662) );
NAND3_X2 inst_676 ( .A2(net_2169), .A3(net_1583), .ZN(net_604), .A1(net_603) );
CLKBUF_X2 inst_3583 ( .A(net_3374), .Z(net_3375) );
CLKBUF_X2 inst_3348 ( .A(net_2764), .Z(net_3140) );
NAND2_X2 inst_1115 ( .ZN(net_2069), .A1(net_2068), .A2(net_1220) );
CLKBUF_X2 inst_4222 ( .A(net_4013), .Z(net_4014) );
NAND2_X2 inst_874 ( .A1(net_1838), .ZN(net_1206), .A2(net_1205) );
CLKBUF_X2 inst_2976 ( .A(net_2767), .Z(net_2768) );
NAND2_X2 inst_1021 ( .A1(net_839), .ZN(net_549), .A2(net_76) );
INV_X2 inst_1681 ( .ZN(net_2051), .A(net_2049) );
INV_X16 inst_1684 ( .ZN(net_1052), .A(net_962) );
CLKBUF_X2 inst_4204 ( .A(net_3995), .Z(net_3996) );
INV_X2 inst_1386 ( .A(net_591), .ZN(x1253) );
AOI22_X2 inst_2255 ( .B2(net_2119), .A1(net_1967), .B1(net_1450), .ZN(net_1375), .A2(net_1201) );
INV_X2 inst_1652 ( .ZN(net_181), .A(x4998) );
OAI22_X2 inst_217 ( .A2(net_2240), .B1(net_1407), .A1(net_1405), .B2(net_232), .ZN(x1794) );
NAND2_X2 inst_1076 ( .A1(net_2104), .ZN(net_1817), .A2(net_1261) );
NOR2_X2 inst_572 ( .A2(net_2334), .A1(net_2328), .ZN(net_314) );
INV_X2 inst_1622 ( .A(net_2287), .ZN(net_319) );
DFF_X2 inst_1735 ( .QN(net_2315), .D(net_1496), .CK(net_3351) );
OAI22_X2 inst_257 ( .B2(net_2250), .A1(net_745), .ZN(net_708), .A2(net_707), .B1(net_534) );
DFF_X1 inst_2050 ( .Q(net_2387), .D(net_528), .CK(net_3368) );
DFF_X1 inst_2000 ( .Q(net_2164), .D(net_1091), .CK(net_3300) );
CLKBUF_X2 inst_3748 ( .A(net_3539), .Z(net_3540) );
AOI22_X2 inst_2213 ( .B2(net_2144), .A1(net_1916), .B1(net_1915), .ZN(net_1467), .A2(net_1160) );
OAI211_X2 inst_485 ( .C2(net_2316), .C1(net_1052), .ZN(net_1023), .A(net_879), .B(net_858) );
INV_X4 inst_1195 ( .A(net_2020), .ZN(net_614) );
NAND3_X2 inst_672 ( .A1(net_1993), .A2(net_1805), .ZN(net_1070), .A3(net_791) );
INV_X2 inst_1471 ( .A(net_1542), .ZN(net_749) );
CLKBUF_X2 inst_3826 ( .A(net_3617), .Z(net_3618) );
INV_X4 inst_1189 ( .ZN(net_1139), .A(net_1107) );
INV_X4 inst_1205 ( .ZN(net_1426), .A(net_1402) );
AOI22_X2 inst_2360 ( .A1(net_783), .B1(net_782), .ZN(net_770), .A2(net_373), .B2(x3699) );
INV_X2 inst_1525 ( .A(net_2360), .ZN(net_322) );
CLKBUF_X2 inst_3230 ( .A(net_3021), .Z(net_3022) );
AOI22_X2 inst_2248 ( .B2(net_2132), .A1(net_1967), .B1(net_1450), .ZN(net_1382), .A2(net_1196) );
AOI222_X2 inst_2453 ( .C1(net_2016), .A2(net_1570), .A1(net_590), .B1(net_589), .ZN(net_583), .B2(net_172), .C2(x5317) );
INV_X4 inst_1312 ( .A(net_1782), .ZN(net_1781) );
CLKBUF_X2 inst_3281 ( .A(net_2624), .Z(net_3073) );
NAND3_X2 inst_703 ( .ZN(net_2058), .A1(net_1799), .A3(net_800), .A2(net_654) );
XNOR2_X2 inst_33 ( .B(net_1845), .ZN(net_657), .A(net_599) );
DFFR_X1 inst_2107 ( .QN(net_2298), .D(net_1600), .RN(net_1347), .CK(net_2527) );
AOI21_X2 inst_2546 ( .ZN(net_535), .B1(net_511), .B2(net_423), .A(net_267) );
OAI22_X2 inst_232 ( .B2(net_2282), .B1(net_1865), .A1(net_1597), .ZN(net_942), .A2(net_703) );
CLKBUF_X2 inst_3419 ( .A(net_2663), .Z(net_3211) );
NAND2_X2 inst_1067 ( .A2(net_2035), .A1(net_1999), .ZN(net_1765) );
CLKBUF_X2 inst_3794 ( .A(net_3585), .Z(net_3586) );
DFF_X2 inst_1824 ( .Q(net_1534), .CK(net_2496), .D(x5507) );
CLKBUF_X2 inst_3716 ( .A(net_3507), .Z(net_3508) );
INV_X4 inst_1214 ( .A(net_2015), .ZN(net_1407) );
OAI22_X2 inst_253 ( .B2(net_2274), .A1(net_745), .ZN(net_717), .A2(net_716), .B1(net_534) );
NAND2_X2 inst_971 ( .A2(net_1563), .A1(net_961), .ZN(net_868) );
INV_X2 inst_1417 ( .A(net_559), .ZN(x1230) );
INV_X4 inst_1219 ( .ZN(net_500), .A(net_470) );
CLKBUF_X2 inst_3652 ( .A(net_3443), .Z(net_3444) );
NOR2_X2 inst_589 ( .A2(net_2277), .ZN(net_1878), .A1(net_520) );
CLKBUF_X2 inst_3459 ( .A(net_3250), .Z(net_3251) );
NOR2_X2 inst_602 ( .A2(net_2269), .ZN(net_1891), .A1(net_520) );
SDFF_X2 inst_59 ( .Q(net_1567), .D(net_1567), .SE(net_498), .CK(net_2931), .SI(x6968) );
DFF_X1 inst_1877 ( .D(net_1329), .QN(net_87), .CK(net_3933) );
AOI22_X2 inst_2367 ( .B2(net_2126), .A1(net_2038), .A2(net_1556), .B1(net_979), .ZN(net_689) );
OR2_X2 inst_135 ( .A1(net_2416), .A2(net_1904), .ZN(net_468) );
CLKBUF_X2 inst_3335 ( .A(net_3126), .Z(net_3127) );
CLKBUF_X2 inst_3256 ( .A(net_2462), .Z(net_3048) );
CLKBUF_X2 inst_3073 ( .A(net_2864), .Z(net_2865) );
DFF_X1 inst_1865 ( .D(net_1357), .QN(net_97), .CK(net_3657) );
XNOR2_X2 inst_37 ( .B(net_1222), .ZN(net_540), .A(net_526) );
DFF_X1 inst_1980 ( .Q(net_2145), .D(net_1041), .CK(net_3233) );
INV_X2 inst_1664 ( .A(net_1756), .ZN(net_1755) );
INV_X2 inst_1447 ( .A(net_1533), .ZN(net_949) );
CLKBUF_X2 inst_3117 ( .A(net_2908), .Z(net_2909) );
CLKBUF_X2 inst_2885 ( .A(net_2676), .Z(net_2677) );
AND2_X2 inst_2632 ( .A1(net_609), .A2(x7241), .ZN(x781) );
AOI22_X2 inst_2221 ( .B2(net_2146), .A1(net_1916), .B1(net_1915), .ZN(net_1459), .A2(net_1174) );
CLKBUF_X2 inst_3770 ( .A(net_3561), .Z(net_3562) );
DFFR_X2 inst_2082 ( .QN(net_1748), .RN(net_1347), .D(net_1137), .CK(net_3915) );
CLKBUF_X2 inst_3286 ( .A(net_3077), .Z(net_3078) );
CLKBUF_X2 inst_4225 ( .A(net_2809), .Z(net_4017) );
CLKBUF_X2 inst_2709 ( .A(net_2463), .Z(net_2501) );
OAI22_X2 inst_224 ( .B2(net_2296), .B1(net_1865), .ZN(net_954), .A2(net_953), .A1(net_951) );
CLKBUF_X2 inst_3635 ( .A(net_2770), .Z(net_3427) );
CLKBUF_X2 inst_3075 ( .A(net_2739), .Z(net_2867) );
CLKBUF_X2 inst_2800 ( .A(net_2528), .Z(net_2592) );
AOI22_X2 inst_2406 ( .B1(net_2197), .ZN(net_1634), .A1(net_1621), .B2(net_1538), .A2(net_1197) );
NAND2_X4 inst_766 ( .ZN(net_2100), .A2(net_1914), .A1(net_1731) );
CLKBUF_X2 inst_4141 ( .A(net_3932), .Z(net_3933) );
CLKBUF_X2 inst_3270 ( .A(net_3061), .Z(net_3062) );
DFF_X1 inst_1908 ( .D(net_1313), .QN(net_133), .CK(net_3445) );
CLKBUF_X2 inst_3273 ( .A(net_3064), .Z(net_3065) );
NAND2_X2 inst_801 ( .ZN(net_1312), .A1(net_1272), .A2(net_1236) );
NAND3_X2 inst_692 ( .A2(net_2428), .A3(net_2423), .ZN(net_1773), .A1(net_301) );
INV_X2 inst_1517 ( .A(net_2243), .ZN(net_275) );
SDFF_X2 inst_70 ( .Q(net_1559), .D(net_1559), .SE(net_396), .CK(net_2675), .SI(x7190) );
NAND2_X2 inst_870 ( .A1(net_1838), .A2(net_1238), .ZN(net_1211) );
XOR2_X1 inst_11 ( .Z(net_2184), .B(net_2105), .A(net_1649) );
OAI22_X2 inst_188 ( .B1(net_1402), .A1(net_529), .B2(net_178), .A2(net_86), .ZN(x1693) );
CLKBUF_X2 inst_3768 ( .A(net_3248), .Z(net_3560) );
INV_X2 inst_1619 ( .ZN(net_302), .A(net_57) );
CLKBUF_X2 inst_4207 ( .A(net_3998), .Z(net_3999) );
CLKBUF_X2 inst_3110 ( .A(net_2871), .Z(net_2902) );
OAI21_X1 inst_441 ( .B2(net_1579), .ZN(net_1252), .B1(net_1250), .A(net_602) );
CLKBUF_X2 inst_3011 ( .A(net_2546), .Z(net_2803) );
AOI22_X2 inst_2276 ( .ZN(net_1695), .A2(net_1553), .A1(net_1000), .B1(net_999), .B2(net_377) );
CLKBUF_X2 inst_2848 ( .A(net_2639), .Z(net_2640) );
AOI22_X2 inst_2301 ( .A2(net_2150), .B1(net_2096), .A1(net_1769), .B2(net_1524), .ZN(net_908) );
NAND2_X2 inst_808 ( .A2(net_1670), .ZN(net_1305), .A1(net_1282) );
INV_X2 inst_1537 ( .A(net_2305), .ZN(net_329) );
NOR2_X2 inst_557 ( .A2(net_2246), .ZN(net_524), .A1(net_461) );
DFF_X1 inst_2041 ( .Q(net_2389), .D(net_649), .CK(net_3557) );
CLKBUF_X2 inst_3859 ( .A(net_3650), .Z(net_3651) );
CLKBUF_X2 inst_3593 ( .A(net_3157), .Z(net_3385) );
INV_X2 inst_1383 ( .ZN(net_635), .A(net_634) );
CLKBUF_X2 inst_3279 ( .A(net_3042), .Z(net_3071) );
NAND2_X2 inst_823 ( .A1(net_1840), .ZN(net_1337), .A2(net_368) );
INV_X2 inst_1461 ( .ZN(net_1056), .A(net_369) );
CLKBUF_X2 inst_2838 ( .A(net_2629), .Z(net_2630) );
CLKBUF_X2 inst_3773 ( .A(net_3564), .Z(net_3565) );
CLKBUF_X2 inst_3423 ( .A(net_3214), .Z(net_3215) );
CLKBUF_X2 inst_3176 ( .A(net_2967), .Z(net_2968) );
CLKBUF_X2 inst_2833 ( .A(net_2624), .Z(net_2625) );
DFF_X1 inst_2042 ( .QN(net_2408), .D(net_679), .CK(net_3965) );
CLKBUF_X2 inst_3325 ( .A(net_3116), .Z(net_3117) );
CLKBUF_X2 inst_4168 ( .A(net_3959), .Z(net_3960) );
OAI22_X2 inst_195 ( .A2(net_2367), .B2(net_1911), .B1(net_1841), .A1(net_1836), .ZN(net_1245) );
DFF_X1 inst_1987 ( .Q(net_2151), .D(net_1046), .CK(net_2970) );
CLKBUF_X2 inst_2796 ( .A(net_2587), .Z(net_2588) );
INV_X8 inst_1150 ( .A(net_1865), .ZN(net_1603) );
CLKBUF_X2 inst_2729 ( .A(net_2520), .Z(net_2521) );
INV_X2 inst_1413 ( .A(net_563), .ZN(x1207) );
DFF_X2 inst_1815 ( .Q(net_1516), .CK(net_2556), .D(x5796) );
CLKBUF_X2 inst_3993 ( .A(net_3784), .Z(net_3785) );
INV_X2 inst_1589 ( .ZN(net_220), .A(x4089) );
INV_X4 inst_1326 ( .ZN(net_1958), .A(net_1957) );
OAI21_X2 inst_335 ( .B2(net_2320), .B1(net_2041), .ZN(net_1495), .A(net_1458) );
CLKBUF_X2 inst_3875 ( .A(net_3666), .Z(net_3667) );
AND2_X2 inst_2629 ( .A1(net_594), .A2(x7466), .ZN(x878) );
NAND3_X2 inst_658 ( .A1(net_2063), .A2(net_1806), .ZN(net_1133), .A3(net_814) );
OAI21_X2 inst_438 ( .ZN(net_2045), .B2(net_1586), .B1(net_592), .A(net_403) );
INV_X4 inst_1341 ( .ZN(net_2070), .A(net_1748) );
DFFR_X1 inst_2154 ( .QN(net_2271), .RN(net_1347), .D(net_723), .CK(net_2747) );
NOR2_X2 inst_587 ( .A2(net_2266), .ZN(net_1876), .A1(net_520) );
NAND3_X2 inst_666 ( .A2(net_1802), .ZN(net_1076), .A1(net_969), .A3(net_805) );
AND2_X4 inst_2602 ( .A1(net_2378), .A2(net_2377), .ZN(net_2200) );
OAI21_X2 inst_324 ( .B2(net_2323), .A(net_1857), .B1(net_1507), .ZN(net_1506) );
DFF_X2 inst_1829 ( .Q(net_1531), .CK(net_2493), .D(x5468) );
CLKBUF_X2 inst_3550 ( .A(net_3341), .Z(net_3342) );
SDFF_X2 inst_109 ( .SE(net_488), .Q(net_166), .D(net_166), .CK(net_2733), .SI(x4502) );
INV_X4 inst_1182 ( .ZN(net_1441), .A(net_1367) );
CLKBUF_X2 inst_4083 ( .A(net_3474), .Z(net_3875) );
CLKBUF_X2 inst_3983 ( .A(net_3774), .Z(net_3775) );
XNOR2_X1 inst_43 ( .ZN(net_1654), .A(net_1653), .B(net_369) );
DFFR_X1 inst_2128 ( .QN(net_2258), .RN(net_1347), .D(net_750), .CK(net_2840) );
INV_X1 inst_1707 ( .A(net_1785), .ZN(net_1784) );
INV_X2 inst_1444 ( .A(net_1517), .ZN(net_941) );
INV_X4 inst_1231 ( .ZN(net_442), .A(net_405) );
OAI21_X2 inst_375 ( .A(net_1759), .B1(net_1744), .ZN(net_1414), .B2(net_399) );
CLKBUF_X2 inst_3490 ( .A(net_3281), .Z(net_3282) );
NAND2_X2 inst_904 ( .A1(net_1760), .ZN(net_1115), .A2(net_328) );
CLKBUF_X2 inst_3315 ( .A(net_3106), .Z(net_3107) );
OAI22_X2 inst_285 ( .A2(net_2442), .A1(net_1615), .B1(net_1407), .B2(net_454), .ZN(x51) );
DFF_X2 inst_1830 ( .QN(net_1757), .Q(net_1659), .CK(net_3123), .D(x6592) );
CLKBUF_X2 inst_3923 ( .A(net_3714), .Z(net_3715) );
NAND2_X4 inst_757 ( .A1(net_2050), .ZN(net_2020), .A2(net_1905) );
OAI21_X2 inst_343 ( .ZN(net_1487), .B2(net_1484), .A(net_1448), .B1(net_1253) );
INV_X2 inst_1627 ( .ZN(net_194), .A(x6439) );
INV_X2 inst_1563 ( .ZN(net_237), .A(x4435) );
NOR2_X2 inst_543 ( .A2(net_2358), .ZN(net_914), .A1(net_913) );
NAND2_X2 inst_1106 ( .ZN(net_2018), .A1(net_2012), .A2(net_399) );
CLKBUF_X2 inst_3242 ( .A(net_3033), .Z(net_3034) );
CLKBUF_X2 inst_3817 ( .A(net_3608), .Z(net_3609) );
CLKBUF_X2 inst_3138 ( .A(net_2929), .Z(net_2930) );
NAND2_X2 inst_982 ( .A2(net_1552), .A1(net_961), .ZN(net_857) );
NAND2_X2 inst_929 ( .A2(net_1633), .ZN(net_1085), .A1(net_830) );
DFFR_X2 inst_2070 ( .QN(net_1592), .RN(net_1347), .D(net_1249), .CK(net_3952) );
INV_X2 inst_1397 ( .A(net_578), .ZN(x1195) );
INV_X4 inst_1256 ( .A(net_2205), .ZN(net_405) );
CLKBUF_X2 inst_2890 ( .A(net_2681), .Z(net_2682) );
OAI22_X2 inst_299 ( .A2(net_2241), .B1(net_1895), .A1(net_1615), .B2(net_216), .ZN(x1768) );
DFF_X2 inst_1798 ( .QN(net_2311), .D(net_382), .CK(net_3992) );
CLKBUF_X2 inst_2927 ( .A(net_2508), .Z(net_2719) );
CLKBUF_X2 inst_3303 ( .A(net_3094), .Z(net_3095) );
DFF_X1 inst_1903 ( .D(net_1303), .QN(net_119), .CK(net_3570) );
CLKBUF_X2 inst_2760 ( .A(net_2551), .Z(net_2552) );
DFF_X1 inst_1938 ( .Q(net_2398), .D(net_1117), .CK(net_3071) );
AOI21_X2 inst_2554 ( .ZN(net_1853), .B1(net_1852), .A(net_1849), .B2(net_48) );
CLKBUF_X2 inst_2745 ( .A(net_2536), .Z(net_2537) );
DFFR_X1 inst_2095 ( .RN(net_1347), .D(net_1135), .QN(net_47), .CK(net_3548) );
AND2_X2 inst_2604 ( .A1(net_2195), .ZN(net_622), .A2(net_376) );
INV_X4 inst_1244 ( .A(net_2316), .ZN(net_1259) );
CLKBUF_X2 inst_3260 ( .A(net_3051), .Z(net_3052) );
CLKBUF_X2 inst_3248 ( .A(net_3039), .Z(net_3040) );
CLKBUF_X2 inst_4190 ( .A(net_3981), .Z(net_3982) );
CLKBUF_X2 inst_3158 ( .A(net_2949), .Z(net_2950) );
NOR2_X2 inst_582 ( .ZN(net_1774), .A2(net_523), .A1(net_348) );
NAND3_X2 inst_683 ( .ZN(net_430), .A1(net_351), .A3(net_272), .A2(net_269) );
CLKBUF_X2 inst_3269 ( .A(net_3060), .Z(net_3061) );
DFF_X1 inst_1944 ( .Q(net_2110), .D(net_1050), .CK(net_3191) );
OAI22_X2 inst_210 ( .A2(net_2216), .A1(net_1408), .B1(net_1407), .B2(net_246), .ZN(x2289) );
CLKBUF_X2 inst_3101 ( .A(net_2554), .Z(net_2893) );
DFFR_X1 inst_2110 ( .QN(net_2301), .D(net_1609), .RN(net_1347), .CK(net_2760) );
DFF_X1 inst_1850 ( .QN(net_2369), .D(net_1444), .CK(net_3616) );
CLKBUF_X2 inst_3477 ( .A(net_3268), .Z(net_3269) );
DFF_X1 inst_1950 ( .Q(net_2116), .D(net_1092), .CK(net_3542) );
CLKBUF_X2 inst_3881 ( .A(net_3672), .Z(net_3673) );
INV_X4 inst_1294 ( .ZN(net_794), .A(net_63) );
HA_X1 inst_1712 ( .B(net_1259), .CO(net_596), .S(net_528), .A(net_473) );
DFF_X1 inst_2057 ( .D(net_493), .CK(net_4025), .Q(x0) );
CLKBUF_X2 inst_3108 ( .A(net_2899), .Z(net_2900) );
NAND2_X4 inst_747 ( .ZN(net_1970), .A2(net_1969), .A1(net_1968) );
NAND2_X2 inst_843 ( .A1(net_1840), .ZN(net_1270), .A2(net_280) );
CLKBUF_X2 inst_3806 ( .A(net_3597), .Z(net_3598) );
CLKBUF_X2 inst_2853 ( .A(net_2608), .Z(net_2645) );
DFF_X2 inst_1779 ( .QN(net_2424), .D(net_758), .CK(net_3667) );
DFFR_X1 inst_2115 ( .QN(net_2306), .D(net_1608), .RN(net_1347), .CK(net_2477) );
CLKBUF_X2 inst_3251 ( .A(net_3042), .Z(net_3043) );
SDFF_X2 inst_112 ( .SE(net_487), .Q(net_151), .D(net_151), .CK(net_2531), .SI(x4926) );
DFF_X2 inst_1728 ( .QN(net_2323), .D(net_1506), .CK(net_3129) );
CLKBUF_X2 inst_2775 ( .A(net_2528), .Z(net_2567) );
NAND2_X2 inst_916 ( .A1(net_974), .A2(net_777), .ZN(x2993) );
DFF_X2 inst_1722 ( .QN(net_2329), .D(net_1492), .CK(net_2983) );
OAI22_X2 inst_305 ( .A2(net_2222), .B1(net_1895), .A1(net_1405), .B2(net_200), .ZN(x2175) );
INV_X2 inst_1595 ( .ZN(net_215), .A(x4629) );
CLKBUF_X2 inst_3665 ( .A(net_3456), .Z(net_3457) );
CLKBUF_X2 inst_2724 ( .A(net_2515), .Z(net_2516) );
AOI21_X2 inst_2525 ( .A(net_1785), .B1(net_910), .ZN(net_808), .B2(net_72) );
CLKBUF_X2 inst_2968 ( .A(net_2759), .Z(net_2760) );
CLKBUF_X2 inst_2964 ( .A(net_2494), .Z(net_2756) );
CLKBUF_X2 inst_3721 ( .A(net_3512), .Z(net_3513) );
AOI22_X2 inst_2349 ( .ZN(net_785), .A1(net_783), .B1(net_782), .A2(net_356), .B2(x3651) );
NAND3_X4 inst_646 ( .A3(net_2168), .ZN(net_1994), .A1(net_1901), .A2(net_82) );
CLKBUF_X2 inst_4032 ( .A(net_3823), .Z(net_3824) );
CLKBUF_X2 inst_3169 ( .A(net_2960), .Z(net_2961) );
NAND2_X2 inst_963 ( .A2(net_1555), .A1(net_961), .ZN(net_877) );
OAI21_X2 inst_382 ( .A(net_1937), .B2(net_1356), .ZN(net_1354), .B1(net_1333) );
AOI22_X2 inst_2329 ( .ZN(net_841), .A1(net_840), .B1(net_839), .A2(net_447), .B2(net_79) );
NAND2_X2 inst_907 ( .A1(net_977), .A2(net_770), .ZN(x2928) );
NAND2_X2 inst_922 ( .A2(net_1636), .ZN(net_1092), .A1(net_694) );
INV_X2 inst_1614 ( .ZN(net_202), .A(x5078) );
INV_X2 inst_1502 ( .A(net_2354), .ZN(net_1222) );
CLKBUF_X2 inst_2788 ( .A(net_2579), .Z(net_2580) );
CLKBUF_X2 inst_4091 ( .A(net_3882), .Z(net_3883) );
NAND2_X2 inst_1049 ( .A1(net_1746), .ZN(net_1676), .A2(net_1201) );
CLKBUF_X2 inst_3907 ( .A(net_3698), .Z(net_3699) );
OAI22_X2 inst_168 ( .A1(net_2013), .B1(net_1406), .B2(net_185), .A2(net_122), .ZN(x476) );
INV_X2 inst_1568 ( .A(net_2286), .ZN(net_337) );
CLKBUF_X2 inst_3692 ( .A(net_3483), .Z(net_3484) );
CLKBUF_X2 inst_3366 ( .A(net_2926), .Z(net_3158) );
NAND2_X2 inst_873 ( .A1(net_1838), .ZN(net_1208), .A2(net_1207) );
NAND2_X2 inst_991 ( .A1(net_1596), .A2(net_958), .ZN(net_850) );
NAND3_X2 inst_653 ( .A2(net_2003), .ZN(net_1192), .A1(net_611), .A3(net_512) );
CLKBUF_X2 inst_3767 ( .A(net_3558), .Z(net_3559) );
NOR2_X2 inst_580 ( .A2(net_2367), .ZN(net_1734), .A1(net_1151) );
OAI22_X2 inst_170 ( .B1(net_1406), .A1(net_1405), .B2(net_258), .A2(net_120), .ZN(x499) );
DFF_X2 inst_1746 ( .QN(net_2360), .D(net_1416), .CK(net_3872) );
CLKBUF_X2 inst_3691 ( .A(net_3482), .Z(net_3483) );
CLKBUF_X2 inst_3371 ( .A(net_3162), .Z(net_3163) );
CLKBUF_X2 inst_3052 ( .A(net_2843), .Z(net_2844) );
CLKBUF_X2 inst_3649 ( .A(net_3440), .Z(net_3441) );
DFF_X1 inst_1857 ( .QN(net_2437), .D(net_1414), .CK(net_3847) );
CLKBUF_X2 inst_2907 ( .A(net_2698), .Z(net_2699) );
CLKBUF_X2 inst_4072 ( .A(net_3863), .Z(net_3864) );
CLKBUF_X2 inst_2656 ( .A(net_2447), .Z(net_2448) );
CLKBUF_X2 inst_3000 ( .A(net_2791), .Z(net_2792) );
INV_X8 inst_1163 ( .A(net_1959), .ZN(net_1916) );
OAI211_X2 inst_468 ( .C2(net_2320), .C1(net_1052), .ZN(net_1043), .A(net_886), .B(net_855) );
NAND2_X2 inst_1099 ( .ZN(net_1952), .A2(net_1951), .A1(net_1949) );
CLKBUF_X2 inst_3616 ( .A(net_3407), .Z(net_3408) );
INV_X2 inst_1604 ( .A(net_2301), .ZN(net_339) );
CLKBUF_X2 inst_3239 ( .A(net_3030), .Z(net_3031) );
AOI22_X2 inst_2314 ( .A2(net_2111), .B1(net_2096), .A1(net_1769), .B2(net_1519), .ZN(net_895) );
OAI21_X2 inst_429 ( .B1(net_1977), .A(net_1904), .ZN(net_1668), .B2(net_358) );
CLKBUF_X2 inst_2692 ( .A(net_2483), .Z(net_2484) );
INV_X2 inst_1599 ( .ZN(net_211), .A(x6389) );
CLKBUF_X2 inst_2812 ( .A(net_2603), .Z(net_2604) );
CLKBUF_X2 inst_3565 ( .A(net_3356), .Z(net_3357) );
CLKBUF_X2 inst_3197 ( .A(net_2988), .Z(net_2989) );
XOR2_X1 inst_7 ( .Z(net_2180), .B(net_1227), .A(net_1151) );
CLKBUF_X2 inst_3977 ( .A(net_3768), .Z(net_3769) );
CLKBUF_X2 inst_3450 ( .A(net_3241), .Z(net_3242) );
CLKBUF_X2 inst_3467 ( .A(net_3258), .Z(net_3259) );
AND2_X4 inst_2593 ( .ZN(net_2166), .A2(net_1747), .A1(net_1726) );
CLKBUF_X2 inst_3064 ( .A(net_2491), .Z(net_2856) );
CLKBUF_X2 inst_3676 ( .A(net_3418), .Z(net_3468) );
NAND2_X2 inst_1083 ( .A1(net_1934), .ZN(net_1824), .A2(net_1217) );
CLKBUF_X2 inst_4073 ( .A(net_3417), .Z(net_3865) );
OAI21_X2 inst_318 ( .B2(net_2327), .B1(net_2041), .ZN(net_1512), .A(net_1477) );
CLKBUF_X2 inst_4033 ( .A(net_3824), .Z(net_3825) );
INV_X8 inst_1136 ( .A(net_1865), .ZN(net_951) );
AOI222_X2 inst_2466 ( .C1(net_2017), .A2(net_1558), .A1(net_590), .B1(net_589), .ZN(net_570), .B2(net_160), .C2(x5581) );
CLKBUF_X2 inst_2899 ( .A(net_2690), .Z(net_2691) );
CLKBUF_X2 inst_4065 ( .A(net_2829), .Z(net_3857) );
INV_X2 inst_1486 ( .A(net_2346), .ZN(net_934) );
AOI22_X2 inst_2281 ( .B1(net_1768), .ZN(net_1710), .A2(net_1552), .B2(net_1513), .A1(net_1000) );
NAND3_X2 inst_696 ( .A1(net_2100), .ZN(net_1934), .A3(net_1812), .A2(net_1760) );
INV_X8 inst_1175 ( .ZN(net_2038), .A(net_2037) );
CLKBUF_X2 inst_3311 ( .A(net_3102), .Z(net_3103) );
CLKBUF_X2 inst_4096 ( .A(net_3887), .Z(net_3888) );
OAI21_X2 inst_395 ( .B1(net_1829), .ZN(net_1112), .B2(net_950), .A(net_929) );
NAND2_X2 inst_841 ( .A1(net_1840), .ZN(net_1272), .A2(net_330) );
CLKBUF_X2 inst_3963 ( .A(net_3754), .Z(net_3755) );
NAND3_X2 inst_689 ( .A3(net_1733), .ZN(net_1723), .A1(net_1657), .A2(net_987) );
CLKBUF_X2 inst_3969 ( .A(net_3760), .Z(net_3761) );
AOI22_X2 inst_2363 ( .B2(net_2116), .A1(net_2038), .A2(net_1547), .B1(net_979), .ZN(net_694) );
CLKBUF_X2 inst_2689 ( .A(net_2480), .Z(net_2481) );
CLKBUF_X2 inst_4029 ( .A(net_3820), .Z(net_3821) );
INV_X2 inst_1629 ( .ZN(net_192), .A(x4107) );
CLKBUF_X2 inst_3896 ( .A(net_3687), .Z(net_3688) );
INV_X2 inst_1558 ( .ZN(net_242), .A(x4353) );
CLKBUF_X2 inst_3679 ( .A(net_3275), .Z(net_3471) );
CLKBUF_X2 inst_2906 ( .A(net_2697), .Z(net_2698) );
CLKBUF_X2 inst_3424 ( .A(net_2729), .Z(net_3216) );
CLKBUF_X2 inst_3886 ( .A(net_3677), .Z(net_3678) );
INV_X2 inst_1615 ( .ZN(net_201), .A(x4206) );
AND2_X4 inst_2580 ( .A2(net_2418), .A1(net_1872), .ZN(net_429) );
CLKBUF_X2 inst_3713 ( .A(net_3504), .Z(net_3505) );
AOI22_X2 inst_2394 ( .B1(net_2197), .ZN(net_1622), .A1(net_1621), .B2(net_1533), .A2(net_322) );
DFFR_X1 inst_2145 ( .QN(net_2251), .RN(net_1347), .D(net_704), .CK(net_2643) );
NAND3_X1 inst_709 ( .A2(net_1953), .ZN(net_1733), .A3(net_1719), .A1(net_1561) );
AOI22_X2 inst_2375 ( .B2(net_2133), .B1(net_1929), .ZN(net_656), .A1(net_655), .A2(net_293) );
NAND2_X2 inst_920 ( .A1(net_1641), .ZN(net_1097), .A2(net_820) );
CLKBUF_X2 inst_3454 ( .A(net_2817), .Z(net_3246) );
DFF_X1 inst_2054 ( .QN(net_2400), .D(net_504), .CK(net_3785) );
INV_X4 inst_1259 ( .A(net_2320), .ZN(net_345) );
DFF_X2 inst_1796 ( .QN(net_2376), .D(net_467), .CK(net_3850) );
NOR2_X2 inst_535 ( .A1(net_1840), .ZN(net_1255), .A2(net_638) );
CLKBUF_X2 inst_2889 ( .A(net_2505), .Z(net_2681) );
INV_X2 inst_1670 ( .ZN(net_1845), .A(net_1843) );
AOI22_X2 inst_2427 ( .B2(net_2147), .B1(net_1974), .ZN(net_1801), .A1(net_1791), .A2(net_339) );
CLKBUF_X2 inst_4198 ( .A(net_2813), .Z(net_3990) );
OAI21_X4 inst_315 ( .A(net_2416), .B2(net_1872), .B1(net_1712), .ZN(net_480) );
CLKBUF_X2 inst_2935 ( .A(net_2726), .Z(net_2727) );
OAI22_X2 inst_216 ( .A2(net_2219), .B1(net_1407), .A1(net_1403), .B2(net_256), .ZN(x2233) );
CLKBUF_X2 inst_3317 ( .A(net_3108), .Z(net_3109) );
CLKBUF_X2 inst_3369 ( .A(net_3160), .Z(net_3161) );
CLKBUF_X2 inst_3113 ( .A(net_2904), .Z(net_2905) );
DFF_X1 inst_2060 ( .QN(net_2373), .D(net_2185), .CK(net_4020) );
CLKBUF_X2 inst_3695 ( .A(net_2974), .Z(net_3487) );
CLKBUF_X2 inst_2680 ( .A(net_2471), .Z(net_2472) );
CLKBUF_X2 inst_3168 ( .A(net_2485), .Z(net_2960) );
AOI22_X2 inst_2336 ( .B2(net_2134), .A1(net_2038), .A2(net_1568), .B1(net_979), .ZN(net_828) );
AOI22_X2 inst_2385 ( .B1(net_1450), .B2(net_909), .ZN(net_636), .A1(net_630), .A2(net_436) );
OAI21_X2 inst_415 ( .B1(net_768), .ZN(net_754), .A(net_648), .B2(net_318) );
CLKBUF_X2 inst_3855 ( .A(net_3646), .Z(net_3647) );
DFF_X2 inst_1795 ( .QN(net_2243), .D(net_452), .CK(net_2820) );
NAND2_X2 inst_828 ( .A2(net_2066), .A1(net_1840), .ZN(net_1287) );
CLKBUF_X2 inst_3318 ( .A(net_3109), .Z(net_3110) );
OAI22_X2 inst_223 ( .B2(net_2295), .B1(net_1865), .A1(net_1597), .ZN(net_955), .A2(net_735) );
CLKBUF_X2 inst_4164 ( .A(net_3955), .Z(net_3956) );
AOI22_X2 inst_2420 ( .B2(net_2155), .B1(net_1974), .ZN(net_1794), .A1(net_1791), .A2(net_292) );
INV_X2 inst_1561 ( .ZN(net_239), .A(x6289) );
CLKBUF_X2 inst_3564 ( .A(net_3355), .Z(net_3356) );
DFFR_X1 inst_2104 ( .QN(net_2294), .D(net_1602), .RN(net_1347), .CK(net_2846) );
CLKBUF_X2 inst_4205 ( .A(net_3922), .Z(net_3997) );
INV_X4 inst_1322 ( .A(net_2053), .ZN(net_1901) );
AND4_X2 inst_2573 ( .A2(net_2050), .ZN(net_1910), .A3(net_1909), .A1(net_522), .A4(net_397) );
DFFR_X1 inst_2096 ( .Q(net_2165), .RN(net_1347), .D(net_1109), .CK(net_3119) );
NOR2_X2 inst_552 ( .A1(net_1971), .A2(net_621), .ZN(net_600) );
CLKBUF_X2 inst_3050 ( .A(net_2841), .Z(net_2842) );
CLKBUF_X2 inst_3493 ( .A(net_3284), .Z(net_3285) );
CLKBUF_X2 inst_3019 ( .A(net_2810), .Z(net_2811) );
AOI22_X2 inst_2327 ( .A2(net_2156), .B1(net_2096), .A1(net_1769), .B2(net_1515), .ZN(net_875) );
CLKBUF_X2 inst_3913 ( .A(net_3704), .Z(net_3705) );
INV_X2 inst_1564 ( .ZN(net_236), .A(x4066) );
CLKBUF_X2 inst_3487 ( .A(net_3278), .Z(net_3279) );
CLKBUF_X2 inst_3597 ( .A(net_3388), .Z(net_3389) );
DFF_X1 inst_1941 ( .Q(net_2107), .D(net_1024), .CK(net_3070) );
AND2_X2 inst_2607 ( .A1(net_609), .A2(x7509), .ZN(x894) );
SDFF_X2 inst_113 ( .SE(net_487), .Q(net_172), .D(net_172), .CK(net_2703), .SI(x4375) );
XOR2_X1 inst_9 ( .Z(net_2182), .B(net_1239), .A(net_541) );
OAI21_X2 inst_356 ( .B2(net_2399), .B1(net_1443), .ZN(net_1438), .A(net_1377) );
CLKBUF_X2 inst_3358 ( .A(net_3149), .Z(net_3150) );
CLKBUF_X2 inst_2690 ( .A(net_2453), .Z(net_2482) );
INV_X2 inst_1594 ( .ZN(net_216), .A(x4303) );
NAND2_X2 inst_902 ( .A1(net_1648), .A2(net_1645), .ZN(net_1117) );
CLKBUF_X2 inst_3489 ( .A(net_2499), .Z(net_3281) );
NAND2_X2 inst_778 ( .ZN(net_1349), .A2(net_1295), .A1(net_1270) );
INV_X2 inst_1544 ( .A(net_2284), .ZN(net_316) );
DFF_X1 inst_1935 ( .D(net_1123), .QN(net_65), .CK(net_3495) );
CLKBUF_X2 inst_4063 ( .A(net_3101), .Z(net_3855) );
AND2_X2 inst_2625 ( .A1(net_609), .A2(x7484), .ZN(x886) );
CLKBUF_X2 inst_3148 ( .A(net_2939), .Z(net_2940) );
DFFR_X1 inst_2140 ( .QN(net_2273), .RN(net_1347), .D(net_719), .CK(net_2473) );
CLKBUF_X2 inst_3329 ( .A(net_2645), .Z(net_3121) );
NAND2_X2 inst_781 ( .A1(net_2106), .ZN(net_1332), .A2(net_1223) );
CLKBUF_X2 inst_4042 ( .A(net_3833), .Z(net_3834) );
CLKBUF_X2 inst_3026 ( .A(net_2468), .Z(net_2818) );
CLKBUF_X2 inst_3696 ( .A(net_3487), .Z(net_3488) );
INV_X2 inst_1442 ( .A(net_1531), .ZN(net_728) );
CLKBUF_X2 inst_2847 ( .A(net_2638), .Z(net_2639) );
OAI21_X2 inst_332 ( .B2(net_2319), .B1(net_2041), .ZN(net_1498), .A(net_1460) );
CLKBUF_X2 inst_3639 ( .A(net_3430), .Z(net_3431) );
INV_X4 inst_1289 ( .A(net_2356), .ZN(net_1197) );
DFFR_X1 inst_2132 ( .QN(net_2263), .RN(net_1347), .D(net_738), .CK(net_2836) );
CLKBUF_X2 inst_4013 ( .A(net_3804), .Z(net_3805) );
INV_X2 inst_1559 ( .ZN(net_241), .A(x4690) );
DFF_X1 inst_1928 ( .D(net_1129), .QN(net_59), .CK(net_3479) );
DFF_X1 inst_1967 ( .Q(net_2133), .D(net_1103), .CK(net_3399) );
NAND2_X2 inst_927 ( .A2(net_1627), .ZN(net_1087), .A1(net_689) );
NAND2_X4 inst_752 ( .ZN(net_1999), .A2(net_1997), .A1(net_1782) );
CLKBUF_X2 inst_3245 ( .A(net_2462), .Z(net_3037) );
SDFF_X2 inst_73 ( .SE(net_488), .Q(net_161), .D(net_161), .CK(net_2491), .SI(x4629) );
INV_X2 inst_1488 ( .A(net_2424), .ZN(net_373) );
DFF_X2 inst_1719 ( .QN(net_2331), .D(net_1493), .CK(net_3177) );
DFF_X1 inst_1947 ( .Q(net_2113), .D(net_1057), .CK(net_3114) );
CLKBUF_X2 inst_3202 ( .A(net_2559), .Z(net_2994) );
OAI21_X2 inst_378 ( .A(net_1938), .ZN(net_1359), .B2(net_1356), .B1(net_1343) );
DFF_X1 inst_1951 ( .Q(net_2117), .D(net_1097), .CK(net_3538) );
INV_X2 inst_1384 ( .A(net_766), .ZN(net_632) );
DFFR_X1 inst_2118 ( .QN(net_2309), .D(net_1606), .RN(net_1347), .CK(net_2755) );
NAND2_X2 inst_890 ( .A2(net_1691), .A1(net_1690), .ZN(net_1130) );
DFF_X1 inst_1851 ( .QN(net_2368), .D(net_1422), .CK(net_3615) );
INV_X8 inst_1168 ( .ZN(net_1984), .A(net_1983) );
OAI22_X2 inst_250 ( .B2(net_2271), .A1(net_745), .ZN(net_723), .A2(net_722), .B1(net_534) );
NAND3_X2 inst_659 ( .A3(net_1722), .A1(net_1658), .ZN(net_1132), .A2(net_984) );
INV_X8 inst_1161 ( .ZN(net_1872), .A(net_1871) );
CLKBUF_X2 inst_3362 ( .A(net_2546), .Z(net_3154) );
INV_X2 inst_1523 ( .ZN(net_263), .A(x5020) );
AOI21_X2 inst_2539 ( .A(net_1785), .B1(net_910), .ZN(net_789), .B2(net_788) );
NAND2_X2 inst_1048 ( .A1(net_1743), .ZN(net_1675), .A2(net_1207) );
CLKBUF_X2 inst_3199 ( .A(net_2990), .Z(net_2991) );
CLKBUF_X2 inst_2797 ( .A(net_2588), .Z(net_2589) );
CLKBUF_X2 inst_3612 ( .A(net_3321), .Z(net_3404) );
CLKBUF_X2 inst_3431 ( .A(net_3061), .Z(net_3223) );
INV_X2 inst_1581 ( .A(net_2337), .ZN(net_397) );
AOI22_X2 inst_2270 ( .ZN(net_1703), .A2(net_1547), .B1(net_1001), .A1(net_1000), .B2(net_796) );
DFFR_X2 inst_2085 ( .RN(net_1347), .D(net_1132), .QN(net_82), .CK(net_3510) );
AOI22_X2 inst_2388 ( .A1(net_1718), .B1(net_1474), .B2(net_660), .ZN(net_628), .A2(net_370) );
AOI22_X2 inst_2401 ( .B1(net_2197), .ZN(net_1629), .A1(net_1621), .B2(net_1526), .A2(net_1228) );
AOI22_X2 inst_2312 ( .A2(net_2145), .B1(net_2096), .A1(net_1769), .B2(net_1531), .ZN(net_897) );
CLKBUF_X2 inst_3500 ( .A(net_2573), .Z(net_3292) );
AND2_X2 inst_2634 ( .A1(net_594), .A2(x7169), .ZN(x748) );
CLKBUF_X2 inst_3711 ( .A(net_3315), .Z(net_3503) );
AOI22_X2 inst_2241 ( .B2(net_2121), .A1(net_1967), .B1(net_1450), .ZN(net_1389), .A2(net_933) );
NOR2_X2 inst_556 ( .ZN(net_547), .A2(net_524), .A1(net_462) );
NAND3_X2 inst_650 ( .A3(net_2371), .A1(net_1738), .ZN(net_1369), .A2(net_1207) );
OAI22_X2 inst_289 ( .A1(net_1615), .B1(net_1406), .B2(net_194), .A2(net_124), .ZN(x450) );
CLKBUF_X2 inst_2667 ( .A(net_2458), .Z(net_2459) );
CLKBUF_X2 inst_3632 ( .A(net_3331), .Z(net_3424) );
CLKBUF_X2 inst_4194 ( .A(net_3528), .Z(net_3986) );
NAND2_X2 inst_987 ( .A2(net_1571), .A1(net_961), .ZN(net_852) );
OAI21_X2 inst_420 ( .B2(net_2377), .B1(net_2194), .ZN(net_634), .A(net_615) );
NAND3_X2 inst_679 ( .A2(net_2417), .A3(net_1752), .ZN(net_469), .A1(net_468) );
CLKBUF_X2 inst_3006 ( .A(net_2728), .Z(net_2798) );
CLKBUF_X2 inst_3992 ( .A(net_3783), .Z(net_3784) );
CLKBUF_X2 inst_3265 ( .A(net_3056), .Z(net_3057) );
CLKBUF_X2 inst_3364 ( .A(net_3155), .Z(net_3156) );
INV_X4 inst_1351 ( .ZN(net_2196), .A(net_2195) );
SDFF_X2 inst_44 ( .QN(net_2438), .SI(net_2053), .SE(net_1935), .D(net_1246), .CK(net_3884) );
CLKBUF_X2 inst_3300 ( .A(net_3091), .Z(net_3092) );
OAI21_X2 inst_371 ( .B2(net_2180), .B1(net_1443), .ZN(net_1418), .A(net_1381) );
INV_X4 inst_1305 ( .A(net_2369), .ZN(net_1735) );
OAI222_X2 inst_314 ( .A2(net_2333), .B1(net_2186), .A1(net_2041), .ZN(net_2021), .C1(net_1965), .B2(net_1959), .C2(net_44) );
OAI21_X2 inst_435 ( .B2(net_2415), .ZN(net_1979), .B1(net_1978), .A(net_1976) );
CLKBUF_X2 inst_3225 ( .A(net_3016), .Z(net_3017) );
CLKBUF_X2 inst_3822 ( .A(net_3613), .Z(net_3614) );
NOR2_X2 inst_597 ( .A2(net_2262), .ZN(net_1886), .A1(net_520) );
CLKBUF_X2 inst_3307 ( .A(net_3098), .Z(net_3099) );
INV_X2 inst_1587 ( .ZN(net_221), .A(x4129) );
INV_X4 inst_1185 ( .ZN(net_1184), .A(net_1173) );
CLKBUF_X2 inst_3787 ( .A(net_2613), .Z(net_3579) );
NOR2_X1 inst_628 ( .ZN(net_1867), .A1(net_1748), .A2(net_361) );
CLKBUF_X2 inst_3684 ( .A(net_3129), .Z(net_3476) );
DFF_X1 inst_1923 ( .QN(net_2442), .D(net_2166), .CK(net_3682) );
CLKBUF_X2 inst_2748 ( .A(net_2539), .Z(net_2540) );
CLKBUF_X2 inst_3013 ( .A(net_2804), .Z(net_2805) );
OAI211_X2 inst_472 ( .C1(net_1054), .ZN(net_1038), .B(net_861), .A(net_838), .C2(net_406) );
OAI21_X1 inst_447 ( .B2(net_2418), .ZN(net_2052), .A(net_2051), .B1(net_1250) );
CLKBUF_X2 inst_3642 ( .A(net_2712), .Z(net_3434) );
OAI211_X2 inst_457 ( .C2(net_2353), .C1(net_1639), .ZN(net_1094), .A(net_818), .B(net_666) );
DFF_X2 inst_1738 ( .QN(net_2334), .D(net_1485), .CK(net_3170) );
AND2_X2 inst_2623 ( .A1(net_594), .A2(x7369), .ZN(x835) );
CLKBUF_X2 inst_2802 ( .A(net_2593), .Z(net_2594) );
CLKBUF_X2 inst_4171 ( .A(net_3962), .Z(net_3963) );
INV_X2 inst_1391 ( .A(net_584), .ZN(x971) );
CLKBUF_X2 inst_3092 ( .A(net_2761), .Z(net_2884) );
NAND3_X2 inst_665 ( .A1(net_1956), .A2(net_1803), .ZN(net_1077), .A3(net_806) );
CLKBUF_X2 inst_2734 ( .A(net_2525), .Z(net_2526) );
CLKBUF_X2 inst_3395 ( .A(net_3186), .Z(net_3187) );
INV_X8 inst_1130 ( .A(net_2044), .ZN(net_1367) );
CLKBUF_X2 inst_3538 ( .A(net_3329), .Z(net_3330) );
NAND2_X2 inst_855 ( .A2(net_1276), .ZN(net_1234), .A1(net_1233) );
DFF_X1 inst_2039 ( .Q(net_2394), .D(net_673), .CK(net_3150) );
CLKBUF_X2 inst_3755 ( .A(net_3001), .Z(net_3547) );
OR2_X1 inst_146 ( .A1(net_1404), .A2(x6157), .ZN(x101) );
CLKBUF_X2 inst_3233 ( .A(net_2561), .Z(net_3025) );
CLKBUF_X2 inst_3999 ( .A(net_3376), .Z(net_3791) );
INV_X4 inst_1196 ( .ZN(net_714), .A(net_534) );
OAI21_X2 inst_326 ( .B1(net_1507), .ZN(net_1504), .A(net_1470), .B2(net_1056) );
NAND2_X2 inst_817 ( .A1(net_1841), .ZN(net_1295), .A2(net_1199) );
CLKBUF_X2 inst_3428 ( .A(net_3219), .Z(net_3220) );
NOR2_X4 inst_518 ( .ZN(net_479), .A1(net_430), .A2(net_355) );
INV_X2 inst_1363 ( .A(net_1022), .ZN(x2483) );
CLKBUF_X2 inst_3336 ( .A(net_2831), .Z(net_3128) );
CLKBUF_X2 inst_3863 ( .A(net_3654), .Z(net_3655) );
CLKBUF_X2 inst_3293 ( .A(net_2520), .Z(net_3085) );
AOI22_X2 inst_2345 ( .B1(net_2197), .A1(net_2038), .A2(net_1549), .B2(net_1516), .ZN(net_819) );
CLKBUF_X2 inst_2837 ( .A(net_2618), .Z(net_2629) );
CLKBUF_X2 inst_3793 ( .A(net_3584), .Z(net_3585) );
SDFF_X2 inst_108 ( .SE(net_488), .Q(net_171), .D(net_171), .CK(net_3019), .SI(x4397) );
DFF_X1 inst_1845 ( .QN(net_2339), .D(net_1483), .CK(net_3192) );
CLKBUF_X2 inst_3778 ( .A(net_3569), .Z(net_3570) );
CLKBUF_X2 inst_3602 ( .A(net_2743), .Z(net_3394) );
CLKBUF_X2 inst_3940 ( .A(net_3731), .Z(net_3732) );
INV_X2 inst_1354 ( .A(net_1413), .ZN(x108) );
INV_X2 inst_1429 ( .ZN(net_444), .A(net_418) );
NAND2_X2 inst_970 ( .A2(net_1562), .A1(net_961), .ZN(net_869) );
INV_X4 inst_1278 ( .A(net_2351), .ZN(net_1240) );
CLKBUF_X2 inst_3763 ( .A(net_3554), .Z(net_3555) );
NAND4_X2 inst_638 ( .ZN(net_1937), .A3(net_1914), .A2(net_1835), .A1(net_1760), .A4(net_537) );
NOR2_X2 inst_586 ( .A2(net_2278), .ZN(net_1875), .A1(net_520) );
NAND2_X4 inst_749 ( .ZN(net_1977), .A2(net_1872), .A1(net_1666) );
NAND2_X2 inst_1030 ( .A1(net_2094), .ZN(net_482), .A2(net_472) );
DFFR_X1 inst_2127 ( .QN(net_2297), .RN(net_1347), .D(net_952), .CK(net_2751) );
AND2_X4 inst_2591 ( .A2(net_2204), .ZN(net_1980), .A1(net_1757) );
AND2_X2 inst_2649 ( .A2(net_2168), .ZN(net_1902), .A1(net_399) );
CLKBUF_X2 inst_3275 ( .A(net_2526), .Z(net_3067) );
INV_X2 inst_1466 ( .ZN(net_395), .A(net_364) );
DFF_X2 inst_1726 ( .QN(net_2322), .D(net_1508), .CK(net_3322) );
CLKBUF_X2 inst_2841 ( .A(net_2490), .Z(net_2633) );
INV_X2 inst_1373 ( .A(net_1011), .ZN(x2661) );
AOI22_X2 inst_2268 ( .ZN(net_1699), .A2(net_1545), .B1(net_1001), .A1(net_1000), .B2(net_909) );
CLKBUF_X2 inst_2652 ( .A(x7552), .Z(net_2444) );
INV_X4 inst_1203 ( .A(net_1719), .ZN(net_552) );
AOI222_X2 inst_2458 ( .C1(net_2014), .A2(net_1549), .A1(net_590), .B1(net_589), .ZN(net_578), .B2(net_151), .C2(x5796) );
CLKBUF_X2 inst_3828 ( .A(net_3619), .Z(net_3620) );
OAI22_X2 inst_296 ( .A1(net_1615), .B1(net_1404), .B2(net_239), .A2(net_140), .ZN(x140) );
NAND2_X2 inst_802 ( .ZN(net_1311), .A1(net_1277), .A2(net_1237) );
NAND2_X2 inst_905 ( .A1(net_1760), .ZN(net_1114), .A2(net_280) );
CLKBUF_X2 inst_3155 ( .A(net_2946), .Z(net_2947) );
CLKBUF_X2 inst_3134 ( .A(net_2925), .Z(net_2926) );
NAND2_X2 inst_1006 ( .A2(net_2122), .A1(net_979), .ZN(net_666) );
DFF_X1 inst_1985 ( .Q(net_2149), .D(net_1049), .CK(net_2994) );
CLKBUF_X2 inst_4214 ( .A(net_4005), .Z(net_4006) );
CLKBUF_X2 inst_3834 ( .A(net_3625), .Z(net_3626) );
CLKBUF_X2 inst_4043 ( .A(net_3834), .Z(net_3835) );
CLKBUF_X2 inst_3943 ( .A(net_3223), .Z(net_3735) );
CLKBUF_X2 inst_3651 ( .A(net_3442), .Z(net_3443) );
DFF_X2 inst_1759 ( .QN(net_2354), .D(net_1433), .CK(net_3734) );
AND2_X2 inst_2615 ( .A1(net_609), .A2(x7033), .ZN(x691) );
AOI21_X2 inst_2532 ( .A(net_1785), .B1(net_910), .ZN(net_801), .B2(net_79) );
AOI222_X2 inst_2463 ( .C1(net_2017), .A2(net_1561), .A1(net_590), .B1(net_589), .ZN(net_573), .B2(net_163), .C2(x5507) );
CLKBUF_X2 inst_3463 ( .A(net_3254), .Z(net_3255) );
CLKBUF_X2 inst_4055 ( .A(net_3846), .Z(net_3847) );
INV_X4 inst_1247 ( .A(net_1775), .ZN(net_402) );
INV_X2 inst_1464 ( .A(net_1538), .ZN(net_739) );
INV_X2 inst_1493 ( .A(net_1577), .ZN(net_334) );
INV_X4 inst_1308 ( .A(net_1746), .ZN(net_1745) );
SDFF_X2 inst_85 ( .Q(net_1570), .D(net_1570), .SE(net_491), .CK(net_2618), .SI(x6880) );
CLKBUF_X2 inst_3070 ( .A(net_2861), .Z(net_2862) );
CLKBUF_X2 inst_2998 ( .A(net_2472), .Z(net_2790) );
AND2_X2 inst_2612 ( .A1(net_609), .A2(x6845), .ZN(x615) );
CLKBUF_X2 inst_4184 ( .A(net_3975), .Z(net_3976) );
CLKBUF_X2 inst_4049 ( .A(net_3840), .Z(net_3841) );
CLKBUF_X2 inst_2702 ( .A(net_2452), .Z(net_2494) );
CLKBUF_X2 inst_2910 ( .A(net_2701), .Z(net_2702) );
CLKBUF_X2 inst_4022 ( .A(net_3813), .Z(net_3814) );
INV_X2 inst_1362 ( .A(net_989), .ZN(x2496) );
CLKBUF_X2 inst_3238 ( .A(net_3029), .Z(net_3030) );
OAI22_X2 inst_290 ( .A1(net_1615), .B1(net_1404), .B2(net_244), .A2(net_125), .ZN(x439) );
OR2_X1 inst_145 ( .A1(net_1404), .A2(x6122), .ZN(x91) );
DFF_X1 inst_1978 ( .Q(net_2143), .D(net_1035), .CK(net_3066) );
OAI22_X2 inst_272 ( .B2(net_2286), .B1(net_1865), .ZN(net_1604), .A1(net_951), .A2(net_938) );
CLKBUF_X2 inst_2854 ( .A(net_2645), .Z(net_2646) );
CLKBUF_X2 inst_3030 ( .A(net_2821), .Z(net_2822) );
DFFR_X1 inst_2112 ( .QN(net_2303), .RN(net_1347), .D(net_946), .CK(net_2725) );
NAND2_X2 inst_814 ( .ZN(net_1299), .A2(net_1258), .A1(net_1221) );
CLKBUF_X2 inst_3036 ( .A(net_2827), .Z(net_2828) );
AOI22_X2 inst_2230 ( .ZN(net_1412), .A2(net_428), .A1(net_143), .B2(x6207), .B1(x5995) );
INV_X2 inst_1458 ( .A(net_2370), .ZN(net_1207) );
CLKBUF_X2 inst_3471 ( .A(net_3262), .Z(net_3263) );
CLKBUF_X2 inst_4133 ( .A(net_2597), .Z(net_3925) );
NAND2_X2 inst_789 ( .A1(net_1818), .ZN(net_1324), .A2(net_1208) );
DFF_X2 inst_1806 ( .QN(net_2209), .CK(net_2867), .D(x6470) );
DFF_X2 inst_1810 ( .Q(net_1532), .CK(net_2558), .D(x5913) );
DFF_X1 inst_1860 ( .QN(net_2441), .D(net_1409), .CK(net_3695) );
AOI22_X2 inst_2275 ( .ZN(net_1711), .B1(net_1001), .A1(net_999), .B2(net_786), .A2(net_681) );
DFF_X1 inst_1885 ( .D(net_1297), .QN(net_92), .CK(net_3875) );
INV_X2 inst_1437 ( .A(net_1535), .ZN(net_953) );
NAND2_X2 inst_822 ( .A1(net_1840), .ZN(net_1339), .A2(net_401) );
NAND2_X1 inst_1125 ( .A1(net_2385), .A2(net_2376), .ZN(net_523) );
NOR2_X2 inst_609 ( .ZN(net_1969), .A2(net_681), .A1(net_356) );
AOI21_X2 inst_2533 ( .A(net_1785), .B1(net_910), .ZN(net_800), .B2(net_80) );
AOI22_X2 inst_2391 ( .A2(net_2200), .A1(net_2195), .B1(net_839), .ZN(net_625), .B2(net_72) );
NAND2_X2 inst_795 ( .A2(net_1678), .ZN(net_1318), .A1(net_1288) );
AOI222_X1 inst_2496 ( .B1(net_1995), .A1(net_1751), .B2(net_1555), .C1(net_1020), .ZN(net_1004), .A2(net_157), .C2(x3580) );
AOI22_X2 inst_2239 ( .B2(net_2128), .A1(net_1967), .B1(net_1450), .ZN(net_1391), .A2(net_1238) );
XNOR2_X2 inst_27 ( .ZN(net_924), .A(net_670), .B(net_366) );
AOI222_X1 inst_2491 ( .B1(net_1995), .A1(net_1751), .B2(net_1560), .C1(net_1020), .ZN(net_1009), .A2(net_162), .C2(x3465) );
INV_X2 inst_1639 ( .ZN(net_184), .A(x4164) );
NOR2_X1 inst_619 ( .A2(net_2434), .A1(net_1748), .ZN(net_1361) );
CLKBUF_X2 inst_2671 ( .A(net_2462), .Z(net_2463) );
INV_X2 inst_1654 ( .ZN(net_179), .A(x4461) );
NAND4_X2 inst_639 ( .ZN(net_1938), .A3(net_1914), .A2(net_1835), .A1(net_1760), .A4(net_1198) );
INV_X2 inst_1355 ( .A(net_1412), .ZN(x116) );
NAND2_X2 inst_877 ( .A1(net_1838), .A2(net_1240), .ZN(net_1200) );
OAI22_X2 inst_155 ( .B1(net_1428), .A1(net_529), .B2(net_213), .A2(net_106), .ZN(x1425) );
CLKBUF_X2 inst_3939 ( .A(net_2986), .Z(net_3731) );
SDFF_X2 inst_55 ( .SE(net_1768), .SI(net_1535), .Q(net_72), .D(net_72), .CK(net_3235) );
AOI22_X2 inst_2280 ( .B1(net_1768), .ZN(net_1706), .A2(net_1550), .B2(net_1515), .A1(net_1000) );
DFFR_X2 inst_2076 ( .D(net_1952), .QN(net_1582), .RN(net_1347), .CK(net_3982) );
INV_X2 inst_1651 ( .A(net_2280), .ZN(net_310) );
CLKBUF_X2 inst_4127 ( .A(net_3918), .Z(net_3919) );
AOI222_X1 inst_2481 ( .B1(net_1995), .A1(net_1751), .B2(net_1570), .C1(net_1020), .ZN(net_1019), .A2(net_172), .C2(x3295) );
INV_X8 inst_1137 ( .A(net_2097), .ZN(net_962) );
OAI21_X2 inst_323 ( .B2(net_2322), .ZN(net_1508), .B1(net_1507), .A(net_1471) );
INV_X8 inst_1162 ( .A(net_1965), .ZN(net_1915) );
INV_X2 inst_1389 ( .A(net_586), .ZN(x957) );
CLKBUF_X2 inst_2973 ( .A(net_2544), .Z(net_2765) );
CLKBUF_X2 inst_3065 ( .A(net_2856), .Z(net_2857) );
NAND2_X4 inst_715 ( .ZN(net_598), .A1(net_541), .A2(net_325) );
NAND2_X2 inst_793 ( .ZN(net_1320), .A1(net_1289), .A2(net_1231) );
INV_X2 inst_1433 ( .A(net_1521), .ZN(net_707) );
INV_X2 inst_1494 ( .A(net_2430), .ZN(net_772) );
DFF_X1 inst_1894 ( .D(net_1342), .QN(net_127), .CK(net_3757) );
CLKBUF_X2 inst_3525 ( .A(net_3316), .Z(net_3317) );
DFF_X1 inst_1999 ( .Q(net_2163), .D(net_1065), .CK(net_3426) );
CLKBUF_X2 inst_3449 ( .A(net_3240), .Z(net_3241) );
INV_X2 inst_1682 ( .A(net_2311), .ZN(net_2091) );
CLKBUF_X2 inst_2733 ( .A(net_2524), .Z(net_2525) );
INV_X4 inst_1340 ( .A(net_2327), .ZN(net_2066) );
INV_X2 inst_1481 ( .A(net_1541), .ZN(net_747) );
OAI211_X2 inst_475 ( .C2(net_2313), .C1(net_1054), .ZN(net_1034), .A(net_895), .B(net_867) );
XNOR2_X2 inst_31 ( .B(net_1197), .ZN(net_679), .A(net_598) );
CLKBUF_X2 inst_2701 ( .A(net_2492), .Z(net_2493) );
CLKBUF_X2 inst_3505 ( .A(net_3296), .Z(net_3297) );
CLKBUF_X2 inst_3165 ( .A(net_2956), .Z(net_2957) );
CLKBUF_X2 inst_3217 ( .A(net_3008), .Z(net_3009) );
NOR2_X2 inst_575 ( .A2(net_2326), .ZN(net_1647), .A1(net_1643) );
CLKBUF_X2 inst_3537 ( .A(net_3328), .Z(net_3329) );
NOR2_X1 inst_627 ( .A2(net_2327), .ZN(net_1646), .A1(net_1644) );
CLKBUF_X2 inst_3352 ( .A(net_3143), .Z(net_3144) );
OAI21_X2 inst_344 ( .ZN(net_1485), .B2(net_1484), .A(net_1452), .B1(net_1254) );
DFF_X2 inst_1833 ( .Q(net_1535), .CK(net_2775), .D(x5527) );
DFFR_X1 inst_2122 ( .QN(net_2286), .D(net_1604), .RN(net_1347), .CK(net_3547) );
CLKBUF_X2 inst_3044 ( .A(net_2835), .Z(net_2836) );
CLKBUF_X2 inst_3520 ( .A(net_3311), .Z(net_3312) );
CLKBUF_X2 inst_3573 ( .A(net_3364), .Z(net_3365) );
NOR2_X1 inst_623 ( .A2(net_2316), .A1(net_2315), .ZN(net_279) );
NAND2_X2 inst_1072 ( .A1(net_2104), .ZN(net_1813), .A2(net_1242) );
CLKBUF_X2 inst_3580 ( .A(net_3371), .Z(net_3372) );
CLKBUF_X2 inst_3818 ( .A(net_3609), .Z(net_3610) );
INV_X2 inst_1621 ( .ZN(net_198), .A(x6623) );
DFF_X1 inst_1993 ( .Q(net_2157), .D(net_1033), .CK(net_3369) );
INV_X4 inst_1338 ( .A(net_2074), .ZN(net_2030) );
AOI22_X2 inst_2430 ( .B2(net_2112), .B1(net_1974), .ZN(net_1804), .A1(net_1791), .A2(net_288) );
CLKBUF_X2 inst_3080 ( .A(net_2871), .Z(net_2872) );
AOI22_X2 inst_2434 ( .B2(net_2142), .B1(net_1974), .ZN(net_1808), .A1(net_1789), .A2(net_290) );
CLKBUF_X2 inst_3226 ( .A(net_3017), .Z(net_3018) );
CLKBUF_X2 inst_3731 ( .A(net_3522), .Z(net_3523) );
NAND2_X2 inst_1107 ( .ZN(net_2019), .A1(net_2012), .A2(net_82) );
CLKBUF_X2 inst_3617 ( .A(net_2668), .Z(net_3409) );
INV_X2 inst_1377 ( .A(net_1007), .ZN(x2722) );
DFF_X1 inst_2028 ( .QN(net_2409), .D(net_2188), .CK(net_3703) );
CLKBUF_X2 inst_3125 ( .A(net_2916), .Z(net_2917) );
AOI22_X4 inst_2201 ( .ZN(net_2072), .B1(net_2071), .A1(net_2070), .B2(x5181), .A2(x3190) );
NAND2_X4 inst_722 ( .A1(net_2200), .A2(net_2173), .ZN(net_492) );
CLKBUF_X2 inst_2776 ( .A(net_2567), .Z(net_2568) );
NAND2_X4 inst_760 ( .ZN(net_2044), .A1(net_2043), .A2(net_1868) );
NAND2_X4 inst_746 ( .ZN(net_1964), .A1(net_1869), .A2(net_417) );
INV_X16 inst_1696 ( .A(net_1991), .ZN(net_1929) );
CLKBUF_X2 inst_4232 ( .A(net_4023), .Z(net_4024) );
AOI22_X2 inst_2267 ( .ZN(net_1693), .A2(net_1544), .A1(net_1000), .B1(net_999), .B2(net_370) );
CLKBUF_X2 inst_3010 ( .A(net_2801), .Z(net_2802) );
CLKBUF_X2 inst_4115 ( .A(net_3906), .Z(net_3907) );
CLKBUF_X2 inst_3133 ( .A(net_2886), .Z(net_2925) );
CLKBUF_X2 inst_3727 ( .A(net_2801), .Z(net_3519) );
INV_X2 inst_1577 ( .A(net_2271), .ZN(net_289) );
INV_X16 inst_1687 ( .ZN(net_910), .A(net_555) );
NAND2_X2 inst_1110 ( .ZN(net_2039), .A2(net_1965), .A1(net_1957) );
DFF_X1 inst_1970 ( .Q(net_2136), .D(net_1101), .CK(net_3393) );
AND2_X4 inst_2588 ( .A1(net_2384), .A2(net_2383), .ZN(net_1775) );
CLKBUF_X2 inst_3989 ( .A(net_3780), .Z(net_3781) );
CLKBUF_X2 inst_2873 ( .A(net_2664), .Z(net_2665) );
AOI22_X2 inst_2442 ( .A1(net_1974), .ZN(net_1920), .A2(net_1919), .B1(net_1789), .B2(net_308) );
CLKBUF_X2 inst_3569 ( .A(net_2840), .Z(net_3361) );
DFF_X1 inst_2066 ( .QN(net_2374), .D(net_2345), .CK(net_4019) );
CLKBUF_X2 inst_3411 ( .A(net_3202), .Z(net_3203) );
AOI21_X2 inst_2524 ( .A(net_1785), .B1(net_910), .ZN(net_809), .B2(net_71) );
INV_X2 inst_1446 ( .A(net_1516), .ZN(net_939) );
OAI21_X2 inst_390 ( .B1(net_1740), .ZN(net_1336), .A(net_1335), .B2(net_359) );
AOI22_X2 inst_2421 ( .B2(net_2154), .B1(net_1974), .ZN(net_1795), .A1(net_1791), .A2(net_340) );
DFF_X2 inst_1742 ( .QN(net_2364), .D(net_1419), .CK(net_3637) );
NAND2_X2 inst_1062 ( .A1(net_1954), .ZN(net_1721), .A2(net_1559) );
CLKBUF_X2 inst_2663 ( .A(net_2448), .Z(net_2455) );
CLKBUF_X2 inst_2875 ( .A(net_2666), .Z(net_2667) );
CLKBUF_X2 inst_3289 ( .A(net_3080), .Z(net_3081) );
OAI21_X2 inst_401 ( .B2(net_2379), .ZN(net_988), .B1(net_920), .A(net_637) );
AOI22_X2 inst_2302 ( .A2(net_2149), .B1(net_2096), .A1(net_1769), .B2(net_1525), .ZN(net_907) );
CLKBUF_X2 inst_3175 ( .A(net_2966), .Z(net_2967) );
CLKBUF_X2 inst_3389 ( .A(net_3180), .Z(net_3181) );
CLKBUF_X2 inst_3210 ( .A(net_2661), .Z(net_3002) );
AOI222_X2 inst_2447 ( .C1(net_2016), .A2(net_1544), .ZN(net_591), .A1(net_590), .B1(net_589), .B2(net_146), .C2(x5913) );
NAND2_X2 inst_782 ( .A1(net_1814), .ZN(net_1331), .A2(net_1211) );
AND2_X2 inst_2642 ( .A1(net_2013), .A2(x6678), .ZN(x550) );
CLKBUF_X2 inst_2869 ( .A(net_2611), .Z(net_2661) );
XOR2_X1 inst_6 ( .B(net_2336), .Z(net_2179), .A(net_1159) );
AOI222_X1 inst_2486 ( .B1(net_1995), .A1(net_1751), .B2(net_1564), .C1(net_1020), .ZN(net_1014), .A2(net_166), .C2(x3396) );
AOI22_X2 inst_2410 ( .B2(net_2135), .ZN(net_1638), .A1(net_1621), .A2(net_1225), .B1(net_979) );
SDFFR_X1 inst_123 ( .SE(net_1829), .D(net_1539), .RN(net_1347), .SI(net_48), .Q(net_48), .CK(net_2860) );
NAND2_X2 inst_930 ( .A2(net_1628), .ZN(net_1084), .A1(net_683) );
NAND2_X2 inst_935 ( .A2(net_1622), .ZN(net_1065), .A1(net_685) );
AOI22_X2 inst_2298 ( .B1(net_1768), .ZN(net_1698), .B2(net_1521), .A1(net_999), .A2(net_357) );
OAI22_X2 inst_167 ( .B1(net_1406), .A1(net_1403), .B2(net_257), .A2(net_126), .ZN(x421) );
CLKBUF_X2 inst_2944 ( .A(net_2735), .Z(net_2736) );
NAND2_X2 inst_1026 ( .A1(net_1931), .A2(net_1577), .ZN(net_539) );
INV_X4 inst_1320 ( .A(net_2015), .ZN(net_1895) );
CLKBUF_X2 inst_3874 ( .A(net_3665), .Z(net_3666) );
INV_X4 inst_1251 ( .A(net_1583), .ZN(net_601) );
SDFF_X2 inst_95 ( .SE(net_487), .Q(net_162), .D(net_162), .CK(net_2770), .SI(x4604) );
CLKBUF_X2 inst_3376 ( .A(net_3167), .Z(net_3168) );
AOI222_X2 inst_2475 ( .C1(net_2017), .A2(net_1547), .A1(net_590), .B1(net_589), .ZN(net_561), .B2(net_149), .C2(x5846) );
CLKBUF_X2 inst_2921 ( .A(net_2661), .Z(net_2713) );
CLKBUF_X2 inst_2862 ( .A(net_2653), .Z(net_2654) );
OAI21_X2 inst_331 ( .B2(net_2317), .B1(net_2041), .ZN(net_1499), .A(net_1462) );
CLKBUF_X2 inst_4009 ( .A(net_3800), .Z(net_3801) );
AOI22_X2 inst_2353 ( .A1(net_783), .B1(net_782), .ZN(net_779), .A2(net_646), .B2(x3733) );
NAND3_X2 inst_667 ( .A2(net_1809), .A1(net_1762), .ZN(net_1075), .A3(net_804) );
CLKBUF_X2 inst_2762 ( .A(net_2453), .Z(net_2554) );
CLKBUF_X2 inst_2896 ( .A(net_2687), .Z(net_2688) );
NAND2_X2 inst_997 ( .A1(net_1790), .ZN(net_834), .A2(net_674) );
NAND2_X2 inst_857 ( .A1(net_1741), .ZN(net_1230), .A2(net_366) );
CLKBUF_X2 inst_2691 ( .A(net_2482), .Z(net_2483) );
CLKBUF_X2 inst_3590 ( .A(net_3381), .Z(net_3382) );
INV_X2 inst_1511 ( .A(net_2420), .ZN(net_370) );
CLKBUF_X2 inst_4179 ( .A(net_2676), .Z(net_3971) );
OAI21_X2 inst_365 ( .B2(net_2409), .B1(net_1441), .ZN(net_1429), .A(net_1391) );
CLKBUF_X2 inst_4006 ( .A(net_3797), .Z(net_3798) );
SDFF_X2 inst_67 ( .Q(net_1544), .D(net_1544), .SE(net_498), .CK(net_2684), .SI(x7509) );
NAND2_X2 inst_954 ( .A2(net_2358), .ZN(net_982), .A1(net_759) );
CLKBUF_X2 inst_3203 ( .A(net_2774), .Z(net_2995) );
INV_X2 inst_1504 ( .A(net_2324), .ZN(net_369) );
AOI222_X2 inst_2476 ( .C1(net_2016), .A2(net_1554), .A1(net_590), .B1(net_589), .ZN(net_560), .B2(net_156), .C2(x5686) );
CLKBUF_X2 inst_3403 ( .A(net_3194), .Z(net_3195) );
DFF_X2 inst_1823 ( .Q(net_1537), .CK(net_2815), .D(x5581) );
OAI22_X2 inst_202 ( .A2(net_2229), .B1(net_1406), .A1(net_1405), .B2(net_266), .ZN(x2016) );
INV_X4 inst_1310 ( .ZN(net_1751), .A(net_1750) );
AOI22_X2 inst_2212 ( .A2(net_2344), .B2(net_2111), .A1(net_1960), .B1(net_1915), .ZN(net_1468) );
CLKBUF_X2 inst_3280 ( .A(net_2548), .Z(net_3072) );
INV_X2 inst_1401 ( .A(net_574), .ZN(x1241) );
CLKBUF_X2 inst_2823 ( .A(net_2614), .Z(net_2615) );
DFF_X1 inst_2030 ( .QN(net_2240), .D(net_834), .CK(net_2993) );
CLKBUF_X2 inst_3807 ( .A(net_3598), .Z(net_3599) );
NAND2_X2 inst_1069 ( .A2(net_1858), .ZN(net_1771), .A1(net_1770) );
XNOR2_X2 inst_30 ( .B(net_1240), .ZN(net_692), .A(net_619) );
OR2_X2 inst_136 ( .ZN(net_451), .A2(net_426), .A1(net_407) );
NOR2_X2 inst_610 ( .ZN(net_1971), .A1(net_514), .A2(net_356) );
CLKBUF_X2 inst_3541 ( .A(net_3257), .Z(net_3333) );
NAND2_X2 inst_1036 ( .ZN(net_381), .A2(net_302), .A1(net_295) );
OAI22_X2 inst_233 ( .B2(net_2285), .B1(net_1865), .A1(net_951), .ZN(net_940), .A2(net_939) );
INV_X2 inst_1526 ( .A(net_2330), .ZN(net_285) );
AOI21_X2 inst_2547 ( .ZN(net_509), .A(net_479), .B1(net_430), .B2(net_355) );
NAND2_X2 inst_1047 ( .A1(net_1746), .ZN(net_1674), .A2(net_367) );
SDFF_X2 inst_60 ( .Q(net_1554), .D(net_1554), .SE(net_396), .CK(net_2926), .SI(x7314) );
CLKBUF_X2 inst_3850 ( .A(net_3641), .Z(net_3642) );
CLKBUF_X2 inst_3700 ( .A(net_2853), .Z(net_3492) );
DFF_X1 inst_1858 ( .QN(net_2436), .D(net_1397), .CK(net_3913) );
DFF_X2 inst_1786 ( .QN(net_2383), .D(net_765), .CK(net_3854) );
AOI22_X2 inst_2376 ( .B2(net_2134), .B1(net_1929), .A1(net_655), .ZN(net_654), .A2(net_300) );
CLKBUF_X2 inst_3846 ( .A(net_2587), .Z(net_3638) );
INV_X4 inst_1334 ( .ZN(net_2014), .A(net_2012) );
NOR3_X2 inst_496 ( .A1(net_462), .ZN(net_460), .A2(net_459), .A3(net_458) );
NAND2_X2 inst_860 ( .A1(net_1741), .ZN(net_1224), .A2(net_1213) );
NOR2_X2 inst_563 ( .A2(net_1825), .ZN(net_438), .A1(net_275) );
CLKBUF_X2 inst_3962 ( .A(net_3429), .Z(net_3754) );
NAND2_X2 inst_943 ( .ZN(net_1039), .A1(net_960), .A2(net_893) );
CLKBUF_X2 inst_3478 ( .A(net_3269), .Z(net_3270) );
CLKBUF_X2 inst_3749 ( .A(net_3540), .Z(net_3541) );
AND2_X2 inst_2620 ( .A1(net_594), .A2(x7297), .ZN(x794) );
CLKBUF_X2 inst_2782 ( .A(net_2573), .Z(net_2574) );
DFF_X1 inst_1964 ( .Q(net_2130), .D(net_1064), .CK(net_3434) );
INV_X2 inst_1633 ( .ZN(net_189), .A(x4008) );
DFF_X2 inst_1765 ( .QN(net_2430), .D(net_990), .CK(net_3627) );
INV_X4 inst_1262 ( .A(net_2279), .ZN(net_332) );
OAI22_X2 inst_265 ( .B2(net_2252), .A1(net_714), .ZN(net_697), .A2(net_696), .B1(net_534) );
CLKBUF_X2 inst_3720 ( .A(net_3511), .Z(net_3512) );
DFF_X1 inst_2005 ( .QN(net_2229), .D(net_1077), .CK(net_3036) );
DFF_X1 inst_2055 ( .D(net_508), .CK(net_4028), .Q(x8) );
CLKBUF_X2 inst_3856 ( .A(net_3647), .Z(net_3648) );
NOR2_X2 inst_544 ( .A1(net_1829), .ZN(net_849), .A2(net_848) );
NAND2_X4 inst_736 ( .ZN(net_1905), .A2(net_1904), .A1(net_1903) );
CLKBUF_X2 inst_3262 ( .A(net_3053), .Z(net_3054) );
OAI22_X2 inst_178 ( .B1(net_1428), .A1(net_1426), .B2(net_192), .A2(net_99), .ZN(x1507) );
NAND2_X4 inst_734 ( .A1(net_2094), .ZN(net_1869), .A2(net_1772) );
INV_X4 inst_1282 ( .A(net_2413), .ZN(net_277) );
NAND2_X2 inst_1077 ( .A1(net_2104), .A2(net_2076), .ZN(net_1818) );
INV_X8 inst_1148 ( .A(net_1904), .ZN(net_396) );
CLKBUF_X2 inst_3919 ( .A(net_3710), .Z(net_3711) );
CLKBUF_X2 inst_3954 ( .A(net_3745), .Z(net_3746) );
CLKBUF_X2 inst_2757 ( .A(net_2548), .Z(net_2549) );
OAI22_X2 inst_222 ( .B2(net_2292), .B1(net_1865), .A1(net_1597), .ZN(net_956), .A2(net_742) );
DFF_X1 inst_1932 ( .D(net_1127), .QN(net_61), .CK(net_3499) );
CLKBUF_X2 inst_3704 ( .A(net_3080), .Z(net_3496) );
CLKBUF_X2 inst_3587 ( .A(net_3173), .Z(net_3379) );
NAND2_X2 inst_1052 ( .A1(net_1743), .ZN(net_1679), .A2(net_322) );
INV_X4 inst_1280 ( .A(net_2312), .ZN(net_280) );
INV_X4 inst_1302 ( .ZN(net_1619), .A(net_1618) );
INV_X2 inst_1648 ( .A(net_2294), .ZN(net_326) );
NAND2_X2 inst_842 ( .A2(net_2076), .A1(net_1840), .ZN(net_1271) );
NAND2_X2 inst_1079 ( .A1(net_2104), .ZN(net_1820), .A2(net_1262) );
DFFS_X2 inst_2068 ( .QN(net_2413), .SN(net_1347), .D(net_1232), .CK(net_3972) );
CLKBUF_X2 inst_3925 ( .A(net_3083), .Z(net_3717) );
NOR2_X2 inst_551 ( .A1(net_621), .ZN(net_605), .A2(net_351) );
AND2_X2 inst_2606 ( .A1(net_609), .A2(x7383), .ZN(x844) );
DFFR_X1 inst_2101 ( .QN(net_2290), .RN(net_1347), .D(net_957), .CK(net_2887) );
AOI21_X2 inst_2523 ( .A(net_1785), .B1(net_910), .ZN(net_810), .B2(net_362) );
NOR2_X4 inst_506 ( .A2(net_2336), .ZN(net_1166), .A1(net_1159) );
OAI21_X2 inst_353 ( .B2(net_2408), .ZN(net_1442), .B1(net_1441), .A(net_1392) );
CLKBUF_X2 inst_3808 ( .A(net_3599), .Z(net_3600) );
DFF_X1 inst_1940 ( .QN(net_2212), .D(net_1131), .CK(net_3302) );
OR2_X2 inst_134 ( .A1(net_2417), .A2(net_1904), .ZN(net_437) );
AOI22_X2 inst_2409 ( .B2(net_2118), .ZN(net_1637), .A1(net_1621), .A2(net_1203), .B1(net_979) );
CLKBUF_X2 inst_3322 ( .A(net_3113), .Z(net_3114) );
NAND2_X2 inst_1085 ( .A2(net_1914), .ZN(net_1840), .A1(net_1788) );
INV_X4 inst_1323 ( .A(net_2010), .ZN(net_1927) );
CLKBUF_X2 inst_3425 ( .A(net_3216), .Z(net_3217) );
AOI22_X2 inst_2328 ( .ZN(net_842), .A1(net_840), .B1(net_839), .A2(net_412), .B2(net_78) );
CLKBUF_X2 inst_2655 ( .A(x7552), .Z(net_2447) );
OAI22_X2 inst_160 ( .A1(net_1408), .B1(net_1407), .B2(net_252), .A2(net_136), .ZN(x234) );
DFF_X2 inst_1720 ( .QN(net_2330), .D(net_1511), .CK(net_3172) );
CLKBUF_X2 inst_4041 ( .A(net_3832), .Z(net_3833) );
CLKBUF_X2 inst_3701 ( .A(net_3492), .Z(net_3493) );
CLKBUF_X2 inst_3357 ( .A(net_3148), .Z(net_3149) );
XOR2_X1 inst_8 ( .Z(net_2181), .A(net_1655), .B(net_327) );
CLKBUF_X2 inst_2912 ( .A(net_2600), .Z(net_2704) );
NAND2_X4 inst_762 ( .ZN(net_2065), .A2(net_2064), .A1(net_1831) );
OAI21_X2 inst_370 ( .B2(net_1443), .ZN(net_1419), .A(net_1382), .B1(net_1185) );
CLKBUF_X2 inst_3025 ( .A(net_2816), .Z(net_2817) );
INV_X4 inst_1265 ( .ZN(net_352), .A(net_327) );
DFFR_X2 inst_2090 ( .RN(net_1347), .D(net_1108), .QN(net_45), .CK(net_3977) );
NAND2_X2 inst_965 ( .A2(net_1557), .A1(net_961), .ZN(net_874) );
CLKBUF_X2 inst_3370 ( .A(net_2937), .Z(net_3162) );
INV_X4 inst_1321 ( .ZN(net_1896), .A(net_1850) );
NAND2_X2 inst_1012 ( .A2(net_1240), .ZN(net_642), .A1(net_618) );
NAND2_X2 inst_901 ( .A2(net_1703), .A1(net_1702), .ZN(net_1118) );
DFF_X1 inst_1956 ( .Q(net_2122), .D(net_1094), .CK(net_3536) );
CLKBUF_X2 inst_3492 ( .A(net_3283), .Z(net_3284) );
NAND2_X4 inst_751 ( .ZN(net_1991), .A2(net_1988), .A1(net_1927) );
CLKBUF_X2 inst_3149 ( .A(net_2940), .Z(net_2941) );
AOI22_X2 inst_2403 ( .B1(net_2197), .ZN(net_1631), .A1(net_1621), .B2(net_1536), .A2(net_366) );
AOI222_X2 inst_2471 ( .C1(net_2016), .A2(net_1552), .A1(net_590), .B1(net_589), .ZN(net_565), .B2(net_154), .C2(x5740) );
CLKBUF_X2 inst_4034 ( .A(net_3825), .Z(net_3826) );
OAI21_X2 inst_377 ( .B2(net_1967), .ZN(net_1401), .B1(net_1362), .A(net_367) );
DFF_X1 inst_1934 ( .D(net_1126), .QN(net_64), .CK(net_3470) );
CLKBUF_X2 inst_3946 ( .A(net_3737), .Z(net_3738) );
CLKBUF_X2 inst_3098 ( .A(net_2689), .Z(net_2890) );
CLKBUF_X2 inst_3244 ( .A(net_3035), .Z(net_3036) );
CLKBUF_X2 inst_3916 ( .A(net_2468), .Z(net_3708) );
CLKBUF_X2 inst_3920 ( .A(net_3711), .Z(net_3712) );
CLKBUF_X2 inst_3821 ( .A(net_2626), .Z(net_3613) );
CLKBUF_X2 inst_3018 ( .A(net_2809), .Z(net_2810) );
CLKBUF_X2 inst_3078 ( .A(net_2869), .Z(net_2870) );
CLKBUF_X2 inst_3835 ( .A(net_3626), .Z(net_3627) );
DFFR_X1 inst_2097 ( .QN(net_2293), .D(net_1601), .RN(net_1347), .CK(net_2889) );
NAND2_X2 inst_928 ( .A2(net_1631), .ZN(net_1086), .A1(net_687) );
SDFF_X2 inst_107 ( .SE(net_488), .Q(net_158), .D(net_158), .CK(net_2532), .SI(x4718) );
DFFR_X1 inst_2117 ( .QN(net_2281), .RN(net_1347), .D(net_943), .CK(net_2883) );
NAND2_X2 inst_990 ( .ZN(net_1657), .A1(net_1596), .A2(net_1519) );
CLKBUF_X2 inst_3140 ( .A(net_2485), .Z(net_2932) );
INV_X2 inst_1539 ( .A(net_2306), .ZN(net_312) );
CLKBUF_X2 inst_2662 ( .A(net_2453), .Z(net_2454) );
CLKBUF_X2 inst_3628 ( .A(net_3134), .Z(net_3420) );
DFF_X2 inst_1718 ( .QN(net_2332), .D(net_1489), .CK(net_2964) );
NAND2_X2 inst_1050 ( .A1(net_1746), .ZN(net_1677), .A2(net_1203) );
AOI22_X2 inst_2366 ( .B2(net_2164), .A1(net_2038), .A2(net_1552), .B1(net_979), .ZN(net_690) );
CLKBUF_X2 inst_3316 ( .A(net_2639), .Z(net_3108) );
INV_X4 inst_1296 ( .A(net_2358), .ZN(net_933) );
DFF_X1 inst_1852 ( .QN(net_2367), .D(net_1418), .CK(net_3614) );
CLKBUF_X2 inst_3671 ( .A(net_3462), .Z(net_3463) );
CLKBUF_X2 inst_3282 ( .A(net_3073), .Z(net_3074) );
CLKBUF_X2 inst_4014 ( .A(net_3805), .Z(net_3806) );
CLKBUF_X2 inst_3694 ( .A(net_3131), .Z(net_3486) );
CLKBUF_X2 inst_4074 ( .A(net_3865), .Z(net_3866) );
CLKBUF_X2 inst_3783 ( .A(net_2598), .Z(net_3575) );
INV_X2 inst_1557 ( .A(net_2384), .ZN(net_243) );
AOI22_X2 inst_2399 ( .B1(net_2197), .A2(net_1845), .ZN(net_1627), .A1(net_1621), .B2(net_1539) );
CLKBUF_X2 inst_2698 ( .A(net_2489), .Z(net_2490) );
INV_X4 inst_1237 ( .A(net_1904), .ZN(net_491) );
CLKBUF_X2 inst_3412 ( .A(net_3203), .Z(net_3204) );
AOI21_X2 inst_2518 ( .A(net_1967), .ZN(net_1368), .B2(net_1367), .B1(net_1194) );
CLKBUF_X2 inst_3460 ( .A(net_3251), .Z(net_3252) );
INV_X2 inst_1616 ( .A(net_2257), .ZN(net_338) );
DFFR_X2 inst_2075 ( .QN(net_1579), .RN(net_1347), .D(net_1252), .CK(net_3984) );
CLKBUF_X2 inst_3062 ( .A(net_2853), .Z(net_2854) );
CLKBUF_X2 inst_3310 ( .A(net_3101), .Z(net_3102) );
DFF_X1 inst_1911 ( .D(net_1307), .Q(net_142), .CK(net_3044) );
CLKBUF_X2 inst_4151 ( .A(net_3942), .Z(net_3943) );
DFF_X2 inst_1825 ( .QN(net_2207), .CK(net_2699), .D(x6530) );
NOR2_X2 inst_585 ( .ZN(net_1868), .A2(net_1867), .A1(net_1866) );
INV_X2 inst_1606 ( .A(net_2273), .ZN(net_300) );
CLKBUF_X2 inst_2851 ( .A(net_2486), .Z(net_2643) );
OAI21_X2 inst_410 ( .ZN(net_764), .B2(net_661), .B1(net_622), .A(net_243) );
OAI21_X4 inst_316 ( .B1(net_2073), .ZN(net_1729), .B2(net_1728), .A(net_931) );
INV_X8 inst_1174 ( .ZN(net_2017), .A(net_2012) );
NAND2_X2 inst_1023 ( .A1(net_1997), .ZN(net_553), .A2(net_527) );
OAI21_X2 inst_383 ( .A(net_1941), .B2(net_1356), .ZN(net_1353), .B1(net_1337) );
AOI22_X2 inst_2428 ( .B2(net_2145), .B1(net_1974), .ZN(net_1802), .A1(net_1791), .A2(net_320) );
CLKBUF_X2 inst_4132 ( .A(net_3923), .Z(net_3924) );
CLKBUF_X2 inst_3186 ( .A(net_2977), .Z(net_2978) );
NAND3_X2 inst_678 ( .A1(net_1918), .ZN(net_538), .A2(net_537), .A3(net_420) );
NAND2_X1 inst_1124 ( .ZN(net_530), .A1(net_529), .A2(x3843) );
CLKBUF_X2 inst_4086 ( .A(net_3877), .Z(net_3878) );
CLKBUF_X2 inst_3762 ( .A(net_3553), .Z(net_3554) );
NAND2_X2 inst_854 ( .A1(net_1741), .ZN(net_1236), .A2(net_1235) );
CLKBUF_X2 inst_3259 ( .A(net_3050), .Z(net_3051) );
AOI21_X2 inst_2555 ( .ZN(net_1951), .A(net_1950), .B2(net_1948), .B1(net_608) );
CLKBUF_X2 inst_3375 ( .A(net_2572), .Z(net_3167) );
OAI22_X2 inst_234 ( .B2(net_2287), .B1(net_1865), .A1(net_951), .ZN(net_937), .A2(net_936) );
CLKBUF_X2 inst_3678 ( .A(net_3469), .Z(net_3470) );
CLKBUF_X2 inst_3979 ( .A(net_3770), .Z(net_3771) );
DFF_X1 inst_1946 ( .Q(net_2112), .D(net_1029), .CK(net_3001) );
CLKBUF_X2 inst_3714 ( .A(net_3505), .Z(net_3506) );
INV_X4 inst_1304 ( .ZN(net_1730), .A(net_1728) );
CLKBUF_X2 inst_3429 ( .A(net_3220), .Z(net_3221) );
INV_X4 inst_1328 ( .A(net_2011), .ZN(net_1962) );
CLKBUF_X2 inst_3457 ( .A(net_3248), .Z(net_3249) );
NAND3_X2 inst_688 ( .A3(net_2105), .ZN(net_1653), .A1(net_1652), .A2(net_1649) );
DFF_X2 inst_1749 ( .QN(net_1843), .D(net_1417), .CK(net_3744) );
AOI21_X2 inst_2549 ( .ZN(net_494), .A(net_453), .B1(net_449), .B2(net_373) );
CLKBUF_X2 inst_3292 ( .A(net_3083), .Z(net_3084) );
DFF_X2 inst_1776 ( .QN(net_2378), .D(net_883), .CK(net_3891) );
CLKBUF_X2 inst_3641 ( .A(net_3432), .Z(net_3433) );
AOI22_X2 inst_2335 ( .B2(net_2132), .A1(net_2038), .A2(net_1566), .B1(net_979), .ZN(net_829) );
AOI22_X2 inst_2387 ( .A1(net_2195), .B1(net_839), .ZN(net_629), .A2(net_471), .B2(net_74) );
NAND2_X2 inst_919 ( .A1(net_1638), .ZN(net_1102), .A2(net_823) );
NOR2_X2 inst_598 ( .A2(net_2251), .ZN(net_1887), .A1(net_520) );
DFF_X1 inst_1916 ( .D(net_1294), .QN(net_86), .CK(net_3685) );
CLKBUF_X2 inst_3156 ( .A(net_2567), .Z(net_2948) );
CLKBUF_X2 inst_2747 ( .A(net_2538), .Z(net_2539) );
NAND2_X2 inst_840 ( .A1(net_1840), .ZN(net_1273), .A2(net_285) );
INV_X2 inst_1624 ( .ZN(net_196), .A(x4524) );
INV_X4 inst_1220 ( .A(net_1874), .ZN(net_499) );
INV_X2 inst_1456 ( .A(net_2363), .ZN(net_1235) );
DFF_X2 inst_1797 ( .QN(net_1581), .D(net_396), .CK(net_3994) );
CLKBUF_X2 inst_3167 ( .A(net_2958), .Z(net_2959) );
CLKBUF_X2 inst_2708 ( .A(net_2499), .Z(net_2500) );
CLKBUF_X2 inst_4195 ( .A(net_3986), .Z(net_3987) );
CLKBUF_X2 inst_3530 ( .A(net_3321), .Z(net_3322) );
AND2_X4 inst_2592 ( .ZN(net_2081), .A2(net_1186), .A1(net_1184) );
OAI21_X2 inst_325 ( .B2(net_2312), .B1(net_1507), .ZN(net_1505), .A(net_1472) );
INV_X4 inst_1197 ( .ZN(net_740), .A(net_534) );
CLKBUF_X2 inst_3116 ( .A(net_2907), .Z(net_2908) );
NAND2_X2 inst_955 ( .A1(net_1829), .ZN(net_930), .A2(net_298) );
CLKBUF_X2 inst_4199 ( .A(net_3990), .Z(net_3991) );
SDFF_X2 inst_114 ( .SE(net_488), .Q(net_173), .D(net_173), .CK(net_2942), .SI(x4353) );
AOI22_X2 inst_2278 ( .ZN(net_1705), .A2(net_1549), .A1(net_1000), .B1(net_999), .B2(net_355) );
NOR2_X2 inst_617 ( .A2(net_2175), .ZN(net_2043), .A1(net_2042) );
CLKBUF_X2 inst_4150 ( .A(net_3712), .Z(net_3942) );
NOR2_X2 inst_534 ( .A2(net_2434), .A1(net_1747), .ZN(net_1360) );
NAND2_X2 inst_1057 ( .A2(net_1914), .A1(net_1729), .ZN(net_1685) );
CLKBUF_X2 inst_2842 ( .A(net_2633), .Z(net_2634) );
DFFR_X2 inst_2084 ( .D(net_1723), .QN(net_1576), .RN(net_1347), .CK(net_3514) );
CLKBUF_X2 inst_2836 ( .A(net_2627), .Z(net_2628) );
CLKBUF_X2 inst_3792 ( .A(net_3466), .Z(net_3584) );
NAND2_X4 inst_748 ( .ZN(net_1973), .A2(net_1927), .A1(net_1665) );
CLKBUF_X2 inst_2839 ( .A(net_2630), .Z(net_2631) );
CLKBUF_X2 inst_2770 ( .A(net_2561), .Z(net_2562) );
CLKBUF_X2 inst_3444 ( .A(net_2540), .Z(net_3236) );
NAND2_X2 inst_803 ( .A2(net_1672), .ZN(net_1310), .A1(net_1280) );
DFF_X1 inst_1986 ( .Q(net_2150), .D(net_1047), .CK(net_2971) );
CLKBUF_X2 inst_2909 ( .A(net_2700), .Z(net_2701) );
DFF_X1 inst_1949 ( .Q(net_2115), .D(net_1083), .CK(net_3400) );
AOI22_X2 inst_2348 ( .B1(net_2197), .A1(net_2038), .A2(net_1561), .B2(net_1534), .ZN(net_816) );
CLKBUF_X2 inst_3135 ( .A(net_2524), .Z(net_2927) );
CLKBUF_X2 inst_4021 ( .A(net_3812), .Z(net_3813) );
NAND3_X2 inst_701 ( .ZN(net_2047), .A1(net_2045), .A2(net_1829), .A3(net_472) );
NAND3_X2 inst_662 ( .A1(net_1986), .A2(net_1808), .ZN(net_1080), .A3(net_809) );
CLKBUF_X2 inst_2911 ( .A(net_2702), .Z(net_2703) );
INV_X2 inst_1533 ( .A(net_2303), .ZN(net_274) );
AOI22_X2 inst_2380 ( .B1(net_1915), .A1(net_1718), .B2(net_794), .ZN(net_645), .A2(net_373) );
CLKBUF_X2 inst_3495 ( .A(net_2742), .Z(net_3287) );
DFF_X1 inst_1859 ( .QN(net_2440), .D(net_1398), .CK(net_3936) );
INV_X2 inst_1465 ( .A(net_2348), .ZN(net_1205) );
SDFF_X2 inst_53 ( .SE(net_1768), .SI(net_1536), .Q(net_71), .D(net_71), .CK(net_3236) );
NAND2_X2 inst_1007 ( .A2(net_2131), .A1(net_979), .ZN(net_665) );
CLKBUF_X2 inst_2815 ( .A(net_2606), .Z(net_2607) );
CLKBUF_X2 inst_4208 ( .A(net_3999), .Z(net_4000) );
CLKBUF_X2 inst_3605 ( .A(net_3396), .Z(net_3397) );
AND2_X2 inst_2614 ( .A1(net_609), .A2(x6968), .ZN(x665) );
CLKBUF_X2 inst_3337 ( .A(net_3128), .Z(net_3129) );
CLKBUF_X2 inst_4215 ( .A(net_3913), .Z(net_4007) );
NAND3_X2 inst_651 ( .ZN(net_1232), .A1(net_1191), .A2(net_611), .A3(net_532) );
CLKBUF_X2 inst_4090 ( .A(net_3881), .Z(net_3882) );
NAND2_X2 inst_999 ( .A1(net_1669), .ZN(net_761), .A2(net_307) );
DFFR_X1 inst_2111 ( .QN(net_2302), .RN(net_1347), .D(net_947), .CK(net_2756) );
CLKBUF_X2 inst_2883 ( .A(net_2674), .Z(net_2675) );
INV_X8 inst_1157 ( .A(net_2009), .ZN(net_1782) );
DFF_X1 inst_1846 ( .QN(net_2341), .D(net_1487), .CK(net_3415) );
DFFR_X1 inst_2139 ( .QN(net_2272), .RN(net_1347), .D(net_721), .CK(net_3013) );
INV_X2 inst_1463 ( .ZN(net_366), .A(net_315) );
OAI22_X2 inst_186 ( .B1(net_1428), .A1(net_529), .B2(net_234), .A2(net_88), .ZN(x1663) );
CLKBUF_X2 inst_3528 ( .A(net_3319), .Z(net_3320) );
NAND2_X4 inst_759 ( .A2(net_2198), .ZN(net_2037), .A1(net_1979) );
CLKBUF_X2 inst_3071 ( .A(net_2862), .Z(net_2863) );
DFF_X1 inst_2061 ( .Q(net_2246), .D(net_460), .CK(net_3604) );
CLKBUF_X2 inst_3685 ( .A(net_3476), .Z(net_3477) );
NAND2_X2 inst_863 ( .A1(net_1838), .ZN(net_1220), .A2(net_933) );
INV_X2 inst_1472 ( .A(net_1526), .ZN(net_718) );
INV_X2 inst_1385 ( .ZN(net_619), .A(net_618) );
INV_X2 inst_1573 ( .A(net_2245), .ZN(net_461) );
INV_X4 inst_1183 ( .ZN(net_1443), .A(net_1367) );
CLKBUF_X2 inst_3784 ( .A(net_3575), .Z(net_3576) );
INV_X2 inst_1390 ( .A(net_585), .ZN(x962) );
CLKBUF_X2 inst_3586 ( .A(net_3377), .Z(net_3378) );
OAI22_X2 inst_229 ( .B2(net_2304), .B1(net_1865), .A1(net_1597), .ZN(net_945), .A2(net_718) );
AOI22_X2 inst_2282 ( .A1(net_1996), .B1(net_1749), .A2(net_1552), .ZN(net_981), .B2(net_154) );
INV_X2 inst_1489 ( .A(net_2317), .ZN(net_1264) );
AOI22_X2 inst_2415 ( .B2(net_2143), .B1(net_1974), .A1(net_1789), .ZN(net_1661), .A2(net_343) );
AOI22_X2 inst_2262 ( .B1(net_1768), .ZN(net_1690), .B2(net_1580), .A1(net_1001), .A2(net_815) );
CLKBUF_X2 inst_3288 ( .A(net_3079), .Z(net_3080) );
INV_X8 inst_1160 ( .ZN(net_1828), .A(net_1827) );
INV_X2 inst_1394 ( .A(net_581), .ZN(x996) );
DFFR_X1 inst_2131 ( .QN(net_2262), .RN(net_1347), .D(net_741), .CK(net_2607) );
DFF_X2 inst_1808 ( .Q(net_1522), .CK(net_2717), .D(x5269) );
NAND2_X2 inst_988 ( .A2(net_1564), .A1(net_961), .ZN(net_851) );
DFF_X1 inst_1876 ( .D(net_1328), .QN(net_91), .CK(net_3718) );
OAI22_X2 inst_169 ( .B1(net_1406), .A1(net_1405), .B2(net_187), .A2(net_121), .ZN(x491) );
OAI21_X2 inst_421 ( .ZN(net_496), .A(net_477), .B1(net_429), .B2(net_396) );
INV_X4 inst_1315 ( .A(net_2065), .ZN(net_1832) );
NOR2_X2 inst_555 ( .A2(net_2291), .A1(net_1848), .ZN(net_557) );
NAND2_X2 inst_816 ( .ZN(net_1297), .A2(net_1256), .A1(net_1214) );
AOI22_X2 inst_2392 ( .B1(net_839), .ZN(net_624), .A1(net_623), .A2(net_374), .B2(net_75) );
CLKBUF_X2 inst_2798 ( .A(net_2589), .Z(net_2590) );
CLKBUF_X2 inst_3667 ( .A(net_3458), .Z(net_3459) );
INV_X4 inst_1184 ( .A(net_1739), .ZN(net_1194) );
NAND3_X2 inst_656 ( .A1(net_1721), .ZN(net_1137), .A3(net_994), .A2(net_985) );
SDFF_X2 inst_45 ( .SE(net_1768), .SI(net_1530), .Q(net_76), .D(net_76), .CK(net_3449) );
NAND2_X2 inst_1108 ( .ZN(net_2027), .A1(net_2025), .A2(net_1777) );
OAI211_X2 inst_458 ( .C2(net_2359), .C1(net_1639), .ZN(net_1093), .A(net_816), .B(net_671) );
CLKBUF_X2 inst_3093 ( .A(net_2884), .Z(net_2885) );
INV_X2 inst_1562 ( .ZN(net_238), .A(x4096) );
CLKBUF_X2 inst_4148 ( .A(net_3939), .Z(net_3940) );
DFF_X1 inst_1922 ( .QN(net_2434), .D(net_1713), .CK(net_3904) );
CLKBUF_X2 inst_3361 ( .A(net_3152), .Z(net_3153) );
NAND2_X4 inst_741 ( .A1(net_1965), .ZN(net_1959), .A2(net_1958) );
CLKBUF_X2 inst_3170 ( .A(net_2690), .Z(net_2962) );
CLKBUF_X2 inst_3232 ( .A(net_3023), .Z(net_3024) );
CLKBUF_X2 inst_3991 ( .A(net_3694), .Z(net_3783) );
CLKBUF_X2 inst_3343 ( .A(net_2684), .Z(net_3135) );
INV_X4 inst_1350 ( .A(net_2412), .ZN(net_2191) );
CLKBUF_X2 inst_4140 ( .A(net_3931), .Z(net_3932) );
CLKBUF_X2 inst_3012 ( .A(net_2803), .Z(net_2804) );
AND2_X2 inst_2635 ( .A1(net_594), .A2(x4283), .ZN(x1739) );
INV_X2 inst_1543 ( .A(net_2304), .ZN(net_283) );
CLKBUF_X2 inst_2828 ( .A(net_2619), .Z(net_2620) );
CLKBUF_X2 inst_4219 ( .A(net_4010), .Z(net_4011) );
CLKBUF_X2 inst_2801 ( .A(net_2592), .Z(net_2593) );
NAND2_X2 inst_1118 ( .ZN(net_2078), .A2(net_2077), .A1(net_1184) );
AOI22_X2 inst_2303 ( .A2(net_2139), .B1(net_2096), .A1(net_1769), .B2(net_1521), .ZN(net_906) );
CLKBUF_X2 inst_3363 ( .A(net_3154), .Z(net_3155) );
CLKBUF_X2 inst_3877 ( .A(net_3668), .Z(net_3669) );
CLKBUF_X2 inst_2666 ( .A(net_2457), .Z(net_2458) );
OAI211_X2 inst_473 ( .C1(net_1052), .ZN(net_1037), .C2(net_1036), .A(net_902), .B(net_872) );
INV_X8 inst_1131 ( .A(net_1760), .ZN(net_1356) );
INV_X2 inst_1357 ( .A(net_1410), .ZN(x132) );
NAND3_X2 inst_691 ( .A1(net_1999), .A3(net_1977), .ZN(net_1766), .A2(net_612) );
AOI22_X2 inst_2211 ( .A2(net_2396), .B2(net_2141), .A1(net_1916), .B1(net_1915), .ZN(net_1469) );
CLKBUF_X2 inst_3771 ( .A(net_2674), .Z(net_3563) );
CLKBUF_X2 inst_3083 ( .A(net_2874), .Z(net_2875) );
INV_X16 inst_1695 ( .A(net_1896), .ZN(net_1863) );
NAND2_X2 inst_770 ( .A2(net_2436), .A1(net_2168), .ZN(x1285) );
NOR2_X2 inst_565 ( .A1(net_537), .ZN(net_421), .A2(net_420) );
NOR2_X1 inst_622 ( .A2(net_2355), .A1(net_1843), .ZN(net_325) );
DFF_X1 inst_1971 ( .Q(net_2137), .D(net_1100), .CK(net_3392) );
INV_X2 inst_1404 ( .A(net_572), .ZN(x1097) );
CLKBUF_X2 inst_2989 ( .A(net_2705), .Z(net_2781) );
CLKBUF_X2 inst_3479 ( .A(net_3270), .Z(net_3271) );
OAI21_X2 inst_409 ( .ZN(net_765), .B1(net_650), .A(net_639), .B2(net_376) );
AOI22_X2 inst_2288 ( .A1(net_1996), .B1(net_1749), .A2(net_1545), .ZN(net_974), .B2(net_147) );
INV_X4 inst_1339 ( .ZN(net_2033), .A(net_2032) );
DFF_X2 inst_1834 ( .Q(net_1520), .CK(net_2712), .D(x5247) );
CLKBUF_X2 inst_3575 ( .A(net_3366), .Z(net_3367) );
CLKBUF_X2 inst_3506 ( .A(net_3297), .Z(net_3298) );
CLKBUF_X2 inst_3654 ( .A(net_2732), .Z(net_3446) );
NAND2_X2 inst_977 ( .A2(net_1570), .A1(net_961), .ZN(net_862) );
AOI22_X2 inst_2228 ( .B2(net_2153), .A1(net_2040), .B1(net_1450), .ZN(net_1448), .A2(net_309) );
CLKBUF_X2 inst_3574 ( .A(net_3290), .Z(net_3366) );
NAND2_X4 inst_768 ( .ZN(net_2168), .A1(net_459), .A2(x3865) );
NAND3_X2 inst_663 ( .A2(net_1661), .ZN(net_1079), .A1(net_971), .A3(net_808) );
DFFR_X1 inst_2121 ( .QN(net_2285), .RN(net_1347), .D(net_940), .CK(net_3117) );
OAI22_X2 inst_297 ( .A2(net_2232), .B1(net_1895), .A1(net_1615), .B2(net_183), .ZN(x1956) );
CLKBUF_X2 inst_3227 ( .A(net_2653), .Z(net_3019) );
INV_X2 inst_1395 ( .A(net_580), .ZN(x1007) );
AOI222_X2 inst_2477 ( .C1(net_2016), .A2(net_1546), .A1(net_590), .B1(net_589), .ZN(net_559), .B2(net_148), .C2(x5868) );
CLKBUF_X2 inst_3436 ( .A(net_3139), .Z(net_3228) );
CLKBUF_X2 inst_3494 ( .A(net_3285), .Z(net_3286) );
CLKBUF_X2 inst_4224 ( .A(net_4015), .Z(net_4016) );
DFF_X1 inst_1875 ( .D(net_1331), .QN(net_98), .CK(net_3690) );
CLKBUF_X2 inst_3351 ( .A(net_3142), .Z(net_3143) );
DFF_X1 inst_1867 ( .D(net_1359), .QN(net_93), .CK(net_3908) );
CLKBUF_X2 inst_3190 ( .A(net_2686), .Z(net_2982) );
OAI22_X2 inst_162 ( .A1(net_1408), .B1(net_1407), .B2(net_208), .A2(net_134), .ZN(x272) );
CLKBUF_X2 inst_3308 ( .A(net_3073), .Z(net_3100) );
AOI22_X2 inst_2290 ( .A1(net_1996), .B1(net_1749), .A2(net_1543), .ZN(net_972), .B2(net_145) );
CLKBUF_X2 inst_3397 ( .A(net_3188), .Z(net_3189) );
CLKBUF_X2 inst_2829 ( .A(net_2620), .Z(net_2621) );
CLKBUF_X2 inst_3819 ( .A(net_3610), .Z(net_3611) );
CLKBUF_X2 inst_4233 ( .A(net_4024), .Z(net_4025) );
CLKBUF_X2 inst_3668 ( .A(net_3459), .Z(net_3460) );
CLKBUF_X2 inst_3968 ( .A(net_3658), .Z(net_3760) );
CLKBUF_X2 inst_3342 ( .A(net_3133), .Z(net_3134) );
NAND2_X2 inst_1098 ( .ZN(net_1945), .A1(net_1834), .A2(net_1777) );
AND2_X2 inst_2621 ( .A1(net_594), .A2(x7314), .ZN(x807) );
CLKBUF_X2 inst_4149 ( .A(net_3940), .Z(net_3941) );
CLKBUF_X2 inst_3895 ( .A(net_3686), .Z(net_3687) );
AOI22_X2 inst_2443 ( .B1(net_2096), .ZN(net_1921), .A2(net_1919), .A1(net_1769), .B2(net_1528) );
NAND2_X4 inst_723 ( .A1(net_1291), .ZN(net_457), .A2(net_365) );
OAI22_X2 inst_303 ( .A2(net_2213), .B1(net_1895), .A1(net_1403), .B2(net_181), .ZN(x2333) );
NOR2_X2 inst_618 ( .ZN(net_2192), .A1(net_2191), .A2(net_1584) );
AOI22_X2 inst_2444 ( .B2(net_2132), .ZN(net_2060), .B1(net_1929), .A1(net_655), .A2(net_289) );
CLKBUF_X2 inst_3893 ( .A(net_3684), .Z(net_3685) );
INV_X2 inst_1647 ( .A(net_2297), .ZN(net_288) );
CLKBUF_X2 inst_3263 ( .A(net_2994), .Z(net_3055) );
CLKBUF_X2 inst_3057 ( .A(net_2848), .Z(net_2849) );
INV_X4 inst_1275 ( .A(net_1575), .ZN(net_303) );
AOI222_X2 inst_2462 ( .C1(net_2016), .A2(net_1545), .A1(net_590), .B1(net_589), .ZN(net_574), .B2(net_147), .C2(x5892) );
OAI211_X2 inst_474 ( .C1(net_1052), .ZN(net_1035), .A(net_901), .B(net_871), .C2(net_287) );
XNOR2_X2 inst_26 ( .B(net_2433), .A(net_2359), .ZN(net_1141) );
DFF_X1 inst_2067 ( .Q(net_2343), .D(net_2312), .CK(net_3139) );
NOR2_X1 inst_626 ( .A1(net_2357), .A2(net_315), .ZN(net_268) );
INV_X2 inst_1376 ( .A(net_1008), .ZN(x2706) );
CLKBUF_X2 inst_2882 ( .A(net_2673), .Z(net_2674) );
CLKBUF_X2 inst_2777 ( .A(net_2568), .Z(net_2569) );
AOI222_X2 inst_2446 ( .C1(net_2016), .A2(net_1560), .ZN(net_610), .A1(net_590), .B1(net_589), .B2(net_162), .C2(x5527) );
CLKBUF_X2 inst_3765 ( .A(net_3556), .Z(net_3557) );
INV_X2 inst_1659 ( .A(net_2368), .ZN(net_1225) );
CLKBUF_X2 inst_4218 ( .A(net_4009), .Z(net_4010) );
NAND2_X2 inst_798 ( .A2(net_1673), .ZN(net_1315), .A1(net_1266) );
OAI21_X2 inst_398 ( .B1(net_1829), .ZN(net_1109), .B2(net_939), .A(net_926) );
OAI21_X2 inst_436 ( .B2(net_2414), .A(net_2174), .B1(net_2074), .ZN(net_2029) );
INV_X2 inst_1434 ( .A(net_1524), .ZN(net_713) );
DFF_X1 inst_1886 ( .D(net_1298), .QN(net_110), .CK(net_3826) );
CLKBUF_X2 inst_3705 ( .A(net_3496), .Z(net_3497) );
AOI22_X2 inst_2231 ( .ZN(net_1411), .A2(net_408), .A1(net_142), .B2(x6236), .B1(x5995) );
OR2_X1 inst_144 ( .A1(net_1404), .A2(x6096), .ZN(x83) );
INV_X2 inst_1457 ( .A(net_2426), .ZN(net_398) );
INV_X2 inst_1438 ( .A(net_1534), .ZN(net_950) );
DFF_X2 inst_1818 ( .Q(net_1514), .CK(net_2596), .D(x5755) );
CLKBUF_X2 inst_3662 ( .A(net_3453), .Z(net_3454) );
DFF_X2 inst_1766 ( .QN(net_2382), .D(net_2199), .CK(net_3895) );
CLKBUF_X2 inst_2670 ( .A(net_2461), .Z(net_2462) );
NAND2_X2 inst_880 ( .ZN(net_1176), .A2(net_1169), .A1(net_767) );
CLKBUF_X2 inst_2974 ( .A(net_2765), .Z(net_2766) );
DFF_X1 inst_1895 ( .D(net_1308), .QN(net_139), .CK(net_3484) );
CLKBUF_X2 inst_2681 ( .A(net_2472), .Z(net_2473) );
CLKBUF_X2 inst_2730 ( .A(net_2521), .Z(net_2522) );
CLKBUF_X2 inst_3445 ( .A(net_2646), .Z(net_3237) );
NAND2_X4 inst_737 ( .A1(net_2024), .ZN(net_1914), .A2(net_84) );
NAND2_X2 inst_876 ( .A1(net_1838), .ZN(net_1202), .A2(net_1201) );
CLKBUF_X2 inst_2979 ( .A(net_2643), .Z(net_2771) );
NOR2_X2 inst_545 ( .ZN(net_920), .A1(net_634), .A2(net_607) );
CLKBUF_X2 inst_3972 ( .A(net_3698), .Z(net_3764) );
INV_X2 inst_1388 ( .A(net_587), .ZN(x950) );
AOI22_X2 inst_2433 ( .B2(net_2159), .B1(net_1974), .ZN(net_1807), .A1(net_1789), .A2(net_344) );
CLKBUF_X2 inst_2699 ( .A(net_2490), .Z(net_2491) );
CLKBUF_X2 inst_3517 ( .A(net_3245), .Z(net_3309) );
NOR2_X2 inst_562 ( .A2(net_1716), .ZN(net_445), .A1(net_377) );
AOI222_X1 inst_2480 ( .B1(net_1995), .A1(net_1749), .B2(net_1571), .ZN(net_1021), .C1(net_1020), .A2(net_173), .C2(x3277) );
INV_X2 inst_1372 ( .A(net_1012), .ZN(x2471) );
CLKBUF_X2 inst_3396 ( .A(net_3187), .Z(net_3188) );
INV_X2 inst_1360 ( .ZN(net_1148), .A(net_1147) );
OAI211_X2 inst_466 ( .C1(net_1054), .ZN(net_1047), .A(net_908), .B(net_862), .C2(net_410) );
CLKBUF_X2 inst_2761 ( .A(net_2552), .Z(net_2553) );
CLKBUF_X2 inst_3981 ( .A(net_3772), .Z(net_3773) );
NAND2_X2 inst_989 ( .ZN(net_1658), .A1(net_1596), .A2(net_1521) );
AOI22_X2 inst_2283 ( .A1(net_1996), .B1(net_1749), .A2(net_1551), .ZN(net_980), .B2(net_153) );
CLKBUF_X2 inst_3038 ( .A(net_2829), .Z(net_2830) );
NAND2_X2 inst_858 ( .A1(net_1741), .ZN(net_1229), .A2(net_933) );
CLKBUF_X2 inst_3659 ( .A(net_3450), .Z(net_3451) );
CLKBUF_X2 inst_3604 ( .A(net_3395), .Z(net_3396) );
NAND2_X2 inst_1109 ( .A1(net_2074), .ZN(net_2028), .A2(net_1870) );
CLKBUF_X2 inst_3864 ( .A(net_2614), .Z(net_3656) );
CLKBUF_X2 inst_4209 ( .A(net_4000), .Z(net_4001) );
CLKBUF_X2 inst_3037 ( .A(net_2538), .Z(net_2829) );
SDFF_X2 inst_54 ( .SE(net_1768), .SI(net_1525), .Q(net_81), .D(net_81), .CK(net_3198) );
AOI222_X2 inst_2468 ( .C1(net_2016), .A2(net_1550), .A1(net_590), .B1(net_589), .ZN(net_568), .B2(net_152), .C2(x5779) );
CLKBUF_X2 inst_2936 ( .A(net_2727), .Z(net_2728) );
INV_X4 inst_1314 ( .A(net_2010), .ZN(net_1826) );
INV_X2 inst_1420 ( .ZN(net_603), .A(net_539) );
INV_X2 inst_1482 ( .A(net_1527), .ZN(net_720) );
INV_X8 inst_1156 ( .A(net_1840), .ZN(net_1746) );
CLKBUF_X2 inst_3378 ( .A(net_3169), .Z(net_3170) );
CLKBUF_X2 inst_3484 ( .A(net_3275), .Z(net_3276) );
CLKBUF_X2 inst_4062 ( .A(net_3853), .Z(net_3854) );
NAND2_X2 inst_942 ( .ZN(net_1044), .A1(net_963), .A2(net_885) );
INV_X4 inst_1295 ( .ZN(net_790), .A(net_65) );
DFF_X1 inst_1880 ( .D(net_1326), .QN(net_102), .CK(net_3827) );
CLKBUF_X2 inst_4108 ( .A(net_2991), .Z(net_3900) );
OAI22_X2 inst_262 ( .B2(net_2255), .A2(net_938), .A1(net_740), .ZN(net_700), .B1(net_534) );
CLKBUF_X2 inst_3829 ( .A(net_3620), .Z(net_3621) );
CLKBUF_X2 inst_3630 ( .A(net_3421), .Z(net_3422) );
NOR3_X2 inst_497 ( .A2(net_2366), .A1(net_2365), .A3(net_2364), .ZN(net_386) );
NAND2_X2 inst_1035 ( .A2(net_2366), .ZN(net_404), .A1(net_364) );
INV_X4 inst_1335 ( .ZN(net_2015), .A(net_2012) );
CLKBUF_X2 inst_3845 ( .A(net_3627), .Z(net_3637) );
CLKBUF_X2 inst_3637 ( .A(net_3428), .Z(net_3429) );
CLKBUF_X2 inst_3128 ( .A(net_2643), .Z(net_2920) );
DFF_X1 inst_1883 ( .D(net_1322), .QN(net_89), .CK(net_3928) );
NAND2_X2 inst_1078 ( .A1(net_2104), .ZN(net_1819), .A2(net_285) );
AOI21_X2 inst_2517 ( .B2(net_2115), .B1(net_1915), .ZN(net_1399), .A(net_1365) );
CLKBUF_X2 inst_3621 ( .A(net_3412), .Z(net_3413) );
NAND2_X2 inst_864 ( .A1(net_1838), .ZN(net_1219), .A2(net_1218) );
OAI21_X2 inst_418 ( .B2(net_1718), .ZN(net_682), .A(net_681), .B1(net_600) );
SDFF_X2 inst_86 ( .Q(net_1564), .D(net_1564), .SE(net_491), .CK(net_2669), .SI(x7061) );
CLKBUF_X2 inst_4183 ( .A(net_3974), .Z(net_3975) );
NAND2_X2 inst_949 ( .ZN(net_990), .A2(net_844), .A1(net_751) );
CLKBUF_X2 inst_3283 ( .A(net_3074), .Z(net_3075) );
CLKBUF_X2 inst_3557 ( .A(net_3348), .Z(net_3349) );
NAND2_X2 inst_1039 ( .A1(net_2198), .A2(net_2035), .ZN(net_1618) );
DFF_X1 inst_1992 ( .Q(net_2156), .D(net_1025), .CK(net_3373) );
CLKBUF_X2 inst_3961 ( .A(net_3752), .Z(net_3753) );
NAND2_X4 inst_714 ( .A1(net_2198), .ZN(net_556), .A2(net_543) );
CLKBUF_X2 inst_3730 ( .A(net_3521), .Z(net_3522) );
CLKBUF_X2 inst_2895 ( .A(net_2686), .Z(net_2687) );
CLKBUF_X2 inst_3005 ( .A(net_2796), .Z(net_2797) );
CLKBUF_X2 inst_3598 ( .A(net_3141), .Z(net_3390) );
CLKBUF_X2 inst_4048 ( .A(net_3777), .Z(net_3840) );
DFF_X2 inst_1826 ( .Q(net_1539), .CK(net_2632), .D(x5628) );
DFFR_X1 inst_2109 ( .QN(net_2299), .RN(net_1347), .D(net_948), .CK(net_2519) );
CLKBUF_X2 inst_4003 ( .A(net_3344), .Z(net_3795) );
DFF_X1 inst_2020 ( .QN(net_2213), .D(net_1060), .CK(net_3327) );
NAND2_X2 inst_1061 ( .A1(net_1954), .ZN(net_1720), .A2(net_1562) );
INV_X8 inst_1177 ( .ZN(net_2102), .A(net_2101) );
AOI22_X2 inst_2326 ( .A2(net_2155), .B1(net_2096), .A1(net_1769), .B2(net_1516), .ZN(net_879) );
CLKBUF_X2 inst_2820 ( .A(net_2611), .Z(net_2612) );
AOI21_X2 inst_2548 ( .B2(net_646), .ZN(net_495), .B1(net_475), .A(net_450) );
SDFF_X2 inst_72 ( .Q(net_1553), .D(net_1553), .SE(net_396), .CK(net_2910), .SI(x7329) );
AOI22_X2 inst_2404 ( .B2(net_2242), .B1(net_2197), .ZN(net_1632), .A1(net_1621), .A2(net_537) );
INV_X2 inst_1578 ( .ZN(net_228), .A(x4375) );
INV_X2 inst_1634 ( .ZN(net_188), .A(x6372) );
INV_X2 inst_1666 ( .ZN(net_1778), .A(x3190) );
CLKBUF_X2 inst_3542 ( .A(net_2974), .Z(net_3334) );
NAND2_X4 inst_735 ( .A2(net_1902), .A1(net_1901), .ZN(net_1750) );
INV_X2 inst_1529 ( .A(net_2302), .ZN(net_308) );
SDFF_X2 inst_115 ( .SE(net_488), .Q(net_163), .D(net_163), .CK(net_2728), .SI(x4578) );
INV_X2 inst_1653 ( .ZN(net_180), .A(x4258) );
CLKBUF_X2 inst_3726 ( .A(net_3517), .Z(net_3518) );
CLKBUF_X2 inst_3045 ( .A(net_2480), .Z(net_2837) );
INV_X2 inst_1582 ( .ZN(net_225), .A(x6367) );
CLKBUF_X2 inst_2984 ( .A(net_2725), .Z(net_2776) );
OAI22_X2 inst_175 ( .B1(net_1428), .A1(net_529), .B2(net_220), .A2(net_101), .ZN(x1474) );
CLKBUF_X2 inst_3258 ( .A(net_3049), .Z(net_3050) );
DFF_X2 inst_1737 ( .QN(net_2317), .D(net_1499), .CK(net_3549) );
DFF_X2 inst_1805 ( .Q(net_1527), .CK(net_2718), .D(x5386) );
DFF_X1 inst_1840 ( .QN(net_2338), .D(net_1491), .CK(net_2979) );
CLKBUF_X2 inst_2995 ( .A(net_2722), .Z(net_2787) );
CLKBUF_X2 inst_3563 ( .A(net_3354), .Z(net_3355) );
OR2_X2 inst_133 ( .A2(net_1904), .A1(net_1579), .ZN(net_439) );
INV_X4 inst_1263 ( .A(net_2323), .ZN(net_331) );
CLKBUF_X2 inst_2752 ( .A(net_2543), .Z(net_2544) );
CLKBUF_X2 inst_3330 ( .A(net_3121), .Z(net_3122) );
INV_X8 inst_1149 ( .A(net_1865), .ZN(net_1597) );
DFF_X2 inst_1721 ( .QN(net_2337), .D(net_1510), .CK(net_2961) );
INV_X2 inst_1445 ( .A(net_1515), .ZN(net_938) );
INV_X4 inst_1281 ( .A(net_2326), .ZN(net_846) );
INV_X2 inst_1509 ( .A(net_2382), .ZN(net_281) );
CLKBUF_X2 inst_3088 ( .A(net_2879), .Z(net_2880) );
CLKBUF_X2 inst_3990 ( .A(net_3781), .Z(net_3782) );
OR4_X4 inst_126 ( .ZN(net_2190), .A1(net_79), .A2(net_76), .A3(net_72), .A4(net_71) );
CLKBUF_X2 inst_3782 ( .A(net_3573), .Z(net_3574) );
INV_X2 inst_1512 ( .A(net_2367), .ZN(net_1227) );
CLKBUF_X2 inst_3887 ( .A(net_3678), .Z(net_3679) );
INV_X2 inst_1631 ( .A(net_2296), .ZN(net_343) );
CLKBUF_X2 inst_3934 ( .A(net_3556), .Z(net_3726) );
NAND2_X2 inst_948 ( .A2(net_1518), .ZN(net_993), .A1(net_992) );
INV_X8 inst_1140 ( .ZN(net_839), .A(net_525) );
NAND2_X2 inst_1086 ( .A1(net_1975), .ZN(net_1847), .A2(net_1846) );
AND2_X2 inst_2643 ( .A2(net_2421), .ZN(net_436), .A1(net_351) );
INV_X16 inst_1688 ( .A(net_1918), .ZN(net_1450) );
AOI22_X2 inst_2299 ( .B1(net_1768), .ZN(net_1702), .B2(net_1518), .A1(net_999), .A2(net_646) );
DFF_X2 inst_1800 ( .Q(net_1513), .CK(net_2563), .D(x5740) );
OAI211_X4 inst_448 ( .A(net_1943), .C1(net_1741), .B(net_1616), .ZN(net_1294), .C2(net_1115) );
NAND2_X2 inst_914 ( .A1(net_976), .A2(net_779), .ZN(x2950) );
DFF_X1 inst_2002 ( .QN(net_2232), .D(net_1074), .CK(net_3227) );
OAI21_X2 inst_384 ( .A(net_2434), .ZN(net_1352), .B1(net_1168), .B2(net_399) );
INV_X2 inst_1642 ( .ZN(net_183), .A(x4476) );
INV_X4 inst_1252 ( .A(net_2415), .ZN(net_531) );
NOR2_X2 inst_608 ( .A2(net_2267), .ZN(net_1955), .A1(net_520) );
INV_X4 inst_1343 ( .ZN(net_2074), .A(net_2072) );
CLKBUF_X2 inst_3800 ( .A(net_2750), .Z(net_3592) );
NAND2_X2 inst_834 ( .A1(net_1840), .A2(net_1812), .ZN(net_1280) );
CLKBUF_X2 inst_2920 ( .A(net_2593), .Z(net_2712) );
CLKBUF_X2 inst_4054 ( .A(net_3845), .Z(net_3846) );
NAND2_X2 inst_966 ( .A2(net_1558), .A1(net_961), .ZN(net_873) );
OAI22_X2 inst_199 ( .A2(net_2220), .A1(net_1408), .B1(net_1407), .B2(net_218), .ZN(x2220) );
INV_X4 inst_1246 ( .A(net_2340), .ZN(net_1284) );
CLKBUF_X2 inst_2961 ( .A(net_2752), .Z(net_2753) );
CLKBUF_X2 inst_3185 ( .A(net_2976), .Z(net_2977) );
AOI22_X2 inst_2209 ( .A2(net_2393), .B2(net_2140), .A1(net_1916), .ZN(net_1471), .B1(net_1450) );
AOI221_X2 inst_2506 ( .B2(net_2162), .B1(net_1929), .A(net_1889), .ZN(net_911), .C1(net_910), .C2(net_909) );
CLKBUF_X2 inst_2722 ( .A(net_2513), .Z(net_2514) );
INV_X4 inst_1238 ( .A(net_1778), .ZN(net_488) );
CLKBUF_X2 inst_3607 ( .A(net_3398), .Z(net_3399) );
DFF_X1 inst_2029 ( .Q(net_2247), .D(net_849), .CK(net_3059) );
CLKBUF_X2 inst_3402 ( .A(net_2719), .Z(net_3194) );
NAND2_X2 inst_1011 ( .ZN(net_651), .A1(net_650), .A2(net_549) );
NOR2_X2 inst_540 ( .A1(net_2432), .A2(net_2328), .ZN(net_1145) );
CLKBUF_X2 inst_4114 ( .A(net_3905), .Z(net_3906) );
OAI21_X2 inst_404 ( .B2(net_2421), .ZN(net_882), .B1(net_880), .A(net_636) );
AOI22_X2 inst_2356 ( .A1(net_783), .ZN(net_776), .B1(net_775), .A2(net_370), .B2(x3796) );
NAND2_X2 inst_998 ( .A1(net_1669), .ZN(net_762), .A2(net_334) );
CLKBUF_X2 inst_3209 ( .A(net_3000), .Z(net_3001) );
CLKBUF_X2 inst_3160 ( .A(net_2951), .Z(net_2952) );
CLKBUF_X2 inst_2861 ( .A(net_2652), .Z(net_2653) );
SDFF_X2 inst_66 ( .Q(net_1565), .D(net_1565), .SE(net_396), .CK(net_2854), .SI(x7033) );
CLKBUF_X2 inst_3615 ( .A(net_3406), .Z(net_3407) );
CLKBUF_X2 inst_3216 ( .A(net_3007), .Z(net_3008) );
OAI22_X2 inst_273 ( .B2(net_2284), .B1(net_1865), .ZN(net_1605), .A1(net_1597), .A2(net_941) );
OAI22_X2 inst_192 ( .B1(net_1428), .A1(net_529), .B2(net_177), .A2(net_107), .ZN(x1415) );
DFF_X1 inst_1965 ( .Q(net_2131), .D(net_1106), .CK(net_3433) );
CLKBUF_X2 inst_3915 ( .A(net_3706), .Z(net_3707) );
OAI21_X2 inst_366 ( .B2(net_2403), .B1(net_1441), .ZN(net_1425), .A(net_1373) );
AOI22_X2 inst_2418 ( .B2(net_2107), .B1(net_1974), .ZN(net_1792), .A1(net_1791), .A2(net_284) );
CLKBUF_X2 inst_2715 ( .A(net_2506), .Z(net_2507) );
CLKBUF_X2 inst_3540 ( .A(net_3331), .Z(net_3332) );
CLKBUF_X2 inst_4126 ( .A(net_3652), .Z(net_3918) );
CLKBUF_X2 inst_4178 ( .A(net_3969), .Z(net_3970) );
CLKBUF_X2 inst_3547 ( .A(net_3338), .Z(net_3339) );
INV_X2 inst_1574 ( .ZN(net_230), .A(x4949) );
AOI22_X2 inst_2413 ( .B1(net_2197), .ZN(net_1642), .A1(net_1619), .B2(net_1528), .A2(net_1196) );
CLKBUF_X2 inst_3285 ( .A(net_3076), .Z(net_3077) );
OAI22_X2 inst_228 ( .B2(net_2303), .B1(net_1865), .A1(net_951), .ZN(net_946), .A2(net_720) );
NOR4_X2 inst_486 ( .A2(net_2190), .ZN(net_467), .A3(net_347), .A1(net_78), .A4(net_75) );
INV_X4 inst_1240 ( .ZN(net_380), .A(net_314) );
NAND2_X2 inst_1025 ( .A2(net_1932), .ZN(net_615), .A1(net_525) );
NAND3_X1 inst_707 ( .A2(net_2028), .A1(net_1918), .ZN(net_1350), .A3(net_537) );
CLKBUF_X2 inst_3670 ( .A(net_2654), .Z(net_3462) );
OAI22_X2 inst_244 ( .B2(net_2266), .A2(net_950), .A1(net_740), .ZN(net_733), .B1(net_534) );
CLKBUF_X2 inst_2804 ( .A(net_2595), .Z(net_2596) );
INV_X2 inst_1521 ( .ZN(net_264), .A(x6326) );
AND2_X4 inst_2576 ( .A2(net_2168), .A1(net_2053), .ZN(net_783) );
CLKBUF_X2 inst_3079 ( .A(net_2870), .Z(net_2871) );
AND2_X2 inst_2631 ( .A1(net_609), .A2(x7007), .ZN(x679) );
INV_X4 inst_1306 ( .ZN(net_1739), .A(net_1737) );
NAND2_X2 inst_772 ( .A1(net_1966), .ZN(net_1423), .A2(net_1364) );
AOI211_X2 inst_2563 ( .C2(net_2137), .C1(net_1929), .A(net_1878), .B(net_1785), .ZN(net_675) );
CLKBUF_X2 inst_3810 ( .A(net_3601), .Z(net_3602) );
INV_X2 inst_1407 ( .A(net_569), .ZN(x1124) );
CLKBUF_X2 inst_3682 ( .A(net_3473), .Z(net_3474) );
AND2_X2 inst_2636 ( .A1(net_609), .A2(x6880), .ZN(x627) );
OAI21_X1 inst_445 ( .ZN(net_1193), .B1(net_1192), .B2(net_496), .A(net_271) );
SDFF_X2 inst_93 ( .SE(net_488), .Q(net_148), .D(net_148), .CK(net_2542), .SI(x4998) );
CLKBUF_X2 inst_3606 ( .A(net_2731), .Z(net_3398) );
NOR2_X2 inst_606 ( .A2(net_2270), .ZN(net_1946), .A1(net_520) );
CLKBUF_X2 inst_2942 ( .A(net_2658), .Z(net_2734) );
CLKBUF_X2 inst_3761 ( .A(net_3404), .Z(net_3553) );
NAND2_X2 inst_853 ( .A1(net_1841), .ZN(net_1237), .A2(net_364) );
OR2_X2 inst_139 ( .A2(net_2320), .A1(net_2319), .ZN(net_294) );
NAND3_X2 inst_657 ( .A1(net_1720), .ZN(net_1136), .A3(net_993), .A2(net_986) );
INV_X2 inst_1675 ( .ZN(net_1904), .A(x5181) );
NOR2_X2 inst_584 ( .ZN(net_1861), .A1(net_1851), .A2(net_1577) );
INV_X4 inst_1316 ( .A(net_2086), .ZN(net_1831) );
CLKBUF_X2 inst_3433 ( .A(net_3224), .Z(net_3225) );
DFFR_X1 inst_2098 ( .QN(net_2287), .RN(net_1347), .D(net_937), .CK(net_3342) );
OAI211_X2 inst_470 ( .C1(net_1052), .ZN(net_1041), .A(net_897), .B(net_868), .C2(net_400) );
CLKBUF_X2 inst_3551 ( .A(net_3180), .Z(net_3343) );
DFF_X1 inst_1921 ( .D(net_1244), .QN(net_105), .CK(net_3811) );
CLKBUF_X2 inst_4237 ( .A(net_3069), .Z(net_4029) );
OR2_X1 inst_148 ( .A1(net_1427), .A2(x3900), .ZN(x1306) );
DFF_X2 inst_1752 ( .QN(net_2356), .D(net_1442), .CK(net_3741) );
NOR2_X2 inst_554 ( .A2(net_2282), .A1(net_1848), .ZN(net_558) );
INV_X4 inst_1187 ( .ZN(net_1154), .A(net_84) );
OAI22_X2 inst_191 ( .B1(net_1428), .A1(net_529), .B2(net_219), .A2(net_109), .ZN(x1387) );
NAND2_X2 inst_1063 ( .A1(net_1954), .ZN(net_1722), .A2(net_1560) );
CLKBUF_X2 inst_2700 ( .A(net_2469), .Z(net_2492) );
DFF_X1 inst_1917 ( .D(net_1293), .QN(net_85), .CK(net_3683) );
AND2_X2 inst_2638 ( .A1(net_775), .A2(x7264), .ZN(x788) );
CLKBUF_X2 inst_3252 ( .A(net_3043), .Z(net_3044) );
CLKBUF_X2 inst_3235 ( .A(net_3026), .Z(net_3027) );
INV_X8 inst_1167 ( .ZN(net_1978), .A(net_1977) );
CLKBUF_X2 inst_3879 ( .A(net_3670), .Z(net_3671) );
DFFR_X2 inst_2087 ( .RN(net_1347), .D(net_1112), .QN(net_53), .CK(net_3052) );
INV_X4 inst_1303 ( .A(net_1917), .ZN(net_1718) );
NAND2_X2 inst_892 ( .A2(net_1695), .A1(net_1694), .ZN(net_1128) );
INV_X2 inst_1623 ( .ZN(net_197), .A(x6358) );
CLKBUF_X2 inst_2665 ( .A(net_2448), .Z(net_2457) );
CLKBUF_X2 inst_4088 ( .A(net_3879), .Z(net_3880) );
INV_X8 inst_1132 ( .A(net_1787), .ZN(net_931) );
NAND2_X2 inst_968 ( .A2(net_1560), .A1(net_961), .ZN(net_871) );
NAND2_X2 inst_819 ( .A1(net_1840), .ZN(net_1290), .A2(net_397) );
CLKBUF_X2 inst_4100 ( .A(net_3748), .Z(net_3892) );
CLKBUF_X2 inst_3320 ( .A(net_2852), .Z(net_3112) );
INV_X2 inst_1468 ( .A(net_1522), .ZN(net_709) );
CLKBUF_X2 inst_3452 ( .A(net_2938), .Z(net_3244) );
DFF_X2 inst_1803 ( .QN(net_2203), .CK(net_2642), .D(x6650) );
INV_X2 inst_1516 ( .ZN(net_266), .A(x4549) );
CLKBUF_X2 inst_3776 ( .A(net_3567), .Z(net_3568) );
CLKBUF_X2 inst_3153 ( .A(net_2944), .Z(net_2945) );
OAI21_X2 inst_386 ( .B2(net_2353), .B1(net_1842), .ZN(net_1344), .A(net_1343) );
CLKBUF_X2 inst_2814 ( .A(net_2605), .Z(net_2606) );
AND2_X2 inst_2617 ( .A1(net_609), .A2(x7120), .ZN(x722) );
NAND2_X2 inst_936 ( .A2(net_1620), .ZN(net_1064), .A1(net_684) );
CLKBUF_X2 inst_3809 ( .A(net_2885), .Z(net_3601) );
CLKBUF_X2 inst_4004 ( .A(net_3795), .Z(net_3796) );
CLKBUF_X2 inst_3942 ( .A(net_2678), .Z(net_3734) );
CLKBUF_X2 inst_3068 ( .A(net_2859), .Z(net_2860) );
AOI22_X2 inst_2277 ( .ZN(net_1701), .A2(net_1546), .A1(net_1000), .B1(net_999), .B2(net_350) );
CLKBUF_X2 inst_2778 ( .A(net_2569), .Z(net_2570) );
CLKBUF_X2 inst_3798 ( .A(net_3589), .Z(net_3590) );
CLKBUF_X2 inst_4109 ( .A(net_3900), .Z(net_3901) );
CLKBUF_X2 inst_4192 ( .A(net_3983), .Z(net_3984) );
CLKBUF_X2 inst_2962 ( .A(net_2753), .Z(net_2754) );
CLKBUF_X2 inst_3004 ( .A(net_2795), .Z(net_2796) );
CLKBUF_X2 inst_3780 ( .A(net_3571), .Z(net_3572) );
AND2_X2 inst_2647 ( .A1(net_2017), .A2(x3145), .ZN(x2435) );
NAND2_X2 inst_811 ( .ZN(net_1302), .A1(net_1281), .A2(net_1241) );
OAI22_X2 inst_208 ( .A2(net_2221), .A1(net_1408), .B1(net_1404), .B2(net_259), .ZN(x2200) );
CLKBUF_X2 inst_4202 ( .A(net_3993), .Z(net_3994) );
AOI222_X2 inst_2456 ( .C1(net_2015), .A2(net_1567), .A1(net_590), .B1(net_589), .ZN(net_580), .B2(net_169), .C2(x5386) );
CLKBUF_X2 inst_3774 ( .A(net_3401), .Z(net_3566) );
CLKBUF_X2 inst_2710 ( .A(net_2501), .Z(net_2502) );
NAND2_X2 inst_1058 ( .ZN(net_1714), .A1(net_1713), .A2(net_1360) );
CLKBUF_X2 inst_2887 ( .A(net_2678), .Z(net_2679) );
CLKBUF_X2 inst_3909 ( .A(net_3700), .Z(net_3701) );
DFF_X1 inst_1869 ( .D(net_1349), .QN(net_115), .CK(net_3583) );
NAND2_X2 inst_897 ( .A2(net_1707), .A1(net_1706), .ZN(net_1123) );
CLKBUF_X2 inst_3360 ( .A(net_3151), .Z(net_3152) );
CLKBUF_X2 inst_3945 ( .A(net_3736), .Z(net_3737) );
INV_X4 inst_1201 ( .ZN(net_630), .A(net_621) );
INV_X2 inst_1473 ( .A(net_1778), .ZN(net_361) );
DFF_X2 inst_1788 ( .QN(net_2443), .D(net_547), .CK(net_3586) );
INV_X4 inst_1272 ( .A(net_2346), .ZN(net_414) );
CLKBUF_X2 inst_4182 ( .A(net_3973), .Z(net_3974) );
NAND4_X2 inst_636 ( .A2(net_2050), .ZN(net_1911), .A3(net_1909), .A1(net_522), .A4(net_363) );
NAND4_X2 inst_632 ( .ZN(net_459), .A1(net_391), .A2(net_390), .A3(net_389), .A4(net_388) );
XOR2_X2 inst_0 ( .A(net_2084), .Z(net_1253), .B(net_309) );
CLKBUF_X2 inst_2852 ( .A(net_2569), .Z(net_2644) );
DFF_X1 inst_1927 ( .D(net_1130), .QN(net_58), .CK(net_3267) );
OAI22_X2 inst_184 ( .B1(net_1428), .A1(net_529), .B2(net_217), .A2(net_90), .ZN(x1628) );
DFF_X1 inst_1847 ( .QN(net_2371), .D(net_1455), .CK(net_3410) );
CLKBUF_X2 inst_3973 ( .A(net_3764), .Z(net_3765) );
DFF_X1 inst_1907 ( .D(net_1306), .Q(net_143), .CK(net_3045) );
OAI21_X2 inst_433 ( .ZN(net_1893), .A(net_520), .B1(net_519), .B2(net_466) );
DFF_X1 inst_1983 ( .D(net_1051), .QN(net_44), .CK(net_3185) );
CLKBUF_X2 inst_3836 ( .A(net_3298), .Z(net_3628) );
DFF_X1 inst_1948 ( .Q(net_2114), .D(net_1099), .CK(net_3403) );
DFFR_X1 inst_2114 ( .QN(net_2305), .RN(net_1347), .D(net_944), .CK(net_2481) );
CLKBUF_X2 inst_2784 ( .A(net_2575), .Z(net_2576) );
CLKBUF_X2 inst_4216 ( .A(net_4007), .Z(net_4008) );
SDFF_X2 inst_106 ( .SE(net_487), .Q(net_156), .D(net_156), .CK(net_2766), .SI(x4790) );
OAI21_X2 inst_422 ( .B2(net_1904), .B1(net_1872), .ZN(net_478), .A(net_477) );
AND2_X4 inst_2583 ( .A1(net_2420), .A2(net_2419), .ZN(net_351) );
AOI22_X2 inst_2243 ( .B2(net_2163), .A1(net_1967), .B1(net_1915), .ZN(net_1387), .A2(net_322) );
INV_X2 inst_1475 ( .A(net_1514), .ZN(net_936) );
INV_X2 inst_1426 ( .ZN(net_1594), .A(net_444) );
CLKBUF_X2 inst_3090 ( .A(net_2881), .Z(net_2882) );
INV_X2 inst_1637 ( .ZN(net_391), .A(x3976) );
CLKBUF_X2 inst_3997 ( .A(net_3788), .Z(net_3789) );
INV_X4 inst_1352 ( .A(net_2198), .ZN(net_2197) );
AOI22_X2 inst_2261 ( .A2(net_2031), .ZN(net_1169), .A1(net_1168), .B1(net_1154), .B2(net_354) );
CLKBUF_X2 inst_4142 ( .A(net_3373), .Z(net_3934) );
CLKBUF_X2 inst_3390 ( .A(net_3181), .Z(net_3182) );
CLKBUF_X2 inst_2930 ( .A(net_2663), .Z(net_2722) );
INV_X2 inst_1410 ( .A(net_566), .ZN(x1155) );
CLKBUF_X2 inst_2859 ( .A(net_2650), .Z(net_2651) );
OAI21_X2 inst_397 ( .B1(net_1829), .ZN(net_1110), .B2(net_941), .A(net_927) );
CLKBUF_X2 inst_3756 ( .A(net_3507), .Z(net_3548) );
NOR2_X4 inst_504 ( .A2(net_1747), .A1(net_1730), .ZN(net_1246) );
CLKBUF_X2 inst_3192 ( .A(net_2787), .Z(net_2984) );
DFF_X2 inst_1733 ( .QN(net_2321), .D(net_1494), .CK(net_3127) );
INV_X4 inst_1297 ( .A(net_2341), .ZN(net_309) );
CLKBUF_X2 inst_3900 ( .A(net_3691), .Z(net_3692) );
CLKBUF_X2 inst_3194 ( .A(net_2985), .Z(net_2986) );
NAND2_X2 inst_918 ( .A1(net_1168), .ZN(net_1107), .A2(net_531) );
CLKBUF_X2 inst_3884 ( .A(net_3675), .Z(net_3676) );
INV_X8 inst_1173 ( .ZN(net_2016), .A(net_2012) );
CLKBUF_X2 inst_3904 ( .A(net_3457), .Z(net_3696) );
CLKBUF_X2 inst_2908 ( .A(net_2592), .Z(net_2700) );
INV_X2 inst_1393 ( .A(net_582), .ZN(x989) );
DFFR_X2 inst_2074 ( .QN(net_2417), .RN(net_1347), .D(net_1251), .CK(net_3985) );
CLKBUF_X2 inst_4035 ( .A(net_3239), .Z(net_3827) );
DFF_X1 inst_1862 ( .D(net_1355), .QN(net_111), .CK(net_3880) );
CLKBUF_X2 inst_3519 ( .A(net_3310), .Z(net_3311) );
INV_X4 inst_1236 ( .ZN(net_411), .A(net_396) );
OAI22_X2 inst_221 ( .B2(net_2290), .B1(net_1865), .A1(net_1597), .ZN(net_957), .A2(net_747) );
CLKBUF_X2 inst_4075 ( .A(net_3430), .Z(net_3867) );
CLKBUF_X2 inst_3313 ( .A(net_3104), .Z(net_3105) );
CLKBUF_X2 inst_3562 ( .A(net_2903), .Z(net_3354) );
AOI22_X2 inst_2334 ( .B2(net_2160), .A1(net_2038), .A2(net_1546), .B1(net_979), .ZN(net_830) );
AOI22_X2 inst_2429 ( .B2(net_2144), .B1(net_1974), .ZN(net_1803), .A1(net_1791), .A2(net_306) );
AOI22_X2 inst_2210 ( .A2(net_2395), .B2(net_2113), .A1(net_1960), .ZN(net_1470), .B1(net_1450) );
NAND2_X4 inst_754 ( .ZN(net_2010), .A1(net_2008), .A2(net_1783) );
CLKBUF_X2 inst_2937 ( .A(net_2543), .Z(net_2729) );
AND2_X4 inst_2590 ( .ZN(net_1954), .A1(net_1953), .A2(net_1719) );
CLKBUF_X2 inst_2913 ( .A(net_2646), .Z(net_2705) );
NAND3_X2 inst_687 ( .A1(net_1935), .A2(net_1901), .ZN(net_1617), .A3(net_478) );
DFF_X2 inst_1774 ( .QN(net_2422), .D(net_881), .CK(net_3676) );
AOI22_X2 inst_2319 ( .A2(net_2154), .B1(net_2096), .A1(net_1769), .B2(net_1518), .ZN(net_890) );
CLKBUF_X2 inst_3295 ( .A(net_3086), .Z(net_3087) );
NAND2_X2 inst_985 ( .A2(net_1550), .A1(net_961), .ZN(net_854) );
AOI22_X2 inst_2225 ( .B2(net_2148), .A1(net_2040), .B1(net_1474), .ZN(net_1452), .A2(net_1276) );
AOI221_X2 inst_2513 ( .B2(net_2163), .ZN(net_1956), .A(net_1955), .B1(net_1929), .C1(net_1863), .C2(net_295) );
CLKBUF_X2 inst_4061 ( .A(net_3852), .Z(net_3853) );
AOI22_X2 inst_2254 ( .B2(net_2118), .A1(net_1967), .B1(net_1450), .ZN(net_1376), .A2(net_1203) );
CLKBUF_X2 inst_2923 ( .A(net_2714), .Z(net_2715) );
CLKBUF_X2 inst_2707 ( .A(net_2451), .Z(net_2499) );
NAND2_X2 inst_1117 ( .ZN(net_2075), .A2(net_2072), .A1(net_2000) );
CLKBUF_X2 inst_4015 ( .A(net_3806), .Z(net_3807) );
CLKBUF_X2 inst_3958 ( .A(net_3749), .Z(net_3750) );
DFF_X1 inst_2007 ( .QN(net_2226), .D(net_1080), .CK(net_3245) );
CLKBUF_X2 inst_2725 ( .A(net_2492), .Z(net_2517) );
CLKBUF_X2 inst_3644 ( .A(net_3435), .Z(net_3436) );
INV_X2 inst_1610 ( .ZN(net_660), .A(net_59) );
OAI21_X2 inst_334 ( .B2(net_2315), .B1(net_2041), .ZN(net_1496), .A(net_1463) );
NAND2_X2 inst_805 ( .A2(net_1671), .ZN(net_1308), .A1(net_1286) );
CLKBUF_X2 inst_3707 ( .A(net_3498), .Z(net_3499) );
OAI21_X2 inst_354 ( .B2(net_2375), .B1(net_1441), .ZN(net_1440), .A(net_1384) );
INV_X8 inst_1145 ( .A(net_1402), .ZN(net_529) );
NAND2_X2 inst_1042 ( .A1(net_1828), .ZN(net_1669), .A2(net_275) );
OAI21_X2 inst_373 ( .B1(net_1441), .ZN(net_1416), .A(net_1387), .B2(net_1152) );
CLKBUF_X2 inst_3056 ( .A(net_2847), .Z(net_2848) );
DFF_X1 inst_1868 ( .D(net_1348), .QN(net_117), .CK(net_3803) );
NOR2_X2 inst_595 ( .A2(net_2259), .ZN(net_1884), .A1(net_520) );
AND2_X2 inst_2609 ( .A1(net_609), .A2(x5143), .ZN(x925) );
XNOR2_X2 inst_22 ( .B(net_1190), .ZN(net_1167), .A(net_1153) );
DFF_X2 inst_1717 ( .QN(net_2333), .D(net_2021), .CK(net_3178) );
AOI21_X2 inst_2556 ( .B2(net_2113), .ZN(net_1975), .B1(net_1974), .A(net_1972) );
CLKBUF_X2 inst_3099 ( .A(net_2890), .Z(net_2891) );
INV_X1 inst_1704 ( .ZN(net_483), .A(net_482) );
CLKBUF_X2 inst_2901 ( .A(net_2658), .Z(net_2693) );
NAND2_X4 inst_767 ( .ZN(net_2101), .A1(net_614), .A2(net_522) );
OAI22_X2 inst_161 ( .B1(net_1614), .A1(net_1408), .B2(net_264), .A2(net_135), .ZN(x255) );
CLKBUF_X2 inst_3356 ( .A(net_3147), .Z(net_3148) );
CLKBUF_X2 inst_3849 ( .A(net_3640), .Z(net_3641) );
NAND2_X4 inst_718 ( .A1(net_1984), .ZN(net_520), .A2(net_507) );
NAND2_X2 inst_1029 ( .A2(net_2381), .ZN(net_510), .A1(net_446) );
CLKBUF_X2 inst_4024 ( .A(net_3815), .Z(net_3816) );
AOI22_X2 inst_2408 ( .B1(net_2197), .ZN(net_1636), .A1(net_1621), .B2(net_1518), .A2(net_1291) );
INV_X4 inst_1324 ( .ZN(net_1933), .A(net_1932) );
OAI21_X2 inst_342 ( .B2(net_2328), .B1(net_2041), .ZN(net_1488), .A(net_1479) );
NOR2_X4 inst_526 ( .ZN(net_1772), .A1(net_1578), .A2(net_191) );
DFFR_X1 inst_2147 ( .QN(net_2253), .RN(net_1347), .D(net_702), .CK(net_3339) );
INV_X8 inst_1178 ( .ZN(net_2195), .A(net_2194) );
OAI211_X2 inst_463 ( .C2(net_2333), .A(net_1921), .C1(net_1052), .ZN(net_1051), .B(net_865) );
DFFR_X2 inst_2091 ( .QN(net_1583), .RN(net_1347), .D(net_995), .CK(net_3725) );
INV_X2 inst_1534 ( .ZN(net_260), .A(x6298) );
CLKBUF_X2 inst_3104 ( .A(net_2895), .Z(net_2896) );
CLKBUF_X2 inst_3820 ( .A(net_3611), .Z(net_3612) );
OAI21_X2 inst_319 ( .B1(net_2041), .ZN(net_1511), .A(net_1476), .B2(net_400) );
INV_X2 inst_1450 ( .A(net_1523), .ZN(net_711) );
AOI22_X2 inst_2422 ( .B2(net_2108), .B1(net_1974), .ZN(net_1796), .A1(net_1791), .A2(net_311) );
CLKBUF_X2 inst_3123 ( .A(net_2634), .Z(net_2915) );
NAND3_X2 inst_649 ( .ZN(net_1453), .A1(net_1399), .A3(net_1363), .A2(net_1195) );
CLKBUF_X2 inst_3725 ( .A(net_3516), .Z(net_3517) );
HA_X1 inst_1711 ( .B(net_1201), .CO(net_618), .S(net_551), .A(net_503) );
AND2_X4 inst_2597 ( .ZN(net_2171), .A2(net_2105), .A1(net_1649) );
CLKBUF_X2 inst_3426 ( .A(net_3217), .Z(net_3218) );
NOR3_X2 inst_500 ( .ZN(net_2063), .A3(net_2062), .A2(net_1926), .A1(net_1724) );
INV_X2 inst_1592 ( .ZN(net_217), .A(x4197) );
DFF_X2 inst_1770 ( .QN(net_2429), .D(net_991), .CK(net_3623) );
INV_X2 inst_1575 ( .A(net_2272), .ZN(net_293) );
NAND2_X2 inst_995 ( .A1(net_1797), .ZN(net_836), .A2(net_676) );
NOR2_X2 inst_550 ( .A1(net_2194), .ZN(net_606), .A2(net_412) );
DFF_X1 inst_2052 ( .Q(net_2392), .D(net_2184), .CK(net_3146) );
CLKBUF_X2 inst_3413 ( .A(net_2573), .Z(net_3205) );
AOI222_X2 inst_2470 ( .C1(net_2014), .A2(net_1553), .A1(net_590), .B1(net_589), .ZN(net_566), .B2(net_155), .C2(x5712) );
INV_X4 inst_1258 ( .ZN(net_448), .A(net_354) );
CLKBUF_X2 inst_3141 ( .A(net_2932), .Z(net_2933) );
CLKBUF_X2 inst_3921 ( .A(net_3402), .Z(net_3713) );
DFF_X1 inst_1957 ( .Q(net_2123), .D(net_1095), .CK(net_3534) );
CLKBUF_X2 inst_3857 ( .A(net_2589), .Z(net_3649) );
NAND2_X2 inst_1060 ( .A2(net_2431), .ZN(net_1716), .A1(net_222) );
INV_X2 inst_1419 ( .ZN(net_623), .A(net_615) );
NAND2_X2 inst_900 ( .A2(net_1699), .A1(net_1698), .ZN(net_1119) );
CLKBUF_X2 inst_2661 ( .A(net_2452), .Z(net_2453) );
AOI221_X2 inst_2501 ( .B2(net_2129), .B1(net_1929), .A(net_1876), .C1(net_1863), .ZN(net_970), .C2(net_276) );
CLKBUF_X2 inst_3548 ( .A(net_3084), .Z(net_3340) );
CLKBUF_X2 inst_2807 ( .A(net_2598), .Z(net_2599) );
NOR2_X2 inst_594 ( .A2(net_2275), .ZN(net_1883), .A1(net_520) );
CLKBUF_X2 inst_2983 ( .A(net_2774), .Z(net_2775) );
INV_X2 inst_1632 ( .ZN(net_190), .A(x4175) );
NAND2_X2 inst_925 ( .A2(net_1630), .ZN(net_1089), .A1(net_688) );
AOI22_X2 inst_2378 ( .A1(net_1718), .B1(net_1450), .B2(net_815), .ZN(net_648), .A2(net_318) );
NAND2_X2 inst_1120 ( .ZN(net_2099), .A1(net_2098), .A2(net_1862) );
INV_X2 inst_1536 ( .ZN(net_258), .A(x6530) );
NAND2_X2 inst_881 ( .A2(net_1196), .ZN(net_1188), .A1(net_1172) );
CLKBUF_X2 inst_3876 ( .A(net_2705), .Z(net_3668) );
CLKBUF_X2 inst_3184 ( .A(net_2975), .Z(net_2976) );
CLKBUF_X2 inst_3848 ( .A(net_3453), .Z(net_3640) );
INV_X4 inst_1225 ( .ZN(net_1687), .A(net_431) );
NAND2_X2 inst_947 ( .A2(net_1532), .ZN(net_994), .A1(net_992) );
NAND2_X4 inst_731 ( .A1(net_2006), .ZN(net_1836), .A2(net_1835) );
CLKBUF_X2 inst_3706 ( .A(net_3497), .Z(net_3498) );
AOI222_X2 inst_2459 ( .C1(net_2016), .A2(net_1564), .A1(net_590), .B1(net_589), .ZN(net_577), .B2(net_166), .C2(x5448) );
OAI22_X2 inst_301 ( .A2(net_2239), .A1(net_2013), .B1(net_1895), .B2(net_229), .ZN(x1811) );
OAI21_X2 inst_363 ( .B1(net_1443), .ZN(net_1431), .A(net_1385), .B2(net_1167) );
DFFR_X1 inst_2141 ( .QN(net_2274), .RN(net_1347), .D(net_717), .CK(net_2469) );
OAI22_X2 inst_247 ( .B2(net_2268), .ZN(net_729), .A2(net_728), .A1(net_714), .B1(net_534) );
OAI21_X2 inst_403 ( .B2(net_2378), .ZN(net_883), .B1(net_635), .A(net_625) );
CLKBUF_X2 inst_3446 ( .A(net_3237), .Z(net_3238) );
CLKBUF_X2 inst_2728 ( .A(net_2498), .Z(net_2520) );
INV_X2 inst_1588 ( .ZN(net_786), .A(net_67) );
CLKBUF_X2 inst_3801 ( .A(net_3592), .Z(net_3593) );
CLKBUF_X2 inst_4177 ( .A(net_3968), .Z(net_3969) );
CLKBUF_X2 inst_2956 ( .A(net_2621), .Z(net_2748) );
CLKBUF_X2 inst_3729 ( .A(net_3520), .Z(net_3521) );
OAI21_X2 inst_412 ( .B1(net_768), .ZN(net_757), .A(net_647), .B2(net_495) );
AOI21_X4 inst_2516 ( .A(net_1935), .ZN(net_1758), .B1(net_1684), .B2(net_82) );
AND2_X2 inst_2650 ( .A2(net_2122), .ZN(net_2062), .A1(net_1928) );
DFFR_X1 inst_2155 ( .QN(net_2249), .RN(net_1347), .D(net_731), .CK(net_2504) );
INV_X2 inst_1506 ( .A(net_2314), .ZN(net_286) );
OAI211_X2 inst_464 ( .C2(net_2335), .C1(net_1052), .ZN(net_1050), .A(net_900), .B(net_864) );
OAI21_X2 inst_341 ( .B2(net_2332), .B1(net_2041), .ZN(net_1489), .A(net_1478) );
CLKBUF_X2 inst_3785 ( .A(net_3576), .Z(net_3577) );
CLKBUF_X2 inst_3189 ( .A(net_2980), .Z(net_2981) );
CLKBUF_X2 inst_3163 ( .A(net_2954), .Z(net_2955) );
AOI221_X2 inst_2504 ( .B2(net_2117), .C2(net_2093), .B1(net_1929), .A(net_1881), .C1(net_1863), .ZN(net_965) );
AOI22_X2 inst_2359 ( .A1(net_783), .B1(net_775), .ZN(net_771), .A2(net_377), .B2(x3618) );
CLKBUF_X2 inst_3702 ( .A(net_3493), .Z(net_3494) );
NAND3_X2 inst_684 ( .A1(net_2439), .ZN(net_455), .A3(x5995), .A2(x5957) );
CLKBUF_X2 inst_3374 ( .A(net_3165), .Z(net_3166) );
CLKBUF_X2 inst_3177 ( .A(net_2675), .Z(net_2969) );
CLKBUF_X2 inst_3438 ( .A(net_3229), .Z(net_3230) );
INV_X2 inst_1361 ( .ZN(net_1144), .A(net_1138) );
CLKBUF_X2 inst_3401 ( .A(net_3169), .Z(net_3193) );
CLKBUF_X2 inst_3811 ( .A(net_3602), .Z(net_3603) );
CLKBUF_X2 inst_3653 ( .A(net_3444), .Z(net_3445) );
AOI22_X2 inst_2208 ( .A2(net_2343), .B2(net_2139), .A1(net_1960), .ZN(net_1472), .B1(net_1450) );
INV_X8 inst_1138 ( .ZN(net_745), .A(net_534) );
CLKBUF_X2 inst_4162 ( .A(net_3953), .Z(net_3954) );
INV_X4 inst_1241 ( .A(net_2315), .ZN(net_1260) );
NAND2_X2 inst_1038 ( .A2(net_2382), .A1(net_2381), .ZN(net_348) );
NAND2_X2 inst_940 ( .A1(net_1860), .ZN(net_1060), .A2(net_918) );
NAND2_X2 inst_1004 ( .A2(net_2136), .A1(net_979), .ZN(net_668) );
CLKBUF_X2 inst_3201 ( .A(net_2992), .Z(net_2993) );
CLKBUF_X2 inst_3595 ( .A(net_3386), .Z(net_3387) );
OAI22_X2 inst_189 ( .B1(net_1428), .A1(net_529), .B2(net_180), .A2(net_85), .ZN(x1701) );
XNOR2_X2 inst_14 ( .B(net_2335), .ZN(net_1346), .A(net_1234) );
AOI222_X2 inst_2450 ( .C1(net_2016), .A2(net_1573), .A1(net_590), .B1(net_589), .ZN(net_586), .B2(net_175), .C2(x5247) );
SDFF_X2 inst_62 ( .Q(net_1546), .D(net_1546), .SE(net_498), .CK(net_2692), .SI(x7466) );
AOI22_X2 inst_2325 ( .A2(net_2109), .B1(net_2096), .A1(net_1769), .B2(net_1517), .ZN(net_884) );
CLKBUF_X2 inst_3743 ( .A(net_3102), .Z(net_3535) );
OAI22_X2 inst_251 ( .B2(net_2272), .A1(net_745), .ZN(net_721), .A2(net_720), .B1(net_534) );
CLKBUF_X2 inst_2860 ( .A(net_2517), .Z(net_2652) );
NAND2_X2 inst_1074 ( .A1(net_2104), .ZN(net_1815), .A2(net_1259) );
NAND2_X2 inst_879 ( .A1(net_2003), .A2(net_1668), .ZN(net_1181) );
CLKBUF_X2 inst_4007 ( .A(net_3798), .Z(net_3799) );
INV_X2 inst_1552 ( .ZN(net_248), .A(x4051) );
INV_X2 inst_1524 ( .A(net_2289), .ZN(net_297) );
INV_X2 inst_1602 ( .A(net_2309), .ZN(net_296) );
NAND2_X2 inst_969 ( .A2(net_1561), .A1(net_961), .ZN(net_870) );
NAND4_X4 inst_629 ( .A4(net_2176), .ZN(net_2090), .A3(net_2089), .A2(net_2088), .A1(net_2087) );
NAND2_X2 inst_1100 ( .ZN(net_1949), .A2(net_1948), .A1(net_1181) );
AOI21_X2 inst_2528 ( .A(net_1785), .B1(net_910), .ZN(net_805), .B2(net_75) );
NAND2_X2 inst_791 ( .A1(net_1815), .ZN(net_1322), .A2(net_1204) );
DFF_X1 inst_2021 ( .QN(net_2211), .D(net_1900), .CK(net_3243) );
NAND2_X2 inst_898 ( .A2(net_1711), .A1(net_1710), .ZN(net_1122) );
CLKBUF_X2 inst_3383 ( .A(net_3174), .Z(net_3175) );
DFF_X1 inst_1977 ( .Q(net_2142), .D(net_1037), .CK(net_3041) );
DFF_X2 inst_1793 ( .QN(net_2245), .D(net_463), .CK(net_3807) );
INV_X4 inst_1191 ( .A(net_1829), .ZN(net_992) );
CLKBUF_X2 inst_4227 ( .A(net_4018), .Z(net_4019) );
NOR2_X4 inst_533 ( .ZN(net_2073), .A1(net_2072), .A2(net_1923) );
AOI222_X2 inst_2478 ( .B2(net_2202), .B1(net_1948), .ZN(net_532), .A1(net_531), .A2(net_500), .C2(net_396), .C1(net_358) );
CLKBUF_X2 inst_2751 ( .A(net_2502), .Z(net_2543) );
DFF_X1 inst_1874 ( .D(net_1330), .QN(net_101), .CK(net_3612) );
DFF_X2 inst_1760 ( .D(net_1682), .QN(net_1589), .CK(net_3903) );
AOI22_X2 inst_2291 ( .A1(net_1996), .B1(net_1749), .A2(net_1553), .ZN(net_968), .B2(net_155) );
AOI22_X2 inst_2343 ( .B1(net_2197), .A1(net_2038), .A2(net_1573), .B2(net_1520), .ZN(net_821) );
AOI21_X2 inst_2538 ( .A(net_1785), .B1(net_910), .ZN(net_791), .B2(net_790) );
DFF_X1 inst_2022 ( .QN(net_2410), .D(net_924), .CK(net_3679) );
CLKBUF_X2 inst_2821 ( .A(net_2612), .Z(net_2613) );
CLKBUF_X2 inst_3132 ( .A(net_2923), .Z(net_2924) );
CLKBUF_X2 inst_3960 ( .A(net_3751), .Z(net_3752) );
NAND2_X2 inst_1095 ( .A1(net_1965), .ZN(net_1917), .A2(net_1716) );
OAI22_X2 inst_176 ( .B1(net_1402), .A1(net_529), .B2(net_238), .A2(net_100), .ZN(x1492) );
AOI22_X2 inst_2439 ( .B2(net_2394), .B1(net_1916), .A1(net_1915), .ZN(net_1857), .A2(net_1855) );
CLKBUF_X2 inst_2826 ( .A(net_2617), .Z(net_2618) );
CLKBUF_X2 inst_3910 ( .A(net_3701), .Z(net_3702) );
INV_X4 inst_1336 ( .ZN(net_2022), .A(net_1834) );
INV_X4 inst_1332 ( .ZN(net_2000), .A(net_1923) );
DFF_X1 inst_1841 ( .QN(net_2327), .D(net_1512), .CK(net_3308) );
INV_X2 inst_1665 ( .A(net_1757), .ZN(net_1756) );
CLKBUF_X2 inst_3345 ( .A(net_3136), .Z(net_3137) );
CLKBUF_X2 inst_3264 ( .A(net_2790), .Z(net_3056) );
NAND2_X2 inst_780 ( .ZN(net_1345), .A2(net_1255), .A1(net_1178) );
AOI22_X2 inst_2332 ( .B2(net_2125), .A1(net_2038), .A2(net_1555), .B1(net_979), .ZN(net_832) );
CLKBUF_X2 inst_3967 ( .A(net_3431), .Z(net_3759) );
AOI22_X2 inst_2310 ( .A2(net_2112), .B1(net_2096), .A1(net_1769), .B2(net_1534), .ZN(net_899) );
NAND2_X2 inst_1089 ( .A1(net_2435), .ZN(net_1866), .A2(net_291) );
CLKBUF_X2 inst_4018 ( .A(net_3809), .Z(net_3810) );
DFF_X2 inst_1767 ( .QN(net_2384), .D(net_997), .CK(net_3871) );
CLKBUF_X2 inst_3669 ( .A(net_3460), .Z(net_3461) );
AOI22_X2 inst_2219 ( .A2(net_2389), .B2(net_2157), .A1(net_1960), .ZN(net_1461), .B1(net_1450) );
INV_X4 inst_1284 ( .A(net_1592), .ZN(net_271) );
NOR2_X2 inst_546 ( .A2(net_1718), .ZN(net_880), .A1(net_605) );
AOI222_X2 inst_2465 ( .C1(net_2015), .A2(net_1565), .A1(net_590), .B1(net_589), .ZN(net_571), .B2(net_167), .C2(x5429) );
AOI22_X2 inst_2361 ( .B1(net_1915), .B2(net_811), .ZN(net_751), .A1(net_640), .A2(net_379) );
INV_X4 inst_1290 ( .A(net_2372), .ZN(net_537) );
NAND3_X2 inst_704 ( .ZN(net_2059), .A1(net_1800), .A3(net_801), .A2(net_656) );
AOI22_X2 inst_2226 ( .B2(net_2110), .A1(net_2040), .A2(net_1812), .ZN(net_1451), .B1(net_1450) );
NAND3_X2 inst_694 ( .A2(net_2203), .ZN(net_1874), .A1(net_444), .A3(net_442) );
DFF_X1 inst_2046 ( .Q(net_2393), .D(net_1651), .CK(net_3084) );
AOI222_X1 inst_2498 ( .B1(net_1995), .A1(net_1751), .B2(net_1572), .C1(net_1020), .ZN(net_989), .A2(net_174), .C2(x3261) );
CLKBUF_X2 inst_4129 ( .A(net_3920), .Z(net_3921) );
CLKBUF_X2 inst_3154 ( .A(net_2945), .Z(net_2946) );
CLKBUF_X2 inst_3861 ( .A(net_3652), .Z(net_3653) );
INV_X4 inst_1342 ( .ZN(net_2071), .A(net_2070) );
CLKBUF_X2 inst_2971 ( .A(net_2762), .Z(net_2763) );
CLKBUF_X2 inst_4196 ( .A(net_3987), .Z(net_3988) );
CLKBUF_X2 inst_3524 ( .A(net_3315), .Z(net_3316) );
NAND2_X2 inst_1014 ( .A1(net_2195), .ZN(net_620), .A2(net_510) );
NAND2_X2 inst_787 ( .A1(net_1820), .ZN(net_1326), .A2(net_1210) );
AOI21_X2 inst_2531 ( .A(net_1785), .B1(net_910), .ZN(net_802), .B2(net_78) );
CLKBUF_X2 inst_3933 ( .A(net_3724), .Z(net_3725) );
INV_X4 inst_1347 ( .ZN(net_2089), .A(net_1773) );
NAND2_X2 inst_825 ( .A1(net_1840), .ZN(net_1333), .A2(net_309) );
INV_X2 inst_1656 ( .ZN(net_178), .A(x4251) );
NOR2_X4 inst_509 ( .ZN(net_555), .A1(net_542), .A2(net_533) );
AND2_X4 inst_2586 ( .A2(net_2424), .A1(net_2422), .ZN(net_269) );
CLKBUF_X2 inst_2687 ( .A(net_2478), .Z(net_2479) );
INV_X2 inst_1680 ( .ZN(net_2025), .A(net_2022) );
DFF_X1 inst_1881 ( .D(net_1327), .QN(net_95), .CK(net_3717) );
INV_X2 inst_1626 ( .ZN(net_195), .A(x4080) );
AND2_X2 inst_2622 ( .A1(net_594), .A2(x7329), .ZN(x817) );
OAI22_X2 inst_153 ( .B1(net_1427), .A1(net_1426), .B2(net_388), .A2(net_114), .ZN(x1337) );
DFF_X1 inst_1892 ( .D(net_1340), .QN(net_134), .CK(net_3448) );
CLKBUF_X2 inst_3034 ( .A(net_2825), .Z(net_2826) );
INV_X2 inst_1459 ( .A(net_2361), .ZN(net_932) );
NAND2_X4 inst_726 ( .A1(net_1746), .A2(net_1730), .ZN(net_1713) );
OAI22_X2 inst_295 ( .B2(net_2292), .A1(net_1973), .ZN(net_1849), .B1(net_1848), .A2(net_43) );
CLKBUF_X2 inst_4094 ( .A(net_3885), .Z(net_3886) );
OAI22_X2 inst_209 ( .A2(net_2218), .A1(net_2017), .B1(net_1406), .B2(net_206), .ZN(x2260) );
CLKBUF_X2 inst_3894 ( .A(net_2611), .Z(net_3686) );
NAND2_X2 inst_1087 ( .ZN(net_1848), .A1(net_1665), .A2(net_499) );
DFF_X2 inst_1781 ( .QN(net_2420), .D(net_753), .CK(net_3452) );
OAI21_X2 inst_320 ( .B2(net_2337), .B1(net_2041), .ZN(net_1510), .A(net_1475) );
NOR2_X2 inst_607 ( .A1(net_2202), .A2(net_2170), .ZN(net_1950) );
CLKBUF_X2 inst_2769 ( .A(net_2560), .Z(net_2561) );
AOI22_X2 inst_2432 ( .B2(net_2158), .B1(net_1974), .ZN(net_1806), .A1(net_1789), .A2(net_297) );
INV_X2 inst_1375 ( .A(net_1009), .ZN(x2690) );
XOR2_X2 inst_1 ( .A(net_2432), .B(net_2328), .Z(net_1150) );
DFF_X1 inst_1891 ( .D(net_1338), .QN(net_136), .CK(net_3653) );
CLKBUF_X2 inst_3982 ( .A(net_3585), .Z(net_3774) );
CLKBUF_X2 inst_3215 ( .A(net_3006), .Z(net_3007) );
OAI22_X2 inst_235 ( .B2(net_2288), .B1(net_1865), .A1(net_951), .ZN(net_935), .A2(net_848) );
CLKBUF_X2 inst_3063 ( .A(net_2526), .Z(net_2855) );
AOI211_X2 inst_2564 ( .C2(net_2114), .C1(net_1929), .A(net_1875), .B(net_1785), .ZN(net_674) );
DFF_X2 inst_1812 ( .Q(net_1523), .CK(net_2715), .D(x5294) );
NAND2_X2 inst_1082 ( .A1(net_2104), .ZN(net_1823), .A2(net_1264) );
CLKBUF_X2 inst_4167 ( .A(net_3958), .Z(net_3959) );
CLKBUF_X2 inst_2677 ( .A(net_2468), .Z(net_2469) );
DFF_X1 inst_1995 ( .Q(net_2159), .D(net_1032), .CK(net_3153) );
SDFF_X2 inst_105 ( .SE(net_487), .Q(net_149), .D(net_149), .CK(net_2811), .SI(x4974) );
CLKBUF_X2 inst_3518 ( .A(net_3309), .Z(net_3310) );
NOR2_X1 inst_625 ( .ZN(net_270), .A2(net_55), .A1(net_52) );
CLKBUF_X2 inst_3367 ( .A(net_3158), .Z(net_3159) );
CLKBUF_X2 inst_2835 ( .A(net_2626), .Z(net_2627) );
NOR2_X2 inst_568 ( .ZN(net_353), .A2(net_249), .A1(x3098) );
INV_X2 inst_1483 ( .A(net_2350), .ZN(net_1201) );
NOR2_X4 inst_523 ( .ZN(net_1649), .A1(net_433), .A2(net_294) );
CLKBUF_X2 inst_2731 ( .A(net_2522), .Z(net_2523) );
AOI22_X2 inst_2207 ( .A2(net_2397), .B2(net_2142), .A1(net_1960), .B1(net_1474), .ZN(net_1473) );
INV_X2 inst_1492 ( .A(net_1197), .ZN(net_336) );
OAI22_X2 inst_181 ( .B1(net_1428), .A1(net_529), .B2(net_233), .A2(net_94), .ZN(x1578) );
CLKBUF_X2 inst_4234 ( .A(net_3847), .Z(net_4026) );
CLKBUF_X2 inst_3892 ( .A(net_2640), .Z(net_3684) );
NAND2_X4 inst_713 ( .A1(net_2195), .ZN(net_650), .A2(net_550) );
CLKBUF_X2 inst_3930 ( .A(net_3721), .Z(net_3722) );
CLKBUF_X2 inst_2867 ( .A(net_2462), .Z(net_2659) );
CLKBUF_X2 inst_2898 ( .A(net_2689), .Z(net_2690) );
OAI211_X2 inst_477 ( .C1(net_1054), .ZN(net_1032), .C2(net_1031), .A(net_887), .B(net_853) );
CLKBUF_X2 inst_3398 ( .A(net_3189), .Z(net_3190) );
INV_X2 inst_1368 ( .A(net_1016), .ZN(x2592) );
CLKBUF_X2 inst_3576 ( .A(net_3367), .Z(net_3368) );
OAI21_X2 inst_423 ( .B2(net_2422), .B1(net_2421), .ZN(net_476), .A(net_475) );
NAND2_X2 inst_835 ( .A1(net_1840), .ZN(net_1279), .A2(net_1264) );
DFFR_X2 inst_2088 ( .RN(net_1347), .D(net_1111), .QN(net_54), .CK(net_2745) );
CLKBUF_X2 inst_3305 ( .A(net_2647), .Z(net_3097) );
CLKBUF_X2 inst_3082 ( .A(net_2873), .Z(net_2874) );
CLKBUF_X2 inst_3208 ( .A(net_2999), .Z(net_3000) );
CLKBUF_X2 inst_4137 ( .A(net_2850), .Z(net_3929) );
NAND2_X2 inst_1112 ( .ZN(net_2046), .A1(net_2045), .A2(net_47) );
CLKBUF_X2 inst_4134 ( .A(net_3925), .Z(net_3926) );
CLKBUF_X2 inst_3507 ( .A(net_3298), .Z(net_3299) );
NAND2_X4 inst_710 ( .ZN(net_1182), .A1(net_1175), .A2(net_330) );
CLKBUF_X2 inst_4081 ( .A(net_2742), .Z(net_3873) );
INV_X2 inst_1379 ( .A(net_1005), .ZN(x2752) );
NAND2_X2 inst_941 ( .ZN(net_1059), .A1(net_967), .A2(net_891) );
OAI22_X2 inst_271 ( .B2(net_2294), .B1(net_1865), .ZN(net_1602), .A1(net_1597), .A2(net_737) );
CLKBUF_X2 inst_3350 ( .A(net_2571), .Z(net_3142) );
DFF_X2 inst_1817 ( .Q(net_1515), .CK(net_2597), .D(x5779) );
SDFF_X2 inst_56 ( .SE(net_1998), .D(net_1537), .SI(net_362), .Q(net_70), .CK(net_3276) );
OAI22_X2 inst_308 ( .B1(net_1895), .A1(net_1408), .B2(net_188), .A2(net_130), .ZN(x361) );
INV_X2 inst_1546 ( .A(net_2249), .ZN(net_305) );
INV_X4 inst_1230 ( .A(net_2076), .ZN(net_406) );
OAI211_X2 inst_455 ( .C1(net_1639), .ZN(net_1099), .C2(net_1098), .A(net_821), .B(net_667) );
CLKBUF_X2 inst_3535 ( .A(net_3326), .Z(net_3327) );
INV_X16 inst_1694 ( .ZN(net_1841), .A(net_1840) );
CLKBUF_X2 inst_2871 ( .A(net_2662), .Z(net_2663) );
AOI21_X2 inst_2540 ( .A(net_1785), .B1(net_910), .ZN(net_787), .B2(net_786) );
CLKBUF_X2 inst_3497 ( .A(net_3288), .Z(net_3289) );
NAND2_X2 inst_1064 ( .A1(net_2002), .A2(net_1732), .ZN(net_1726) );
CLKBUF_X2 inst_3629 ( .A(net_3420), .Z(net_3421) );
CLKBUF_X2 inst_3599 ( .A(net_3390), .Z(net_3391) );
CLKBUF_X2 inst_3024 ( .A(net_2673), .Z(net_2816) );
NOR2_X2 inst_583 ( .ZN(net_1859), .A1(net_1851), .A2(net_1576) );
DFF_X1 inst_1904 ( .D(net_1304), .QN(net_118), .CK(net_3799) );
CLKBUF_X2 inst_3581 ( .A(net_3372), .Z(net_3373) );
DFF_X1 inst_2065 ( .Q(net_1586), .D(net_353), .CK(net_3917) );
AOI22_X2 inst_2251 ( .B2(net_2136), .A1(net_1967), .A2(net_1735), .B1(net_1450), .ZN(net_1379) );
CLKBUF_X2 inst_3085 ( .A(net_2444), .Z(net_2877) );
CLKBUF_X2 inst_3987 ( .A(net_3778), .Z(net_3779) );
CLKBUF_X2 inst_3951 ( .A(net_3742), .Z(net_3743) );
DFF_X1 inst_1899 ( .D(net_1300), .QN(net_122), .CK(net_3580) );
CLKBUF_X2 inst_2943 ( .A(net_2495), .Z(net_2735) );
INV_X2 inst_1593 ( .ZN(net_389), .A(x3954) );
AND4_X4 inst_2569 ( .A3(net_2418), .A4(net_2415), .A1(net_1754), .A2(net_1592), .ZN(net_384) );
NAND2_X4 inst_724 ( .A1(net_1655), .ZN(net_1643), .A2(net_327) );
CLKBUF_X2 inst_2716 ( .A(net_2507), .Z(net_2508) );
AOI222_X2 inst_2449 ( .C1(net_2017), .A2(net_1574), .A1(net_590), .B1(net_589), .ZN(net_587), .B2(net_176), .C2(x5224) );
CLKBUF_X2 inst_3228 ( .A(net_2611), .Z(net_3020) );
NAND2_X2 inst_975 ( .A2(net_1568), .A1(net_961), .ZN(net_864) );
DFFR_X1 inst_2124 ( .QN(net_2283), .D(net_1598), .RN(net_1347), .CK(net_2844) );
CLKBUF_X2 inst_2789 ( .A(net_2580), .Z(net_2581) );
CLKBUF_X2 inst_3191 ( .A(net_2982), .Z(net_2983) );
AOI22_X2 inst_2289 ( .A1(net_1996), .B1(net_1749), .A2(net_1544), .ZN(net_973), .B2(net_146) );
INV_X2 inst_1435 ( .A(net_1186), .ZN(net_1045) );
INV_X2 inst_1431 ( .A(net_2331), .ZN(net_401) );
CLKBUF_X2 inst_3760 ( .A(net_3551), .Z(net_3552) );
INV_X2 inst_1398 ( .A(net_577), .ZN(x1036) );
CLKBUF_X2 inst_3746 ( .A(net_3537), .Z(net_3538) );
DFF_X2 inst_1804 ( .Q(net_1541), .CK(net_2817), .D(x5686) );
CLKBUF_X2 inst_2750 ( .A(net_2541), .Z(net_2542) );
CLKBUF_X2 inst_2849 ( .A(net_2640), .Z(net_2641) );
AOI22_X2 inst_2440 ( .ZN(net_1858), .A1(net_1852), .B1(net_1789), .A2(net_472), .B2(net_332) );
CLKBUF_X2 inst_4121 ( .A(net_3912), .Z(net_3913) );
INV_X2 inst_1467 ( .ZN(net_362), .A(net_301) );
AND2_X2 inst_2640 ( .A1(net_775), .A2(x6773), .ZN(x596) );
CLKBUF_X2 inst_3327 ( .A(net_2618), .Z(net_3119) );
CLKBUF_X2 inst_2659 ( .A(net_2450), .Z(net_2451) );
DFFR_X1 inst_2134 ( .QN(net_2266), .RN(net_1347), .D(net_733), .CK(net_2797) );
DFF_X2 inst_1744 ( .QN(net_2362), .D(net_1431), .CK(net_3591) );
CLKBUF_X2 inst_2834 ( .A(net_2625), .Z(net_2626) );
INV_X2 inst_1513 ( .A(net_2422), .ZN(net_350) );
INV_X8 inst_1155 ( .A(net_1840), .ZN(net_1743) );
CLKBUF_X2 inst_4117 ( .A(net_3604), .Z(net_3909) );
OAI22_X2 inst_207 ( .A2(net_2223), .B1(net_1614), .A1(net_1405), .B2(net_261), .ZN(x2149) );
CLKBUF_X2 inst_3321 ( .A(net_3112), .Z(net_3113) );
CLKBUF_X2 inst_4080 ( .A(net_3322), .Z(net_3872) );
INV_X2 inst_1545 ( .ZN(net_253), .A(x4184) );
OAI21_X2 inst_333 ( .B2(net_2318), .B1(net_2041), .ZN(net_1497), .A(net_1461) );
CLKBUF_X2 inst_3338 ( .A(net_2600), .Z(net_3130) );
NAND2_X4 inst_712 ( .A2(net_2036), .A1(net_1963), .ZN(net_633) );
INV_X4 inst_1215 ( .A(net_1984), .ZN(net_516) );
OR2_X4 inst_131 ( .ZN(net_1834), .A2(net_1833), .A1(net_82) );
OAI21_X2 inst_406 ( .ZN(net_798), .B2(net_768), .A(net_643), .B1(net_595) );
OAI21_X2 inst_328 ( .B2(net_2313), .B1(net_1507), .ZN(net_1502), .A(net_1468) );
CLKBUF_X2 inst_3111 ( .A(net_2902), .Z(net_2903) );
DFF_X1 inst_2035 ( .QN(net_2241), .D(net_912), .CK(net_3210) );
SDFF_X2 inst_47 ( .SE(net_1768), .SI(net_1534), .Q(net_73), .D(net_73), .CK(net_3423) );
CLKBUF_X2 inst_4217 ( .A(net_4008), .Z(net_4009) );
CLKBUF_X2 inst_2764 ( .A(net_2555), .Z(net_2556) );
NAND2_X2 inst_818 ( .A1(net_1841), .ZN(net_1292), .A2(net_1291) );
DFF_X1 inst_1984 ( .Q(net_2148), .D(net_1039), .CK(net_3183) );
CLKBUF_X2 inst_4101 ( .A(net_3892), .Z(net_3893) );
CLKBUF_X2 inst_3178 ( .A(net_2969), .Z(net_2970) );
CLKBUF_X2 inst_3274 ( .A(net_3065), .Z(net_3066) );
CLKBUF_X2 inst_4203 ( .A(net_3798), .Z(net_3995) );
CLKBUF_X2 inst_2840 ( .A(net_2631), .Z(net_2632) );
NOR2_X4 inst_525 ( .A1(net_1780), .A2(net_1756), .ZN(net_1665) );
CLKBUF_X2 inst_2781 ( .A(net_2552), .Z(net_2573) );
OAI21_X2 inst_434 ( .B2(net_2414), .ZN(net_1925), .A(net_1727), .B1(net_632) );
CLKBUF_X2 inst_3455 ( .A(net_3246), .Z(net_3247) );
NAND2_X2 inst_1032 ( .A2(net_2176), .ZN(net_475), .A1(net_351) );
NAND2_X2 inst_906 ( .A1(net_973), .A2(net_776), .ZN(x3020) );
INV_X4 inst_1248 ( .A(net_2322), .ZN(net_1265) );
AND2_X4 inst_2598 ( .ZN(net_2172), .A1(net_1734), .A2(net_1225) );
AOI22_X2 inst_2402 ( .B1(net_2197), .ZN(net_1630), .A1(net_1621), .B2(net_1535), .A2(net_933) );
INV_X2 inst_1392 ( .A(net_583), .ZN(x981) );
AND2_X2 inst_2616 ( .A1(net_609), .A2(x7087), .ZN(x711) );
CLKBUF_X2 inst_4044 ( .A(net_3445), .Z(net_3836) );
INV_X2 inst_1476 ( .A(net_1536), .ZN(net_735) );
AOI22_X2 inst_2249 ( .B2(net_2124), .A1(net_1967), .B1(net_1474), .ZN(net_1381), .A2(net_1227) );
CLKBUF_X2 inst_3998 ( .A(net_3789), .Z(net_3790) );
DFFR_X1 inst_2113 ( .QN(net_2304), .RN(net_1347), .D(net_945), .CK(net_2486) );
DFF_X2 inst_1820 ( .Q(net_1518), .CK(net_2591), .D(x5846) );
AOI22_X2 inst_2269 ( .B1(net_1768), .ZN(net_1700), .B2(net_1519), .A1(net_1001), .A2(net_917) );
DFF_X2 inst_1780 ( .QN(net_2419), .D(net_754), .CK(net_3457) );
AOI22_X2 inst_2390 ( .B1(net_839), .ZN(net_626), .A1(net_623), .A2(net_313), .B2(net_71) );
INV_X2 inst_1436 ( .A(net_1903), .ZN(net_383) );
OAI22_X2 inst_183 ( .B1(net_1427), .A1(net_529), .B2(net_253), .A2(net_91), .ZN(x1613) );
NAND2_X2 inst_852 ( .A1(net_1841), .ZN(net_1241), .A2(net_1240) );
CLKBUF_X2 inst_3871 ( .A(net_3662), .Z(net_3663) );
INV_X2 inst_1474 ( .A(net_1525), .ZN(net_716) );
AOI22_X2 inst_2271 ( .ZN(net_1689), .A2(net_1548), .B1(net_1001), .A1(net_1000), .B2(net_794) );
DFF_X1 inst_2045 ( .Q(net_2388), .D(net_617), .CK(net_3555) );
DFF_X1 inst_1920 ( .D(net_1243), .QN(net_107), .CK(net_3605) );
CLKBUF_X2 inst_3779 ( .A(net_3364), .Z(net_3571) );
DFF_X1 inst_1848 ( .QN(net_2370), .D(net_1454), .CK(net_3408) );
INV_X4 inst_1311 ( .A(net_2204), .ZN(net_1779) );
NAND3_X2 inst_697 ( .ZN(net_1936), .A2(net_1914), .A1(net_1835), .A3(net_1190) );
CLKBUF_X2 inst_3415 ( .A(net_3206), .Z(net_3207) );
NOR4_X2 inst_487 ( .ZN(net_463), .A1(net_462), .A2(net_461), .A3(net_459), .A4(x3884) );
INV_X2 inst_1640 ( .ZN(net_909), .A(net_60) );
CLKBUF_X2 inst_4143 ( .A(net_3934), .Z(net_3935) );
CLKBUF_X2 inst_3234 ( .A(net_3025), .Z(net_3026) );
AND2_X2 inst_2639 ( .A1(net_775), .A2(x7061), .ZN(x702) );
DFFR_X1 inst_2133 ( .QN(net_2265), .RN(net_1347), .D(net_734), .CK(net_3081) );
AOI221_X2 inst_2509 ( .B2(net_2128), .B1(net_1929), .A(net_1877), .C1(net_1863), .ZN(net_1763), .C2(net_50) );
AOI21_X2 inst_2542 ( .ZN(net_843), .B1(net_680), .A(net_536), .B2(net_445) );
CLKBUF_X2 inst_3091 ( .A(net_2882), .Z(net_2883) );
CLKBUF_X2 inst_4197 ( .A(net_2630), .Z(net_3989) );
OAI21_X2 inst_417 ( .B1(net_768), .ZN(net_752), .A(net_644), .B2(net_509) );
DFF_X1 inst_1861 ( .D(net_1354), .QN(net_114), .CK(net_3844) );
NAND3_X2 inst_671 ( .A2(net_1794), .ZN(net_1071), .A1(net_966), .A3(net_793) );
XNOR2_X2 inst_21 ( .A(net_1734), .B(net_1225), .ZN(net_1170) );
CLKBUF_X2 inst_3570 ( .A(net_3361), .Z(net_3362) );
DFF_X1 inst_2004 ( .QN(net_2230), .D(net_1076), .CK(net_3249) );
AOI22_X2 inst_2311 ( .A2(net_2144), .B1(net_2096), .A1(net_1769), .B2(net_1533), .ZN(net_898) );
CLKBUF_X2 inst_3885 ( .A(net_3648), .Z(net_3677) );
CLKBUF_X2 inst_2857 ( .A(net_2648), .Z(net_2649) );
OAI22_X2 inst_220 ( .B2(net_2279), .B1(net_1865), .ZN(net_959), .A2(net_958), .A1(net_951) );
INV_X2 inst_1585 ( .ZN(net_223), .A(x4974) );
INV_X4 inst_1317 ( .ZN(net_1842), .A(net_1841) );
CLKBUF_X2 inst_3683 ( .A(net_3474), .Z(net_3475) );
CLKBUF_X2 inst_2941 ( .A(net_2732), .Z(net_2733) );
OAI22_X2 inst_245 ( .B2(net_2267), .A2(net_949), .ZN(net_732), .A1(net_714), .B1(net_534) );
DFF_X1 inst_1873 ( .D(net_1332), .QN(net_94), .CK(net_3719) );
CLKBUF_X2 inst_4111 ( .A(net_3902), .Z(net_3903) );
NOR2_X1 inst_624 ( .A2(net_2417), .ZN(net_1712), .A1(net_1579) );
OR2_X1 inst_147 ( .A1(net_1404), .A2(x6063), .ZN(x75) );
OAI22_X1 inst_313 ( .B2(net_2443), .A1(net_2168), .A2(net_1904), .B1(net_529), .ZN(x934) );
INV_X2 inst_1676 ( .ZN(net_1919), .A(net_44) );
CLKBUF_X2 inst_4170 ( .A(net_3478), .Z(net_3962) );
NAND2_X2 inst_1041 ( .A2(net_2327), .ZN(net_1648), .A1(net_1647) );
DFFR_X2 inst_2086 ( .RN(net_1347), .D(net_1113), .QN(net_52), .CK(net_3075) );
CLKBUF_X2 inst_3114 ( .A(net_2712), .Z(net_2906) );
CLKBUF_X2 inst_3577 ( .A(net_2572), .Z(net_3369) );
AND2_X2 inst_2637 ( .A1(net_775), .A2(x7345), .ZN(x828) );
CLKBUF_X2 inst_3624 ( .A(net_2628), .Z(net_3416) );
OAI22_X2 inst_236 ( .B2(net_2258), .ZN(net_750), .A2(net_749), .A1(net_745), .B1(net_534) );
NOR2_X2 inst_553 ( .ZN(net_592), .A1(net_535), .A2(net_409) );
CLKBUF_X2 inst_3878 ( .A(net_3669), .Z(net_3670) );
CLKBUF_X2 inst_3331 ( .A(net_3001), .Z(net_3123) );
OAI22_X2 inst_242 ( .B2(net_2264), .ZN(net_736), .A2(net_735), .A1(net_714), .B1(net_534) );
NAND2_X2 inst_986 ( .A2(net_1554), .A1(net_961), .ZN(net_853) );
CLKBUF_X2 inst_3172 ( .A(net_2963), .Z(net_2964) );
INV_X2 inst_1422 ( .ZN(net_517), .A(net_516) );
CLKBUF_X2 inst_3508 ( .A(net_3299), .Z(net_3300) );
INV_X4 inst_1186 ( .A(net_1914), .ZN(net_1158) );
DFF_X2 inst_1753 ( .QN(net_2346), .D(net_1440), .CK(net_4011) );
DFF_X2 inst_1727 ( .QN(net_2324), .D(net_1504), .CK(net_3318) );
INV_X4 inst_1221 ( .ZN(net_453), .A(net_430) );
INV_X8 inst_1166 ( .ZN(net_1965), .A(net_1964) );
DFF_X2 inst_1739 ( .QN(net_2366), .D(net_1486), .CK(net_3600) );
SDFF_X2 inst_116 ( .SE(net_487), .Q(net_160), .D(net_160), .CK(net_2764), .SI(x4658) );
INV_X8 inst_1133 ( .A(net_1767), .ZN(net_1001) );
OAI211_X2 inst_471 ( .C2(net_2332), .C1(net_1054), .ZN(net_1040), .A(net_894), .B(net_866) );
CLKBUF_X2 inst_4087 ( .A(net_2593), .Z(net_3879) );
DFFR_X1 inst_2103 ( .QN(net_2292), .RN(net_1347), .D(net_956), .CK(net_2647) );
CLKBUF_X2 inst_3609 ( .A(net_2779), .Z(net_3401) );
NAND2_X2 inst_896 ( .A2(net_1697), .A1(net_1696), .ZN(net_1124) );
OAI21_X2 inst_339 ( .B1(net_1507), .ZN(net_1491), .A(net_1456), .B2(net_1045) );
CLKBUF_X2 inst_2664 ( .A(net_2455), .Z(net_2456) );
OAI21_X2 inst_351 ( .B2(net_2406), .ZN(net_1445), .B1(net_1441), .A(net_1394) );
AND2_X2 inst_2608 ( .A1(net_594), .A2(x5118), .ZN(x910) );
AOI21_X2 inst_2557 ( .ZN(net_2056), .B2(net_2055), .B1(net_2054), .A(net_515) );
AOI21_X2 inst_2521 ( .A(net_1785), .B1(net_910), .ZN(net_814), .B2(net_813) );
OAI21_X2 inst_385 ( .A(net_2434), .ZN(net_1351), .B1(net_1168), .B2(net_82) );
CLKBUF_X2 inst_3319 ( .A(net_3110), .Z(net_3111) );
CLKBUF_X2 inst_2653 ( .A(net_2444), .Z(net_2445) );
AOI21_X2 inst_2550 ( .B2(net_1904), .A(net_1753), .ZN(net_477), .B1(net_375) );
INV_X2 inst_1560 ( .ZN(net_240), .A(x6303) );
CLKBUF_X2 inst_3932 ( .A(net_3723), .Z(net_3724) );
NOR2_X2 inst_596 ( .A2(net_2265), .ZN(net_1885), .A1(net_520) );
CLKBUF_X2 inst_2771 ( .A(net_2562), .Z(net_2563) );
DFFR_X1 inst_2142 ( .QN(net_2276), .RN(net_1347), .D(net_712), .CK(net_2464) );
INV_X1 inst_1705 ( .A(net_83), .ZN(x15) );
NAND2_X2 inst_847 ( .A1(net_1840), .ZN(net_1266), .A2(net_1263) );
CLKBUF_X2 inst_2720 ( .A(net_2511), .Z(net_2512) );
DFF_X1 inst_1942 ( .Q(net_2108), .D(net_1038), .CK(net_2974) );
HA_X1 inst_1716 ( .A(net_2171), .S(net_1651), .CO(net_1650), .B(net_1265) );
CLKBUF_X2 inst_3253 ( .A(net_2615), .Z(net_3045) );
AND2_X2 inst_2648 ( .A1(net_2017), .A2(x3134), .ZN(x2416) );
INV_X8 inst_1146 ( .ZN(net_1402), .A(net_1020) );
NAND4_X2 inst_637 ( .A2(net_2050), .ZN(net_1912), .A4(net_1909), .A3(net_1284), .A1(net_522) );
CLKBUF_X2 inst_3708 ( .A(net_2537), .Z(net_3500) );
NOR2_X2 inst_547 ( .A1(net_1970), .ZN(net_640), .A2(net_621) );
CLKBUF_X2 inst_4023 ( .A(net_3814), .Z(net_3815) );
CLKBUF_X2 inst_3105 ( .A(net_2624), .Z(net_2897) );
CLKBUF_X2 inst_3673 ( .A(net_3464), .Z(net_3465) );
CLKBUF_X2 inst_3781 ( .A(net_3572), .Z(net_3573) );
CLKBUF_X2 inst_3539 ( .A(net_2566), .Z(net_3331) );
AOI222_X2 inst_2457 ( .C1(net_2017), .A2(net_1566), .A1(net_590), .B1(net_589), .ZN(net_579), .B2(net_168), .C2(x5413) );
CLKBUF_X2 inst_3552 ( .A(net_3343), .Z(net_3344) );
INV_X16 inst_1702 ( .ZN(net_2104), .A(net_2103) );
OAI22_X2 inst_274 ( .B2(net_2309), .B1(net_1865), .ZN(net_1606), .A1(net_951), .A2(net_705) );
INV_X2 inst_1607 ( .ZN(net_206), .A(x4866) );
INV_X4 inst_1277 ( .ZN(net_298), .A(net_52) );
CLKBUF_X2 inst_2817 ( .A(net_2608), .Z(net_2609) );
CLKBUF_X2 inst_4076 ( .A(net_3867), .Z(net_3868) );
DFFR_X2 inst_2092 ( .D(net_2048), .RN(net_1347), .QN(net_56), .CK(net_3272) );
OAI22_X2 inst_164 ( .B1(net_1407), .A1(net_1405), .B2(net_197), .A2(net_132), .ZN(x317) );
CLKBUF_X2 inst_3207 ( .A(net_2998), .Z(net_2999) );
CLKBUF_X2 inst_3143 ( .A(net_2934), .Z(net_2935) );
DFF_X1 inst_1854 ( .QN(net_2358), .D(net_1430), .CK(net_3941) );
CLKBUF_X2 inst_2696 ( .A(net_2487), .Z(net_2488) );
INV_X1 inst_1710 ( .ZN(net_2026), .A(net_2025) );
AOI22_X2 inst_2407 ( .B1(net_2197), .ZN(net_1635), .A1(net_1621), .B2(net_1513), .A2(net_1213) );
DFF_X2 inst_1771 ( .QN(net_2380), .D(net_921), .CK(net_3864) );
CLKBUF_X2 inst_2880 ( .A(net_2671), .Z(net_2672) );
INV_X2 inst_1440 ( .A(net_1532), .ZN(net_730) );
CLKBUF_X2 inst_2660 ( .A(net_2450), .Z(net_2452) );
CLKBUF_X2 inst_3142 ( .A(net_2933), .Z(net_2934) );
AOI22_X2 inst_2305 ( .A2(net_2113), .B1(net_2096), .A1(net_1769), .B2(net_1538), .ZN(net_904) );
CLKBUF_X2 inst_3355 ( .A(net_2929), .Z(net_3147) );
NAND2_X4 inst_753 ( .ZN(net_2007), .A2(net_419), .A1(net_405) );
DFFR_X1 inst_2150 ( .QN(net_2257), .RN(net_1347), .D(net_698), .CK(net_2789) );
AOI22_X2 inst_2389 ( .A1(net_1718), .B1(net_1450), .B2(net_790), .ZN(net_627), .A2(net_398) );
CLKBUF_X2 inst_3427 ( .A(net_2687), .Z(net_3219) );
NAND2_X2 inst_946 ( .ZN(net_996), .A1(net_841), .A2(net_662) );
DFF_X1 inst_1954 ( .Q(net_2120), .D(net_1067), .CK(net_3559) );
AOI22_X2 inst_2260 ( .B2(net_2134), .B1(net_1915), .ZN(net_1370), .A2(net_1367), .A1(net_1189) );
DFFR_X1 inst_2148 ( .QN(net_2255), .RN(net_1347), .D(net_700), .CK(net_3335) );
CLKBUF_X2 inst_3941 ( .A(net_3732), .Z(net_3733) );
CLKBUF_X2 inst_2900 ( .A(net_2691), .Z(net_2692) );
INV_X2 inst_1591 ( .ZN(net_218), .A(x4821) );
CLKBUF_X2 inst_3247 ( .A(net_3038), .Z(net_3039) );
CLKBUF_X2 inst_3697 ( .A(net_2881), .Z(net_3489) );
CLKBUF_X2 inst_3858 ( .A(net_3649), .Z(net_3650) );
OAI21_X2 inst_379 ( .A(net_1940), .B1(net_1839), .ZN(net_1358), .B2(net_1356) );
NAND2_X2 inst_926 ( .A2(net_1634), .ZN(net_1088), .A1(net_831) );
CLKBUF_X2 inst_3922 ( .A(net_3713), .Z(net_3714) );
DFF_X1 inst_2053 ( .D(net_521), .QN(net_46), .CK(net_3699) );
INV_X4 inst_1325 ( .ZN(net_1948), .A(net_1582) );
AND4_X4 inst_2570 ( .A4(net_2427), .A1(net_2426), .A3(net_2425), .A2(net_2424), .ZN(net_2087) );
CLKBUF_X2 inst_4153 ( .A(net_3944), .Z(net_3945) );
CLKBUF_X2 inst_3312 ( .A(net_2532), .Z(net_3104) );
CLKBUF_X2 inst_3646 ( .A(net_3437), .Z(net_3438) );
CLKBUF_X2 inst_3719 ( .A(net_3431), .Z(net_3511) );
NAND2_X2 inst_891 ( .A2(net_1693), .A1(net_1692), .ZN(net_1129) );
CLKBUF_X2 inst_4095 ( .A(net_3886), .Z(net_3887) );
SDFF_X2 inst_74 ( .Q(net_1561), .D(net_1561), .SE(net_491), .CK(net_2905), .SI(x7145) );
INV_X4 inst_1235 ( .A(net_531), .ZN(net_409) );
AOI22_X2 inst_2244 ( .B2(net_2130), .A1(net_1967), .B1(net_1450), .ZN(net_1386), .A2(net_932) );
CLKBUF_X2 inst_3561 ( .A(net_3352), .Z(net_3353) );
OAI22_X2 inst_288 ( .A1(net_1615), .B1(net_1404), .B2(net_205), .A2(net_123), .ZN(x461) );
CLKBUF_X2 inst_3284 ( .A(net_2599), .Z(net_3076) );
CLKBUF_X2 inst_3046 ( .A(net_2837), .Z(net_2838) );
CLKBUF_X2 inst_3626 ( .A(net_3417), .Z(net_3418) );
CLKBUF_X2 inst_4036 ( .A(net_3361), .Z(net_3828) );
INV_X4 inst_1298 ( .A(net_2357), .ZN(net_1238) );
CLKBUF_X2 inst_3757 ( .A(net_3471), .Z(net_3549) );
NAND2_X2 inst_917 ( .A1(net_972), .A2(net_774), .ZN(x3041) );
CLKBUF_X2 inst_3712 ( .A(net_3096), .Z(net_3504) );
DFF_X2 inst_1743 ( .QN(net_2363), .D(net_1421), .CK(net_3636) );
OAI21_X2 inst_372 ( .B2(net_2407), .B1(net_1443), .ZN(net_1417), .A(net_1393) );
INV_X2 inst_1600 ( .ZN(net_210), .A(x6400) );
OAI22_X2 inst_215 ( .A2(net_2233), .B1(net_1406), .A1(net_1405), .B2(net_179), .ZN(x1937) );
CLKBUF_X2 inst_2850 ( .A(net_2641), .Z(net_2642) );
AND2_X2 inst_2624 ( .A1(net_594), .A2(x7442), .ZN(x870) );
NAND2_X2 inst_849 ( .A2(net_1910), .A1(net_1840), .ZN(net_1257) );
DFF_X2 inst_1775 ( .QN(net_2421), .D(net_882), .CK(net_3461) );
AOI22_X2 inst_2397 ( .B1(net_2197), .ZN(net_1625), .A1(net_1621), .B2(net_1514), .A2(net_1240) );
XOR2_X2 inst_3 ( .A(net_2313), .B(net_2312), .Z(net_392) );
INV_X8 inst_1172 ( .ZN(net_2008), .A(net_2007) );
NAND2_X2 inst_1090 ( .A2(net_2417), .ZN(net_1871), .A1(net_1579) );
CLKBUF_X2 inst_3060 ( .A(net_2851), .Z(net_2852) );
CLKBUF_X2 inst_3903 ( .A(net_3694), .Z(net_3695) );
AOI22_X2 inst_2372 ( .B2(net_2130), .A1(net_2038), .A2(net_1563), .B1(net_979), .ZN(net_684) );
AND3_X2 inst_2575 ( .ZN(net_2067), .A3(net_2066), .A2(net_614), .A1(net_522) );
NOR2_X2 inst_566 ( .A1(net_2165), .A2(net_601), .ZN(net_403) );
INV_X2 inst_1399 ( .A(net_576), .ZN(x1044) );
INV_X4 inst_1239 ( .ZN(net_1048), .A(net_363) );
CLKBUF_X2 inst_3126 ( .A(net_2917), .Z(net_2918) );
NOR2_X4 inst_503 ( .A2(net_2333), .ZN(net_1233), .A1(net_1182) );
AOI22_X2 inst_2333 ( .B2(net_2127), .A1(net_2038), .A2(net_1557), .B1(net_979), .ZN(net_831) );
DFF_X1 inst_1936 ( .D(net_1125), .QN(net_66), .CK(net_3494) );
CLKBUF_X2 inst_3193 ( .A(net_2944), .Z(net_2985) );
CLKBUF_X2 inst_4193 ( .A(net_3043), .Z(net_3985) );
DFFR_X1 inst_2099 ( .QN(net_2279), .RN(net_1347), .D(net_959), .CK(net_3340) );
CLKBUF_X2 inst_4069 ( .A(net_3860), .Z(net_3861) );
NAND2_X2 inst_1097 ( .ZN(net_1932), .A2(net_1588), .A1(net_226) );
NAND3_X2 inst_686 ( .A1(net_1935), .A2(net_1901), .ZN(net_1616), .A3(net_469) );
CLKBUF_X2 inst_4016 ( .A(net_2816), .Z(net_3808) );
DFF_X2 inst_1732 ( .QN(net_2320), .D(net_1495), .CK(net_3317) );
CLKBUF_X2 inst_2914 ( .A(net_2705), .Z(net_2706) );
CLKBUF_X2 inst_2888 ( .A(net_2679), .Z(net_2680) );
CLKBUF_X2 inst_3294 ( .A(net_3085), .Z(net_3086) );
CLKBUF_X2 inst_2741 ( .A(net_2519), .Z(net_2533) );
CLKBUF_X2 inst_3643 ( .A(net_2688), .Z(net_3435) );
NAND2_X2 inst_967 ( .A2(net_1559), .A1(net_961), .ZN(net_872) );
DFFR_X1 inst_2119 ( .QN(net_2282), .RN(net_1347), .D(net_942), .CK(net_2609) );
DFF_X1 inst_1929 ( .D(net_1128), .QN(net_68), .CK(net_3265) );
INV_X2 inst_1522 ( .ZN(net_390), .A(x3961) );
CLKBUF_X2 inst_3391 ( .A(net_3182), .Z(net_3183) );
DFF_X2 inst_1794 ( .QN(net_2244), .D(net_456), .CK(net_2824) );
INV_X4 inst_1227 ( .A(net_1716), .ZN(net_413) );
AOI22_X2 inst_2324 ( .A2(net_2152), .B1(net_2096), .A1(net_1769), .B2(net_1520), .ZN(net_885) );
CLKBUF_X2 inst_3069 ( .A(net_2445), .Z(net_2861) );
CLKBUF_X2 inst_3631 ( .A(net_3422), .Z(net_3423) );
NAND2_X2 inst_1101 ( .A2(net_2209), .A1(net_2206), .ZN(net_1981) );
CLKBUF_X2 inst_3047 ( .A(net_2838), .Z(net_2839) );
CLKBUF_X2 inst_2950 ( .A(net_2741), .Z(net_2742) );
CLKBUF_X2 inst_3847 ( .A(net_3638), .Z(net_3639) );
CLKBUF_X2 inst_2897 ( .A(net_2546), .Z(net_2689) );
NAND2_X2 inst_861 ( .A1(net_1838), .ZN(net_1223), .A2(net_1222) );
AOI21_X2 inst_2529 ( .A(net_1785), .B1(net_910), .ZN(net_804), .B2(net_76) );
DFF_X2 inst_1787 ( .QN(net_2426), .D(net_769), .CK(net_3661) );
CLKBUF_X2 inst_2990 ( .A(net_2781), .Z(net_2782) );
INV_X4 inst_1283 ( .ZN(net_276), .A(net_53) );
AOI222_X2 inst_2451 ( .C1(net_2016), .A2(net_1572), .A1(net_590), .B1(net_589), .ZN(net_585), .B2(net_174), .C2(x5269) );
INV_X4 inst_1202 ( .A(net_2015), .ZN(net_1404) );
INV_X2 inst_1540 ( .ZN(net_256), .A(x4843) );
AOI22_X2 inst_2227 ( .B2(net_2152), .A1(net_2040), .B1(net_1450), .ZN(net_1449), .A2(net_1284) );
INV_X2 inst_1660 ( .A(net_1840), .ZN(net_1744) );
CLKBUF_X2 inst_2742 ( .A(net_2533), .Z(net_2534) );
CLKBUF_X2 inst_3536 ( .A(net_3068), .Z(net_3328) );
NAND3_X2 inst_660 ( .A2(net_1807), .A1(net_1761), .ZN(net_1082), .A3(net_812) );
AOI222_X1 inst_2490 ( .B1(net_1995), .A1(net_1751), .B2(net_1561), .C1(net_1020), .ZN(net_1010), .A2(net_163), .C2(x3447) );
NOR2_X4 inst_517 ( .ZN(net_486), .A1(net_457), .A2(net_424) );
INV_X2 inst_1576 ( .ZN(net_229), .A(x4336) );
AOI22_X2 inst_2346 ( .B1(net_2197), .A1(net_2038), .A2(net_1553), .B2(net_1542), .ZN(net_818) );
INV_X4 inst_1261 ( .A(net_2385), .ZN(net_333) );
CLKBUF_X2 inst_3462 ( .A(net_3253), .Z(net_3254) );
OAI22_X2 inst_310 ( .B1(net_1895), .A1(net_1403), .B2(net_260), .A2(net_139), .ZN(x169) );
NAND2_X2 inst_794 ( .A2(net_1680), .ZN(net_1319), .A1(net_1275) );
CLKBUF_X2 inst_2754 ( .A(net_2545), .Z(net_2546) );
NAND2_X2 inst_1005 ( .A2(net_2114), .A1(net_979), .ZN(net_667) );
CLKBUF_X2 inst_2759 ( .A(net_2451), .Z(net_2551) );
INV_X8 inst_1147 ( .A(net_2168), .ZN(net_1020) );
DFF_X2 inst_1768 ( .QN(net_2385), .D(net_996), .CK(net_3866) );
INV_X2 inst_1580 ( .A(net_1589), .ZN(net_226) );
DFF_X1 inst_1842 ( .QN(net_2326), .D(net_1509), .CK(net_3047) );
CLKBUF_X2 inst_2688 ( .A(net_2479), .Z(net_2480) );
CLKBUF_X2 inst_2917 ( .A(net_2578), .Z(net_2709) );
AOI22_X2 inst_2423 ( .B2(net_2151), .B1(net_1974), .ZN(net_1797), .A1(net_1791), .A2(net_299) );
INV_X2 inst_1408 ( .A(net_568), .ZN(x1187) );
NAND2_X2 inst_996 ( .A1(net_1796), .ZN(net_835), .A2(net_675) );
AOI22_X2 inst_2351 ( .A1(net_783), .B1(net_782), .ZN(net_781), .A2(net_398), .B2(x3669) );
DFF_X1 inst_1853 ( .D(net_1432), .QN(net_315), .CK(net_3696) );
DFF_X1 inst_1889 ( .D(net_1344), .QN(net_123), .CK(net_3758) );
INV_X2 inst_1527 ( .A(net_2308), .ZN(net_311) );
DFF_X1 inst_2011 ( .QN(net_2217), .D(net_1070), .CK(net_3485) );
DFF_X2 inst_1761 ( .Q(net_2412), .D(net_1840), .CK(net_3899) );
NAND2_X4 inst_740 ( .A1(net_2094), .ZN(net_1930), .A2(net_1772) );
OAI22_X2 inst_264 ( .B2(net_2257), .A2(net_848), .A1(net_714), .ZN(net_698), .B1(net_534) );
CLKBUF_X2 inst_3703 ( .A(net_2553), .Z(net_3495) );
CLKBUF_X2 inst_4189 ( .A(net_3980), .Z(net_3981) );
SDFF_X2 inst_84 ( .Q(net_1558), .D(net_1558), .SE(net_491), .CK(net_2901), .SI(x7215) );
INV_X4 inst_1333 ( .ZN(net_2013), .A(net_2012) );
DFF_X1 inst_1937 ( .D(net_1122), .QN(net_67), .CK(net_3261) );
OAI22_X2 inst_173 ( .A1(net_1426), .B1(net_1402), .B2(net_189), .A2(net_108), .ZN(x1402) );
CLKBUF_X2 inst_3710 ( .A(net_3501), .Z(net_3502) );
NOR2_X2 inst_611 ( .A2(net_2264), .ZN(net_1985), .A1(net_520) );
CLKBUF_X2 inst_3953 ( .A(net_2547), .Z(net_3745) );
AOI222_X1 inst_2487 ( .B1(net_1995), .A1(net_1751), .B2(net_1563), .C1(net_1020), .ZN(net_1013), .A2(net_165), .C2(x3411) );
INV_X2 inst_1551 ( .ZN(net_249), .A(x3067) );
INV_X4 inst_1260 ( .A(net_2085), .ZN(net_372) );
NAND2_X2 inst_1088 ( .ZN(net_1854), .A2(net_1853), .A1(net_678) );
DFF_X1 inst_1943 ( .Q(net_2109), .D(net_1026), .CK(net_3379) );
NOR3_X4 inst_490 ( .A1(net_1780), .A3(net_1755), .ZN(net_533), .A2(net_515) );
CLKBUF_X2 inst_3332 ( .A(net_2480), .Z(net_3124) );
CLKBUF_X2 inst_2717 ( .A(net_2508), .Z(net_2509) );
AOI22_X2 inst_2218 ( .A2(net_2388), .B2(net_2156), .A1(net_1960), .B1(net_1915), .ZN(net_1462) );
CLKBUF_X2 inst_4176 ( .A(net_3967), .Z(net_3968) );
OR3_X2 inst_129 ( .ZN(net_347), .A3(net_77), .A1(net_74), .A2(net_73) );
INV_X4 inst_1309 ( .A(net_1750), .ZN(net_1749) );
CLKBUF_X2 inst_2740 ( .A(net_2515), .Z(net_2532) );
DFF_X2 inst_1754 ( .QN(net_2347), .D(net_1439), .CK(net_4006) );
INV_X2 inst_1531 ( .A(net_2300), .ZN(net_335) );
CLKBUF_X2 inst_2931 ( .A(net_2722), .Z(net_2723) );
AOI21_X2 inst_2530 ( .A(net_1785), .B1(net_910), .ZN(net_803), .B2(net_77) );
CLKBUF_X2 inst_2727 ( .A(net_2518), .Z(net_2519) );
CLKBUF_X2 inst_2922 ( .A(net_2713), .Z(net_2714) );
CLKBUF_X2 inst_3803 ( .A(net_3594), .Z(net_3595) );
CLKBUF_X2 inst_3183 ( .A(net_2532), .Z(net_2975) );
INV_X2 inst_1503 ( .A(net_2428), .ZN(net_681) );
NAND2_X2 inst_777 ( .A2(net_1367), .ZN(net_1364), .A1(net_1188) );
CLKBUF_X2 inst_3802 ( .A(net_3593), .Z(net_3594) );
NAND2_X2 inst_1037 ( .A1(net_2414), .A2(net_1575), .ZN(net_354) );
NAND2_X2 inst_933 ( .A2(net_1625), .ZN(net_1067), .A1(net_691) );
OAI22_X2 inst_300 ( .B2(net_2439), .B1(net_2017), .A1(net_1895), .A2(net_1778), .ZN(x2451) );
CLKBUF_X2 inst_3596 ( .A(net_2813), .Z(net_3388) );
CLKBUF_X2 inst_3724 ( .A(net_3515), .Z(net_3516) );
INV_X4 inst_1250 ( .A(net_2328), .ZN(net_1263) );
INV_X4 inst_1226 ( .ZN(net_419), .A(net_418) );
NAND2_X2 inst_1013 ( .A2(net_1592), .ZN(net_638), .A1(net_604) );
OAI21_X1 inst_446 ( .B2(net_2380), .B1(net_2379), .A(net_492), .ZN(net_471) );
DFF_X1 inst_1979 ( .Q(net_2144), .D(net_1028), .CK(net_2997) );
OAI21_X2 inst_364 ( .B2(net_2411), .B1(net_1441), .ZN(net_1430), .A(net_1389) );
CLKBUF_X2 inst_3613 ( .A(net_3313), .Z(net_3405) );
AOI22_X2 inst_2354 ( .A1(net_783), .ZN(net_778), .B1(net_775), .A2(net_350), .B2(x3758) );
NAND2_X2 inst_824 ( .A1(net_1840), .ZN(net_1335), .A2(net_1186) );
CLKBUF_X2 inst_2997 ( .A(net_2788), .Z(net_2789) );
CLKBUF_X2 inst_3533 ( .A(net_3324), .Z(net_3325) );
OAI21_X2 inst_411 ( .B1(net_768), .ZN(net_758), .A(net_645), .B2(net_494) );
SDFFR_X1 inst_124 ( .SE(net_1829), .D(net_1536), .RN(net_1347), .SI(net_51), .Q(net_51), .CK(net_3024) );
CLKBUF_X2 inst_3515 ( .A(net_3306), .Z(net_3307) );
CLKBUF_X2 inst_3750 ( .A(net_3541), .Z(net_3542) );
CLKBUF_X2 inst_4026 ( .A(net_3817), .Z(net_3818) );
CLKBUF_X2 inst_4056 ( .A(net_3456), .Z(net_3848) );
CLKBUF_X2 inst_3430 ( .A(net_3221), .Z(net_3222) );
CLKBUF_X2 inst_3869 ( .A(net_3660), .Z(net_3661) );
CLKBUF_X2 inst_3488 ( .A(net_3279), .Z(net_3280) );
INV_X4 inst_1270 ( .ZN(net_317), .A(net_56) );
CLKBUF_X2 inst_3448 ( .A(net_3239), .Z(net_3240) );
CLKBUF_X2 inst_3439 ( .A(net_3230), .Z(net_3231) );
SDFF_X2 inst_61 ( .Q(net_1557), .D(net_1557), .SE(net_498), .CK(net_2924), .SI(x7241) );
OAI22_X2 inst_203 ( .A2(net_2228), .A1(net_1408), .B1(net_1407), .B2(net_231), .ZN(x2050) );
INV_X8 inst_1139 ( .ZN(net_655), .A(net_520) );
INV_X2 inst_1519 ( .A(net_1576), .ZN(net_291) );
DFFR_X1 inst_2156 ( .QN(net_2264), .RN(net_1347), .D(net_736), .CK(net_2786) );
INV_X2 inst_1571 ( .ZN(net_454), .A(x6039) );
OAI211_X2 inst_456 ( .C2(net_2354), .C1(net_1639), .ZN(net_1095), .A(net_817), .B(net_672) );
NAND2_X2 inst_832 ( .A1(net_1840), .ZN(net_1282), .A2(net_328) );
AOI221_X2 inst_2515 ( .B2(net_2119), .ZN(net_1993), .A(net_1992), .B1(net_1929), .C1(net_1863), .C2(net_601) );
INV_X2 inst_1491 ( .A(net_2318), .ZN(net_1242) );
INV_X2 inst_1402 ( .A(net_573), .ZN(x1071) );
OAI22_X2 inst_275 ( .B2(net_2308), .B1(net_1865), .ZN(net_1607), .A1(net_951), .A2(net_709) );
SDFF_X2 inst_117 ( .Q(net_1556), .D(net_1556), .SE(net_491), .CK(net_2660), .SI(x7264) );
CLKBUF_X2 inst_2676 ( .A(net_2467), .Z(net_2468) );
CLKBUF_X2 inst_3106 ( .A(net_2897), .Z(net_2898) );
CLKBUF_X2 inst_3728 ( .A(net_3466), .Z(net_3520) );
OAI22_X2 inst_154 ( .B1(net_1428), .A1(net_529), .B2(net_391), .A2(net_111), .ZN(x1371) );
AOI22_X2 inst_2416 ( .B2(net_2141), .B1(net_1974), .A1(net_1789), .ZN(net_1662), .A2(net_326) );
CLKBUF_X2 inst_3812 ( .A(net_3603), .Z(net_3604) );
CLKBUF_X2 inst_4106 ( .A(net_3897), .Z(net_3898) );
OAI211_X2 inst_465 ( .C1(net_1054), .ZN(net_1049), .C2(net_1048), .A(net_907), .B(net_863) );
AOI22_X2 inst_2304 ( .A2(net_2140), .B1(net_2096), .A1(net_1769), .B2(net_1540), .ZN(net_905) );
CLKBUF_X2 inst_3959 ( .A(net_3362), .Z(net_3751) );
AOI221_X2 inst_2503 ( .C2(net_2165), .B2(net_2118), .B1(net_1929), .A(net_1879), .C1(net_1863), .ZN(net_966) );
DFF_X2 inst_1790 ( .QN(net_1590), .D(net_483), .CK(net_3996) );
SDFF_X2 inst_94 ( .SE(net_488), .Q(net_170), .D(net_170), .CK(net_2711), .SI(x4416) );
CLKBUF_X2 inst_3214 ( .A(net_3005), .Z(net_3006) );
DFF_X1 inst_1905 ( .D(net_1312), .QN(net_135), .CK(net_3446) );
AOI22_X2 inst_2264 ( .B1(net_1768), .ZN(net_1694), .B2(net_1542), .A1(net_1001), .A2(net_813) );
INV_X2 inst_1378 ( .A(net_1006), .ZN(x2739) );
OAI22_X2 inst_243 ( .B2(net_2265), .A2(net_953), .A1(net_740), .ZN(net_734), .B1(net_534) );
OAI21_X2 inst_424 ( .ZN(net_428), .B1(net_426), .B2(x6188), .A(x5995) );
NOR2_X2 inst_591 ( .A2(net_2256), .ZN(net_1880), .A1(net_520) );
CLKBUF_X2 inst_2697 ( .A(net_2488), .Z(net_2489) );
CLKBUF_X2 inst_3166 ( .A(net_2957), .Z(net_2958) );
XNOR2_X2 inst_15 ( .B(net_1276), .ZN(net_1254), .A(net_1233) );
CLKBUF_X2 inst_3747 ( .A(net_3267), .Z(net_3539) );
CLKBUF_X2 inst_3656 ( .A(net_3128), .Z(net_3448) );
AOI22_X2 inst_2237 ( .B2(net_2126), .A1(net_1967), .A2(net_1845), .B1(net_1474), .ZN(net_1393) );
CLKBUF_X2 inst_3496 ( .A(net_3287), .Z(net_3288) );
DFFR_X1 inst_2123 ( .QN(net_2288), .RN(net_1347), .D(net_935), .CK(net_2806) );
CLKBUF_X2 inst_3229 ( .A(net_3020), .Z(net_3021) );
CLKBUF_X2 inst_2706 ( .A(net_2489), .Z(net_2498) );
OAI211_X2 inst_476 ( .C2(net_2318), .C1(net_1054), .ZN(net_1033), .A(net_889), .B(net_856) );
CLKBUF_X2 inst_4135 ( .A(net_3926), .Z(net_3927) );
CLKBUF_X2 inst_3742 ( .A(net_3533), .Z(net_3534) );
AOI221_X2 inst_2499 ( .B2(net_2120), .B1(net_1929), .A(net_1880), .C1(net_1863), .ZN(net_983), .C2(net_324) );
CLKBUF_X2 inst_2827 ( .A(net_2527), .Z(net_2619) );
XNOR2_X2 inst_20 ( .ZN(net_1174), .A(net_1171), .B(net_401) );
AOI222_X2 inst_2448 ( .C1(net_2017), .A2(net_1543), .A1(net_590), .B1(net_589), .ZN(net_588), .B2(net_145), .C2(x5934) );
INV_X2 inst_1369 ( .A(net_1015), .ZN(x2611) );
CLKBUF_X2 inst_3988 ( .A(net_3779), .Z(net_3780) );
OAI21_X2 inst_349 ( .B2(net_2370), .ZN(net_1454), .A(net_1400), .B1(net_1368) );
AOI21_X2 inst_2541 ( .A(net_2382), .ZN(net_763), .B1(net_620), .B2(net_615) );
NOR2_X2 inst_576 ( .A1(net_2323), .A2(net_2322), .ZN(net_1652) );
INV_X16 inst_1693 ( .ZN(net_1838), .A(net_1836) );
CLKBUF_X2 inst_4235 ( .A(net_4026), .Z(net_4027) );
AOI211_X2 inst_2561 ( .C2(net_2135), .C1(net_1929), .A(net_1883), .B(net_1785), .ZN(net_677) );
CLKBUF_X2 inst_3306 ( .A(net_3097), .Z(net_3098) );
NAND2_X2 inst_1020 ( .A2(net_2169), .ZN(net_611), .A1(net_539) );
CLKBUF_X2 inst_2876 ( .A(net_2667), .Z(net_2668) );
CLKBUF_X2 inst_3055 ( .A(net_2602), .Z(net_2847) );
NAND2_X2 inst_976 ( .A2(net_1569), .A1(net_961), .ZN(net_863) );
CLKBUF_X2 inst_3952 ( .A(net_3743), .Z(net_3744) );
CLKBUF_X2 inst_4226 ( .A(net_4017), .Z(net_4018) );
INV_X4 inst_1279 ( .A(net_1735), .ZN(net_359) );
AOI22_X2 inst_2252 ( .B2(net_2116), .A1(net_1967), .B1(net_1474), .ZN(net_1378), .A2(net_1291) );
CLKBUF_X2 inst_3588 ( .A(net_2886), .Z(net_3380) );
NAND2_X2 inst_1096 ( .ZN(net_1923), .A1(net_1922), .A2(net_84) );
CLKBUF_X2 inst_4229 ( .A(net_3218), .Z(net_4021) );
AOI22_X2 inst_2238 ( .B2(net_2127), .A1(net_1967), .B1(net_1474), .ZN(net_1392), .A2(net_1197) );
CLKBUF_X2 inst_2763 ( .A(net_2554), .Z(net_2555) );
DFF_X2 inst_1839 ( .Q(net_1538), .CK(net_2581), .D(x5605) );
CLKBUF_X2 inst_3151 ( .A(net_2842), .Z(net_2943) );
NAND2_X4 inst_761 ( .A2(net_2418), .ZN(net_2053), .A1(net_2051) );
CLKBUF_X2 inst_3399 ( .A(net_2772), .Z(net_3191) );
CLKBUF_X2 inst_3414 ( .A(net_3205), .Z(net_3206) );
CLKBUF_X2 inst_2803 ( .A(net_2594), .Z(net_2595) );
INV_X2 inst_1432 ( .A(net_1190), .ZN(net_1105) );
NAND2_X4 inst_725 ( .A2(net_1914), .A1(net_1729), .ZN(net_1684) );
CLKBUF_X2 inst_4120 ( .A(net_3911), .Z(net_3912) );
CLKBUF_X2 inst_3084 ( .A(net_2875), .Z(net_2876) );
AOI22_X2 inst_2259 ( .B2(net_2123), .A1(net_1967), .B1(net_1450), .ZN(net_1371), .A2(net_1222) );
INV_X4 inst_1337 ( .ZN(net_2023), .A(net_1777) );
AOI222_X2 inst_2464 ( .C1(net_2016), .A2(net_1559), .A1(net_590), .B1(net_589), .ZN(net_572), .B2(net_161), .C2(x5556) );
AND2_X2 inst_2641 ( .A1(net_2013), .A2(x6706), .ZN(x564) );
CLKBUF_X2 inst_3096 ( .A(net_2509), .Z(net_2888) );
CLKBUF_X2 inst_3015 ( .A(net_2772), .Z(net_2807) );
CLKBUF_X2 inst_4010 ( .A(net_2894), .Z(net_3802) );
INV_X2 inst_1638 ( .ZN(net_185), .A(x6470) );
CLKBUF_X2 inst_3328 ( .A(net_2850), .Z(net_3120) );
AOI22_X2 inst_2441 ( .ZN(net_1897), .A1(net_1789), .B1(net_655), .A2(net_310), .B2(net_305) );
NAND2_X2 inst_1111 ( .ZN(net_2042), .A2(net_1869), .A1(net_417) );
CLKBUF_X2 inst_3220 ( .A(net_3011), .Z(net_3012) );
CLKBUF_X2 inst_2658 ( .A(net_2449), .Z(net_2450) );
NAND2_X2 inst_878 ( .ZN(net_1191), .A1(net_1180), .A2(net_277) );
OAI211_X2 inst_480 ( .C2(net_2329), .C1(net_1052), .ZN(net_1028), .A(net_898), .B(net_869) );
DFF_X1 inst_1926 ( .QN(net_2201), .D(net_1139), .CK(net_3970) );
NOR2_X2 inst_564 ( .A2(net_2348), .A1(net_457), .ZN(net_435) );
CLKBUF_X2 inst_2986 ( .A(net_2777), .Z(net_2778) );
AOI22_X2 inst_2206 ( .B2(net_2150), .A1(net_1960), .ZN(net_1475), .B1(net_1474), .A2(net_1179) );
CLKBUF_X2 inst_2792 ( .A(net_2583), .Z(net_2584) );
NAND2_X4 inst_739 ( .ZN(net_1931), .A1(net_1930), .A2(net_1591) );
CLKBUF_X2 inst_3862 ( .A(net_3056), .Z(net_3654) );
SDFF_X2 inst_46 ( .SE(net_1768), .SI(net_1526), .Q(net_80), .D(net_80), .CK(net_3166) );
NAND2_X2 inst_934 ( .A2(net_1624), .ZN(net_1066), .A1(net_833) );
AOI21_X2 inst_2537 ( .A(net_1785), .B1(net_910), .ZN(net_793), .B2(net_792) );
NAND2_X2 inst_1000 ( .A1(net_1669), .ZN(net_760), .A2(net_317) );
NAND2_X1 inst_1126 ( .A1(net_1977), .A2(net_1904), .ZN(net_1667) );
CLKBUF_X2 inst_3470 ( .A(net_3149), .Z(net_3262) );
NAND2_X2 inst_796 ( .ZN(net_1317), .A1(net_1283), .A2(net_1230) );
AND2_X4 inst_2585 ( .A2(net_2423), .A1(net_2421), .ZN(net_272) );
NAND4_X2 inst_633 ( .A2(net_2200), .A4(net_2173), .ZN(net_1776), .A3(net_1775), .A1(net_1774) );
AOI22_X2 inst_2364 ( .B2(net_2119), .A1(net_2038), .A2(net_1550), .B1(net_979), .ZN(net_693) );
NOR2_X4 inst_524 ( .A2(net_2324), .ZN(net_1655), .A1(net_1653) );
DFF_X1 inst_1882 ( .D(net_1321), .QN(net_90), .CK(net_3716) );
SDFF_X2 inst_104 ( .SE(net_488), .Q(net_167), .D(net_167), .CK(net_2734), .SI(x4476) );
CLKBUF_X2 inst_4060 ( .A(net_3851), .Z(net_3852) );
AOI22_X2 inst_2285 ( .A1(net_1996), .B1(net_1749), .A2(net_1548), .ZN(net_977), .B2(net_150) );
AOI22_X2 inst_2331 ( .B2(net_2162), .A1(net_2038), .A2(net_1545), .B1(net_979), .ZN(net_833) );
CLKBUF_X2 inst_3344 ( .A(net_3135), .Z(net_3136) );
CLKBUF_X2 inst_3447 ( .A(net_2798), .Z(net_3239) );
INV_X2 inst_1499 ( .A(net_2366), .ZN(net_1228) );
AOI22_X2 inst_2377 ( .B2(net_2124), .B1(net_1929), .A1(net_655), .ZN(net_653), .A2(net_304) );
AOI21_X2 inst_2522 ( .A(net_1785), .B1(net_910), .ZN(net_812), .B2(net_811) );
CLKBUF_X2 inst_2972 ( .A(net_2763), .Z(net_2764) );
NAND2_X4 inst_727 ( .A1(net_2002), .A2(net_1732), .ZN(net_1728) );
NAND2_X2 inst_882 ( .ZN(net_1173), .A1(net_1166), .A2(net_397) );
CLKBUF_X2 inst_2874 ( .A(net_2606), .Z(net_2666) );
AOI22_X2 inst_2431 ( .B2(net_2156), .B1(net_1974), .ZN(net_1805), .A1(net_1789), .A2(net_337) );
CLKBUF_X2 inst_3297 ( .A(net_2973), .Z(net_3089) );
CLKBUF_X2 inst_2938 ( .A(net_2729), .Z(net_2730) );
INV_X4 inst_1346 ( .A(net_2244), .ZN(net_2085) );
NAND3_X1 inst_708 ( .A1(net_2139), .A3(net_1927), .A2(net_1665), .ZN(net_1663) );
CLKBUF_X2 inst_3523 ( .A(net_3314), .Z(net_3315) );
INV_X2 inst_1374 ( .A(net_1010), .ZN(x2674) );
NAND2_X2 inst_953 ( .A1(net_1830), .ZN(net_984), .A2(net_399) );
AOI221_X2 inst_2510 ( .C2(net_2193), .B2(net_2116), .B1(net_1929), .A(net_1888), .C1(net_1863), .ZN(net_1764) );
CLKBUF_X2 inst_3510 ( .A(net_3301), .Z(net_3302) );
NAND2_X2 inst_1071 ( .A1(net_2090), .ZN(net_1787), .A2(net_1776) );
INV_X2 inst_1421 ( .A(net_1918), .ZN(net_536) );
CLKBUF_X2 inst_3373 ( .A(net_3164), .Z(net_3165) );
DFF_X1 inst_1994 ( .Q(net_2158), .D(net_1043), .CK(net_3103) );
CLKBUF_X2 inst_3664 ( .A(net_3455), .Z(net_3456) );
CLKBUF_X2 inst_3486 ( .A(net_2553), .Z(net_3278) );
OAI21_X2 inst_392 ( .B2(net_2001), .ZN(net_1178), .B1(net_766), .A(net_303) );
SDFF_X2 inst_120 ( .Q(net_1562), .D(net_1562), .SE(net_491), .CK(net_2655), .SI(x7120) );
OAI22_X2 inst_294 ( .B2(net_1912), .ZN(net_1837), .A1(net_1836), .B1(net_1743), .A2(net_1098) );
CLKBUF_X2 inst_4165 ( .A(net_3250), .Z(net_3957) );
INV_X2 inst_1514 ( .A(net_1578), .ZN(net_472) );
CLKBUF_X2 inst_3384 ( .A(net_3175), .Z(net_3176) );
AOI22_X2 inst_2272 ( .B1(net_1768), .ZN(net_1704), .B2(net_1516), .A1(net_1001), .A2(net_792) );
INV_X2 inst_1608 ( .ZN(net_815), .A(net_58) );
NOR2_X2 inst_567 ( .ZN(net_387), .A1(net_341), .A2(net_270) );
CLKBUF_X2 inst_3200 ( .A(net_2991), .Z(net_2992) );
NAND2_X2 inst_810 ( .A2(net_1677), .ZN(net_1303), .A1(net_1268) );
OAI22_X2 inst_230 ( .B2(net_2305), .B1(net_1865), .A1(net_1597), .ZN(net_944), .A2(net_716) );
INV_X2 inst_1601 ( .ZN(net_209), .A(x4118) );
INV_X2 inst_1484 ( .ZN(net_349), .A(net_348) );
CLKBUF_X2 inst_3035 ( .A(net_2826), .Z(net_2827) );
CLKBUF_X2 inst_3526 ( .A(net_3005), .Z(net_3318) );
NAND2_X2 inst_856 ( .A1(net_1741), .ZN(net_1231), .A2(net_1222) );
DFF_X1 inst_1893 ( .D(net_1336), .Q(net_141), .CK(net_3004) );

endmodule
