module c5315 (
n562,
n123,
n315,
n293,
n34,
n351,
n94,
n556,
n4,
n61,
n188,
n53,
n3552,
n120,
n46,
n1690,
n136,
n272,
n27,
n149,
n113,
n422,
n254,
n323,
n146,
n1,
n14,
n3546,
n128,
n80,
n4092,
n245,
n411,
n226,
n116,
n503,
n43,
n341,
n210,
n49,
n264,
n119,
n109,
n3548,
n114,
n374,
n176,
n11,
n400,
n3550,
n141,
n83,
n3173,
n545,
n361,
n103,
n4090,
n155,
n197,
n81,
n40,
n372,
n251,
n25,
n366,
n76,
n131,
n4089,
n446,
n288,
n308,
n67,
n191,
n20,
n234,
n206,
n97,
n145,
n126,
n534,
n4115,
n122,
n1497,
n2174,
n490,
n73,
n173,
n52,
n91,
n87,
n129,
n23,
n1694,
n130,
n3724,
n479,
n127,
n137,
n299,
n273,
n179,
n2358,
n118,
n457,
n161,
n307,
n88,
n54,
n4087,
n1691,
n64,
n82,
n1689,
n242,
n292,
n4091,
n140,
n112,
n167,
n435,
n302,
n514,
n369,
n17,
n135,
n332,
n164,
n281,
n132,
n117,
n289,
n324,
n549,
n265,
n37,
n185,
n203,
n152,
n331,
n170,
n348,
n523,
n100,
n552,
n115,
n217,
n4088,
n209,
n26,
n218,
n182,
n257,
n86,
n468,
n373,
n158,
n31,
n121,
n386,
n79,
n194,
n335,
n2824,
n248,
n106,
n24,
n3717,
n338,
n559,
n280,
n70,
n233,
n358,
n225,
n241,
n200,
n316,
n389,
n651,
n826,
n688,
n602,
n593,
n693,
n611,
n797,
n658,
n699,
n676,
n656,
n1002,
n615,
n594,
n863,
n632,
n591,
n599,
n939,
n802,
n673,
n889,
n871,
n712,
n690,
n849,
n732,
n865,
n722,
n685,
n737,
n815,
n824,
n604,
n854,
n834,
n807,
n923,
n877,
n813,
n601,
n702,
n873,
n667,
n828,
n850,
n777,
n704,
n600,
n1004,
n838,
n882,
n598,
n818,
n629,
n993,
n727,
n747,
n626,
n978,
n845,
n820,
n634,
n636,
n682,
n623,
n887,
n861,
n847,
n867,
n998,
n822,
n782,
n772,
n606,
n949,
n851,
n298,
n612,
n717,
n859,
n707,
n921,
n588,
n645,
n654,
n661,
n926,
n830,
n575,
n642,
n670,
n144,
n648,
n875,
n836,
n843,
n603,
n639,
n973,
n767,
n679,
n809,
n810,
n715,
n621,
n762,
n585,
n1000,
n832,
n696,
n664,
n787,
n869,
n848,
n792,
n752,
n610,
n892,
n618,
n757,
n742);

// Start PIs
input n562;
input n123;
input n315;
input n293;
input n34;
input n351;
input n94;
input n556;
input n4;
input n61;
input n188;
input n53;
input n3552;
input n120;
input n46;
input n1690;
input n136;
input n272;
input n27;
input n149;
input n113;
input n422;
input n254;
input n323;
input n146;
input n1;
input n14;
input n3546;
input n128;
input n80;
input n4092;
input n245;
input n411;
input n226;
input n116;
input n503;
input n43;
input n341;
input n210;
input n49;
input n264;
input n119;
input n109;
input n3548;
input n114;
input n374;
input n176;
input n11;
input n400;
input n3550;
input n141;
input n83;
input n3173;
input n545;
input n361;
input n103;
input n4090;
input n155;
input n197;
input n81;
input n40;
input n372;
input n251;
input n25;
input n366;
input n76;
input n131;
input n4089;
input n446;
input n288;
input n308;
input n67;
input n191;
input n20;
input n234;
input n206;
input n97;
input n145;
input n126;
input n534;
input n4115;
input n122;
input n1497;
input n2174;
input n490;
input n73;
input n173;
input n52;
input n91;
input n87;
input n129;
input n23;
input n1694;
input n130;
input n3724;
input n479;
input n127;
input n137;
input n299;
input n273;
input n179;
input n2358;
input n118;
input n457;
input n161;
input n307;
input n88;
input n54;
input n4087;
input n1691;
input n64;
input n82;
input n1689;
input n242;
input n292;
input n4091;
input n140;
input n112;
input n167;
input n435;
input n302;
input n514;
input n369;
input n17;
input n135;
input n332;
input n164;
input n281;
input n132;
input n117;
input n289;
input n324;
input n549;
input n265;
input n37;
input n185;
input n203;
input n152;
input n331;
input n170;
input n348;
input n523;
input n100;
input n552;
input n115;
input n217;
input n4088;
input n209;
input n26;
input n218;
input n182;
input n257;
input n86;
input n468;
input n373;
input n158;
input n31;
input n121;
input n386;
input n79;
input n194;
input n335;
input n2824;
input n248;
input n106;
input n24;
input n3717;
input n338;
input n559;
input n280;
input n70;
input n233;
input n358;
input n225;
input n241;
input n200;
input n316;
input n389;

// Start POs
output n651;
output n826;
output n688;
output n602;
output n593;
output n693;
output n611;
output n797;
output n658;
output n699;
output n676;
output n656;
output n1002;
output n615;
output n594;
output n863;
output n632;
output n591;
output n599;
output n939;
output n802;
output n673;
output n889;
output n871;
output n712;
output n690;
output n849;
output n732;
output n865;
output n722;
output n685;
output n737;
output n815;
output n824;
output n604;
output n854;
output n834;
output n807;
output n923;
output n877;
output n813;
output n601;
output n702;
output n873;
output n667;
output n828;
output n850;
output n777;
output n704;
output n600;
output n1004;
output n838;
output n882;
output n598;
output n818;
output n629;
output n993;
output n727;
output n747;
output n626;
output n978;
output n845;
output n820;
output n634;
output n636;
output n682;
output n623;
output n887;
output n861;
output n847;
output n867;
output n998;
output n822;
output n782;
output n772;
output n606;
output n949;
output n851;
output n298;
output n612;
output n717;
output n859;
output n707;
output n921;
output n588;
output n645;
output n654;
output n661;
output n926;
output n830;
output n575;
output n642;
output n670;
output n144;
output n648;
output n875;
output n836;
output n843;
output n603;
output n639;
output n973;
output n767;
output n679;
output n809;
output n810;
output n715;
output n621;
output n762;
output n585;
output n1000;
output n832;
output n696;
output n664;
output n787;
output n869;
output n848;
output n792;
output n752;
output n610;
output n892;
output n618;
output n757;
output n742;

// Start wires
wire net_416;
wire net_215;
wire net_54;
wire net_526;
wire net_429;
wire net_694;
wire net_129;
wire net_648;
wire net_373;
wire net_98;
wire net_739;
wire net_151;
wire net_356;
wire net_53;
wire net_452;
wire net_545;
wire net_284;
wire net_560;
wire net_774;
wire net_439;
wire net_259;
wire net_548;
wire n146;
wire net_501;
wire net_187;
wire net_111;
wire net_264;
wire net_225;
wire n116;
wire net_636;
wire net_263;
wire net_252;
wire net_124;
wire net_343;
wire n119;
wire net_160;
wire n141;
wire net_322;
wire net_511;
wire net_420;
wire net_665;
wire net_447;
wire n4090;
wire net_410;
wire net_508;
wire net_390;
wire net_35;
wire net_586;
wire net_703;
wire net_239;
wire net_193;
wire net_310;
wire net_120;
wire n308;
wire net_292;
wire net_201;
wire net_109;
wire net_80;
wire n234;
wire n206;
wire net_96;
wire net_167;
wire net_651;
wire net_682;
wire net_280;
wire net_744;
wire net_495;
wire net_34;
wire net_458;
wire net_108;
wire net_598;
wire net_685;
wire n87;
wire n129;
wire n130;
wire net_789;
wire n618;
wire net_593;
wire net_617;
wire net_672;
wire net_777;
wire net_554;
wire n658;
wire net_490;
wire net_742;
wire net_46;
wire net_584;
wire n939;
wire net_632;
wire net_538;
wire net_165;
wire net_464;
wire n604;
wire net_366;
wire net_13;
wire net_747;
wire net_446;
wire n549;
wire n850;
wire n170;
wire net_248;
wire net_384;
wire net_198;
wire n26;
wire n845;
wire net_209;
wire net_3;
wire net_634;
wire net_294;
wire net_371;
wire n859;
wire n31;
wire n588;
wire n575;
wire net_485;
wire n194;
wire n335;
wire net_503;
wire net_256;
wire n3717;
wire net_82;
wire n621;
wire n280;
wire net_64;
wire net_726;
wire net_679;
wire n241;
wire n664;
wire net_308;
wire net_75;
wire net_515;
wire net_600;
wire net_757;
wire net_701;
wire net_206;
wire net_125;
wire net_397;
wire n757;
wire n562;
wire net_223;
wire net_715;
wire net_235;
wire n123;
wire n293;
wire n315;
wire net_606;
wire net_623;
wire n188;
wire net_663;
wire net_320;
wire net_579;
wire n863;
wire net_250;
wire net_769;
wire net_312;
wire net_130;
wire net_572;
wire net_286;
wire net_147;
wire net_787;
wire net_481;
wire net_369;
wire net_403;
wire net_32;
wire n80;
wire net_282;
wire net_645;
wire net_426;
wire n3548;
wire net_780;
wire net_609;
wire net_541;
wire net_414;
wire n83;
wire net_794;
wire net_528;
wire n197;
wire net_456;
wire net_155;
wire net_705;
wire net_335;
wire net_506;
wire net_181;
wire n76;
wire n4089;
wire n782;
wire net_349;
wire net_39;
wire net_245;
wire n446;
wire net_395;
wire net_331;
wire net_493;
wire net_386;
wire net_641;
wire net_277;
wire net_89;
wire net_290;
wire n832;
wire n52;
wire net_680;
wire n23;
wire net_338;
wire n137;
wire net_721;
wire net_243;
wire net_400;
wire n179;
wire n2358;
wire net_759;
wire n602;
wire net_602;
wire n693;
wire net_175;
wire net_657;
wire net_106;
wire net_140;
wire net_740;
wire net_247;
wire net_329;
wire net_279;
wire net_698;
wire net_25;
wire net_70;
wire net_691;
wire n112;
wire net_194;
wire net_730;
wire net_615;
wire n369;
wire net_478;
wire n685;
wire net_441;
wire n815;
wire net_596;
wire net_138;
wire net_749;
wire net_333;
wire net_639;
wire net_728;
wire n289;
wire n324;
wire net_719;
wire n667;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_77;
wire net_20;
wire net_49;
wire net_518;
wire net_15;
wire net_57;
wire net_71;
wire net_771;
wire net_1;
wire net_708;
wire net_696;
wire n707;
wire net_537;
wire net_180;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire n648;
wire net_432;
wire n875;
wire net_513;
wire net_204;
wire n248;
wire net_232;
wire n338;
wire net_604;
wire net_163;
wire net_67;
wire net_268;
wire net_459;
wire net_483;
wire net_48;
wire net_8;
wire net_737;
wire net_203;
wire net_505;
wire net_176;
wire net_296;
wire net_137;
wire net_613;
wire net_237;
wire n94;
wire net_782;
wire n53;
wire n656;
wire n3552;
wire net_614;
wire net_532;
wire net_93;
wire net_578;
wire n673;
wire n272;
wire net_786;
wire net_302;
wire n871;
wire n254;
wire net_127;
wire net_348;
wire net_753;
wire n1;
wire n3546;
wire net_626;
wire net_101;
wire net_388;
wire net_326;
wire net_707;
wire net_589;
wire net_100;
wire net_655;
wire net_686;
wire net_652;
wire net_536;
wire net_455;
wire n374;
wire net_221;
wire net_115;
wire net_689;
wire net_751;
wire net_393;
wire n3173;
wire net_442;
wire net_542;
wire net_575;
wire net_595;
wire net_378;
wire net_408;
wire net_724;
wire net_423;
wire net_328;
wire n131;
wire n717;
wire net_157;
wire net_42;
wire n926;
wire n67;
wire n191;
wire net_66;
wire net_466;
wire net_765;
wire net_675;
wire n122;
wire n973;
wire net_443;
wire n1000;
wire net_522;
wire net_270;
wire net_183;
wire net_668;
wire n479;
wire net_150;
wire net_304;
wire net_352;
wire net_644;
wire n307;
wire net_30;
wire net_643;
wire net_436;
wire net_24;
wire net_622;
wire net_186;
wire n167;
wire n690;
wire net_792;
wire n732;
wire net_767;
wire net_219;
wire net_18;
wire net_309;
wire net_659;
wire net_131;
wire net_196;
wire net_29;
wire net_358;
wire n203;
wire n152;
wire n600;
wire net_516;
wire net_31;
wire n115;
wire n4088;
wire net_713;
wire n623;
wire net_693;
wire net_360;
wire n887;
wire net_213;
wire net_729;
wire n921;
wire net_260;
wire net_438;
wire net_732;
wire net_580;
wire net_314;
wire n2824;
wire net_341;
wire n679;
wire net_468;
wire net_58;
wire net_488;
wire net_73;
wire net_86;
wire n869;
wire n651;
wire net_179;
wire net_159;
wire net_61;
wire n34;
wire net_449;
wire net_383;
wire net_62;
wire net_6;
wire n120;
wire net_553;
wire net_534;
wire net_217;
wire net_733;
wire n46;
wire net_763;
wire net_427;
wire net_486;
wire net_135;
wire net_473;
wire net_406;
wire n422;
wire n737;
wire net_633;
wire net_324;
wire net_113;
wire net_710;
wire net_497;
wire n4092;
wire net_454;
wire net_462;
wire net_418;
wire net_40;
wire n411;
wire n264;
wire net_709;
wire n109;
wire n873;
wire net_161;
wire net_300;
wire net_748;
wire net_677;
wire net_95;
wire n103;
wire net_173;
wire net_78;
wire n372;
wire net_514;
wire n636;
wire net_376;
wire net_22;
wire net_354;
wire net_524;
wire n661;
wire n654;
wire net_646;
wire net_363;
wire n830;
wire net_445;
wire net_573;
wire net_776;
wire n126;
wire net_44;
wire net_784;
wire net_520;
wire net_422;
wire net_561;
wire n810;
wire n715;
wire net_567;
wire net_45;
wire net_381;
wire net_591;
wire net_746;
wire net_272;
wire n848;
wire net_178;
wire n127;
wire net_762;
wire net_695;
wire n611;
wire n797;
wire n88;
wire net_556;
wire n699;
wire net_629;
wire n1691;
wire net_55;
wire net_559;
wire net_635;
wire net_255;
wire net_266;
wire n594;
wire net_345;
wire n1689;
wire net_620;
wire net_619;
wire net_350;
wire net_398;
wire net_306;
wire n435;
wire net_500;
wire n17;
wire n164;
wire n117;
wire net_631;
wire net_11;
wire net_123;
wire n828;
wire net_527;
wire net_362;
wire net_262;
wire net_318;
wire net_68;
wire n682;
wire net_316;
wire net_84;
wire net_670;
wire net_611;
wire net_231;
wire net_103;
wire net_226;
wire net_228;
wire n670;
wire net_143;
wire net_190;
wire net_391;
wire net_533;
wire net_145;
wire net_37;
wire n233;
wire net_582;
wire net_188;
wire net_755;
wire net_509;
wire net_661;
wire net_211;
wire net_133;
wire net_568;
wire net_47;
wire n556;
wire n61;
wire n676;
wire net_557;
wire net_119;
wire net_210;
wire net_168;
wire n136;
wire n27;
wire net_741;
wire net_477;
wire n849;
wire net_385;
wire n865;
wire net_269;
wire net_469;
wire n14;
wire net_727;
wire net_90;
wire net_671;
wire n43;
wire n503;
wire net_283;
wire n702;
wire net_85;
wire net_778;
wire net_770;
wire n176;
wire net_404;
wire net_240;
wire n838;
wire net_4;
wire n882;
wire net_295;
wire n81;
wire n626;
wire net_307;
wire n251;
wire net_344;
wire n366;
wire net_16;
wire net_712;
wire n612;
wire net_257;
wire net_233;
wire net_474;
wire net_472;
wire net_65;
wire net_484;
wire net_136;
wire net_207;
wire net_700;
wire net_126;
wire n173;
wire n73;
wire n585;
wire net_278;
wire n1694;
wire n752;
wire net_571;
wire net_63;
wire net_274;
wire net_601;
wire n118;
wire n826;
wire net_321;
wire net_425;
wire n457;
wire net_287;
wire net_189;
wire net_720;
wire net_99;
wire n64;
wire net_480;
wire net_216;
wire net_433;
wire n632;
wire net_544;
wire net_717;
wire net_368;
wire net_224;
wire net_684;
wire net_52;
wire net_608;
wire n332;
wire net_370;
wire net_510;
wire n807;
wire net_413;
wire net_716;
wire net_114;
wire n777;
wire n331;
wire net_36;
wire n727;
wire net_253;
wire net_637;
wire net_276;
wire net_311;
wire net_760;
wire n978;
wire net_494;
wire n634;
wire net_547;
wire net_154;
wire n257;
wire net_666;
wire n86;
wire net_507;
wire net_616;
wire n158;
wire n645;
wire net_238;
wire net_28;
wire net_529;
wire net_704;
wire n79;
wire net_587;
wire net_97;
wire net_192;
wire net_793;
wire n843;
wire net_649;
wire n767;
wire net_460;
wire net_650;
wire net_291;
wire net_457;
wire net_735;
wire net_772;
wire net_121;
wire net_200;
wire net_597;
wire n787;
wire net_743;
wire n200;
wire net_396;
wire n316;
wire net_195;
wire net_107;
wire net_166;
wire net_530;
wire n351;
wire n4;
wire n1002;
wire net_594;
wire net_603;
wire net_23;
wire net_271;
wire net_117;
wire net_74;
wire net_673;
wire net_401;
wire net_642;
wire net_205;
wire net_699;
wire net_242;
wire net_359;
wire net_440;
wire n722;
wire n323;
wire net_758;
wire net_26;
wire net_470;
wire net_334;
wire n923;
wire net_430;
wire n813;
wire net_365;
wire net_718;
wire net_380;
wire n11;
wire net_141;
wire n3550;
wire net_467;
wire net_83;
wire net_372;
wire n993;
wire net_437;
wire net_56;
wire net_566;
wire net_336;
wire net_624;
wire net_555;
wire net_2;
wire net_9;
wire n642;
wire net_298;
wire net_790;
wire net_688;
wire net_697;
wire net_475;
wire n145;
wire net_563;
wire n603;
wire net_605;
wire net_199;
wire net_502;
wire net_431;
wire n91;
wire n3724;
wire net_638;
wire net_222;
wire net_152;
wire net_313;
wire net_489;
wire net_714;
wire net_683;
wire net_258;
wire net_607;
wire net_148;
wire n242;
wire net_419;
wire n802;
wire n140;
wire net_251;
wire n302;
wire n514;
wire net_244;
wire net_664;
wire net_128;
wire net_585;
wire n824;
wire net_549;
wire net_785;
wire net_374;
wire n265;
wire n37;
wire net_411;
wire net_788;
wire net_214;
wire n1004;
wire net_249;
wire n100;
wire n552;
wire net_706;
wire n209;
wire net_156;
wire net_92;
wire net_112;
wire net_394;
wire net_139;
wire n851;
wire net_551;
wire net_332;
wire net_409;
wire net_463;
wire net_492;
wire net_656;
wire net_88;
wire net_197;
wire n639;
wire net_766;
wire n106;
wire n24;
wire net_81;
wire n809;
wire net_402;
wire net_202;
wire n225;
wire net_110;
wire net_379;
wire net_722;
wire net_33;
wire n892;
wire n389;
wire net_289;
wire net_450;
wire net_621;
wire net_435;
wire net_132;
wire net_105;
wire n615;
wire net_12;
wire n591;
wire n113;
wire net_569;
wire net_768;
wire net_327;
wire net_357;
wire net_630;
wire net_76;
wire n128;
wire net_353;
wire n601;
wire net_519;
wire net_412;
wire n400;
wire net_17;
wire n598;
wire n545;
wire net_319;
wire n361;
wire net_453;
wire net_581;
wire net_164;
wire n155;
wire net_731;
wire net_377;
wire net_87;
wire net_0;
wire net_288;
wire n820;
wire n25;
wire net_658;
wire net_734;
wire net_540;
wire net_512;
wire net_779;
wire net_662;
wire net_50;
wire n97;
wire net_234;
wire net_38;
wire net_342;
wire net_612;
wire net_19;
wire n490;
wire net_738;
wire net_504;
wire n696;
wire net_674;
wire net_618;
wire net_303;
wire n742;
wire n273;
wire n161;
wire net_491;
wire net_681;
wire net_783;
wire n4087;
wire net_392;
wire net_118;
wire n82;
wire net_754;
wire net_421;
wire net_146;
wire net_764;
wire net_550;
wire net_122;
wire net_417;
wire net_7;
wire net_172;
wire n834;
wire n281;
wire net_428;
wire net_94;
wire net_246;
wire net_461;
wire n877;
wire n132;
wire net_640;
wire net_482;
wire net_775;
wire net_149;
wire net_142;
wire net_752;
wire n348;
wire n523;
wire net_387;
wire net_654;
wire net_330;
wire net_498;
wire net_535;
wire net_158;
wire n818;
wire n629;
wire net_676;
wire net_41;
wire n747;
wire net_577;
wire n861;
wire net_570;
wire n182;
wire net_444;
wire net_525;
wire n822;
wire n772;
wire n468;
wire net_325;
wire net_301;
wire n121;
wire net_299;
wire n144;
wire net_182;
wire net_60;
wire net_521;
wire net_337;
wire net_590;
wire net_267;
wire net_273;
wire net_424;
wire net_576;
wire net_690;
wire net_465;
wire net_177;
wire n792;
wire net_523;
wire net_407;
wire net_476;
wire net_564;
wire net_382;
wire n593;
wire n688;
wire net_725;
wire net_583;
wire net_351;
wire n1690;
wire n599;
wire net_340;
wire net_265;
wire net_517;
wire n149;
wire net_434;
wire net_628;
wire net_791;
wire n889;
wire n712;
wire net_14;
wire net_220;
wire net_293;
wire n854;
wire n245;
wire n226;
wire n210;
wire n341;
wire n49;
wire net_69;
wire net_543;
wire n114;
wire net_625;
wire n704;
wire net_339;
wire net_361;
wire net_27;
wire net_317;
wire net_305;
wire n40;
wire net_191;
wire net_261;
wire net_558;
wire n867;
wire n606;
wire net_660;
wire net_144;
wire net_102;
wire net_227;
wire net_59;
wire n288;
wire net_162;
wire n20;
wire net_781;
wire net_230;
wire net_653;
wire n4115;
wire n534;
wire net_134;
wire n1497;
wire net_678;
wire net_546;
wire n2174;
wire n762;
wire net_185;
wire net_702;
wire net_588;
wire n610;
wire net_667;
wire net_208;
wire net_236;
wire net_212;
wire net_315;
wire net_487;
wire n299;
wire net_552;
wire net_415;
wire net_116;
wire n54;
wire net_347;
wire net_756;
wire net_91;
wire net_297;
wire net_346;
wire net_104;
wire net_448;
wire net_72;
wire n292;
wire net_229;
wire n4091;
wire net_627;
wire net_241;
wire net_687;
wire net_5;
wire net_405;
wire n135;
wire net_355;
wire net_184;
wire net_599;
wire net_711;
wire net_610;
wire net_723;
wire n185;
wire net_389;
wire net_451;
wire net_323;
wire net_750;
wire net_736;
wire net_275;
wire net_399;
wire net_539;
wire n217;
wire net_692;
wire net_153;
wire n847;
wire net_218;
wire net_174;
wire n218;
wire n998;
wire net_375;
wire net_562;
wire n949;
wire n298;
wire net_364;
wire net_43;
wire n373;
wire net_10;
wire n386;
wire net_592;
wire net_21;
wire net_79;
wire net_647;
wire n836;
wire net_773;
wire net_285;
wire net_281;
wire net_669;
wire n559;
wire net_254;
wire n70;
wire n358;
wire net_761;
wire net_496;
wire net_479;
wire net_574;
wire net_745;

// Start cells
NAND2_X1 inst_537 ( .ZN(net_455), .A2(net_441), .A1(net_392) );
MUX2_X2 inst_696 ( .A(net_634), .B(net_41), .Z(n863), .S(n4092) );
INV_X1 inst_826 ( .ZN(net_405), .A(net_404) );
NAND2_X1 inst_481 ( .ZN(net_195), .A2(net_194), .A1(n91) );
NAND2_X1 inst_551 ( .A2(net_460), .ZN(net_442), .A1(net_441) );
NOR2_X1 inst_228 ( .ZN(net_31), .A2(n3548), .A1(n218) );
XNOR2_X1 inst_125 ( .ZN(net_711), .B(net_645), .A(net_551) );
NAND2_X1 inst_486 ( .A2(net_203), .ZN(net_201), .A1(n64) );
NAND2_X1 inst_506 ( .ZN(net_421), .A2(net_286), .A1(n534) );
NAND2_X1 inst_495 ( .A2(net_217), .ZN(net_212), .A1(n185) );
NAND3_X1 inst_353 ( .ZN(net_92), .A1(n1694), .A3(n1691), .A2(n161) );
NOR3_X1 inst_207 ( .A2(net_482), .A1(net_437), .A3(net_418), .ZN(n598) );
AND3_X4 inst_872 ( .ZN(net_666), .A2(net_665), .A3(net_661), .A1(n2174) );
OR2_X2 inst_159 ( .A1(net_519), .ZN(net_429), .A2(net_428) );
MUX2_X2 inst_707 ( .A(net_644), .B(net_67), .Z(n826), .S(n4092) );
INV_X1 inst_779 ( .ZN(n604), .A(n545) );
NAND3_X1 inst_395 ( .A3(net_677), .A2(net_200), .A1(net_120), .ZN(n797) );
INV_X1 inst_841 ( .A(net_716), .ZN(n867) );
XNOR2_X1 inst_134 ( .ZN(net_762), .B(net_744), .A(net_656) );
NOR2_X1 inst_244 ( .ZN(net_54), .A1(net_53), .A2(n3546) );
NOR2_X1 inst_333 ( .ZN(net_520), .A1(net_519), .A2(net_473) );
MUX2_X2 inst_712 ( .Z(net_696), .B(net_694), .A(net_693), .S(net_541) );
NAND2_X1 inst_452 ( .ZN(net_398), .A1(net_164), .A2(n809) );
MUX2_X2 inst_689 ( .A(net_649), .B(net_648), .Z(net_646), .S(n4089) );
NAND2_X1 inst_430 ( .ZN(net_32), .A2(n257), .A1(n242) );
XNOR2_X1 inst_131 ( .ZN(net_744), .A(net_688), .B(net_536) );
NAND3_X1 inst_406 ( .A3(net_724), .A2(net_195), .A1(net_123), .ZN(n742) );
NOR2_X1 inst_214 ( .ZN(net_9), .A2(n251), .A1(n218) );
NAND2_X1 inst_462 ( .A2(net_178), .ZN(net_172), .A1(n182) );
OR2_X2 inst_160 ( .A1(net_756), .ZN(net_496), .A2(net_495) );
AND4_X1 inst_869 ( .A4(net_601), .ZN(n854), .A3(n562), .A2(n556), .A1(n552) );
NOR2_X1 inst_328 ( .A1(net_526), .A2(net_501), .ZN(n626) );
XNOR2_X1 inst_47 ( .ZN(net_296), .A(net_295), .B(net_290) );
XOR2_X1 inst_19 ( .Z(net_656), .B(net_295), .A(n514) );
NAND2_X1 inst_548 ( .ZN(net_490), .A1(net_421), .A2(net_362) );
NAND2_X1 inst_515 ( .ZN(net_269), .A1(net_225), .A2(net_103) );
XOR2_X1 inst_8 ( .Z(net_284), .A(net_283), .B(net_282) );
INV_X1 inst_772 ( .ZN(n848), .A(n245) );
INV_X1 inst_818 ( .A(net_630), .ZN(net_331) );
MUX2_X2 inst_728 ( .Z(net_719), .A(net_717), .B(net_716), .S(n1691) );
INV_X1 inst_762 ( .ZN(net_2), .A(n446) );
NAND3_X1 inst_370 ( .ZN(net_161), .A3(net_160), .A1(n4092), .A2(n120) );
NAND2_X1 inst_573 ( .A1(net_738), .ZN(net_685), .A2(net_669) );
XNOR2_X1 inst_100 ( .ZN(net_770), .B(net_538), .A(net_499) );
MUX2_X2 inst_642 ( .Z(net_152), .B(n3552), .A(n3550), .S(n257) );
NAND2_X1 inst_459 ( .A2(net_181), .ZN(net_169), .A1(n197) );
NOR2_X1 inst_279 ( .ZN(net_268), .A1(net_227), .A2(net_111) );
NAND2_X1 inst_445 ( .ZN(net_86), .A2(net_38), .A1(n254) );
CLKBUF_X1 inst_850 ( .Z(n978), .A(n1) );
MUX2_X2 inst_709 ( .Z(net_689), .A(net_673), .B(net_132), .S(n1694) );
XNOR2_X1 inst_93 ( .A(net_602), .ZN(net_552), .B(net_551) );
MUX2_X2 inst_700 ( .Z(net_674), .A(net_672), .B(net_671), .S(n1689) );
XNOR2_X1 inst_81 ( .ZN(net_529), .B(net_524), .A(net_454) );
MUX2_X2 inst_612 ( .Z(net_107), .B(n3552), .A(n3550), .S(n218) );
MUX2_X2 inst_606 ( .Z(net_97), .A(n254), .B(n242), .S(n234) );
NAND3_X1 inst_367 ( .ZN(net_153), .A1(n1694), .A3(n1691), .A2(n164) );
NAND2_X1 inst_525 ( .ZN(net_319), .A2(net_318), .A1(n25) );
CLKBUF_X1 inst_853 ( .Z(n939), .A(n1) );
AND2_X2 inst_901 ( .A2(net_676), .ZN(n664), .A1(n137) );
OR3_X4 inst_139 ( .A1(net_729), .A2(net_630), .ZN(net_453), .A3(net_452) );
MUX2_X2 inst_657 ( .Z(net_559), .B(n861), .A(n822), .S(n1691) );
NAND2_X1 inst_559 ( .A2(net_524), .ZN(net_515), .A1(net_442) );
NAND2_X1 inst_584 ( .ZN(net_781), .A2(net_779), .A1(net_774) );
NAND2_X1 inst_521 ( .ZN(net_313), .A2(net_312), .A1(n24) );
INV_X1 inst_790 ( .ZN(net_136), .A(n4088) );
NAND2_X1 inst_434 ( .ZN(net_58), .A2(net_57), .A1(n3550) );
NAND2_X1 inst_470 ( .ZN(net_182), .A2(net_181), .A1(n203) );
AND2_X2 inst_906 ( .A2(net_689), .ZN(n702), .A1(n137) );
INV_X1 inst_751 ( .ZN(n849), .A(n552) );
INV_X1 inst_845 ( .A(net_700), .ZN(n832) );
NAND2_X1 inst_535 ( .ZN(net_372), .A2(net_363), .A1(net_359) );
NAND2_X1 inst_450 ( .A2(net_160), .ZN(net_150), .A1(n129) );
MUX2_X2 inst_745 ( .Z(net_785), .A(net_780), .B(n97), .S(n4092) );
NAND2_X1 inst_520 ( .A2(net_312), .ZN(net_311), .A1(n79) );
NOR2_X1 inst_237 ( .A1(net_774), .ZN(net_184), .A2(n4091) );
OR2_X4 inst_148 ( .A2(net_519), .ZN(net_378), .A1(net_377) );
NAND2_X1 inst_554 ( .A1(net_454), .ZN(net_448), .A2(net_447) );
MUX2_X2 inst_733 ( .Z(net_737), .A(net_735), .B(net_734), .S(n4089) );
NAND3_X1 inst_377 ( .ZN(net_303), .A3(net_58), .A1(net_12), .A2(n422) );
NOR3_X1 inst_191 ( .ZN(net_236), .A2(net_235), .A1(net_145), .A3(net_33) );
INV_X1 inst_813 ( .ZN(net_729), .A(net_441) );
XNOR2_X1 inst_51 ( .ZN(net_322), .A(net_321), .B(net_128) );
OR3_X2 inst_142 ( .A1(net_76), .A3(net_14), .A2(n809), .ZN(n636) );
NOR2_X1 inst_315 ( .A2(net_679), .A1(net_630), .ZN(net_460) );
XNOR2_X1 inst_80 ( .ZN(net_569), .A(net_519), .B(net_471) );
INV_X1 inst_836 ( .A(net_649), .ZN(n836) );
NOR2_X1 inst_216 ( .ZN(net_14), .A2(n86), .A1(n2358) );
XNOR2_X1 inst_78 ( .ZN(net_507), .A(net_433), .B(net_347) );
NOR2_X1 inst_241 ( .ZN(net_49), .A1(net_48), .A2(n3546) );
OR2_X2 inst_177 ( .ZN(net_728), .A2(net_704), .A1(n1694) );
AND2_X4 inst_885 ( .A1(net_364), .ZN(net_350), .A2(net_349) );
INV_X1 inst_783 ( .ZN(net_6), .A(n242) );
CLKBUF_X1 inst_862 ( .A(n604), .Z(n603) );
NOR4_X1 inst_183 ( .ZN(net_747), .A2(net_713), .A4(net_712), .A1(net_666), .A3(net_664) );
CLKBUF_X1 inst_852 ( .Z(n949), .A(n1) );
OR2_X4 inst_151 ( .ZN(net_495), .A1(net_447), .A2(net_426) );
XNOR2_X1 inst_64 ( .ZN(net_531), .B(net_412), .A(net_253) );
MUX2_X2 inst_743 ( .Z(net_779), .A(net_777), .B(net_776), .S(n4091) );
NAND3_X1 inst_415 ( .A2(net_782), .A3(net_775), .A1(net_161), .ZN(n843) );
MUX2_X2 inst_615 ( .Z(net_110), .B(n3552), .A(n3550), .S(n234) );
NAND3_X1 inst_393 ( .A3(net_653), .A2(net_210), .A1(net_191), .ZN(n762) );
XNOR2_X1 inst_107 ( .ZN(net_600), .B(net_573), .A(net_572) );
INV_X1 inst_828 ( .ZN(net_462), .A(net_461) );
AND2_X4 inst_892 ( .ZN(net_665), .A2(net_662), .A1(net_501) );
XNOR2_X1 inst_92 ( .A(net_656), .ZN(net_586), .B(net_518) );
NAND4_X1 inst_345 ( .ZN(net_437), .A1(net_436), .A2(net_435), .A3(net_434), .A4(net_352) );
NOR2_X1 inst_223 ( .ZN(net_25), .A2(n351), .A1(n251) );
NAND3_X1 inst_402 ( .A3(net_721), .A2(net_198), .A1(net_112), .ZN(n782) );
INV_X1 inst_819 ( .A(net_575), .ZN(net_332) );
NAND4_X1 inst_340 ( .A2(net_399), .A3(net_398), .ZN(net_396), .A4(net_317), .A1(net_314) );
MUX2_X2 inst_643 ( .Z(net_417), .S(n302), .A(n251), .B(n248) );
MUX2_X2 inst_697 ( .A(net_672), .B(net_671), .Z(net_669), .S(n4089) );
NAND2_X1 inst_494 ( .A2(net_217), .ZN(net_211), .A1(n170) );
NAND2_X1 inst_487 ( .A2(net_203), .ZN(net_202), .A1(n61) );
NOR2_X1 inst_329 ( .A1(net_503), .A2(net_502), .ZN(n588) );
NAND2_X1 inst_574 ( .A1(net_740), .ZN(net_686), .A2(net_670) );
NAND3_X1 inst_386 ( .A3(net_592), .A2(net_202), .A1(net_156), .ZN(n859) );
OR2_X2 inst_158 ( .ZN(net_263), .A2(net_90), .A1(n479) );
OR3_X4 inst_141 ( .ZN(net_517), .A1(net_466), .A3(net_465), .A2(net_310) );
NOR3_X1 inst_200 ( .ZN(net_247), .A1(net_54), .A3(net_27), .A2(n435) );
NAND2_X1 inst_507 ( .A2(net_289), .ZN(net_257), .A1(n435) );
NAND2_X1 inst_571 ( .A1(net_740), .ZN(net_678), .A2(net_647) );
XNOR2_X1 inst_57 ( .ZN(net_384), .B(net_299), .A(net_83) );
NOR2_X1 inst_338 ( .ZN(net_662), .A2(net_528), .A1(net_422) );
AND2_X4 inst_884 ( .ZN(net_379), .A1(net_343), .A2(net_342) );
MUX2_X2 inst_711 ( .Z(net_695), .A(net_694), .B(net_693), .S(net_540) );
INV_X1 inst_827 ( .ZN(net_419), .A(net_391) );
NAND2_X1 inst_552 ( .ZN(net_444), .A2(net_443), .A1(net_376) );
MUX2_X2 inst_599 ( .Z(net_89), .S(n351), .A(n254), .B(n242) );
NAND3_X1 inst_417 ( .A3(net_790), .A2(net_201), .A1(net_157), .ZN(n807) );
MUX2_X2 inst_671 ( .Z(net_648), .A(net_580), .B(net_140), .S(n4092) );
NAND2_X1 inst_579 ( .A1(net_748), .ZN(net_745), .A2(net_715) );
XOR2_X1 inst_21 ( .Z(net_324), .B(net_287), .A(net_285) );
NAND2_X1 inst_469 ( .ZN(net_180), .A2(net_178), .A1(n200) );
NOR2_X1 inst_281 ( .ZN(net_272), .A1(net_271), .A2(net_152) );
NAND2_X1 inst_585 ( .ZN(net_789), .A2(net_787), .A1(net_750) );
MUX2_X2 inst_698 ( .A(net_672), .B(net_671), .Z(net_670), .S(n4088) );
XOR2_X1 inst_18 ( .A(net_602), .Z(net_390), .B(n132) );
AND2_X2 inst_915 ( .A2(net_758), .ZN(n642), .A1(n137) );
AND2_X2 inst_893 ( .ZN(n634), .A1(n373), .A2(n1) );
INV_X1 inst_811 ( .ZN(net_756), .A(net_394) );
NAND2_X1 inst_541 ( .ZN(net_375), .A1(net_364), .A2(net_363) );
NAND3_X1 inst_410 ( .ZN(net_760), .A1(net_745), .A3(net_169), .A2(net_121) );
NOR3_X1 inst_208 ( .ZN(net_562), .A1(net_514), .A3(net_406), .A2(net_360) );
XNOR2_X1 inst_88 ( .ZN(net_537), .B(net_536), .A(net_497) );
NOR2_X1 inst_316 ( .ZN(net_424), .A2(net_423), .A1(net_402) );
NOR2_X1 inst_220 ( .ZN(net_20), .A2(n3548), .A1(n351) );
CLKBUF_X1 inst_851 ( .Z(n973), .A(n3173) );
XOR2_X1 inst_9 ( .Z(net_358), .B(net_283), .A(n411) );
XNOR2_X1 inst_113 ( .ZN(net_614), .A(net_585), .B(net_564) );
INV_X1 inst_831 ( .ZN(net_527), .A(net_513) );
NAND2_X1 inst_505 ( .ZN(net_454), .A2(net_282), .A1(n374) );
NAND3_X1 inst_356 ( .ZN(net_114), .A1(n1694), .A3(n1691), .A2(n167) );
NAND3_X1 inst_383 ( .ZN(net_501), .A3(net_468), .A1(net_404), .A2(net_363) );
NAND3_X1 inst_360 ( .ZN(net_119), .A1(n1690), .A3(n1689), .A2(n161) );
INV_X1 inst_773 ( .ZN(net_280), .A(n523) );
NOR3_X1 inst_198 ( .ZN(net_245), .A1(net_146), .A3(net_26), .A2(n457) );
XNOR2_X1 inst_50 ( .ZN(net_299), .A(net_147), .B(net_85) );
NOR2_X1 inst_245 ( .ZN(net_56), .A1(net_55), .A2(n3546) );
AND2_X2 inst_897 ( .A2(net_400), .ZN(n639), .A1(n141) );
NAND2_X1 inst_569 ( .ZN(net_716), .A2(net_635), .A1(net_186) );
MUX2_X2 inst_678 ( .Z(net_618), .B(n877), .A(n838), .S(n4088) );
MUX2_X2 inst_624 ( .Z(net_321), .S(n335), .B(n209), .A(n206) );
NOR2_X1 inst_260 ( .ZN(net_141), .A1(net_50), .A2(n3546) );
CLKBUF_X1 inst_854 ( .Z(n926), .A(n137) );
INV_X1 inst_784 ( .ZN(net_7), .A(n3552) );
MUX2_X2 inst_721 ( .Z(net_707), .B(n865), .A(n826), .S(n4088) );
AND2_X2 inst_902 ( .A2(net_675), .ZN(n696), .A1(n137) );
INV_X1 inst_837 ( .ZN(net_621), .A(net_611) );
OR2_X4 inst_147 ( .A2(net_679), .A1(net_454), .ZN(net_374) );
MUX2_X2 inst_744 ( .Z(net_786), .A(net_773), .B(n94), .S(n4092) );
NOR2_X1 inst_313 ( .A2(net_729), .ZN(net_463), .A1(net_446) );
NOR2_X1 inst_293 ( .ZN(net_380), .A1(net_272), .A2(net_242) );
INV_X1 inst_778 ( .ZN(net_278), .A(n422) );
MUX2_X2 inst_636 ( .Z(net_293), .S(n335), .B(n233), .A(n226) );
MUX2_X2 inst_632 ( .Z(net_130), .S(n1689), .A(n149), .B(n146) );
NAND2_X1 inst_549 ( .ZN(net_430), .A2(net_369), .A1(net_257) );
NOR2_X1 inst_234 ( .A1(net_740), .ZN(net_194), .A2(n4088) );
XOR2_X1 inst_0 ( .Z(net_79), .A(n302), .B(n293) );
NAND2_X1 inst_522 ( .ZN(net_314), .A2(net_312), .A1(n82) );
NOR3_X1 inst_184 ( .ZN(net_222), .A2(net_221), .A1(net_51), .A3(net_19) );
MUX2_X2 inst_690 ( .A(net_649), .B(net_648), .Z(net_647), .S(n4088) );
NOR2_X1 inst_236 ( .A2(net_748), .ZN(net_215), .A1(net_4) );
NAND2_X1 inst_433 ( .A2(net_160), .ZN(net_44), .A1(n131) );
NAND2_X1 inst_553 ( .ZN(net_488), .A1(net_446), .A2(net_374) );
NAND2_X1 inst_478 ( .A2(net_194), .ZN(net_191), .A1(n67) );
XNOR2_X1 inst_65 ( .ZN(net_596), .B(net_412), .A(net_383) );
NAND2_X1 inst_536 ( .A2(net_578), .ZN(net_485), .A1(net_348) );
NOR2_X1 inst_242 ( .ZN(net_51), .A1(net_50), .A2(n248) );
MUX2_X2 inst_688 ( .Z(net_644), .B(net_643), .A(net_417), .S(n4091) );
INV_X1 inst_781 ( .ZN(net_271), .A(n389) );
MUX2_X2 inst_732 ( .Z(net_736), .A(net_735), .B(net_734), .S(n4088) );
NAND2_X1 inst_516 ( .ZN(net_274), .A1(net_229), .A2(net_95) );
XNOR2_X1 inst_98 ( .ZN(net_579), .A(net_578), .B(net_533) );
INV_X1 inst_804 ( .ZN(net_165), .A(n809) );
NOR2_X1 inst_263 ( .ZN(net_318), .A1(net_164), .A2(n809) );
NOR3_X1 inst_190 ( .ZN(net_234), .A2(net_233), .A1(net_115), .A3(net_35) );
NOR3_X1 inst_185 ( .ZN(net_224), .A2(net_223), .A1(net_127), .A3(net_34) );
XOR2_X1 inst_13 ( .Z(net_363), .B(net_288), .A(n523) );
XNOR2_X1 inst_75 ( .B(net_519), .ZN(net_505), .A(net_470) );
NOR2_X1 inst_332 ( .ZN(net_518), .A2(net_517), .A1(net_477) );
OR2_X2 inst_166 ( .ZN(net_653), .A2(net_618), .A1(n4087) );
XNOR2_X1 inst_116 ( .ZN(net_632), .B(net_599), .A(net_575) );
MUX2_X2 inst_598 ( .Z(net_436), .S(n361), .A(n251), .B(n248) );
NAND3_X1 inst_416 ( .A2(net_782), .A3(net_781), .A1(net_162), .ZN(n882) );
AND4_X1 inst_868 ( .ZN(net_601), .A2(net_556), .A4(n559), .A3(n386), .A1(n245) );
OR2_X2 inst_163 ( .ZN(net_594), .A2(net_559), .A1(n1694) );
NAND2_X1 inst_471 ( .ZN(net_183), .A2(net_181), .A1(n188) );
NAND3_X1 inst_394 ( .A3(net_652), .A2(net_206), .A1(net_188), .ZN(n802) );
XNOR2_X1 inst_79 ( .ZN(net_571), .A(net_547), .B(net_521) );
INV_X1 inst_799 ( .ZN(net_158), .A(n514) );
XNOR2_X1 inst_106 ( .ZN(net_599), .B(net_570), .A(net_547) );
MUX2_X2 inst_738 ( .Z(net_767), .B(net_762), .A(net_657), .S(n2174) );
NAND2_X1 inst_422 ( .ZN(net_782), .A2(n4092), .A1(n4091) );
NOR2_X1 inst_219 ( .ZN(net_19), .A2(n281), .A1(n251) );
INV_X1 inst_840 ( .ZN(net_634), .A(net_620) );
MUX2_X2 inst_719 ( .Z(net_705), .B(n865), .A(n826), .S(n1689) );
NOR3_X1 inst_201 ( .A3(net_656), .ZN(net_422), .A2(net_421), .A1(net_372) );
MUX2_X2 inst_605 ( .Z(net_96), .S(n316), .A(n254), .B(n242) );
NOR2_X1 inst_304 ( .A2(net_547), .A1(net_377), .ZN(net_365) );
INV_X1 inst_752 ( .ZN(n593), .A(n299) );
NAND2_X1 inst_542 ( .A2(net_392), .ZN(net_369), .A1(net_368) );
NOR2_X1 inst_255 ( .ZN(net_102), .A1(net_101), .A2(n3546) );
NAND2_X1 inst_453 ( .ZN(net_399), .A2(n809), .A1(n2358) );
XNOR2_X1 inst_128 ( .ZN(net_692), .B(net_691), .A(net_680) );
XNOR2_X1 inst_73 ( .ZN(net_498), .B(net_436), .A(net_411) );
NAND2_X1 inst_493 ( .ZN(net_210), .A2(net_208), .A1(n70) );
AND2_X2 inst_896 ( .A2(net_401), .ZN(n673), .A1(n141) );
NAND3_X1 inst_378 ( .ZN(net_304), .A2(net_278), .A3(net_135), .A1(net_23) );
XOR2_X1 inst_23 ( .Z(net_578), .B(net_327), .A(n490) );
NOR2_X1 inst_339 ( .A2(net_662), .ZN(net_576), .A1(net_526) );
NAND3_X1 inst_351 ( .ZN(net_40), .A1(n1690), .A3(n1689), .A2(n158) );
AND2_X4 inst_890 ( .ZN(net_532), .A1(net_486), .A2(net_485) );
NAND3_X1 inst_361 ( .ZN(net_120), .A1(n4090), .A3(n4089), .A2(n17) );
NAND3_X1 inst_408 ( .ZN(net_758), .A3(net_743), .A1(net_214), .A2(net_170) );
NOR2_X1 inst_325 ( .ZN(net_475), .A2(net_464), .A1(net_463) );
NAND2_X1 inst_461 ( .A2(net_178), .ZN(net_171), .A1(n188) );
INV_X1 inst_829 ( .ZN(net_484), .A(net_483) );
NAND3_X1 inst_385 ( .ZN(net_551), .A1(net_493), .A2(net_492), .A3(net_485) );
INV_X1 inst_812 ( .ZN(net_583), .A(net_357) );
NOR3_X1 inst_197 ( .ZN(net_244), .A1(net_141), .A3(net_15), .A2(n374) );
MUX2_X2 inst_659 ( .A(net_527), .B(net_150), .Z(n838), .S(n4092) );
NOR2_X1 inst_250 ( .A1(net_750), .ZN(net_178), .A2(n1691) );
INV_X1 inst_848 ( .ZN(net_780), .A(net_778) );
NOR4_X1 inst_179 ( .ZN(net_541), .A3(net_459), .A4(net_456), .A2(net_430), .A1(net_395) );
XOR2_X1 inst_24 ( .Z(net_328), .A(net_327), .B(net_325) );
XNOR2_X1 inst_114 ( .ZN(net_625), .B(net_604), .A(net_469) );
INV_X1 inst_786 ( .ZN(n851), .A(n559) );
MUX2_X2 inst_617 ( .Z(net_113), .S(n4088), .A(n109), .B(n106) );
XNOR2_X1 inst_76 ( .ZN(net_504), .A(net_431), .B(net_409) );
NAND3_X1 inst_397 ( .A3(net_685), .A2(net_196), .A1(net_116), .ZN(n792) );
NAND2_X1 inst_504 ( .ZN(net_256), .A2(net_88), .A1(n523) );
OR2_X4 inst_150 ( .ZN(net_526), .A2(net_485), .A1(net_316) );
OR2_X2 inst_172 ( .ZN(net_723), .A2(net_706), .A1(n4090) );
NAND3_X1 inst_362 ( .ZN(net_121), .A1(n1690), .A3(n1689), .A2(n167) );
NOR2_X1 inst_277 ( .ZN(net_266), .A2(net_100), .A1(n411) );
XNOR2_X1 inst_83 ( .B(net_479), .A(net_388), .ZN(n1000) );
AND2_X4 inst_887 ( .A2(net_460), .ZN(net_445), .A1(n4) );
XNOR2_X1 inst_121 ( .ZN(net_660), .A(net_630), .B(net_614) );
NAND2_X1 inst_534 ( .ZN(net_457), .A1(net_363), .A2(net_357) );
NAND2_X1 inst_440 ( .A2(net_160), .ZN(net_70), .A1(n123) );
NOR2_X1 inst_306 ( .A1(net_656), .A2(net_583), .ZN(net_443) );
XOR2_X1 inst_2 ( .Z(net_81), .A(n210), .B(n206) );
MUX2_X2 inst_644 ( .Z(net_154), .S(n4089), .B(n103), .A(n100) );
MUX2_X2 inst_596 ( .Z(net_87), .S(n257), .A(n251), .B(n248) );
NAND2_X1 inst_578 ( .A1(net_748), .ZN(net_743), .A2(net_701) );
AND2_X4 inst_888 ( .A2(net_468), .ZN(net_449), .A1(n54) );
XNOR2_X1 inst_52 ( .ZN(net_547), .B(net_321), .A(n446) );
XNOR2_X1 inst_90 ( .ZN(net_544), .B(net_515), .A(net_249) );
INV_X1 inst_847 ( .ZN(net_773), .A(net_771) );
NOR2_X1 inst_267 ( .A2(net_282), .ZN(net_249), .A1(n374) );
OR3_X4 inst_140 ( .A1(net_656), .ZN(net_458), .A3(net_457), .A2(net_349) );
MUX2_X2 inst_668 ( .Z(net_637), .S(net_607), .A(net_596), .B(net_531) );
NOR2_X1 inst_221 ( .ZN(net_22), .A2(n251), .A1(n206) );
MUX2_X2 inst_748 ( .Z(net_787), .A(net_786), .B(net_785), .S(n1691) );
MUX2_X2 inst_716 ( .Z(net_702), .A(net_700), .B(net_699), .S(n1691) );
NAND2_X1 inst_556 ( .ZN(net_451), .A2(net_450), .A1(net_315) );
MUX2_X2 inst_650 ( .Z(net_481), .B(net_480), .A(net_438), .S(n4091) );
MUX2_X2 inst_637 ( .Z(net_134), .S(n4089), .A(n109), .B(n106) );
NOR2_X1 inst_289 ( .ZN(net_339), .A2(net_250), .A1(net_232) );
INV_X1 inst_792 ( .ZN(net_231), .A(n468) );
NAND2_X1 inst_547 ( .ZN(net_407), .A2(net_406), .A1(net_359) );
NAND2_X1 inst_530 ( .ZN(net_434), .A1(net_300), .A2(net_269) );
MUX2_X2 inst_720 ( .Z(net_706), .B(n865), .A(n826), .S(n4089) );
NAND2_X1 inst_432 ( .A2(net_160), .ZN(net_41), .A1(n115) );
MUX2_X2 inst_679 ( .Z(net_671), .A(net_589), .B(net_149), .S(n4092) );
NAND3_X1 inst_420 ( .ZN(net_794), .A3(net_789), .A2(net_219), .A1(net_173) );
NOR2_X1 inst_282 ( .ZN(net_273), .A1(net_221), .A2(net_108) );
NAND3_X1 inst_368 ( .ZN(net_156), .A3(net_155), .A1(n4090), .A2(n11) );
NAND2_X1 inst_513 ( .ZN(net_446), .A2(net_283), .A1(n411) );
INV_X1 inst_803 ( .ZN(net_229), .A(n411) );
INV_X1 inst_754 ( .ZN(net_59), .A(n324) );
INV_X1 inst_769 ( .ZN(net_124), .A(n248) );
XNOR2_X1 inst_44 ( .ZN(net_630), .B(net_282), .A(n374) );
NOR2_X1 inst_274 ( .A2(net_602), .A1(net_534), .ZN(net_315) );
OR2_X2 inst_174 ( .ZN(net_725), .A2(net_707), .A1(n4087) );
NAND3_X1 inst_371 ( .ZN(net_162), .A3(net_160), .A1(n4092), .A2(n118) );
MUX2_X2 inst_701 ( .Z(net_699), .A(net_627), .B(net_71), .S(n4092) );
MUX2_X2 inst_662 ( .Z(net_580), .B(net_542), .A(net_381), .S(n4091) );
NOR2_X1 inst_314 ( .ZN(net_403), .A1(net_402), .A2(net_332) );
CLKBUF_X1 inst_867 ( .Z(n144), .A(n141) );
NAND2_X1 inst_435 ( .ZN(net_60), .A2(net_59), .A1(n3550) );
OR2_X2 inst_164 ( .ZN(net_595), .A2(net_560), .A1(n1690) );
INV_X1 inst_820 ( .ZN(net_335), .A(net_334) );
XOR2_X1 inst_5 ( .Z(net_84), .A(n351), .B(n341) );
MUX2_X2 inst_597 ( .Z(net_88), .S(n341), .A(n251), .B(n248) );
MUX2_X2 inst_729 ( .Z(net_731), .A(net_696), .B(net_695), .S(n1497) );
OR2_X2 inst_157 ( .ZN(net_261), .A2(net_96), .A1(n490) );
MUX2_X2 inst_687 ( .Z(net_642), .B(net_638), .A(net_414), .S(n4091) );
INV_X1 inst_774 ( .ZN(net_227), .A(n534) );
MUX2_X2 inst_621 ( .Z(net_286), .B(n358), .A(n351), .S(n332) );
XNOR2_X1 inst_68 ( .ZN(net_478), .B(net_386), .A(net_333) );
NOR3_X1 inst_213 ( .ZN(net_713), .A3(net_711), .A2(net_662), .A1(n2174) );
MUX2_X2 inst_604 ( .Z(net_95), .A(n3548), .B(n3546), .S(n273) );
INV_X1 inst_838 ( .A(net_671), .ZN(n873) );
XNOR2_X1 inst_53 ( .ZN(net_326), .B(net_292), .A(net_291) );
MUX2_X2 inst_628 ( .Z(net_283), .S(n335), .B(n280), .A(n273) );
INV_X1 inst_753 ( .ZN(net_663), .A(n2174) );
NOR3_X1 inst_205 ( .ZN(net_524), .A1(net_464), .A3(net_463), .A2(net_393) );
INV_X1 inst_815 ( .ZN(net_691), .A(net_392) );
NAND2_X1 inst_472 ( .ZN(net_185), .A2(net_184), .A1(n52) );
NAND2_X1 inst_447 ( .ZN(net_125), .A2(net_124), .A1(n316) );
NAND3_X1 inst_380 ( .ZN(net_306), .A2(net_271), .A3(net_86), .A1(net_32) );
NAND2_X1 inst_457 ( .A2(net_181), .ZN(net_167), .A1(n176) );
AND2_X4 inst_875 ( .A2(net_124), .ZN(net_66), .A1(n206) );
MUX2_X2 inst_651 ( .A(net_420), .B(net_44), .Z(n822), .S(n4092) );
MUX2_X2 inst_665 ( .Z(net_589), .B(net_588), .A(net_380), .S(n4091) );
NOR2_X1 inst_292 ( .ZN(net_341), .A2(net_255), .A1(net_228) );
NAND3_X1 inst_379 ( .ZN(net_305), .A2(net_280), .A3(net_151), .A1(net_30) );
XNOR2_X1 inst_127 ( .ZN(net_688), .A(net_668), .B(net_605) );
CLKBUF_X1 inst_855 ( .Z(n923), .A(n141) );
NOR3_X1 inst_186 ( .ZN(net_226), .A2(net_225), .A1(net_122), .A3(net_13) );
XOR2_X1 inst_17 ( .Z(net_575), .B(net_293), .A(n422) );
MUX2_X2 inst_706 ( .A(net_642), .B(net_75), .Z(n830), .S(n4092) );
INV_X1 inst_759 ( .ZN(net_50), .A(n281) );
NAND3_X1 inst_413 ( .ZN(net_764), .A1(net_749), .A3(net_174), .A2(net_119) );
OR2_X4 inst_146 ( .A2(net_547), .ZN(net_425), .A1(net_402) );
NOR2_X1 inst_249 ( .A1(net_0), .ZN(n815), .A2(n3173) );
NOR2_X1 inst_334 ( .ZN(net_546), .A2(net_521), .A1(net_424) );
CLKBUF_X1 inst_859 ( .Z(n887), .A(n299) );
NOR3_X1 inst_187 ( .ZN(net_228), .A2(net_227), .A1(net_52), .A3(net_25) );
NOR3_X1 inst_206 ( .ZN(net_483), .A2(net_469), .A3(net_457), .A1(net_405) );
INV_X1 inst_805 ( .A(net_469), .ZN(net_364) );
XNOR2_X1 inst_122 ( .ZN(net_693), .B(net_632), .A(net_546) );
CLKBUF_X1 inst_863 ( .A(n606), .Z(n602) );
XOR2_X1 inst_25 ( .Z(net_329), .B(net_293), .A(net_289) );
INV_X1 inst_839 ( .ZN(net_672), .A(n834) );
NAND3_X1 inst_354 ( .ZN(net_98), .A1(n4088), .A3(n4087), .A2(n17) );
NAND3_X1 inst_405 ( .A3(net_741), .A2(net_193), .A1(net_37), .ZN(n747) );
NAND2_X1 inst_492 ( .ZN(net_209), .A2(net_208), .A1(n61) );
NOR2_X1 inst_240 ( .A1(net_748), .ZN(net_181), .A2(n1689) );
INV_X1 inst_817 ( .ZN(net_519), .A(net_330) );
NOR2_X1 inst_326 ( .A1(net_488), .ZN(net_487), .A2(net_460) );
XNOR2_X1 inst_110 ( .ZN(net_609), .B(net_584), .A(net_577) );
AND2_X4 inst_891 ( .ZN(net_525), .A2(net_524), .A1(net_495) );
NAND2_X1 inst_518 ( .A1(net_534), .ZN(net_307), .A2(net_163) );
XNOR2_X1 inst_74 ( .ZN(net_499), .A(net_410), .B(net_336) );
NOR2_X1 inst_288 ( .ZN(net_338), .A2(net_248), .A1(net_224) );
NAND3_X1 inst_396 ( .A3(net_678), .A2(net_199), .A1(net_98), .ZN(n757) );
NOR2_X1 inst_229 ( .ZN(net_33), .A2(n265), .A1(n251) );
XNOR2_X1 inst_99 ( .ZN(net_584), .B(net_583), .A(net_537) );
XNOR2_X1 inst_69 ( .B(net_384), .A(net_294), .ZN(n1004) );
NAND3_X1 inst_373 ( .ZN(net_239), .A1(net_65), .A3(net_21), .A2(n479) );
XNOR2_X1 inst_82 ( .B(net_478), .A(net_413), .ZN(n998) );
MUX2_X2 inst_669 ( .Z(net_636), .S(net_607), .A(net_606), .B(net_552) );
XNOR2_X1 inst_108 ( .ZN(net_604), .B(net_563), .A(net_545) );
INV_X1 inst_844 ( .ZN(net_717), .A(n828) );
MUX2_X2 inst_664 ( .Z(net_587), .B(net_586), .A(net_435), .S(n4091) );
MUX2_X2 inst_595 ( .Z(net_64), .A(n251), .B(n248), .S(n226) );
NOR2_X1 inst_283 ( .ZN(net_275), .A1(net_233), .A2(net_110) );
XOR2_X1 inst_22 ( .Z(net_348), .B(net_325), .A(n479) );
NOR2_X1 inst_311 ( .ZN(net_382), .A1(net_381), .A2(net_380) );
AND2_X2 inst_917 ( .A2(net_764), .ZN(n654), .A1(n137) );
NAND2_X1 inst_460 ( .A2(net_181), .ZN(net_170), .A1(n200) );
NAND3_X1 inst_372 ( .ZN(net_237), .A1(net_125), .A3(net_10), .A2(n490) );
OR2_X2 inst_169 ( .ZN(net_659), .A2(net_629), .A1(n4092) );
NOR2_X1 inst_215 ( .ZN(net_13), .A2(n324), .A1(n251) );
NOR2_X1 inst_307 ( .A1(net_656), .A2(net_605), .ZN(net_404) );
INV_X1 inst_767 ( .ZN(net_57), .A(n226) );
MUX2_X2 inst_638 ( .Z(net_602), .S(n332), .B(n299), .A(n293) );
NAND2_X1 inst_421 ( .ZN(n847), .A2(n556), .A1(n386) );
OR2_X2 inst_161 ( .ZN(net_592), .A2(net_557), .A1(n4090) );
NAND2_X1 inst_560 ( .ZN(net_522), .A2(net_483), .A1(n54) );
MUX2_X2 inst_749 ( .Z(net_788), .A(net_786), .B(net_785), .S(n4089) );
NAND2_X1 inst_586 ( .ZN(net_790), .A2(net_788), .A1(net_738) );
CLKBUF_X1 inst_849 ( .Z(n993), .A(n1) );
MUX2_X2 inst_702 ( .Z(net_681), .A(net_650), .B(net_131), .S(n1694) );
NAND2_X1 inst_555 ( .ZN(net_492), .A2(net_450), .A1(net_343) );
XOR2_X1 inst_16 ( .Z(net_330), .B(net_292), .A(n457) );
INV_X1 inst_816 ( .ZN(net_605), .A(net_359) );
MUX2_X2 inst_717 ( .Z(net_703), .B(n869), .A(n830), .S(n1689) );
NOR2_X1 inst_276 ( .ZN(net_265), .A2(net_99), .A1(n374) );
MUX2_X2 inst_718 ( .Z(net_704), .B(n869), .A(n830), .S(n1691) );
NAND2_X1 inst_431 ( .A2(net_8), .ZN(n845), .A1(n27) );
NAND4_X1 inst_348 ( .ZN(net_639), .A3(net_638), .A4(net_637), .A2(net_628), .A1(net_586) );
XOR2_X1 inst_3 ( .Z(net_82), .A(n226), .B(n218) );
OR2_X2 inst_156 ( .ZN(net_21), .A2(n308), .A1(n251) );
AND2_X4 inst_889 ( .ZN(net_477), .A2(net_476), .A1(n54) );
NAND2_X1 inst_577 ( .A1(net_750), .ZN(net_742), .A2(net_702) );
AND2_X4 inst_886 ( .A2(net_394), .A1(net_393), .ZN(net_370) );
INV_X1 inst_802 ( .ZN(net_8), .A(n2824) );
NAND2_X1 inst_566 ( .ZN(net_566), .A2(net_565), .A1(net_496) );
NOR2_X1 inst_296 ( .ZN(net_509), .A1(net_276), .A2(net_245) );
XNOR2_X1 inst_91 ( .ZN(net_545), .A(net_516), .B(net_472) );
AND2_X2 inst_905 ( .A2(net_682), .ZN(n667), .A1(n137) );
XNOR2_X1 inst_132 ( .ZN(net_755), .A(net_729), .B(net_720) );
NAND4_X1 inst_342 ( .ZN(net_400), .A2(net_399), .A3(net_398), .A4(net_319), .A1(net_313) );
NAND2_X1 inst_526 ( .ZN(net_320), .A2(net_318), .A1(n81) );
XOR2_X1 inst_36 ( .B(net_756), .Z(net_588), .A(net_525) );
MUX2_X2 inst_656 ( .Z(net_558), .B(n861), .A(n822), .S(n4088) );
MUX2_X2 inst_645 ( .Z(net_159), .S(net_158), .A(net_124), .B(n242) );
NAND2_X1 inst_463 ( .A2(net_178), .ZN(net_173), .A1(n176) );
NAND2_X1 inst_503 ( .ZN(net_366), .A2(net_292), .A1(n457) );
XNOR2_X1 inst_96 ( .ZN(net_570), .A(net_569), .B(net_568) );
XNOR2_X1 inst_45 ( .B(net_469), .ZN(net_334), .A(n54) );
NAND2_X1 inst_451 ( .ZN(net_151), .A2(net_55), .A1(n254) );
XNOR2_X1 inst_101 ( .ZN(net_585), .A(net_544), .B(net_487) );
NOR2_X1 inst_319 ( .A1(net_583), .ZN(net_476), .A2(net_375) );
NOR2_X1 inst_269 ( .A2(net_327), .ZN(net_253), .A1(n490) );
NAND2_X1 inst_458 ( .A2(net_181), .ZN(net_168), .A1(n194) );
NAND2_X1 inst_444 ( .A2(net_160), .ZN(net_75), .A1(n112) );
NAND3_X1 inst_400 ( .ZN(net_753), .A1(net_726), .A2(net_216), .A3(net_182) );
INV_X1 inst_797 ( .ZN(n611), .A(n338) );
MUX2_X2 inst_614 ( .Z(net_109), .B(n3552), .A(n3550), .S(n341) );
MUX2_X2 inst_686 ( .Z(net_641), .B(net_637), .A(net_415), .S(n4091) );
MUX2_X2 inst_649 ( .A(net_436), .Z(net_420), .B(net_335), .S(n4091) );
INV_X1 inst_821 ( .ZN(net_412), .A(net_348) );
MUX2_X2 inst_741 ( .Z(net_772), .A(net_770), .B(net_769), .S(n4091) );
NOR2_X1 inst_261 ( .ZN(net_145), .A1(net_101), .A2(n248) );
NAND2_X1 inst_514 ( .ZN(net_264), .A2(net_87), .A1(n389) );
NAND2_X1 inst_500 ( .ZN(net_219), .A2(net_217), .A1(n179) );
NAND2_X1 inst_510 ( .ZN(net_389), .A2(net_293), .A1(n422) );
NOR2_X1 inst_268 ( .ZN(net_250), .A2(net_91), .A1(n468) );
MUX2_X2 inst_685 ( .Z(net_640), .B(net_636), .S(n3724), .A(n123) );
NAND3_X1 inst_369 ( .ZN(net_157), .A3(net_155), .A1(n4090), .A2(n14) );
NAND2_X1 inst_550 ( .ZN(net_470), .A2(net_428), .A1(net_377) );
XNOR2_X1 inst_63 ( .ZN(net_411), .A(net_340), .B(net_159) );
XNOR2_X1 inst_119 ( .ZN(net_645), .B(net_608), .A(net_602) );
INV_X1 inst_830 ( .ZN(net_506), .A(net_505) );
MUX2_X2 inst_603 ( .Z(net_94), .A(n254), .B(n242), .S(n206) );
NOR2_X1 inst_327 ( .A1(net_503), .A2(net_462), .ZN(n632) );
MUX2_X2 inst_676 ( .Z(net_616), .B(n877), .A(n838), .S(n1689) );
XNOR2_X1 inst_85 ( .ZN(net_581), .A(net_536), .B(net_491) );
NOR2_X1 inst_291 ( .ZN(net_340), .A2(net_254), .A1(net_226) );
NOR2_X1 inst_266 ( .ZN(net_248), .A2(net_45), .A1(n457) );
INV_X1 inst_776 ( .ZN(net_5), .A(n1691) );
AND2_X2 inst_900 ( .A2(net_624), .ZN(n661), .A1(n137) );
AND3_X2 inst_874 ( .A1(net_683), .A2(net_643), .A3(n623), .ZN(n585) );
NAND2_X1 inst_473 ( .ZN(net_186), .A2(net_184), .A1(n53) );
CLKBUF_X1 inst_866 ( .Z(n298), .A(n293) );
NOR2_X1 inst_217 ( .ZN(net_15), .A2(n3548), .A1(n281) );
NAND2_X1 inst_572 ( .ZN(net_700), .A2(net_659), .A1(net_185) );
MUX2_X2 inst_742 ( .Z(net_778), .A(net_777), .B(net_776), .S(n4091) );
XNOR2_X1 inst_77 ( .ZN(net_549), .B(net_534), .A(net_486) );
OR2_X2 inst_171 ( .ZN(net_722), .A2(net_705), .A1(n1690) );
MUX2_X2 inst_691 ( .Z(net_650), .A(net_649), .B(net_648), .S(n1691) );
NAND2_X1 inst_558 ( .ZN(net_500), .A2(net_461), .A1(n4) );
NAND2_X1 inst_427 ( .ZN(n809), .A2(n31), .A1(n27) );
NOR2_X1 inst_257 ( .ZN(net_122), .A1(net_59), .A2(n248) );
MUX2_X2 inst_594 ( .Z(net_45), .A(n254), .B(n242), .S(n210) );
OR2_X4 inst_145 ( .ZN(net_428), .A2(net_402), .A1(net_389) );
NOR2_X1 inst_290 ( .ZN(net_351), .A1(net_268), .A2(net_240) );
NAND3_X1 inst_374 ( .ZN(net_300), .A3(net_60), .A1(net_16), .A2(n503) );
NOR2_X1 inst_272 ( .ZN(net_259), .A2(net_94), .A1(n446) );
NAND2_X1 inst_502 ( .ZN(net_251), .A2(net_64), .A1(n422) );
XNOR2_X1 inst_103 ( .ZN(net_597), .A(net_596), .B(net_550) );
NAND2_X1 inst_485 ( .ZN(net_200), .A2(net_197), .A1(n73) );
INV_X1 inst_814 ( .ZN(net_536), .A(net_363) );
INV_X1 inst_770 ( .ZN(net_48), .A(n351) );
NAND2_X1 inst_565 ( .A2(net_565), .ZN(net_564), .A1(net_453) );
NOR2_X1 inst_248 ( .A2(net_750), .ZN(net_217), .A1(net_5) );
CLKBUF_X1 inst_861 ( .A(n629), .Z(n618) );
MUX2_X2 inst_672 ( .Z(net_649), .A(net_582), .B(net_69), .S(n4092) );
MUX2_X2 inst_622 ( .Z(net_288), .B(n348), .A(n341), .S(n332) );
OR4_X1 inst_138 ( .A1(net_539), .A2(net_520), .A4(net_367), .A3(net_252), .ZN(n621) );
NAND3_X1 inst_389 ( .ZN(net_624), .A3(net_595), .A2(net_220), .A1(net_166) );
INV_X1 inst_789 ( .ZN(net_225), .A(n503) );
NAND3_X1 inst_357 ( .ZN(net_116), .A1(n4090), .A3(n4089), .A2(n20) );
NAND3_X1 inst_409 ( .ZN(net_759), .A3(net_742), .A1(net_211), .A2(net_180) );
AND2_X2 inst_899 ( .A2(net_623), .ZN(n693), .A1(n137) );
INV_X1 inst_809 ( .ZN(net_316), .A(net_315) );
AND2_X4 inst_881 ( .ZN(net_368), .A2(net_285), .A1(n389) );
INV_X1 inst_822 ( .ZN(net_352), .A(net_351) );
AND2_X2 inst_913 ( .A2(net_759), .ZN(n676), .A1(n137) );
NOR4_X1 inst_180 ( .ZN(net_556), .A3(n998), .A2(n1004), .A1(n1002), .A4(n1000) );
MUX2_X2 inst_703 ( .Z(net_682), .A(net_651), .B(net_129), .S(n1690) );
XOR2_X1 inst_33 ( .Z(net_432), .A(net_354), .B(net_341) );
NOR2_X1 inst_312 ( .ZN(net_450), .A2(net_412), .A1(net_383) );
MUX2_X2 inst_660 ( .Z(net_612), .S(net_574), .A(net_573), .B(net_568) );
AND2_X2 inst_912 ( .A2(net_763), .ZN(n679), .A1(n137) );
MUX2_X2 inst_731 ( .A(net_735), .B(net_734), .Z(net_733), .S(n1691) );
MUX2_X2 inst_609 ( .Z(net_103), .A(n3548), .B(n3546), .S(n324) );
NAND2_X1 inst_517 ( .ZN(net_279), .A1(net_278), .A2(net_105) );
NOR2_X1 inst_309 ( .A2(net_536), .ZN(net_465), .A1(net_421) );
NOR2_X1 inst_232 ( .ZN(net_36), .A2(n3548), .A1(n341) );
NAND4_X1 inst_347 ( .ZN(net_528), .A1(net_467), .A2(net_407), .A4(net_361), .A3(net_258) );
INV_X1 inst_768 ( .ZN(net_3), .A(n332) );
INV_X1 inst_795 ( .ZN(n599), .A(n348) );
MUX2_X2 inst_663 ( .Z(net_582), .B(net_581), .A(net_482), .S(n4091) );
NOR2_X1 inst_301 ( .ZN(net_346), .A2(net_266), .A1(net_230) );
NAND3_X1 inst_363 ( .ZN(net_123), .A1(n4088), .A3(n4087), .A2(n40) );
INV_X1 inst_755 ( .ZN(net_155), .A(n4089) );
XOR2_X1 inst_27 ( .Z(net_568), .A(net_402), .B(net_260) );
NOR2_X1 inst_247 ( .A1(net_740), .ZN(net_208), .A2(net_136) );
NOR2_X1 inst_297 ( .ZN(net_510), .A2(net_259), .A1(net_238) );
NAND3_X1 inst_403 ( .A3(net_739), .A2(net_187), .A1(net_117), .ZN(n787) );
NOR2_X1 inst_302 ( .ZN(net_347), .A2(net_265), .A1(net_222) );
NOR2_X1 inst_310 ( .A1(net_534), .ZN(net_493), .A2(net_379) );
NOR2_X1 inst_322 ( .A2(net_490), .ZN(net_472), .A1(net_468) );
MUX2_X2 inst_673 ( .Z(net_611), .B(net_610), .A(net_509), .S(n4091) );
NOR2_X1 inst_253 ( .ZN(net_295), .A1(net_3), .A2(n338) );
NOR3_X1 inst_211 ( .A1(net_667), .A3(net_619), .A2(net_610), .ZN(n575) );
MUX2_X2 inst_619 ( .Z(net_325), .S(n332), .B(n315), .A(n308) );
MUX2_X2 inst_681 ( .Z(net_620), .B(net_619), .A(net_510), .S(n4091) );
OR2_X2 inst_162 ( .ZN(net_593), .A2(net_558), .A1(n4087) );
NAND2_X1 inst_589 ( .A2(net_794), .ZN(n690), .A1(n137) );
NAND2_X1 inst_561 ( .A2(net_541), .ZN(net_540), .A1(net_502) );
INV_X1 inst_794 ( .ZN(net_738), .A(n4090) );
NAND3_X1 inst_412 ( .ZN(net_763), .A3(net_728), .A2(net_218), .A1(net_179) );
NAND2_X1 inst_449 ( .ZN(net_142), .A2(net_77), .A1(n3550) );
MUX2_X2 inst_639 ( .Z(net_469), .B(n366), .A(n361), .S(n332) );
AND2_X4 inst_877 ( .A2(net_160), .ZN(net_71), .A1(n122) );
OR2_X2 inst_155 ( .ZN(net_10), .A2(n316), .A1(n251) );
NAND2_X1 inst_464 ( .A2(net_181), .ZN(net_174), .A1(n191) );
AND3_X4 inst_871 ( .ZN(net_664), .A1(net_663), .A2(net_662), .A3(net_661) );
MUX2_X2 inst_602 ( .Z(net_93), .S(n265), .A(n254), .B(n242) );
XNOR2_X1 inst_59 ( .ZN(net_386), .A(net_323), .B(net_296) );
XNOR2_X1 inst_135 ( .ZN(net_766), .B(net_756), .A(net_755) );
NAND4_X1 inst_341 ( .A2(net_399), .A3(net_398), .ZN(net_397), .A1(net_311), .A4(net_301) );
NOR3_X1 inst_196 ( .ZN(net_243), .A1(net_102), .A3(net_17), .A2(n400) );
NAND2_X1 inst_532 ( .ZN(net_439), .A1(net_302), .A2(net_274) );
XNOR2_X1 inst_55 ( .B(net_417), .A(net_416), .ZN(net_336) );
XOR2_X1 inst_37 ( .Z(net_548), .A(net_547), .B(net_546) );
MUX2_X2 inst_641 ( .Z(net_148), .B(n3552), .A(n3550), .S(n210) );
NAND2_X1 inst_498 ( .ZN(net_216), .A2(net_215), .A1(n173) );
MUX2_X2 inst_740 ( .Z(net_771), .A(net_770), .B(net_769), .S(n4091) );
MUX2_X2 inst_684 ( .Z(net_629), .B(net_628), .A(net_434), .S(n4091) );
NOR2_X1 inst_264 ( .ZN(net_312), .A2(n809), .A1(n2358) );
XNOR2_X1 inst_84 ( .A(net_729), .ZN(net_542), .B(net_489) );
MUX2_X2 inst_723 ( .Z(net_709), .B(n869), .A(n830), .S(n4089) );
OR2_X2 inst_173 ( .ZN(net_724), .A2(net_710), .A1(n4087) );
NOR2_X1 inst_298 ( .ZN(net_355), .A1(net_277), .A2(net_246) );
NOR2_X1 inst_303 ( .A2(net_656), .ZN(net_406), .A1(net_309) );
MUX2_X2 inst_611 ( .Z(net_106), .B(n3552), .A(n3550), .S(n265) );
NOR2_X1 inst_224 ( .ZN(net_26), .A2(n3548), .A1(n210) );
XNOR2_X1 inst_42 ( .ZN(net_43), .A(n369), .B(n361) );
NOR2_X1 inst_287 ( .ZN(net_482), .A1(net_281), .A2(net_241) );
NOR2_X1 inst_323 ( .ZN(net_473), .A2(net_427), .A1(net_365) );
MUX2_X2 inst_618 ( .Z(net_290), .S(n332), .B(n331), .A(n324) );
NAND2_X1 inst_426 ( .ZN(net_18), .A2(n3552), .A1(n273) );
NAND2_X1 inst_588 ( .ZN(net_792), .A2(net_784), .A1(net_748) );
MUX2_X2 inst_648 ( .A(net_416), .Z(net_391), .B(net_390), .S(n3724) );
NAND3_X1 inst_350 ( .ZN(net_37), .A1(n4088), .A3(n4087), .A2(n37) );
NOR2_X1 inst_231 ( .ZN(net_35), .A2(n251), .A1(n234) );
NOR2_X1 inst_270 ( .ZN(net_254), .A2(net_42), .A1(n503) );
NAND2_X1 inst_474 ( .A2(net_197), .ZN(net_187), .A1(n43) );
INV_X1 inst_793 ( .ZN(n606), .A(n549) );
INV_X1 inst_766 ( .ZN(net_46), .A(n218) );
MUX2_X2 inst_715 ( .Z(net_701), .A(net_700), .B(net_699), .S(n1689) );
XOR2_X1 inst_26 ( .A(net_630), .Z(net_480), .B(n4) );
NAND2_X1 inst_437 ( .A2(net_124), .ZN(net_65), .A1(n308) );
NAND2_X1 inst_490 ( .ZN(net_206), .A2(net_203), .A1(n70) );
INV_X1 inst_801 ( .ZN(net_221), .A(n374) );
MUX2_X2 inst_626 ( .Z(net_291), .S(n335), .B(n225), .A(n218) );
MUX2_X2 inst_692 ( .Z(net_651), .A(net_649), .B(net_648), .S(n1689) );
XNOR2_X1 inst_70 ( .B(net_387), .A(net_298), .ZN(n1002) );
AND3_X4 inst_870 ( .ZN(net_395), .A1(net_394), .A2(net_393), .A3(net_392) );
XNOR2_X1 inst_129 ( .ZN(net_720), .B(net_691), .A(net_687) );
NOR3_X1 inst_189 ( .ZN(net_232), .A2(net_231), .A1(net_61), .A3(net_9) );
XOR2_X1 inst_11 ( .Z(net_357), .B(net_286), .A(n534) );
MUX2_X2 inst_631 ( .Z(net_129), .S(n1689), .A(n155), .B(n152) );
NOR3_X1 inst_188 ( .ZN(net_230), .A2(net_229), .A1(net_78), .A3(net_29) );
XOR2_X1 inst_14 ( .Z(net_392), .B(net_289), .A(n435) );
NAND2_X1 inst_475 ( .A2(net_197), .ZN(net_188), .A1(n67) );
NAND2_X1 inst_441 ( .A2(net_160), .ZN(net_72), .A1(n126) );
XOR2_X1 inst_31 ( .Z(net_431), .A(net_353), .B(net_339) );
NAND2_X1 inst_528 ( .ZN(net_414), .A2(net_261), .A1(net_237) );
CLKBUF_X1 inst_865 ( .A(n621), .Z(n591) );
NOR2_X1 inst_252 ( .ZN(net_78), .A1(net_77), .A2(n248) );
AND2_X2 inst_903 ( .A2(net_684), .A1(net_11), .ZN(n818) );
INV_X1 inst_798 ( .ZN(n850), .A(n562) );
XNOR2_X1 inst_62 ( .ZN(net_408), .B(net_346), .A(net_345) );
INV_X1 inst_808 ( .ZN(net_310), .A(net_309) );
INV_X1 inst_777 ( .ZN(net_235), .A(n400) );
NAND2_X1 inst_557 ( .ZN(net_494), .A1(net_493), .A2(net_492) );
NOR2_X1 inst_251 ( .A1(net_164), .ZN(net_76), .A2(n87) );
NAND3_X1 inst_352 ( .ZN(net_62), .A1(n1690), .A3(n1689), .A2(n164) );
NAND2_X1 inst_575 ( .ZN(net_739), .A1(net_738), .A2(net_697) );
NAND3_X1 inst_398 ( .A3(net_686), .A2(net_192), .A1(net_143), .ZN(n752) );
INV_X1 inst_846 ( .ZN(net_735), .A(n824) );
NOR2_X1 inst_286 ( .ZN(net_281), .A1(net_280), .A2(net_109) );
NAND2_X1 inst_436 ( .A2(net_160), .ZN(net_63), .A1(n113) );
AND2_X4 inst_879 ( .A2(net_160), .ZN(net_149), .A1(n128) );
INV_X1 inst_823 ( .ZN(net_356), .A(net_355) );
NAND2_X1 inst_484 ( .ZN(net_199), .A2(net_194), .A1(n73) );
MUX2_X2 inst_627 ( .Z(net_282), .S(n335), .B(n288), .A(n281) );
NOR2_X1 inst_300 ( .ZN(net_345), .A2(net_267), .A1(net_236) );
XNOR2_X1 inst_102 ( .ZN(net_777), .B(net_553), .A(net_504) );
XOR2_X1 inst_32 ( .B(net_583), .Z(net_512), .A(net_350) );
NAND4_X1 inst_344 ( .ZN(net_418), .A1(net_417), .A2(net_416), .A3(net_415), .A4(net_414) );
NAND2_X1 inst_428 ( .ZN(net_23), .A2(n242), .A1(n226) );
NAND2_X1 inst_446 ( .A2(net_160), .ZN(net_104), .A1(n117) );
NAND3_X1 inst_364 ( .ZN(net_137), .A1(net_136), .A3(n4087), .A2(n11) );
OR2_X4 inst_144 ( .ZN(net_438), .A1(net_273), .A2(net_244) );
MUX2_X2 inst_629 ( .Z(net_292), .S(n335), .B(n217), .A(n210) );
NOR3_X1 inst_195 ( .ZN(net_242), .A1(net_39), .A3(net_28), .A2(n389) );
NAND3_X1 inst_407 ( .A3(net_725), .A2(net_205), .A1(net_189), .ZN(n732) );
INV_X1 inst_824 ( .ZN(net_373), .A(net_372) );
INV_X1 inst_791 ( .ZN(net_750), .A(n1694) );
MUX2_X2 inst_623 ( .Z(net_287), .S(n335), .B(n272), .A(n265) );
NAND3_X1 inst_411 ( .ZN(net_761), .A1(net_746), .A3(net_177), .A2(net_114) );
XNOR2_X1 inst_97 ( .ZN(net_577), .A(net_562), .B(net_517) );
MUX2_X2 inst_616 ( .Z(net_111), .B(n3552), .A(n3550), .S(n351) );
AND2_X2 inst_898 ( .A2(net_396), .ZN(n715), .A1(n141) );
AND2_X4 inst_880 ( .A2(net_321), .ZN(net_252), .A1(n446) );
INV_X1 inst_775 ( .ZN(net_4), .A(n1689) );
XNOR2_X1 inst_124 ( .ZN(net_680), .A(net_679), .B(net_631) );
NAND2_X1 inst_533 ( .ZN(net_530), .A1(net_303), .A2(net_279) );
MUX2_X2 inst_620 ( .Z(net_289), .S(n335), .B(n241), .A(n234) );
MUX2_X2 inst_652 ( .Z(net_513), .B(net_512), .A(net_351), .S(n4091) );
MUX2_X2 inst_680 ( .A(net_587), .B(net_74), .Z(n834), .S(n4092) );
INV_X1 inst_785 ( .ZN(net_233), .A(n435) );
MUX2_X2 inst_737 ( .A(net_737), .B(net_134), .Z(n712), .S(n4090) );
AND2_X4 inst_876 ( .A2(net_160), .ZN(net_69), .A1(n119) );
XNOR2_X1 inst_137 ( .ZN(net_776), .B(net_768), .A(net_731) );
MUX2_X2 inst_677 ( .Z(net_617), .B(n877), .A(n838), .S(n4089) );
NAND2_X1 inst_425 ( .ZN(net_16), .A2(n3552), .A1(n324) );
NAND2_X1 inst_545 ( .A1(net_575), .ZN(net_423), .A2(net_330) );
XNOR2_X1 inst_130 ( .ZN(net_730), .B(net_729), .A(net_692) );
MUX2_X2 inst_722 ( .Z(net_708), .B(n865), .A(n826), .S(n1691) );
NOR2_X1 inst_227 ( .ZN(net_29), .A2(n273), .A1(n251) );
NAND3_X1 inst_399 ( .ZN(net_752), .A1(net_722), .A3(net_168), .A2(net_62) );
INV_X1 inst_760 ( .ZN(net_1), .A(n254) );
MUX2_X2 inst_746 ( .A(net_786), .B(net_785), .Z(net_783), .S(n4088) );
NAND2_X1 inst_527 ( .ZN(net_415), .A2(net_263), .A1(net_239) );
NOR2_X1 inst_226 ( .ZN(net_28), .A2(n3548), .A1(n257) );
OR2_X2 inst_176 ( .ZN(net_727), .A2(net_708), .A1(n1694) );
XNOR2_X1 inst_58 ( .ZN(net_385), .A(net_329), .B(net_322) );
NAND3_X1 inst_414 ( .ZN(net_765), .A1(net_751), .A3(net_175), .A2(net_92) );
XNOR2_X1 inst_87 ( .ZN(net_535), .B(net_534), .A(net_532) );
XNOR2_X1 inst_61 ( .ZN(net_388), .B(net_324), .A(net_284) );
NAND2_X1 inst_562 ( .ZN(net_574), .A2(net_541), .A1(net_500) );
NAND2_X1 inst_531 ( .ZN(net_354), .A2(net_305), .A1(net_256) );
NOR3_X1 inst_203 ( .ZN(net_456), .A1(net_455), .A2(net_454), .A3(net_452) );
NOR3_X1 inst_212 ( .ZN(net_712), .A3(net_711), .A2(net_665), .A1(net_663) );
NAND2_X1 inst_499 ( .ZN(net_218), .A2(net_217), .A1(n173) );
NOR2_X1 inst_335 ( .A1(net_756), .ZN(net_523), .A2(net_475) );
MUX2_X2 inst_674 ( .Z(net_613), .B(net_612), .A(net_355), .S(n4091) );
INV_X1 inst_800 ( .ZN(net_748), .A(n1690) );
NAND2_X1 inst_466 ( .A2(net_178), .ZN(net_176), .A1(n194) );
INV_X1 inst_780 ( .ZN(net_160), .A(n4091) );
MUX2_X2 inst_658 ( .Z(net_560), .B(n861), .A(n822), .S(n1689) );
XOR2_X1 inst_10 ( .Z(net_394), .B(net_285), .A(n389) );
XOR2_X1 inst_4 ( .Z(net_83), .A(n273), .B(n265) );
INV_X1 inst_832 ( .ZN(net_543), .A(net_542) );
NAND2_X1 inst_456 ( .A2(net_181), .ZN(net_166), .A1(n182) );
NAND2_X1 inst_581 ( .ZN(net_749), .A1(net_748), .A2(net_732) );
MUX2_X2 inst_600 ( .Z(net_90), .S(n308), .A(n254), .B(n242) );
XOR2_X1 inst_28 ( .Z(net_573), .A(net_402), .B(net_389) );
NOR2_X1 inst_275 ( .ZN(net_262), .A2(net_97), .A1(n435) );
CLKBUF_X1 inst_858 ( .Z(n889), .A(n299) );
XNOR2_X1 inst_117 ( .ZN(net_694), .A(net_600), .B(net_506) );
NAND2_X1 inst_438 ( .A2(net_160), .ZN(net_67), .A1(n121) );
NAND2_X1 inst_501 ( .ZN(net_220), .A2(net_215), .A1(n185) );
XNOR2_X1 inst_49 ( .ZN(net_298), .A(net_80), .B(net_79) );
NOR3_X1 inst_204 ( .A1(net_756), .ZN(net_459), .A3(net_455), .A2(net_446) );
NAND2_X1 inst_587 ( .ZN(net_791), .A2(net_783), .A1(net_740) );
MUX2_X2 inst_666 ( .A(net_555), .B(net_72), .Z(n877), .S(n4092) );
OR2_X4 inst_154 ( .ZN(net_491), .A2(net_490), .A1(net_449) );
MUX2_X2 inst_592 ( .Z(net_534), .S(n332), .B(n307), .A(n302) );
NAND2_X1 inst_546 ( .ZN(net_447), .A2(net_331), .A1(n4) );
NOR2_X1 inst_324 ( .ZN(net_474), .A2(net_466), .A1(net_465) );
AND2_X2 inst_910 ( .A2(net_753), .ZN(n645), .A1(n137) );
NAND2_X1 inst_465 ( .A2(net_178), .ZN(net_175), .A1(n191) );
MUX2_X2 inst_704 ( .Z(net_684), .B(net_640), .A(net_419), .S(n3717) );
XNOR2_X1 inst_109 ( .ZN(net_608), .B(net_579), .A(net_534) );
XNOR2_X1 inst_54 ( .A(net_364), .ZN(net_333), .B(net_144) );
MUX2_X2 inst_693 ( .S(net_774), .B(net_621), .A(net_68), .Z(n865) );
NAND2_X1 inst_570 ( .A1(net_738), .ZN(net_677), .A2(net_646) );
NAND3_X1 inst_390 ( .A3(net_603), .A1(net_451), .A2(net_307), .ZN(n629) );
MUX2_X2 inst_640 ( .Z(net_144), .B(n372), .A(n369), .S(n332) );
XNOR2_X1 inst_43 ( .ZN(net_402), .B(net_291), .A(n468) );
NAND3_X1 inst_359 ( .ZN(net_118), .A1(n1694), .A3(n1691), .A2(n158) );
INV_X1 inst_765 ( .ZN(net_38), .A(n257) );
NOR2_X1 inst_256 ( .ZN(net_115), .A1(net_53), .A2(n248) );
MUX2_X2 inst_694 ( .S(net_774), .B(net_622), .A(net_63), .Z(n869) );
XNOR2_X1 inst_94 ( .ZN(net_553), .B(net_507), .A(net_408) );
NAND2_X1 inst_454 ( .A2(net_165), .ZN(n656), .A1(n140) );
MUX2_X2 inst_630 ( .Z(net_128), .S(n335), .B(n292), .A(n289) );
NAND3_X1 inst_375 ( .ZN(net_301), .A3(net_165), .A1(n2358), .A2(n23) );
AND2_X2 inst_904 ( .A2(net_681), .ZN(n699), .A1(n137) );
NAND3_X1 inst_401 ( .ZN(net_754), .A1(net_727), .A3(net_176), .A2(net_153) );
NOR2_X1 inst_262 ( .ZN(net_146), .A1(net_126), .A2(n3546) );
NAND2_X1 inst_512 ( .ZN(net_377), .A2(net_291), .A1(n468) );
AND2_X2 inst_908 ( .A2(net_754), .ZN(n685), .A1(n137) );
NAND3_X1 inst_355 ( .ZN(net_112), .A1(n4090), .A3(n4089), .A2(n40) );
NOR2_X1 inst_243 ( .ZN(net_52), .A1(net_48), .A2(n248) );
NOR2_X1 inst_285 ( .ZN(net_277), .A1(net_231), .A2(net_107) );
MUX2_X2 inst_591 ( .Z(net_327), .S(n332), .B(n323), .A(n316) );
NAND2_X1 inst_424 ( .ZN(net_12), .A2(n3552), .A1(n226) );
INV_X1 inst_782 ( .ZN(net_164), .A(n2358) );
NAND2_X1 inst_497 ( .A2(net_215), .ZN(net_214), .A1(n170) );
NOR2_X1 inst_218 ( .ZN(net_17), .A2(n3548), .A1(n265) );
XOR2_X1 inst_15 ( .Z(net_359), .B(net_290), .A(n503) );
INV_X1 inst_757 ( .ZN(net_740), .A(n4087) );
MUX2_X2 inst_647 ( .Z(net_435), .B(net_7), .S(n514), .A(n3546) );
NAND4_X1 inst_343 ( .ZN(net_401), .A2(net_399), .A3(net_398), .A4(net_320), .A1(net_308) );
XOR2_X1 inst_6 ( .Z(net_85), .A(n289), .B(n281) );
NOR3_X1 inst_194 ( .ZN(net_241), .A1(net_56), .A3(net_36), .A2(n523) );
NAND2_X1 inst_543 ( .ZN(net_452), .A1(net_394), .A2(net_358) );
NOR2_X1 inst_337 ( .A2(net_541), .ZN(net_539), .A1(net_503) );
INV_X1 inst_787 ( .ZN(net_53), .A(n234) );
INV_X1 inst_825 ( .ZN(net_376), .A(net_375) );
INV_X1 inst_833 ( .ZN(net_591), .A(net_590) );
MUX2_X2 inst_670 ( .Z(net_643), .S(net_607), .A(net_549), .B(net_535) );
XNOR2_X1 inst_123 ( .ZN(net_668), .A(net_625), .B(net_583) );
NAND2_X1 inst_509 ( .A2(net_290), .ZN(net_258), .A1(n503) );
NOR2_X1 inst_299 ( .ZN(net_344), .A2(net_262), .A1(net_234) );
MUX2_X2 inst_699 ( .Z(net_673), .A(net_672), .B(net_671), .S(n1691) );
CLKBUF_X1 inst_864 ( .A(n604), .Z(n594) );
NAND3_X1 inst_418 ( .A3(net_791), .A2(net_207), .A1(net_138), .ZN(n767) );
NAND2_X1 inst_476 ( .A2(net_194), .ZN(net_189), .A1(n46) );
XNOR2_X1 inst_118 ( .A(net_636), .B(net_390), .ZN(n813) );
XNOR2_X1 inst_86 ( .ZN(net_606), .A(net_602), .B(net_494) );
OR2_X4 inst_153 ( .ZN(net_489), .A1(net_488), .A2(net_445) );
XOR2_X1 inst_20 ( .Z(net_323), .A(net_288), .B(net_286) );
NAND2_X1 inst_442 ( .A2(net_160), .ZN(net_73), .A1(n116) );
MUX2_X2 inst_613 ( .Z(net_108), .B(n3552), .A(n3550), .S(n281) );
XOR2_X1 inst_38 ( .A(net_578), .Z(net_550), .B(net_549) );
MUX2_X2 inst_714 ( .A(net_700), .B(net_699), .Z(net_698), .S(n4088) );
NAND3_X1 inst_381 ( .ZN(net_440), .A2(net_439), .A3(net_438), .A1(net_382) );
MUX2_X2 inst_726 ( .A(net_717), .B(net_716), .Z(net_715), .S(n1689) );
NOR2_X1 inst_295 ( .ZN(net_508), .A1(net_275), .A2(net_247) );
NAND4_X1 inst_349 ( .ZN(net_667), .A4(net_633), .A1(net_554), .A2(net_543), .A3(net_480) );
NAND2_X1 inst_483 ( .ZN(net_198), .A2(net_197), .A1(n91) );
NAND2_X1 inst_576 ( .ZN(net_741), .A1(net_740), .A2(net_698) );
AND2_X4 inst_883 ( .ZN(net_342), .A2(net_325), .A1(n479) );
NOR3_X1 inst_209 ( .ZN(net_565), .A1(net_523), .A3(net_370), .A2(net_368) );
NOR2_X1 inst_259 ( .A1(net_164), .ZN(net_139), .A2(n34) );
XOR2_X1 inst_40 ( .Z(net_590), .A(net_575), .B(net_574) );
NOR2_X1 inst_320 ( .ZN(net_427), .A2(net_425), .A1(net_389) );
OR2_X2 inst_167 ( .ZN(net_654), .A2(net_615), .A1(n1694) );
MUX2_X2 inst_607 ( .Z(net_99), .S(n281), .A(n254), .B(n242) );
NOR2_X1 inst_246 ( .ZN(net_61), .A1(net_46), .A2(n248) );
INV_X1 inst_756 ( .ZN(net_223), .A(n457) );
MUX2_X2 inst_635 ( .Z(net_133), .S(n4088), .B(n103), .A(n100) );
INV_X1 inst_807 ( .A(net_534), .ZN(net_343) );
XNOR2_X1 inst_95 ( .ZN(net_567), .B(net_529), .A(net_488) );
MUX2_X2 inst_705 ( .A(net_641), .B(net_73), .Z(n828), .S(n4092) );
XOR2_X1 inst_1 ( .Z(net_80), .A(n316), .B(n308) );
AND2_X2 inst_911 ( .A2(net_761), .ZN(n682), .A1(n137) );
XNOR2_X1 inst_72 ( .B(net_605), .ZN(net_497), .A(net_490) );
NAND2_X1 inst_519 ( .A2(net_312), .ZN(net_308), .A1(n26) );
NAND2_X1 inst_439 ( .A2(net_160), .ZN(net_68), .A1(n114) );
AND2_X2 inst_909 ( .A2(net_752), .ZN(n651), .A1(n137) );
NOR2_X1 inst_331 ( .A2(net_517), .ZN(net_516), .A1(net_476) );
NAND2_X1 inst_582 ( .ZN(net_751), .A1(net_750), .A2(net_733) );
MUX2_X2 inst_735 ( .A(net_714), .B(net_154), .Z(n777), .S(n4090) );
MUX2_X2 inst_683 ( .Z(net_627), .B(net_626), .A(net_508), .S(n4091) );
XNOR2_X1 inst_115 ( .ZN(net_631), .A(net_630), .B(net_598) );
NOR2_X1 inst_235 ( .ZN(net_39), .A1(net_38), .A2(n3546) );
INV_X1 inst_750 ( .ZN(net_55), .A(n341) );
NOR3_X1 inst_210 ( .ZN(net_603), .A2(net_602), .A1(net_576), .A3(net_379) );
NOR2_X1 inst_317 ( .ZN(net_464), .A1(net_454), .A2(net_426) );
AND2_X2 inst_894 ( .ZN(n810), .A2(n145), .A1(n141) );
MUX2_X2 inst_667 ( .Z(net_619), .S(net_574), .A(net_571), .B(net_548) );
NOR2_X1 inst_278 ( .ZN(net_267), .A2(net_93), .A1(n400) );
NAND2_X1 inst_467 ( .A2(net_178), .ZN(net_177), .A1(n197) );
INV_X1 inst_761 ( .ZN(net_774), .A(n4092) );
NOR2_X1 inst_239 ( .A1(net_738), .ZN(net_197), .A2(n4089) );
XNOR2_X1 inst_105 ( .ZN(net_598), .B(net_567), .A(net_565) );
NAND2_X1 inst_488 ( .ZN(net_204), .A2(net_203), .A1(n49) );
NAND3_X1 inst_387 ( .A3(net_593), .A2(net_209), .A1(net_137), .ZN(n722) );
MUX2_X2 inst_725 ( .A(net_717), .B(net_716), .Z(net_714), .S(n4089) );
MUX2_X2 inst_593 ( .Z(net_42), .S(n324), .A(n254), .B(n242) );
OR2_X2 inst_175 ( .ZN(net_726), .A2(net_703), .A1(n1690) );
CLKBUF_X1 inst_857 ( .Z(n892), .A(n549) );
MUX2_X2 inst_747 ( .A(net_786), .B(net_785), .Z(net_784), .S(n1689) );
NOR2_X1 inst_254 ( .A2(n850), .A1(n849), .ZN(n601) );
INV_X1 inst_843 ( .A(net_699), .ZN(n871) );
MUX2_X2 inst_654 ( .Z(net_555), .B(net_554), .A(net_439), .S(n4091) );
MUX2_X2 inst_625 ( .Z(net_285), .S(n335), .B(n264), .A(n257) );
NOR2_X1 inst_225 ( .ZN(net_27), .A2(n3548), .A1(n234) );
MUX2_X2 inst_601 ( .Z(net_91), .A(n254), .B(n242), .S(n218) );
XNOR2_X1 inst_133 ( .ZN(net_757), .B(net_756), .A(net_730) );
NAND2_X1 inst_508 ( .ZN(net_309), .A2(net_288), .A1(n523) );
NAND2_X1 inst_568 ( .A1(net_774), .ZN(net_635), .A2(net_613) );
XNOR2_X1 inst_112 ( .ZN(net_661), .A(net_606), .B(net_597) );
NAND2_X1 inst_523 ( .A2(net_364), .ZN(net_349), .A1(n54) );
AND2_X2 inst_916 ( .A2(net_765), .ZN(n688), .A1(n137) );
NAND3_X1 inst_365 ( .ZN(net_138), .A1(net_136), .A3(n4087), .A2(n14) );
INV_X1 inst_764 ( .ZN(net_126), .A(n210) );
XNOR2_X1 inst_67 ( .ZN(net_433), .B(net_371), .A(net_344) );
NOR4_X1 inst_181 ( .ZN(net_633), .A2(net_626), .A4(net_612), .A3(net_590), .A1(net_588) );
NOR2_X1 inst_305 ( .A2(net_547), .ZN(net_367), .A1(net_366) );
NAND2_X1 inst_479 ( .A2(net_194), .ZN(net_192), .A1(n76) );
XOR2_X1 inst_29 ( .B(net_510), .Z(net_409), .A(net_338) );
INV_X1 inst_771 ( .ZN(n612), .A(n358) );
NAND3_X1 inst_391 ( .ZN(net_675), .A1(net_654), .A3(net_171), .A2(net_118) );
MUX2_X2 inst_661 ( .Z(net_610), .S(net_574), .B(net_569), .A(net_505) );
NAND2_X1 inst_590 ( .A2(net_793), .ZN(n658), .A1(n137) );
AND2_X4 inst_878 ( .A2(net_160), .ZN(net_140), .A1(n127) );
MUX2_X2 inst_713 ( .A(net_700), .B(net_699), .Z(net_697), .S(n4089) );
NOR3_X1 inst_202 ( .A1(net_630), .ZN(net_461), .A2(net_455), .A3(net_452) );
XNOR2_X1 inst_126 ( .ZN(net_687), .A(net_679), .B(net_660) );
NAND2_X1 inst_480 ( .A2(net_194), .ZN(net_193), .A1(n43) );
MUX2_X2 inst_634 ( .Z(net_132), .S(n1691), .A(n149), .B(n146) );
NAND3_X1 inst_419 ( .ZN(net_793), .A3(net_792), .A2(net_213), .A1(net_167) );
NAND2_X1 inst_477 ( .A2(net_197), .ZN(net_190), .A1(n46) );
MUX2_X2 inst_646 ( .Z(net_416), .B(net_6), .A(net_1), .S(n293) );
NAND2_X1 inst_564 ( .ZN(net_563), .A2(net_562), .A1(net_444) );
NAND2_X1 inst_538 ( .A2(net_441), .ZN(net_426), .A1(net_358) );
NAND2_X1 inst_423 ( .ZN(net_11), .A2(n4115), .A1(n135) );
MUX2_X2 inst_739 ( .Z(net_768), .B(net_766), .A(net_757), .S(n1497) );
XOR2_X1 inst_35 ( .Z(net_533), .A(net_532), .B(net_531) );
NAND3_X1 inst_382 ( .A2(net_469), .ZN(net_467), .A3(net_443), .A1(net_373) );
AND2_X2 inst_907 ( .A2(net_690), .ZN(n670), .A1(n137) );
INV_X1 inst_835 ( .A(net_648), .ZN(n875) );
XNOR2_X1 inst_48 ( .ZN(net_297), .A(net_43), .B(n324) );
NAND3_X1 inst_358 ( .ZN(net_117), .A1(n4090), .A3(n4089), .A2(n37) );
XNOR2_X1 inst_46 ( .ZN(net_294), .B(net_82), .A(net_81) );
XNOR2_X1 inst_136 ( .ZN(net_769), .B(net_767), .A(net_747) );
XOR2_X1 inst_30 ( .A(net_415), .B(net_414), .Z(net_410) );
NOR2_X1 inst_330 ( .A1(net_656), .ZN(net_514), .A2(net_474) );
MUX2_X2 inst_610 ( .Z(net_105), .A(n3548), .B(n3546), .S(n226) );
NOR2_X1 inst_233 ( .A2(net_738), .ZN(net_203), .A1(net_155) );
MUX2_X2 inst_710 ( .Z(net_690), .A(net_674), .B(net_130), .S(n1690) );
OR2_X2 inst_165 ( .ZN(net_652), .A2(net_617), .A1(n4090) );
INV_X1 inst_796 ( .ZN(net_77), .A(n273) );
NOR2_X1 inst_271 ( .ZN(net_255), .A2(net_89), .A1(n534) );
NAND2_X1 inst_443 ( .A2(net_160), .ZN(net_74), .A1(n130) );
MUX2_X2 inst_633 ( .Z(net_131), .S(n1691), .A(n155), .B(n152) );
XOR2_X1 inst_34 ( .A(net_679), .Z(net_554), .B(net_448) );
XOR2_X1 inst_12 ( .Z(net_441), .B(net_287), .A(n400) );
NAND2_X1 inst_529 ( .ZN(net_353), .A2(net_304), .A1(net_251) );
NAND2_X1 inst_524 ( .A2(net_318), .ZN(net_317), .A1(n80) );
XNOR2_X1 inst_56 ( .B(net_602), .A(net_343), .ZN(net_337) );
XNOR2_X1 inst_71 ( .ZN(net_479), .B(net_385), .A(net_326) );
MUX2_X2 inst_655 ( .Z(net_557), .B(n861), .A(n822), .S(n4089) );
NOR2_X1 inst_308 ( .A2(net_583), .A1(net_469), .ZN(net_468) );
XNOR2_X1 inst_104 ( .B(net_691), .ZN(net_626), .A(net_566) );
NAND2_X1 inst_448 ( .ZN(net_135), .A2(net_57), .A1(n254) );
XNOR2_X1 inst_60 ( .ZN(net_387), .B(net_297), .A(net_84) );
NAND2_X1 inst_455 ( .A2(net_165), .ZN(n820), .A1(n83) );
OR2_X2 inst_168 ( .ZN(net_655), .A2(net_616), .A1(n1690) );
AND2_X2 inst_914 ( .A2(net_760), .ZN(n648), .A1(n137) );
MUX2_X2 inst_695 ( .Z(net_658), .A(net_416), .B(n623), .S(n4091) );
MUX2_X2 inst_730 ( .A(net_735), .B(net_734), .Z(net_732), .S(n1689) );
AND3_X2 inst_873 ( .A2(net_530), .A1(net_511), .A3(net_356), .ZN(n610) );
MUX2_X2 inst_727 ( .Z(net_718), .A(net_717), .B(net_716), .S(n4088) );
MUX2_X2 inst_675 ( .Z(net_615), .B(n877), .A(n838), .S(n1691) );
NAND3_X1 inst_384 ( .ZN(net_521), .A1(net_429), .A3(net_378), .A2(net_366) );
INV_X1 inst_758 ( .ZN(net_0), .A(n136) );
NOR2_X1 inst_321 ( .ZN(net_486), .A2(net_450), .A1(net_342) );
NAND2_X1 inst_496 ( .A2(net_215), .ZN(net_213), .A1(n179) );
MUX2_X2 inst_653 ( .S(net_774), .B(net_481), .A(net_104), .Z(n861) );
CLKBUF_X1 inst_860 ( .A(n717), .Z(n704) );
MUX2_X2 inst_608 ( .Z(net_100), .S(n273), .A(n254), .B(n242) );
NOR2_X1 inst_336 ( .A1(net_526), .A2(net_484), .ZN(n615) );
AND2_X4 inst_882 ( .ZN(net_393), .A2(net_287), .A1(n400) );
INV_X1 inst_834 ( .A(net_636), .ZN(n623) );
NAND2_X1 inst_563 ( .A2(net_562), .ZN(net_561), .A1(net_458) );
NAND2_X1 inst_583 ( .ZN(net_775), .A1(net_774), .A2(net_772) );
NAND2_X1 inst_580 ( .A1(net_750), .ZN(net_746), .A2(net_719) );
OR2_X2 inst_170 ( .ZN(net_721), .A2(net_709), .A1(n4090) );
NOR2_X1 inst_258 ( .ZN(net_127), .A1(net_126), .A2(n248) );
NAND3_X1 inst_376 ( .ZN(net_302), .A3(net_142), .A1(net_18), .A2(n411) );
NOR3_X1 inst_199 ( .ZN(net_246), .A1(net_47), .A3(net_31), .A2(n468) );
XOR2_X1 inst_41 ( .Z(net_628), .A(net_605), .B(net_561) );
NAND2_X1 inst_511 ( .ZN(net_383), .A2(net_327), .A1(n490) );
OR3_X2 inst_143 ( .A1(net_139), .A3(net_24), .A2(n809), .ZN(n717) );
MUX2_X2 inst_708 ( .A(net_658), .B(net_70), .Z(n824), .S(n4092) );
OR2_X4 inst_152 ( .ZN(net_471), .A1(net_470), .A2(net_403) );
NOR2_X1 inst_265 ( .ZN(net_360), .A2(net_295), .A1(net_158) );
NAND2_X1 inst_482 ( .A2(net_197), .ZN(net_196), .A1(n76) );
NAND2_X1 inst_468 ( .ZN(net_179), .A2(net_178), .A1(n203) );
MUX2_X2 inst_682 ( .Z(net_622), .B(net_591), .A(net_530), .S(n4091) );
MUX2_X2 inst_736 ( .A(net_736), .B(net_113), .Z(n727), .S(n4087) );
NAND2_X1 inst_544 ( .ZN(net_371), .A2(net_306), .A1(net_264) );
NOR2_X1 inst_238 ( .ZN(net_47), .A1(net_46), .A2(n3546) );
NAND2_X1 inst_540 ( .A1(net_469), .ZN(net_362), .A2(net_357) );
NAND2_X1 inst_539 ( .ZN(net_361), .A1(net_360), .A2(net_359) );
NAND2_X1 inst_429 ( .ZN(net_30), .A2(n341), .A1(n242) );
MUX2_X2 inst_724 ( .Z(net_710), .B(n869), .A(n830), .S(n4088) );
NAND3_X1 inst_404 ( .A3(net_723), .A2(net_204), .A1(net_190), .ZN(n772) );
AND2_X2 inst_895 ( .A2(net_397), .ZN(n707), .A1(n141) );
NOR4_X1 inst_178 ( .ZN(net_511), .A1(net_510), .A2(net_509), .A3(net_508), .A4(net_440) );
XNOR2_X1 inst_89 ( .ZN(net_538), .B(net_498), .A(net_432) );
XNOR2_X1 inst_111 ( .ZN(net_638), .B(net_607), .A(net_578) );
XNOR2_X1 inst_66 ( .ZN(net_413), .B(net_337), .A(net_328) );
NAND3_X1 inst_388 ( .ZN(net_623), .A3(net_594), .A2(net_212), .A1(net_172) );
MUX2_X2 inst_734 ( .A(net_718), .B(net_133), .Z(n737), .S(n4087) );
XOR2_X1 inst_7 ( .Z(net_147), .A(n257), .B(n234) );
NOR4_X1 inst_182 ( .ZN(net_683), .A4(net_639), .A2(net_581), .A1(net_512), .A3(net_334) );
NAND3_X1 inst_392 ( .ZN(net_676), .A1(net_655), .A3(net_183), .A2(net_40) );
XNOR2_X1 inst_120 ( .ZN(net_657), .A(net_656), .B(net_609) );
NOR2_X1 inst_273 ( .A2(net_293), .ZN(net_260), .A1(n422) );
INV_X1 inst_788 ( .ZN(net_101), .A(n265) );
NOR2_X1 inst_294 ( .ZN(net_381), .A1(net_270), .A2(net_243) );
NOR2_X1 inst_222 ( .ZN(net_24), .A2(n88), .A1(n2358) );
NOR2_X1 inst_284 ( .ZN(net_276), .A1(net_223), .A2(net_148) );
NAND2_X1 inst_489 ( .A2(net_208), .ZN(net_205), .A1(n49) );
INV_X1 inst_806 ( .A(net_602), .ZN(net_163) );
NOR3_X1 inst_192 ( .ZN(net_238), .A1(net_66), .A3(net_22), .A2(net_2) );
NOR2_X1 inst_280 ( .ZN(net_270), .A1(net_235), .A2(net_106) );
INV_X1 inst_763 ( .ZN(n600), .A(n366) );
NAND3_X1 inst_366 ( .ZN(net_143), .A1(n4088), .A3(n4087), .A2(n20) );
NAND4_X1 inst_346 ( .ZN(net_502), .A4(net_460), .A2(net_441), .A1(net_394), .A3(net_392) );
NAND2_X1 inst_491 ( .A2(net_208), .ZN(net_207), .A1(n64) );
NAND2_X1 inst_567 ( .A2(net_662), .ZN(net_607), .A1(net_522) );
NOR3_X1 inst_193 ( .ZN(net_240), .A1(net_49), .A3(net_20), .A2(n534) );
OR2_X4 inst_149 ( .ZN(net_503), .A2(net_425), .A1(net_423) );
INV_X1 inst_810 ( .ZN(net_679), .A(net_358) );
NOR2_X1 inst_318 ( .ZN(net_466), .A2(net_457), .A1(net_364) );
XOR2_X1 inst_39 ( .A(net_575), .Z(net_572), .B(net_571) );
NOR2_X1 inst_230 ( .ZN(net_34), .A2(n251), .A1(n210) );
CLKBUF_X1 inst_856 ( .Z(n921), .A(n1) );
INV_X1 inst_842 ( .ZN(net_734), .A(n863) );

endmodule
