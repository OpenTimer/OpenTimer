module c3540 (
n317,
n179,
n223,
n329,
n238,
n169,
n143,
n190,
n257,
n311,
n1698,
n213,
n283,
n68,
n58,
n244,
n322,
n41,
n20,
n97,
n274,
n232,
n77,
n326,
n1,
n107,
n128,
n50,
n125,
n330,
n132,
n45,
n116,
n159,
n226,
n250,
n150,
n270,
n294,
n264,
n222,
n87,
n343,
n2897,
n33,
n303,
n13,
n200,
n137,
n124,
n399,
n361,
n369,
n364,
n407,
n367,
n409,
n384,
n351,
n372,
n375,
n358,
n387,
n381,
n390,
n355,
n393,
n378,
n402,
n405,
n396,
n353);

// Start PIs
input n317;
input n179;
input n223;
input n329;
input n238;
input n169;
input n143;
input n190;
input n257;
input n311;
input n1698;
input n213;
input n283;
input n68;
input n58;
input n244;
input n322;
input n41;
input n20;
input n97;
input n274;
input n232;
input n77;
input n326;
input n1;
input n107;
input n128;
input n50;
input n125;
input n330;
input n132;
input n45;
input n116;
input n159;
input n226;
input n250;
input n150;
input n270;
input n294;
input n264;
input n222;
input n87;
input n343;
input n2897;
input n33;
input n303;
input n13;
input n200;
input n137;
input n124;

// Start POs
output n399;
output n361;
output n369;
output n364;
output n407;
output n367;
output n409;
output n384;
output n351;
output n372;
output n375;
output n358;
output n387;
output n381;
output n390;
output n355;
output n393;
output n378;
output n402;
output n405;
output n396;
output n353;

// Start wires
wire net_568;
wire net_47;
wire net_416;
wire net_215;
wire net_54;
wire net_526;
wire net_429;
wire net_557;
wire net_129;
wire net_648;
wire net_373;
wire net_119;
wire net_98;
wire net_151;
wire net_356;
wire net_53;
wire net_452;
wire net_210;
wire net_545;
wire net_284;
wire net_168;
wire net_560;
wire net_477;
wire net_439;
wire net_385;
wire net_259;
wire net_269;
wire net_548;
wire net_469;
wire net_501;
wire net_187;
wire net_111;
wire net_264;
wire net_90;
wire net_225;
wire n116;
wire net_283;
wire n150;
wire net_636;
wire net_85;
wire net_263;
wire net_252;
wire net_124;
wire net_343;
wire net_404;
wire net_240;
wire net_160;
wire net_322;
wire n378;
wire net_511;
wire net_4;
wire n124;
wire net_420;
wire net_665;
wire net_447;
wire net_295;
wire net_410;
wire net_508;
wire net_390;
wire net_307;
wire net_35;
wire net_586;
wire net_344;
wire net_16;
wire net_239;
wire net_193;
wire net_257;
wire net_310;
wire net_233;
wire net_474;
wire net_120;
wire net_292;
wire net_201;
wire net_472;
wire net_109;
wire net_80;
wire net_65;
wire net_96;
wire net_484;
wire net_167;
wire net_207;
wire net_136;
wire net_651;
wire net_280;
wire net_126;
wire n159;
wire net_495;
wire net_278;
wire net_34;
wire net_458;
wire net_108;
wire net_598;
wire n390;
wire n87;
wire net_571;
wire n303;
wire net_63;
wire net_593;
wire net_617;
wire net_601;
wire net_274;
wire net_554;
wire net_425;
wire net_321;
wire net_287;
wire net_189;
wire net_490;
wire net_99;
wire net_46;
wire net_480;
wire net_216;
wire net_433;
wire net_584;
wire n355;
wire net_544;
wire net_368;
wire net_224;
wire net_632;
wire net_52;
wire net_538;
wire net_165;
wire net_608;
wire net_510;
wire net_370;
wire net_464;
wire net_366;
wire net_13;
wire net_413;
wire net_446;
wire net_114;
wire n343;
wire net_248;
wire net_384;
wire net_36;
wire net_198;
wire net_637;
wire net_253;
wire net_311;
wire net_276;
wire net_494;
wire net_209;
wire net_3;
wire net_547;
wire net_634;
wire net_294;
wire net_154;
wire net_666;
wire n257;
wire net_507;
wire net_616;
wire net_371;
wire net_238;
wire net_529;
wire net_28;
wire n58;
wire net_587;
wire net_485;
wire net_97;
wire n364;
wire net_192;
wire net_649;
wire net_503;
wire net_256;
wire net_460;
wire net_82;
wire net_650;
wire net_64;
wire net_457;
wire net_291;
wire n250;
wire net_121;
wire net_597;
wire net_200;
wire net_308;
wire net_75;
wire net_515;
wire net_600;
wire net_396;
wire n200;
wire net_206;
wire net_195;
wire net_125;
wire net_397;
wire net_107;
wire net_166;
wire net_223;
wire net_235;
wire net_530;
wire n351;
wire net_606;
wire net_623;
wire net_663;
wire net_603;
wire net_594;
wire net_320;
wire net_271;
wire net_23;
wire net_117;
wire net_74;
wire net_642;
wire net_579;
wire net_401;
wire net_250;
wire net_205;
wire net_242;
wire net_312;
wire net_130;
wire net_572;
wire net_359;
wire net_440;
wire net_286;
wire net_147;
wire net_481;
wire net_369;
wire n367;
wire net_470;
wire net_26;
wire net_403;
wire net_334;
wire net_32;
wire net_430;
wire n330;
wire net_365;
wire net_282;
wire net_645;
wire net_426;
wire net_380;
wire net_141;
wire net_467;
wire net_83;
wire net_609;
wire net_541;
wire net_414;
wire net_372;
wire n407;
wire net_437;
wire net_528;
wire net_56;
wire net_566;
wire net_456;
wire net_155;
wire net_335;
wire net_506;
wire net_181;
wire net_336;
wire n381;
wire net_624;
wire net_349;
wire net_39;
wire net_555;
wire net_245;
wire net_2;
wire n283;
wire net_9;
wire net_395;
wire net_331;
wire net_298;
wire net_493;
wire net_475;
wire net_563;
wire net_386;
wire net_641;
wire net_605;
wire net_277;
wire net_199;
wire n107;
wire n50;
wire net_502;
wire net_431;
wire net_89;
wire n45;
wire n387;
wire net_290;
wire net_338;
wire n137;
wire net_638;
wire net_243;
wire net_400;
wire n399;
wire n179;
wire net_222;
wire net_602;
wire net_313;
wire n329;
wire net_152;
wire net_489;
wire net_175;
wire net_657;
wire net_106;
wire net_607;
wire net_258;
wire net_140;
wire net_247;
wire net_329;
wire net_279;
wire net_148;
wire n1698;
wire net_419;
wire net_25;
wire net_70;
wire net_251;
wire net_194;
wire net_615;
wire n369;
wire net_478;
wire net_244;
wire net_664;
wire net_585;
wire net_441;
wire net_128;
wire net_596;
wire net_138;
wire net_333;
wire net_639;
wire net_549;
wire net_374;
wire net_411;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_214;
wire net_77;
wire net_249;
wire net_20;
wire net_49;
wire net_518;
wire net_15;
wire net_57;
wire net_71;
wire net_156;
wire net_394;
wire net_1;
wire net_92;
wire net_112;
wire net_139;
wire net_551;
wire net_537;
wire net_332;
wire net_180;
wire net_409;
wire n68;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire net_492;
wire net_463;
wire net_656;
wire net_432;
wire net_88;
wire net_197;
wire n77;
wire net_513;
wire net_204;
wire net_81;
wire net_232;
wire net_604;
wire net_163;
wire net_402;
wire net_67;
wire net_202;
wire net_268;
wire n270;
wire net_110;
wire net_379;
wire net_459;
wire net_483;
wire net_48;
wire net_33;
wire net_8;
wire net_203;
wire net_450;
wire net_289;
wire net_505;
wire net_621;
wire net_435;
wire net_176;
wire net_137;
wire net_296;
wire net_132;
wire net_613;
wire net_237;
wire net_105;
wire net_614;
wire net_532;
wire net_12;
wire net_93;
wire net_578;
wire net_302;
wire net_569;
wire net_127;
wire net_327;
wire net_357;
wire net_348;
wire n1;
wire net_630;
wire n128;
wire net_76;
wire net_626;
wire net_101;
wire net_388;
wire net_326;
wire net_353;
wire net_589;
wire net_519;
wire net_100;
wire net_412;
wire net_655;
wire net_652;
wire net_536;
wire net_455;
wire net_221;
wire net_115;
wire net_393;
wire net_442;
wire net_17;
wire net_319;
wire n361;
wire net_542;
wire net_453;
wire net_575;
wire net_595;
wire net_581;
wire n223;
wire net_378;
wire net_164;
wire net_408;
wire net_377;
wire net_87;
wire net_0;
wire net_288;
wire net_423;
wire net_658;
wire n143;
wire n190;
wire net_328;
wire net_157;
wire net_540;
wire net_512;
wire net_42;
wire net_662;
wire net_50;
wire n97;
wire net_234;
wire net_38;
wire net_66;
wire net_466;
wire n409;
wire net_342;
wire net_612;
wire net_19;
wire net_443;
wire net_504;
wire net_522;
wire net_270;
wire net_183;
wire net_668;
wire net_618;
wire net_150;
wire n405;
wire net_303;
wire net_304;
wire net_352;
wire net_491;
wire n238;
wire net_644;
wire net_30;
wire net_643;
wire n375;
wire net_436;
wire net_24;
wire net_392;
wire net_622;
wire net_186;
wire net_118;
wire net_421;
wire net_146;
wire net_550;
wire net_122;
wire net_417;
wire net_7;
wire net_172;
wire n384;
wire net_428;
wire net_461;
wire net_94;
wire net_246;
wire n132;
wire net_219;
wire net_640;
wire net_18;
wire net_482;
wire n294;
wire net_309;
wire net_659;
wire n222;
wire net_131;
wire n2897;
wire net_196;
wire net_29;
wire net_358;
wire net_142;
wire net_149;
wire net_516;
wire net_654;
wire net_31;
wire net_387;
wire net_330;
wire net_535;
wire net_498;
wire net_158;
wire net_41;
wire net_577;
wire net_360;
wire net_570;
wire net_525;
wire net_444;
wire net_213;
wire net_325;
wire net_301;
wire net_260;
wire net_299;
wire net_438;
wire n322;
wire net_580;
wire net_314;
wire net_182;
wire net_521;
wire net_60;
wire net_590;
wire net_337;
wire net_341;
wire net_267;
wire net_273;
wire net_424;
wire net_468;
wire net_58;
wire net_576;
wire net_488;
wire net_73;
wire net_465;
wire net_86;
wire net_177;
wire net_523;
wire n13;
wire net_476;
wire net_407;
wire net_564;
wire net_382;
wire net_179;
wire net_159;
wire net_61;
wire net_583;
wire net_449;
wire net_383;
wire net_62;
wire net_6;
wire net_553;
wire net_534;
wire net_217;
wire net_351;
wire n311;
wire n213;
wire net_427;
wire net_486;
wire net_135;
wire net_340;
wire net_265;
wire net_517;
wire net_628;
wire net_434;
wire net_473;
wire net_406;
wire net_14;
wire net_220;
wire net_633;
wire net_293;
wire net_324;
wire net_113;
wire net_497;
wire net_454;
wire net_462;
wire net_418;
wire net_40;
wire n226;
wire net_69;
wire net_543;
wire n264;
wire net_161;
wire net_625;
wire net_300;
wire net_339;
wire net_95;
wire net_173;
wire n317;
wire net_361;
wire net_78;
wire net_27;
wire net_317;
wire net_305;
wire n372;
wire net_514;
wire net_191;
wire net_261;
wire net_22;
wire net_376;
wire net_558;
wire net_354;
wire net_660;
wire net_524;
wire net_144;
wire net_102;
wire net_227;
wire net_59;
wire net_646;
wire net_363;
wire n244;
wire net_445;
wire net_573;
wire n396;
wire net_162;
wire n20;
wire net_44;
wire net_230;
wire net_653;
wire n232;
wire net_520;
wire n326;
wire net_422;
wire net_134;
wire net_546;
wire net_561;
wire net_567;
wire net_45;
wire net_381;
wire net_591;
wire net_185;
wire net_588;
wire net_272;
wire net_178;
wire net_667;
wire n393;
wire n402;
wire net_208;
wire net_236;
wire net_487;
wire net_212;
wire net_315;
wire net_552;
wire net_415;
wire net_116;
wire net_556;
wire net_347;
wire net_91;
wire n169;
wire net_297;
wire net_346;
wire net_629;
wire net_55;
wire net_559;
wire net_635;
wire net_255;
wire net_266;
wire net_345;
wire net_104;
wire net_620;
wire net_448;
wire net_619;
wire net_72;
wire net_350;
wire net_229;
wire net_398;
wire net_627;
wire net_306;
wire net_241;
wire net_5;
wire net_405;
wire net_500;
wire net_355;
wire net_184;
wire net_599;
wire net_631;
wire net_11;
wire net_610;
wire net_123;
wire net_527;
wire net_262;
wire net_362;
wire net_389;
wire net_68;
wire net_318;
wire net_451;
wire net_323;
wire net_275;
wire net_539;
wire net_399;
wire net_153;
wire net_316;
wire net_84;
wire net_218;
wire net_174;
wire net_611;
wire net_231;
wire net_562;
wire net_103;
wire net_375;
wire net_226;
wire net_364;
wire net_43;
wire net_10;
wire net_228;
wire net_592;
wire net_21;
wire net_647;
wire net_79;
wire n41;
wire net_143;
wire net_190;
wire n274;
wire net_391;
wire net_533;
wire net_145;
wire net_285;
wire net_281;
wire n125;
wire net_254;
wire net_37;
wire net_582;
wire n358;
wire net_188;
wire net_496;
wire net_509;
wire net_574;
wire net_479;
wire net_661;
wire net_211;
wire net_133;
wire n33;
wire n353;

// Start cells
NAND2_X1 inst_537 ( .ZN(net_456), .A1(net_455), .A2(net_423) );
NAND2_X1 inst_481 ( .A1(net_350), .ZN(net_279), .A2(net_278) );
NAND2_X1 inst_551 ( .ZN(net_493), .A1(net_451), .A2(net_427) );
NAND3_X1 inst_228 ( .ZN(net_141), .A1(net_94), .A3(net_63), .A2(net_16) );
NOR2_X1 inst_125 ( .ZN(net_125), .A1(net_73), .A2(net_53) );
NAND2_X1 inst_486 ( .A2(net_305), .ZN(net_287), .A1(n68) );
NAND2_X1 inst_506 ( .A2(net_324), .ZN(net_323), .A1(net_296) );
NAND2_X1 inst_495 ( .ZN(net_306), .A2(net_305), .A1(n303) );
NAND2_X1 inst_353 ( .A2(net_97), .ZN(net_93), .A1(n238) );
NAND4_X1 inst_207 ( .ZN(net_544), .A2(net_526), .A1(net_525), .A4(net_522), .A3(net_519) );
NOR2_X1 inst_159 ( .ZN(net_478), .A1(net_477), .A2(net_436) );
NAND2_X1 inst_395 ( .A2(net_165), .ZN(net_158), .A1(n326) );
NOR2_X1 inst_134 ( .ZN(net_280), .A1(net_111), .A2(net_108) );
NAND3_X1 inst_244 ( .ZN(net_395), .A2(net_373), .A3(net_316), .A1(net_237) );
NAND2_X1 inst_333 ( .A2(net_61), .ZN(net_60), .A1(n232) );
NAND2_X1 inst_452 ( .ZN(net_236), .A2(net_235), .A1(n264) );
AND2_X4 inst_689 ( .ZN(net_603), .A2(net_588), .A1(net_587) );
NAND2_X1 inst_430 ( .A2(net_265), .ZN(net_209), .A1(n283) );
NOR2_X1 inst_131 ( .ZN(net_168), .A1(net_111), .A2(net_89) );
NAND2_X1 inst_406 ( .A2(net_254), .ZN(net_178), .A1(n159) );
NAND4_X1 inst_214 ( .A1(net_574), .ZN(net_566), .A4(net_536), .A2(net_509), .A3(net_457) );
NAND2_X1 inst_462 ( .A2(net_283), .ZN(net_247), .A1(n322) );
NOR2_X1 inst_160 ( .ZN(net_480), .A1(net_479), .A2(net_437) );
NAND2_X1 inst_328 ( .A2(net_549), .ZN(net_76), .A1(net_73) );
XNOR2_X1 inst_47 ( .ZN(net_664), .A(net_657), .B(net_655) );
XNOR2_X1 inst_19 ( .ZN(net_278), .A(net_91), .B(net_47) );
NAND2_X1 inst_548 ( .ZN(net_490), .A1(net_453), .A2(net_440) );
NAND2_X1 inst_515 ( .ZN(net_347), .A1(net_333), .A2(net_308) );
XOR2_X1 inst_8 ( .Z(net_666), .B(net_664), .A(net_663) );
NAND2_X1 inst_370 ( .A1(net_298), .ZN(net_127), .A2(net_125) );
NAND2_X1 inst_573 ( .A1(net_549), .ZN(net_548), .A2(net_547) );
NOR3_X1 inst_100 ( .ZN(net_171), .A3(net_170), .A2(net_17), .A1(net_3) );
INV_X1 inst_642 ( .ZN(net_305), .A(net_197) );
NAND2_X1 inst_459 ( .A2(net_283), .ZN(net_244), .A1(n326) );
NAND3_X1 inst_279 ( .ZN(net_630), .A1(net_620), .A3(net_538), .A2(net_502) );
NAND2_X1 inst_445 ( .A2(net_265), .ZN(net_228), .A1(n150) );
OR2_X2 inst_93 ( .ZN(net_604), .A2(net_603), .A1(n1) );
OR2_X4 inst_81 ( .A2(net_542), .ZN(net_532), .A1(net_76) );
INV_X1 inst_612 ( .ZN(net_363), .A(n33) );
MUX2_X2 inst_606 ( .Z(net_437), .S(net_413), .B(n200), .A(n190) );
NAND2_X1 inst_367 ( .A1(net_201), .A2(net_125), .ZN(net_123) );
NAND2_X1 inst_525 ( .ZN(net_391), .A2(net_389), .A1(n107) );
NOR2_X1 inst_139 ( .ZN(net_265), .A1(net_114), .A2(net_108) );
AND4_X1 inst_657 ( .ZN(net_349), .A2(net_208), .A4(net_164), .A3(net_151), .A1(n33) );
NAND2_X1 inst_559 ( .A1(net_513), .ZN(net_510), .A2(net_492) );
NAND2_X1 inst_584 ( .ZN(net_609), .A1(net_603), .A2(net_602) );
NAND2_X1 inst_521 ( .ZN(net_386), .A2(net_384), .A1(n77) );
NAND2_X1 inst_434 ( .ZN(net_344), .A2(net_220), .A1(n58) );
NAND2_X1 inst_470 ( .ZN(net_256), .A2(net_254), .A1(n132) );
NAND2_X1 inst_535 ( .A2(net_447), .ZN(net_432), .A1(n179) );
NAND2_X1 inst_450 ( .ZN(net_233), .A2(net_231), .A1(n244) );
NAND2_X1 inst_520 ( .ZN(net_385), .A2(net_384), .A1(n58) );
NAND3_X1 inst_237 ( .ZN(net_272), .A1(net_106), .A3(net_105), .A2(net_78) );
NOR2_X1 inst_148 ( .ZN(net_200), .A1(net_199), .A2(net_197) );
NAND2_X1 inst_554 ( .A1(net_558), .ZN(net_555), .A2(net_501) );
NAND2_X1 inst_377 ( .ZN(net_135), .A2(net_133), .A1(n159) );
NAND4_X1 inst_191 ( .A2(net_363), .ZN(net_352), .A1(net_218), .A3(net_190), .A4(net_188) );
XNOR2_X1 inst_51 ( .A(net_668), .B(net_667), .ZN(n405) );
NOR2_X1 inst_142 ( .ZN(net_333), .A2(net_83), .A1(net_44) );
NAND2_X1 inst_315 ( .ZN(net_114), .A2(net_1), .A1(n20) );
OR2_X4 inst_80 ( .ZN(net_476), .A1(net_475), .A2(net_435) );
NAND4_X1 inst_216 ( .A2(net_574), .ZN(net_572), .A4(net_548), .A3(net_511), .A1(net_202) );
OR2_X4 inst_78 ( .ZN(net_458), .A1(net_424), .A2(net_397) );
NAND3_X1 inst_241 ( .ZN(net_331), .A1(net_219), .A2(net_163), .A3(net_150) );
NOR2_X1 inst_177 ( .ZN(net_579), .A1(net_578), .A2(net_560) );
NOR2_X1 inst_183 ( .ZN(net_639), .A1(net_637), .A2(net_636) );
NOR2_X1 inst_151 ( .A2(net_295), .ZN(net_290), .A1(net_289) );
OR2_X4 inst_64 ( .A1(net_298), .A2(net_51), .ZN(n355) );
NAND2_X1 inst_415 ( .A2(net_254), .ZN(net_191), .A1(n116) );
INV_X1 inst_615 ( .ZN(net_289), .A(n116) );
NAND2_X1 inst_393 ( .A2(net_165), .ZN(net_156), .A1(n132) );
NOR2_X1 inst_107 ( .ZN(net_7), .A2(n58), .A1(n50) );
OR2_X2 inst_92 ( .A1(net_591), .A2(net_579), .ZN(n369) );
NAND2_X1 inst_345 ( .ZN(net_81), .A2(net_79), .A1(n283) );
NAND3_X1 inst_223 ( .ZN(net_136), .A1(net_90), .A3(net_59), .A2(net_19) );
NAND2_X1 inst_402 ( .ZN(net_167), .A2(net_165), .A1(n143) );
NAND2_X1 inst_340 ( .A2(net_79), .ZN(net_72), .A1(n97) );
INV_X1 inst_643 ( .ZN(net_392), .A(net_183) );
NAND2_X1 inst_494 ( .A2(net_305), .ZN(net_303), .A1(n294) );
NAND2_X1 inst_487 ( .A2(net_305), .ZN(net_291), .A1(n50) );
NAND2_X1 inst_329 ( .ZN(net_89), .A1(net_52), .A2(net_40) );
NAND2_X1 inst_574 ( .ZN(net_550), .A1(net_549), .A2(net_530) );
NAND2_X1 inst_386 ( .A2(net_165), .ZN(net_149), .A1(n159) );
NOR2_X1 inst_158 ( .ZN(net_474), .A1(net_473), .A2(net_434) );
NOR2_X1 inst_141 ( .A1(net_118), .ZN(net_116), .A2(net_68) );
NAND4_X1 inst_200 ( .ZN(net_372), .A1(net_371), .A3(net_359), .A4(net_354), .A2(net_149) );
NAND2_X1 inst_507 ( .ZN(net_325), .A2(net_324), .A1(net_298) );
NAND2_X1 inst_571 ( .A2(net_617), .A1(net_593), .ZN(net_576) );
OR3_X2 inst_57 ( .ZN(net_427), .A1(net_369), .A3(net_338), .A2(n33) );
NAND2_X1 inst_338 ( .A2(net_79), .ZN(net_65), .A1(n107) );
NAND2_X1 inst_552 ( .A1(net_513), .ZN(net_494), .A2(net_458) );
MUX2_X2 inst_599 ( .Z(net_104), .S(net_82), .A(n274), .B(n250) );
NAND2_X1 inst_417 ( .ZN(net_354), .A2(net_220), .A1(n107) );
AND3_X4 inst_671 ( .ZN(net_506), .A2(net_477), .A1(net_411), .A3(net_408) );
NAND2_X1 inst_579 ( .A2(net_597), .ZN(net_586), .A1(n330) );
XNOR2_X1 inst_21 ( .A(net_317), .B(net_278), .ZN(n351) );
NAND2_X1 inst_469 ( .ZN(net_255), .A2(net_254), .A1(n137) );
NAND3_X1 inst_281 ( .A2(net_652), .ZN(net_629), .A3(net_625), .A1(net_623) );
NAND2_X1 inst_585 ( .ZN(net_616), .A2(net_594), .A1(net_498) );
XNOR2_X1 inst_18 ( .ZN(net_317), .A(net_55), .B(net_32) );
NAND2_X1 inst_541 ( .A2(net_481), .A1(net_465), .ZN(net_462) );
NAND2_X1 inst_410 ( .A2(net_254), .ZN(net_186), .A1(n50) );
NAND4_X1 inst_208 ( .ZN(net_578), .A3(net_524), .A4(net_523), .A2(net_520), .A1(net_518) );
OR2_X4 inst_88 ( .A2(net_636), .ZN(net_634), .A1(net_633) );
NAND2_X1 inst_316 ( .ZN(net_656), .A2(net_2), .A1(n213) );
NAND3_X1 inst_220 ( .A1(net_73), .ZN(net_33), .A2(n45), .A3(n13) );
XNOR2_X1 inst_9 ( .ZN(net_32), .B(n58), .A(n50) );
NOR2_X1 inst_113 ( .ZN(net_24), .A2(n68), .A1(n50) );
NAND2_X1 inst_505 ( .A2(net_324), .ZN(net_322), .A1(net_289) );
NAND2_X1 inst_356 ( .ZN(net_98), .A2(net_97), .A1(n223) );
NAND2_X1 inst_383 ( .ZN(net_361), .A2(net_168), .A1(n87) );
NAND2_X1 inst_360 ( .ZN(net_105), .A2(net_95), .A1(n20) );
NAND4_X1 inst_198 ( .ZN(net_369), .A4(net_293), .A2(net_227), .A3(net_187), .A1(net_178) );
XNOR2_X1 inst_50 ( .A(net_667), .B(net_662), .ZN(n402) );
NAND3_X1 inst_245 ( .ZN(net_403), .A2(net_374), .A3(net_309), .A1(net_232) );
NAND2_X1 inst_569 ( .A1(net_549), .ZN(net_540), .A2(net_539) );
AND2_X4 inst_678 ( .ZN(net_220), .A2(net_113), .A1(net_111) );
INV_X1 inst_624 ( .ZN(net_3), .A(n250) );
NAND3_X1 inst_260 ( .ZN(net_468), .A1(net_388), .A3(net_321), .A2(net_127) );
NOR2_X1 inst_147 ( .A1(net_296), .ZN(net_198), .A2(net_197) );
NAND2_X1 inst_313 ( .ZN(net_31), .A1(n264), .A2(n107) );
NAND2_X1 inst_293 ( .ZN(net_40), .A1(n20), .A2(n179) );
INV_X1 inst_636 ( .ZN(net_314), .A(net_172) );
INV_X1 inst_632 ( .A(net_114), .ZN(net_111) );
NAND2_X1 inst_549 ( .ZN(net_491), .A1(net_454), .A2(net_441) );
NAND3_X1 inst_234 ( .ZN(net_181), .A1(net_132), .A3(net_81), .A2(net_29) );
XOR2_X1 inst_0 ( .Z(net_41), .A(n244), .B(n238) );
NAND2_X1 inst_522 ( .A2(net_389), .ZN(net_387), .A1(n116) );
NOR2_X1 inst_184 ( .A2(net_644), .ZN(net_643), .A1(net_636) );
AND2_X4 inst_690 ( .A1(net_617), .A2(net_616), .ZN(net_614) );
NAND3_X1 inst_236 ( .ZN(net_271), .A1(net_131), .A3(net_85), .A2(net_65) );
NAND2_X1 inst_433 ( .A2(net_280), .ZN(net_216), .A1(n159) );
NAND2_X1 inst_553 ( .A1(net_558), .A2(net_507), .ZN(net_498) );
NAND2_X1 inst_478 ( .ZN(net_266), .A2(net_265), .A1(n311) );
OR2_X4 inst_65 ( .A2(net_269), .ZN(net_170), .A1(net_73) );
NAND2_X1 inst_536 ( .A2(net_447), .ZN(net_433), .A1(net_5) );
NAND3_X1 inst_242 ( .ZN(net_346), .A3(net_344), .A2(net_337), .A1(net_148) );
AND2_X4 inst_688 ( .ZN(net_524), .A1(net_505), .A2(net_476) );
NAND2_X1 inst_516 ( .ZN(net_367), .A1(net_350), .A2(net_318) );
NOR4_X1 inst_98 ( .ZN(net_485), .A2(net_444), .A3(net_443), .A4(net_442), .A1(net_432) );
NAND3_X1 inst_263 ( .ZN(net_475), .A1(net_383), .A3(net_334), .A2(net_119) );
NAND4_X1 inst_190 ( .A2(net_363), .ZN(net_348), .A1(net_284), .A4(net_281), .A3(net_185) );
NAND4_X1 inst_185 ( .ZN(net_75), .A2(net_31), .A4(net_27), .A1(net_18), .A3(net_13) );
XNOR2_X1 inst_13 ( .ZN(net_46), .A(n232), .B(n226) );
OR2_X4 inst_75 ( .A2(net_409), .ZN(net_408), .A1(n179) );
NAND2_X1 inst_332 ( .A2(net_61), .ZN(net_59), .A1(n223) );
NOR2_X1 inst_166 ( .ZN(net_519), .A1(net_501), .A2(net_472) );
NOR2_X1 inst_116 ( .A1(net_363), .ZN(net_79), .A2(n20) );
NAND2_X1 inst_598 ( .ZN(net_657), .A1(net_656), .A2(n375) );
NAND2_X1 inst_416 ( .A2(net_220), .ZN(net_192), .A1(n116) );
NOR2_X1 inst_163 ( .ZN(net_487), .A1(net_486), .A2(net_448) );
NAND2_X1 inst_471 ( .A2(net_280), .ZN(net_257), .A1(n116) );
NAND2_X1 inst_394 ( .A2(net_165), .ZN(net_157), .A1(n294) );
OR2_X4 inst_79 ( .ZN(net_469), .A1(net_468), .A2(net_396) );
NOR3_X1 inst_106 ( .ZN(net_590), .A3(net_563), .A1(net_554), .A2(net_499) );
NAND2_X1 inst_422 ( .A2(net_265), .ZN(net_195), .A1(n97) );
NAND4_X1 inst_219 ( .ZN(net_577), .A2(net_574), .A4(net_550), .A3(net_514), .A1(net_206) );
NAND4_X1 inst_201 ( .ZN(net_376), .A2(net_371), .A4(net_257), .A1(net_195), .A3(net_193) );
MUX2_X2 inst_605 ( .Z(net_436), .S(net_409), .B(n200), .A(n190) );
NAND2_X1 inst_304 ( .ZN(net_21), .A2(n50), .A1(n226) );
NAND2_X1 inst_542 ( .A2(net_471), .A1(net_465), .ZN(net_463) );
NAND3_X1 inst_255 ( .ZN(net_445), .A1(net_444), .A2(net_443), .A3(net_442) );
NAND2_X1 inst_453 ( .ZN(net_237), .A2(net_235), .A1(n257) );
NOR2_X1 inst_128 ( .ZN(net_83), .A2(net_35), .A1(n13) );
OR2_X4 inst_73 ( .A2(net_403), .ZN(net_402), .A1(n179) );
NAND2_X1 inst_493 ( .A2(net_305), .ZN(net_301), .A1(n159) );
NAND2_X1 inst_378 ( .ZN(net_337), .A2(net_168), .A1(n68) );
XNOR2_X1 inst_23 ( .ZN(net_617), .A(net_520), .B(net_460) );
NAND2_X1 inst_339 ( .A2(net_79), .ZN(net_66), .A1(n87) );
NAND2_X1 inst_351 ( .A2(net_97), .ZN(net_88), .A1(n264) );
NAND2_X1 inst_361 ( .A2(net_133), .ZN(net_106), .A1(n150) );
NAND2_X1 inst_408 ( .ZN(net_342), .A2(net_220), .A1(n68) );
NAND2_X1 inst_325 ( .A2(net_61), .ZN(net_50), .A1(n250) );
NAND2_X1 inst_461 ( .A2(net_283), .ZN(net_246), .A1(n311) );
NAND2_X1 inst_385 ( .A2(net_165), .ZN(net_148), .A1(n283) );
NAND4_X1 inst_197 ( .ZN(net_368), .A4(net_287), .A2(net_216), .A3(net_189), .A1(net_186) );
AND4_X1 inst_659 ( .ZN(net_355), .A4(net_354), .A3(net_155), .A2(net_145), .A1(n33) );
NAND3_X1 inst_250 ( .ZN(net_444), .A2(net_373), .A3(net_315), .A1(net_236) );
NOR2_X1 inst_179 ( .A2(net_587), .ZN(net_585), .A1(net_547) );
XNOR2_X1 inst_24 ( .ZN(net_593), .A(net_518), .B(net_461) );
NOR2_X1 inst_114 ( .ZN(net_51), .A2(n97), .A1(n107) );
INV_X1 inst_617 ( .ZN(net_296), .A(n107) );
OR2_X4 inst_76 ( .A2(net_413), .ZN(net_412), .A1(n179) );
NAND2_X1 inst_397 ( .A2(net_165), .ZN(net_161), .A1(n128) );
NAND2_X1 inst_504 ( .A1(net_333), .ZN(net_321), .A2(net_273) );
NOR2_X1 inst_150 ( .A1(net_289), .ZN(net_288), .A2(net_143) );
NOR2_X1 inst_172 ( .ZN(net_554), .A1(net_553), .A2(net_545) );
NAND2_X1 inst_362 ( .ZN(net_197), .A1(net_114), .A2(net_113) );
NAND3_X1 inst_277 ( .A3(net_604), .A1(net_275), .A2(net_215), .ZN(n364) );
OR2_X4 inst_83 ( .ZN(net_543), .A2(net_542), .A1(n330) );
NOR2_X1 inst_121 ( .ZN(net_97), .A2(net_61), .A1(n33) );
NAND2_X1 inst_534 ( .A1(net_455), .ZN(net_431), .A2(net_393) );
NAND2_X1 inst_440 ( .A2(net_254), .ZN(net_223), .A1(n294) );
NAND2_X1 inst_306 ( .ZN(net_23), .A2(n77), .A1(n244) );
XOR2_X1 inst_2 ( .Z(net_533), .B(net_525), .A(net_466) );
INV_X1 inst_644 ( .A(net_333), .ZN(net_176) );
NAND2_X1 inst_596 ( .ZN(net_653), .A1(net_652), .A2(net_647) );
NAND2_X1 inst_578 ( .A2(net_569), .A1(net_565), .ZN(n396) );
OR4_X1 inst_52 ( .ZN(net_658), .A3(n396), .A4(n390), .A1(n384), .A2(n378) );
OR2_X4 inst_90 ( .ZN(net_650), .A2(net_643), .A1(net_637) );
NAND3_X1 inst_267 ( .ZN(net_452), .A1(net_419), .A3(net_261), .A2(net_238) );
NOR2_X1 inst_140 ( .A1(net_319), .A2(net_214), .ZN(net_115) );
AND3_X4 inst_668 ( .ZN(net_343), .A3(net_342), .A1(net_156), .A2(net_146) );
NAND3_X1 inst_221 ( .ZN(net_483), .A3(net_73), .A1(net_54), .A2(n213) );
NAND2_X1 inst_556 ( .A2(net_504), .ZN(net_502), .A1(net_483) );
INV_X1 inst_650 ( .A(net_617), .ZN(net_530) );
INV_X1 inst_637 ( .ZN(net_633), .A(net_626) );
NAND3_X1 inst_289 ( .A3(net_653), .A1(net_645), .A2(net_575), .ZN(n378) );
NAND2_X1 inst_547 ( .ZN(net_489), .A1(net_450), .A2(net_428) );
NAND2_X1 inst_530 ( .A1(net_410), .ZN(net_407), .A2(net_406) );
NAND2_X1 inst_432 ( .A2(net_280), .ZN(net_211), .A1(n283) );
AND2_X4 inst_679 ( .A2(net_165), .ZN(net_160), .A1(n124) );
NAND2_X1 inst_420 ( .ZN(net_356), .A2(net_220), .A1(n97) );
NAND3_X1 inst_282 ( .A3(net_624), .A1(net_613), .A2(net_573), .ZN(n390) );
NAND2_X1 inst_368 ( .A1(net_296), .A2(net_125), .ZN(net_124) );
NAND2_X1 inst_513 ( .A1(net_333), .ZN(net_332), .A2(net_271) );
XNOR2_X1 inst_44 ( .ZN(net_647), .A(net_644), .B(net_639) );
NAND3_X1 inst_274 ( .ZN(net_569), .A1(net_568), .A2(net_567), .A3(net_543) );
NOR2_X1 inst_174 ( .A1(net_568), .ZN(net_562), .A2(net_561) );
NAND2_X1 inst_371 ( .A2(net_133), .ZN(net_128), .A1(n68) );
AND4_X1 inst_662 ( .ZN(net_375), .A2(net_363), .A4(net_301), .A1(net_248), .A3(net_228) );
NAND2_X1 inst_314 ( .ZN(net_82), .A2(net_44), .A1(n45) );
NAND2_X1 inst_435 ( .A2(net_265), .ZN(net_217), .A1(n159) );
NOR2_X1 inst_164 ( .ZN(net_497), .A2(net_485), .A1(net_470) );
XOR2_X1 inst_5 ( .Z(net_618), .A(net_617), .B(net_616) );
NAND2_X1 inst_597 ( .A1(net_656), .ZN(net_655), .A2(n378) );
NOR2_X1 inst_157 ( .ZN(net_472), .A1(net_471), .A2(net_438) );
AND2_X4 inst_687 ( .A1(net_558), .A2(net_503), .ZN(net_499) );
INV_X1 inst_621 ( .ZN(net_1), .A(n190) );
OR2_X4 inst_68 ( .ZN(net_174), .A2(net_173), .A1(net_0) );
NAND4_X1 inst_213 ( .A1(net_574), .ZN(net_565), .A4(net_532), .A2(net_508), .A3(net_456) );
MUX2_X2 inst_604 ( .Z(net_435), .S(net_406), .B(n200), .A(n190) );
OR3_X4 inst_53 ( .A3(net_661), .ZN(n407), .A1(n393), .A2(n387) );
INV_X1 inst_628 ( .ZN(net_5), .A(n179) );
NAND4_X1 inst_205 ( .ZN(net_429), .A1(net_375), .A2(net_345), .A4(net_263), .A3(net_253) );
NAND2_X1 inst_472 ( .A2(net_280), .ZN(net_258), .A1(n143) );
NAND2_X1 inst_447 ( .A2(net_231), .ZN(net_229), .A1(n238) );
NAND2_X1 inst_380 ( .A2(net_168), .ZN(net_145), .A1(n116) );
NAND2_X1 inst_457 ( .A2(net_283), .ZN(net_242), .A1(n317) );
INV_X1 inst_651 ( .A(net_593), .ZN(net_547) );
AND4_X1 inst_665 ( .ZN(net_420), .A4(net_357), .A2(net_294), .A3(net_246), .A1(net_209) );
NAND2_X1 inst_292 ( .ZN(net_9), .A2(n33), .A1(n107) );
NAND2_X1 inst_379 ( .A2(net_168), .ZN(net_144), .A1(n50) );
NOR2_X1 inst_127 ( .ZN(net_107), .A2(net_82), .A1(n41) );
NAND4_X1 inst_186 ( .ZN(net_84), .A3(net_28), .A2(net_26), .A1(net_23), .A4(net_21) );
XNOR2_X1 inst_17 ( .ZN(net_173), .B(net_46), .A(net_41) );
NAND2_X1 inst_413 ( .A2(net_265), .ZN(net_189), .A1(n58) );
NOR2_X1 inst_146 ( .A1(net_350), .ZN(net_324), .A2(net_183) );
NAND3_X1 inst_249 ( .ZN(net_413), .A2(net_374), .A3(net_313), .A1(net_233) );
NAND2_X1 inst_334 ( .ZN(net_62), .A2(net_61), .A1(n244) );
NAND4_X1 inst_187 ( .A4(net_274), .ZN(net_268), .A1(net_25), .A2(net_12), .A3(n58) );
NAND4_X1 inst_206 ( .A4(net_524), .A2(net_523), .ZN(net_521), .A3(net_520), .A1(net_507) );
NOR2_X1 inst_122 ( .ZN(net_109), .A2(net_8), .A1(n1) );
XNOR2_X1 inst_25 ( .ZN(net_619), .A(net_523), .B(net_464) );
NAND2_X1 inst_354 ( .A2(net_97), .ZN(net_94), .A1(n232) );
NAND2_X1 inst_405 ( .ZN(net_558), .A2(net_177), .A1(n343) );
NAND2_X1 inst_492 ( .A2(net_305), .ZN(net_300), .A1(n283) );
NAND3_X1 inst_240 ( .ZN(net_308), .A3(net_135), .A1(net_86), .A2(net_77) );
NAND2_X1 inst_326 ( .ZN(net_172), .A2(net_58), .A1(net_10) );
NOR2_X1 inst_110 ( .ZN(net_549), .A2(n33), .A1(n13) );
NAND2_X1 inst_518 ( .A2(net_384), .ZN(net_382), .A1(n68) );
OR2_X4 inst_74 ( .A2(net_406), .ZN(net_405), .A1(n179) );
NAND3_X1 inst_288 ( .A3(net_651), .A2(net_270), .A1(net_92), .ZN(n367) );
NAND2_X1 inst_396 ( .A2(net_165), .ZN(net_159), .A1(n311) );
NAND3_X1 inst_229 ( .ZN(net_142), .A1(net_88), .A3(net_48), .A2(net_14) );
NOR3_X1 inst_99 ( .ZN(net_71), .A1(net_70), .A3(net_69), .A2(n50) );
OR2_X4 inst_69 ( .ZN(net_215), .A1(net_214), .A2(net_213) );
NAND2_X1 inst_373 ( .A2(net_133), .ZN(net_130), .A1(n58) );
OR2_X4 inst_82 ( .A2(net_556), .A1(net_555), .ZN(net_541) );
AND3_X4 inst_669 ( .ZN(net_345), .A3(net_344), .A1(net_161), .A2(net_144) );
NOR2_X1 inst_108 ( .ZN(net_8), .A2(n45), .A1(n41) );
AND4_X1 inst_664 ( .ZN(net_419), .A4(net_355), .A2(net_300), .A3(net_242), .A1(net_224) );
NAND2_X1 inst_595 ( .ZN(net_649), .A2(net_648), .A1(net_626) );
NAND3_X1 inst_283 ( .A3(net_629), .A1(net_627), .A2(net_564), .ZN(n387) );
XNOR2_X1 inst_22 ( .ZN(net_539), .B(net_524), .A(net_484) );
NAND2_X1 inst_311 ( .ZN(net_29), .A2(n20), .A1(n116) );
NAND2_X1 inst_460 ( .A2(net_283), .ZN(net_245), .A1(n143) );
NAND2_X1 inst_372 ( .A2(net_133), .ZN(net_129), .A1(n50) );
NOR2_X1 inst_169 ( .ZN(net_520), .A1(net_506), .A2(net_478) );
NAND4_X1 inst_215 ( .A2(net_574), .ZN(net_571), .A4(net_540), .A3(net_515), .A1(net_203) );
NAND2_X1 inst_307 ( .ZN(net_25), .A2(n77), .A1(n68) );
INV_X1 inst_638 ( .A(net_125), .ZN(net_100) );
NAND2_X1 inst_421 ( .ZN(net_339), .A2(net_220), .A1(n87) );
NOR2_X1 inst_161 ( .ZN(net_482), .A1(net_481), .A2(net_439) );
NAND2_X1 inst_560 ( .A1(net_513), .ZN(net_511), .A2(net_489) );
NAND2_X1 inst_586 ( .ZN(net_637), .A2(net_605), .A1(net_586) );
NAND2_X1 inst_555 ( .A1(net_558), .ZN(net_553), .A2(net_500) );
XNOR2_X1 inst_16 ( .ZN(net_276), .A(net_45), .B(net_42) );
NAND3_X1 inst_276 ( .A2(net_652), .ZN(net_610), .A3(net_609), .A1(net_601) );
NAND2_X1 inst_431 ( .A2(net_254), .ZN(net_210), .A1(n283) );
NAND2_X1 inst_348 ( .ZN(net_86), .A2(net_67), .A1(n20) );
XOR2_X1 inst_3 ( .Z(net_556), .B(net_522), .A(net_462) );
NOR2_X1 inst_156 ( .ZN(net_389), .A2(net_335), .A1(net_38) );
NAND2_X1 inst_577 ( .ZN(net_588), .A2(net_559), .A1(net_558) );
NAND2_X1 inst_566 ( .A1(net_535), .ZN(net_534), .A2(net_533) );
NAND2_X1 inst_296 ( .ZN(net_13), .A2(n97), .A1(n257) );
OR2_X2 inst_91 ( .A1(net_582), .A2(net_581), .ZN(n399) );
NOR2_X1 inst_132 ( .ZN(net_274), .A2(net_101), .A1(n116) );
NAND2_X1 inst_342 ( .A2(net_79), .ZN(net_77), .A1(n68) );
NAND2_X1 inst_526 ( .A2(net_444), .A1(net_410), .ZN(net_398) );
XNOR2_X1 inst_36 ( .ZN(net_636), .A(net_618), .B(net_585) );
INV_X1 inst_656 ( .ZN(net_640), .A(net_639) );
INV_X1 inst_645 ( .ZN(net_652), .A(net_213) );
NAND2_X1 inst_463 ( .A2(net_283), .ZN(net_248), .A1(n132) );
NAND2_X1 inst_503 ( .ZN(net_316), .A1(net_314), .A2(net_138) );
NOR4_X1 inst_96 ( .ZN(net_417), .A4(net_362), .A1(net_297), .A3(net_285), .A2(net_200) );
XNOR2_X1 inst_45 ( .ZN(net_667), .A(net_646), .B(net_638) );
NAND2_X1 inst_451 ( .A2(net_235), .ZN(net_234), .A1(n270) );
NOR3_X1 inst_101 ( .A1(net_320), .A3(net_171), .A2(net_115), .ZN(n361) );
NAND2_X1 inst_319 ( .A2(net_410), .ZN(net_39), .A1(n20) );
NAND3_X1 inst_269 ( .ZN(net_454), .A1(net_418), .A3(net_262), .A2(net_251) );
NAND2_X1 inst_458 ( .A2(net_283), .ZN(net_243), .A1(n137) );
NAND2_X1 inst_444 ( .A2(net_280), .ZN(net_227), .A1(n150) );
NAND2_X1 inst_400 ( .A2(net_165), .ZN(net_164), .A1(n329) );
INV_X1 inst_614 ( .ZN(net_118), .A(n50) );
AND2_X4 inst_686 ( .A1(net_558), .ZN(net_537), .A2(net_506) );
INV_X1 inst_649 ( .A(net_475), .ZN(net_459) );
NAND3_X1 inst_261 ( .ZN(net_486), .A1(net_390), .A3(net_332), .A2(net_126) );
NAND2_X1 inst_514 ( .ZN(net_334), .A1(net_333), .A2(net_272) );
NAND2_X1 inst_500 ( .A1(net_314), .ZN(net_312), .A2(net_142) );
NAND2_X1 inst_510 ( .A1(net_333), .ZN(net_328), .A2(net_181) );
NAND3_X1 inst_268 ( .ZN(net_453), .A1(net_421), .A3(net_260), .A2(net_252) );
AND2_X4 inst_685 ( .ZN(net_525), .A2(net_496), .A1(net_469) );
NAND2_X1 inst_369 ( .A1(net_199), .ZN(net_126), .A2(net_125) );
NAND2_X1 inst_550 ( .ZN(net_492), .A1(net_452), .A2(net_426) );
OR2_X4 inst_63 ( .ZN(net_269), .A1(net_44), .A2(n13) );
NOR2_X1 inst_119 ( .A2(net_363), .A1(net_73), .ZN(net_35) );
MUX2_X2 inst_603 ( .Z(net_434), .S(net_403), .B(n200), .A(n190) );
NAND2_X1 inst_327 ( .A1(net_298), .ZN(net_101), .A2(net_51) );
AND2_X4 inst_676 ( .ZN(net_58), .A2(n13), .A1(n1) );
OR2_X4 inst_85 ( .ZN(net_587), .A2(net_570), .A1(net_4) );
NAND3_X1 inst_291 ( .A1(net_660), .ZN(n409), .A3(n407), .A2(n213) );
NAND3_X1 inst_266 ( .ZN(net_451), .A1(net_420), .A3(net_241), .A2(net_223) );
NAND2_X1 inst_473 ( .A2(net_280), .ZN(net_260), .A1(n322) );
NAND4_X1 inst_217 ( .A1(net_574), .ZN(net_573), .A2(net_546), .A4(net_510), .A3(net_430) );
NAND2_X1 inst_572 ( .ZN(net_546), .A2(net_545), .A1(net_535) );
OR2_X4 inst_77 ( .A2(net_444), .ZN(net_415), .A1(n179) );
NOR2_X1 inst_171 ( .A2(net_578), .A1(net_544), .ZN(n372) );
NAND2_X1 inst_558 ( .A1(net_513), .ZN(net_509), .A2(net_491) );
NAND2_X1 inst_427 ( .ZN(net_206), .A1(net_205), .A2(net_204) );
NAND3_X1 inst_257 ( .ZN(net_477), .A1(net_382), .A3(net_327), .A2(net_117) );
NAND2_X1 inst_594 ( .A1(net_637), .A2(net_636), .ZN(net_635) );
NOR2_X1 inst_145 ( .A1(net_549), .A2(net_513), .ZN(net_204) );
NAND3_X1 inst_290 ( .A3(net_654), .A1(net_649), .A2(net_571), .ZN(n375) );
NAND2_X1 inst_374 ( .A2(net_133), .ZN(net_131), .A1(n77) );
NAND3_X1 inst_272 ( .ZN(net_528), .A1(net_524), .A3(net_523), .A2(net_506) );
NAND2_X1 inst_502 ( .ZN(net_315), .A1(net_314), .A2(net_139) );
NOR3_X1 inst_103 ( .ZN(net_425), .A1(net_370), .A3(net_366), .A2(net_160) );
NAND2_X1 inst_485 ( .ZN(net_335), .A2(net_176), .A1(net_100) );
NAND2_X1 inst_565 ( .A2(net_525), .ZN(net_517), .A1(net_503) );
NAND3_X1 inst_248 ( .ZN(net_409), .A2(net_374), .A3(net_311), .A1(net_229) );
AND3_X4 inst_672 ( .ZN(net_507), .A2(net_479), .A1(net_414), .A3(net_412) );
INV_X1 inst_622 ( .ZN(net_2), .A(n343) );
NOR2_X1 inst_138 ( .ZN(net_183), .A2(net_170), .A1(n33) );
NAND2_X1 inst_389 ( .A2(net_168), .ZN(net_152), .A1(n283) );
NAND2_X1 inst_357 ( .ZN(net_99), .A2(net_97), .A1(n244) );
NAND2_X1 inst_409 ( .A2(net_254), .ZN(net_185), .A1(n68) );
NOR2_X1 inst_180 ( .ZN(net_589), .A2(net_588), .A1(net_578) );
XNOR2_X1 inst_33 ( .ZN(net_607), .B(net_590), .A(net_533) );
NAND2_X1 inst_312 ( .ZN(net_30), .A2(n33), .A1(n116) );
AND4_X1 inst_660 ( .ZN(net_357), .A4(net_356), .A3(net_153), .A2(net_147), .A1(n33) );
MUX2_X2 inst_609 ( .Z(net_448), .S(net_447), .A(n200), .B(n190) );
NAND2_X1 inst_517 ( .A2(net_443), .A1(net_410), .ZN(net_381) );
NAND2_X1 inst_309 ( .ZN(net_27), .A2(n87), .A1(n250) );
NAND3_X1 inst_232 ( .ZN(net_179), .A1(net_129), .A3(net_80), .A2(net_43) );
NAND2_X1 inst_347 ( .A2(net_91), .ZN(net_85), .A1(n20) );
AND4_X1 inst_663 ( .ZN(net_418), .A4(net_353), .A2(net_303), .A3(net_247), .A1(net_239) );
NAND2_X1 inst_301 ( .ZN(net_19), .A2(n87), .A1(n33) );
NAND2_X1 inst_363 ( .A1(net_205), .A2(net_125), .ZN(net_117) );
XNOR2_X1 inst_27 ( .ZN(net_542), .A(net_519), .B(net_463) );
NAND3_X1 inst_247 ( .ZN(net_442), .A2(net_373), .A3(net_312), .A1(net_234) );
NAND2_X1 inst_297 ( .ZN(net_14), .A2(n33), .A1(n303) );
NAND2_X1 inst_403 ( .ZN(net_169), .A2(net_168), .A1(n150) );
NAND2_X1 inst_302 ( .ZN(net_52), .A2(n200), .A1(n20) );
NAND2_X1 inst_310 ( .ZN(net_28), .A2(n58), .A1(n232) );
NAND2_X1 inst_322 ( .A1(net_205), .ZN(net_95), .A2(net_7) );
AND3_X4 inst_673 ( .ZN(net_500), .A2(net_481), .A3(net_415), .A1(net_398) );
NAND3_X1 inst_253 ( .ZN(net_422), .A3(net_351), .A1(net_323), .A2(net_302) );
NAND4_X1 inst_211 ( .ZN(net_559), .A3(net_529), .A4(net_527), .A1(net_517), .A2(net_496) );
INV_X1 inst_619 ( .ZN(net_410), .A(n169) );
AND2_X4 inst_681 ( .A2(net_283), .ZN(net_240), .A1(n303) );
NOR2_X1 inst_162 ( .ZN(net_484), .A1(net_483), .A2(net_459) );
NAND2_X1 inst_589 ( .ZN(net_621), .A2(net_606), .A1(net_567) );
NAND2_X1 inst_561 ( .A1(net_513), .ZN(net_512), .A2(net_493) );
NAND2_X1 inst_412 ( .A2(net_280), .ZN(net_188), .A1(n50) );
NAND2_X1 inst_449 ( .ZN(net_232), .A2(net_231), .A1(n232) );
INV_X1 inst_639 ( .A(net_483), .ZN(net_177) );
NOR2_X1 inst_155 ( .ZN(net_384), .A2(net_335), .A1(net_34) );
NAND2_X1 inst_464 ( .A2(net_283), .ZN(net_249), .A1(n128) );
MUX2_X2 inst_602 ( .S(net_443), .Z(net_396), .B(n200), .A(n190) );
OR3_X2 inst_59 ( .ZN(net_441), .A3(net_378), .A1(net_352), .A2(net_286) );
NOR2_X1 inst_135 ( .A2(net_314), .ZN(net_231), .A1(net_109) );
NAND2_X1 inst_341 ( .A2(net_79), .ZN(net_74), .A1(n116) );
NAND4_X1 inst_196 ( .ZN(net_366), .A4(net_282), .A3(net_256), .A1(net_250), .A2(net_69) );
NAND2_X1 inst_532 ( .ZN(net_414), .A2(net_413), .A1(net_410) );
OR3_X2 inst_55 ( .ZN(net_270), .A2(net_269), .A1(net_116), .A3(net_24) );
XNOR2_X1 inst_37 ( .ZN(net_628), .B(net_622), .A(net_619) );
INV_X1 inst_641 ( .A(net_283), .ZN(net_143) );
NAND2_X1 inst_498 ( .A1(net_314), .ZN(net_310), .A2(net_137) );
AND2_X4 inst_684 ( .A2(net_305), .ZN(net_304), .A1(n150) );
NAND3_X1 inst_264 ( .ZN(net_449), .A1(net_417), .A3(net_211), .A2(net_191) );
OR2_X4 inst_84 ( .ZN(net_561), .A1(net_556), .A2(net_545) );
NOR2_X1 inst_173 ( .ZN(net_581), .A2(net_568), .A1(net_556) );
NAND2_X1 inst_298 ( .ZN(net_15), .A2(n77), .A1(n33) );
NAND2_X1 inst_303 ( .ZN(net_20), .A2(n33), .A1(n294) );
MUX2_X2 inst_611 ( .Z(net_668), .A(net_666), .B(net_665), .S(net_103) );
NAND3_X1 inst_224 ( .ZN(net_137), .A1(net_98), .A3(net_57), .A2(net_15) );
XNOR2_X1 inst_42 ( .ZN(net_648), .A(net_631), .B(net_595) );
NAND3_X1 inst_287 ( .ZN(net_654), .A2(net_652), .A1(net_650), .A3(net_648) );
NAND2_X1 inst_323 ( .A2(net_61), .ZN(net_48), .A1(n257) );
INV_X1 inst_618 ( .ZN(net_0), .A(n45) );
NAND2_X1 inst_426 ( .A2(net_204), .ZN(net_203), .A1(net_118) );
NAND2_X1 inst_588 ( .A1(net_626), .ZN(net_613), .A2(net_612) );
INV_X1 inst_648 ( .ZN(net_447), .A(net_395) );
NAND2_X1 inst_350 ( .A2(net_97), .ZN(net_87), .A1(n250) );
NAND3_X1 inst_231 ( .ZN(net_175), .A1(net_99), .A3(net_49), .A2(net_30) );
NAND3_X1 inst_270 ( .ZN(net_505), .A2(net_475), .A1(net_407), .A3(net_405) );
NAND2_X1 inst_474 ( .A2(net_280), .ZN(net_261), .A1(n311) );
XNOR2_X1 inst_26 ( .ZN(net_531), .A(net_526), .B(net_467) );
NAND2_X1 inst_437 ( .A2(net_220), .ZN(net_219), .A1(n50) );
NAND2_X1 inst_490 ( .ZN(net_377), .A2(net_305), .A1(n77) );
INV_X1 inst_626 ( .ZN(net_4), .A(n330) );
OR2_X4 inst_70 ( .A1(net_392), .ZN(net_302), .A2(net_274) );
NOR2_X1 inst_129 ( .ZN(net_165), .A1(net_114), .A2(net_89) );
NAND4_X1 inst_189 ( .ZN(net_341), .A3(net_340), .A4(net_339), .A1(net_222), .A2(net_167) );
XNOR2_X1 inst_11 ( .ZN(net_67), .A(n68), .B(n58) );
INV_X1 inst_631 ( .ZN(net_64), .A(net_40) );
NAND4_X1 inst_188 ( .ZN(net_338), .A3(net_337), .A4(net_336), .A1(net_245), .A2(net_154) );
XNOR2_X1 inst_14 ( .A(net_298), .ZN(net_47), .B(n116) );
NAND2_X1 inst_475 ( .A2(net_280), .ZN(net_262), .A1(n317) );
NAND2_X1 inst_441 ( .A2(net_265), .ZN(net_224), .A1(n294) );
XNOR2_X1 inst_31 ( .ZN(net_612), .B(net_583), .A(net_581) );
NAND2_X1 inst_528 ( .A1(net_410), .ZN(net_400), .A2(net_395) );
NAND3_X1 inst_252 ( .ZN(net_394), .A2(net_392), .A3(net_326), .A1(net_279) );
OR3_X2 inst_62 ( .ZN(net_661), .A1(net_658), .A3(n381), .A2(n375) );
NAND2_X1 inst_557 ( .A1(net_513), .ZN(net_508), .A2(net_490) );
NAND3_X1 inst_251 ( .ZN(net_393), .A1(net_392), .A2(net_325), .A3(net_277) );
NAND2_X1 inst_352 ( .A2(net_97), .ZN(net_90), .A1(n226) );
NAND2_X1 inst_575 ( .ZN(net_552), .A2(net_551), .A1(net_549) );
NAND2_X1 inst_398 ( .A2(net_165), .ZN(net_162), .A1(n303) );
NAND3_X1 inst_286 ( .A3(net_642), .A1(net_634), .A2(net_577), .ZN(n381) );
NAND2_X1 inst_436 ( .A2(net_283), .ZN(net_218), .A1(n159) );
NAND2_X1 inst_484 ( .ZN(net_284), .A2(net_283), .A1(n50) );
INV_X1 inst_627 ( .ZN(net_73), .A(n20) );
NAND2_X1 inst_300 ( .ZN(net_18), .A1(n270), .A2(n116) );
NOR3_X1 inst_102 ( .ZN(net_424), .A1(net_376), .A3(net_365), .A2(net_212) );
XNOR2_X1 inst_32 ( .ZN(net_606), .B(net_600), .A(net_587) );
NAND2_X1 inst_344 ( .ZN(net_80), .A2(net_79), .A1(n77) );
NAND2_X1 inst_428 ( .ZN(net_207), .A2(net_204), .A1(net_120) );
NAND2_X1 inst_446 ( .ZN(net_336), .A2(net_220), .A1(n77) );
NAND2_X1 inst_364 ( .A2(net_125), .ZN(net_119), .A1(net_118) );
NOR2_X1 inst_144 ( .ZN(net_254), .A1(net_114), .A2(net_110) );
INV_X1 inst_629 ( .ZN(net_199), .A(n97) );
NAND4_X1 inst_195 ( .ZN(net_365), .A4(net_342), .A3(net_340), .A2(net_157), .A1(n33) );
NAND2_X1 inst_407 ( .ZN(net_184), .A2(net_183), .A1(n355) );
INV_X1 inst_623 ( .ZN(net_205), .A(n68) );
NAND2_X1 inst_411 ( .A2(net_265), .ZN(net_187), .A1(n50) );
NOR4_X1 inst_97 ( .ZN(net_446), .A4(net_379), .A2(net_346), .A3(net_299), .A1(net_288) );
INV_X1 inst_616 ( .ZN(net_120), .A(n58) );
NOR2_X1 inst_124 ( .ZN(net_133), .A2(net_79), .A1(n20) );
NAND2_X1 inst_533 ( .A1(net_455), .ZN(net_430), .A2(net_394) );
INV_X1 inst_620 ( .ZN(net_201), .A(n77) );
INV_X1 inst_652 ( .A(net_619), .ZN(net_551) );
AND2_X4 inst_680 ( .A2(net_283), .ZN(net_212), .A1(n283) );
NOR2_X1 inst_137 ( .ZN(net_283), .A1(net_111), .A2(net_110) );
AND2_X4 inst_677 ( .ZN(net_513), .A1(net_58), .A2(net_39) );
NAND2_X1 inst_425 ( .A2(net_204), .ZN(net_202), .A1(net_201) );
NAND2_X1 inst_545 ( .A2(net_486), .ZN(net_467), .A1(net_465) );
NOR2_X1 inst_130 ( .A2(net_95), .ZN(n353), .A1(n77) );
NAND3_X1 inst_227 ( .ZN(net_140), .A1(net_93), .A3(net_60), .A2(net_9) );
NAND2_X1 inst_399 ( .A2(net_168), .ZN(net_163), .A1(n159) );
NAND2_X1 inst_527 ( .A2(net_442), .A1(net_410), .ZN(net_399) );
NAND3_X1 inst_226 ( .ZN(net_139), .A1(net_96), .A3(net_50), .A2(net_20) );
NOR2_X1 inst_176 ( .ZN(net_597), .A1(net_578), .A2(net_570) );
OR3_X2 inst_58 ( .ZN(net_440), .A3(net_372), .A1(net_348), .A2(net_292) );
NAND2_X1 inst_414 ( .A2(net_254), .ZN(net_190), .A1(n58) );
OR2_X4 inst_87 ( .A1(net_603), .A2(net_602), .ZN(net_601) );
OR3_X2 inst_61 ( .ZN(net_660), .A2(net_656), .A1(n378), .A3(n375) );
NAND2_X1 inst_562 ( .ZN(net_514), .A1(net_513), .A2(net_488) );
NAND2_X1 inst_531 ( .ZN(net_411), .A1(net_410), .A2(net_409) );
NAND4_X1 inst_203 ( .ZN(net_379), .A1(net_377), .A2(net_196), .A4(net_194), .A3(net_70) );
NAND4_X1 inst_212 ( .A1(net_574), .ZN(net_564), .A4(net_534), .A3(net_512), .A2(net_431) );
NAND2_X1 inst_499 ( .A1(net_314), .ZN(net_311), .A2(net_141) );
NAND2_X1 inst_335 ( .ZN(net_63), .A2(net_61), .A1(n226) );
AND3_X4 inst_674 ( .ZN(net_501), .A2(net_471), .A3(net_401), .A1(net_399) );
NAND2_X1 inst_466 ( .A2(net_254), .ZN(net_251), .A1(n311) );
AND4_X1 inst_658 ( .ZN(net_353), .A4(net_192), .A2(net_158), .A3(net_152), .A1(n33) );
XNOR2_X1 inst_10 ( .ZN(net_42), .A(n257), .B(n250) );
XOR2_X1 inst_4 ( .Z(net_557), .A(net_556), .B(net_555) );
NAND2_X1 inst_456 ( .A2(net_280), .ZN(net_241), .A1(n303) );
NAND2_X1 inst_581 ( .ZN(net_594), .A1(net_593), .A2(net_580) );
MUX2_X2 inst_600 ( .Z(net_318), .B(net_317), .A(net_214), .S(n45) );
XNOR2_X1 inst_28 ( .ZN(net_602), .A(net_568), .B(net_557) );
NAND3_X1 inst_275 ( .ZN(net_608), .A1(net_599), .A3(net_598), .A2(n330) );
NOR2_X1 inst_117 ( .A1(net_363), .ZN(net_70), .A2(n41) );
NAND2_X1 inst_438 ( .ZN(net_221), .A2(net_220), .A1(n159) );
NAND2_X1 inst_501 ( .A1(net_314), .ZN(net_313), .A2(net_140) );
XNOR2_X1 inst_49 ( .ZN(net_665), .A(net_664), .B(net_663) );
NAND4_X1 inst_204 ( .ZN(net_428), .A1(net_358), .A2(net_343), .A4(net_291), .A3(net_217) );
NAND2_X1 inst_587 ( .A2(net_612), .ZN(net_611), .A1(net_602) );
AND4_X1 inst_666 ( .ZN(net_421), .A4(net_349), .A2(net_306), .A1(net_266), .A3(net_244) );
NOR2_X1 inst_154 ( .ZN(net_299), .A1(net_298), .A2(net_295) );
NAND2_X1 inst_592 ( .A2(net_621), .A1(net_572), .ZN(n384) );
NAND2_X1 inst_546 ( .ZN(net_488), .A1(net_449), .A2(net_429) );
NAND2_X1 inst_324 ( .A2(net_61), .ZN(net_49), .A1(n238) );
NAND2_X1 inst_465 ( .A2(net_283), .ZN(net_250), .A1(n125) );
NOR2_X1 inst_109 ( .ZN(net_12), .A2(n50), .A1(n45) );
OR3_X2 inst_54 ( .A1(net_319), .A2(net_289), .ZN(net_92), .A3(net_91) );
NAND2_X1 inst_570 ( .ZN(net_568), .A2(net_542), .A1(n330) );
NAND2_X1 inst_390 ( .A2(net_165), .ZN(net_153), .A1(n317) );
INV_X1 inst_640 ( .ZN(net_295), .A(net_265) );
XNOR2_X1 inst_43 ( .ZN(net_641), .B(net_632), .A(net_608) );
NAND2_X1 inst_359 ( .ZN(net_103), .A2(net_56), .A1(n2897) );
NAND3_X1 inst_256 ( .ZN(net_471), .A1(net_387), .A3(net_328), .A2(net_122) );
NOR4_X1 inst_94 ( .ZN(net_397), .A1(net_364), .A2(net_331), .A4(net_304), .A3(net_259) );
NAND2_X1 inst_454 ( .A2(net_254), .ZN(net_238), .A1(n303) );
INV_X1 inst_630 ( .ZN(net_6), .A(n200) );
NAND2_X1 inst_375 ( .A2(net_133), .ZN(net_132), .A1(n97) );
NAND2_X1 inst_401 ( .ZN(net_166), .A2(net_165), .A1(n150) );
NAND3_X1 inst_262 ( .ZN(net_473), .A1(net_385), .A3(net_347), .A2(net_121) );
NAND2_X1 inst_512 ( .A1(net_333), .ZN(net_330), .A2(net_182) );
NAND2_X1 inst_355 ( .A2(net_97), .ZN(net_96), .A1(n257) );
NAND3_X1 inst_243 ( .ZN(net_351), .A1(net_350), .A2(net_268), .A3(net_174) );
NAND3_X1 inst_285 ( .ZN(net_651), .A3(net_641), .A2(net_319), .A1(net_269) );
NAND2_X1 inst_591 ( .A1(net_652), .ZN(net_624), .A2(net_615) );
NAND2_X1 inst_424 ( .A1(net_633), .ZN(net_567), .A2(net_213) );
NAND2_X1 inst_497 ( .A1(net_314), .ZN(net_309), .A2(net_136) );
NAND4_X1 inst_218 ( .ZN(net_575), .A1(net_574), .A4(net_552), .A3(net_494), .A2(net_207) );
XNOR2_X1 inst_15 ( .A(net_201), .ZN(net_55), .B(n68) );
INV_X1 inst_647 ( .ZN(net_574), .A(net_567) );
NAND2_X1 inst_343 ( .A2(net_79), .ZN(net_78), .A1(n58) );
XOR2_X1 inst_6 ( .Z(net_646), .B(n390), .A(n387) );
NAND4_X1 inst_194 ( .ZN(net_364), .A2(net_363), .A4(net_264), .A3(net_255), .A1(net_249) );
NAND2_X1 inst_543 ( .A2(net_473), .ZN(net_464), .A1(net_177) );
NAND2_X1 inst_337 ( .ZN(net_108), .A2(net_64), .A1(net_6) );
AND3_X4 inst_670 ( .ZN(net_504), .A2(net_473), .A1(net_404), .A3(net_402) );
NOR2_X1 inst_123 ( .A1(net_201), .ZN(net_68), .A2(net_67) );
NAND2_X1 inst_509 ( .A1(net_333), .ZN(net_327), .A2(net_179) );
NAND2_X1 inst_299 ( .ZN(net_16), .A2(n97), .A1(n33) );
NAND2_X1 inst_418 ( .A2(net_254), .ZN(net_193), .A1(n107) );
NAND2_X1 inst_476 ( .A2(net_280), .ZN(net_263), .A1(n137) );
NOR2_X1 inst_118 ( .A1(net_73), .ZN(net_34), .A2(n1) );
OR2_X4 inst_86 ( .ZN(net_599), .A1(net_597), .A2(net_596) );
NOR2_X1 inst_153 ( .ZN(net_297), .A1(net_296), .A2(net_295) );
XNOR2_X1 inst_20 ( .A(net_276), .B(net_173), .ZN(n358) );
NAND2_X1 inst_442 ( .A2(net_254), .ZN(net_225), .A1(n150) );
INV_X1 inst_613 ( .ZN(net_298), .A(n87) );
XNOR2_X1 inst_38 ( .ZN(net_631), .B(net_630), .A(net_539) );
NAND2_X1 inst_381 ( .A2(net_168), .ZN(net_146), .A1(n58) );
NAND2_X1 inst_295 ( .ZN(net_11), .A2(n33), .A1(n283) );
NAND2_X1 inst_349 ( .ZN(net_626), .A2(net_33), .A1(n1) );
NAND2_X1 inst_483 ( .ZN(net_282), .A2(net_280), .A1(n128) );
NAND2_X1 inst_576 ( .ZN(net_582), .A1(net_553), .A2(net_541) );
NAND4_X1 inst_209 ( .ZN(net_527), .A2(net_526), .A3(net_525), .A4(net_522), .A1(net_501) );
NAND3_X1 inst_259 ( .ZN(net_481), .A1(net_391), .A3(net_330), .A2(net_124) );
XNOR2_X1 inst_40 ( .ZN(net_638), .A(n396), .B(n393) );
NAND2_X1 inst_320 ( .ZN(net_53), .A2(net_44), .A1(n13) );
NOR2_X1 inst_167 ( .ZN(net_526), .A1(net_503), .A2(net_487) );
MUX2_X2 inst_607 ( .S(net_442), .Z(net_438), .B(n200), .A(n190) );
NAND3_X1 inst_246 ( .ZN(net_406), .A2(net_374), .A3(net_310), .A1(net_230) );
INV_X1 inst_635 ( .ZN(net_535), .A(net_76) );
NOR4_X1 inst_95 ( .ZN(net_416), .A4(net_360), .A1(net_290), .A3(net_240), .A2(net_198) );
XOR2_X1 inst_1 ( .Z(net_45), .A(n270), .B(n264) );
OR2_X4 inst_72 ( .A2(net_442), .ZN(net_401), .A1(n179) );
NAND2_X1 inst_519 ( .A2(net_384), .ZN(net_383), .A1(n50) );
NAND2_X1 inst_439 ( .A2(net_283), .ZN(net_222), .A1(n150) );
NAND2_X1 inst_331 ( .ZN(net_319), .A2(net_58), .A1(n20) );
NAND2_X1 inst_582 ( .A2(net_596), .ZN(net_595), .A1(n330) );
AND2_X4 inst_683 ( .ZN(net_285), .A2(net_283), .A1(n294) );
NOR2_X1 inst_115 ( .ZN(net_61), .A2(n33), .A1(n1698) );
NAND3_X1 inst_235 ( .ZN(net_182), .A1(net_134), .A3(net_74), .A2(net_37) );
NAND4_X1 inst_210 ( .ZN(net_591), .A3(net_528), .A4(net_521), .A1(net_516), .A2(net_505) );
NAND2_X1 inst_317 ( .A2(net_205), .A1(net_120), .ZN(net_36) );
AND3_X4 inst_667 ( .ZN(net_320), .A2(net_319), .A1(net_170), .A3(net_112) );
NAND3_X1 inst_278 ( .ZN(net_620), .A2(net_619), .A1(net_617), .A3(net_616) );
NAND2_X1 inst_467 ( .A2(net_254), .ZN(net_252), .A1(n317) );
NAND3_X1 inst_239 ( .ZN(net_275), .A3(net_274), .A1(net_213), .A2(n1) );
NOR3_X1 inst_105 ( .ZN(net_596), .A2(net_576), .A3(net_570), .A1(net_551) );
NAND2_X1 inst_488 ( .A2(net_305), .ZN(net_293), .A1(n58) );
NAND2_X1 inst_387 ( .A2(net_165), .ZN(net_150), .A1(n125) );
NAND2_X1 inst_593 ( .ZN(net_627), .A1(net_626), .A2(net_625) );
NOR2_X1 inst_175 ( .ZN(net_563), .A2(net_561), .A1(net_555) );
NAND3_X1 inst_254 ( .ZN(net_423), .A3(net_367), .A1(net_322), .A2(net_184) );
INV_X1 inst_654 ( .ZN(net_560), .A(net_559) );
INV_X1 inst_625 ( .ZN(net_44), .A(n1) );
NAND3_X1 inst_225 ( .ZN(net_138), .A1(net_87), .A3(net_62), .A2(net_11) );
MUX2_X2 inst_601 ( .Z(net_443), .A(net_175), .S(net_172), .B(net_104) );
NOR2_X1 inst_133 ( .A2(net_314), .ZN(net_235), .A1(net_107) );
NAND2_X1 inst_508 ( .ZN(net_326), .A2(net_324), .A1(net_199) );
NAND2_X1 inst_568 ( .A2(net_619), .ZN(net_538), .A1(net_537) );
NOR2_X1 inst_112 ( .ZN(net_69), .A2(n41), .A1(n33) );
NAND2_X1 inst_523 ( .A2(net_389), .ZN(net_388), .A1(n87) );
NAND2_X1 inst_365 ( .A2(net_125), .ZN(net_121), .A1(net_120) );
OR2_X4 inst_67 ( .ZN(net_213), .A2(net_170), .A1(n41) );
NOR2_X1 inst_181 ( .ZN(net_605), .A1(net_591), .A2(net_589) );
NAND2_X1 inst_305 ( .ZN(net_22), .A2(n77), .A1(n20) );
NAND2_X1 inst_479 ( .ZN(net_267), .A2(net_265), .A1(n137) );
XNOR2_X1 inst_29 ( .ZN(net_583), .B(net_582), .A(net_531) );
NAND2_X1 inst_391 ( .A2(net_165), .ZN(net_154), .A1(n137) );
AND4_X1 inst_661 ( .A2(net_363), .ZN(net_358), .A4(net_258), .A1(net_243), .A3(net_225) );
NAND2_X1 inst_590 ( .ZN(net_623), .A2(net_611), .A1(net_603) );
NAND4_X1 inst_202 ( .ZN(net_378), .A1(net_377), .A3(net_361), .A4(net_356), .A2(net_166) );
NOR2_X1 inst_126 ( .ZN(net_113), .A1(net_64), .A2(net_52) );
NAND2_X1 inst_480 ( .A1(net_350), .ZN(net_277), .A2(net_276) );
INV_X1 inst_634 ( .A(net_656), .ZN(net_56) );
NAND2_X1 inst_419 ( .A2(net_280), .ZN(net_194), .A1(n107) );
NAND2_X1 inst_477 ( .A2(net_280), .ZN(net_264), .A1(n132) );
INV_X1 inst_646 ( .A(net_558), .ZN(net_465) );
NAND2_X1 inst_564 ( .A2(net_524), .ZN(net_516), .A1(net_504) );
NAND2_X1 inst_538 ( .ZN(net_457), .A1(net_455), .A2(net_422) );
NAND2_X1 inst_423 ( .A2(net_254), .ZN(net_196), .A1(n97) );
XNOR2_X1 inst_35 ( .ZN(net_625), .A(net_607), .B(net_562) );
NAND2_X1 inst_382 ( .ZN(net_359), .A2(net_168), .A1(n97) );
XNOR2_X1 inst_48 ( .B(net_663), .ZN(net_662), .A(net_659) );
NAND2_X1 inst_358 ( .ZN(net_102), .A2(net_101), .A1(n20) );
XNOR2_X1 inst_46 ( .ZN(net_659), .B(n378), .A(n375) );
NOR2_X1 inst_136 ( .A1(net_363), .ZN(net_350), .A2(net_170) );
XNOR2_X1 inst_30 ( .ZN(net_600), .A(net_593), .B(net_588) );
NAND2_X1 inst_330 ( .A2(net_61), .ZN(net_57), .A1(n222) );
MUX2_X2 inst_610 ( .Z(net_570), .S(net_558), .B(net_544), .A(net_497) );
NAND3_X1 inst_233 ( .ZN(net_180), .A1(net_130), .A3(net_66), .A2(net_22) );
NOR2_X1 inst_165 ( .ZN(net_522), .A1(net_500), .A2(net_482) );
NAND3_X1 inst_271 ( .ZN(net_496), .A3(net_468), .A1(net_381), .A2(net_380) );
NAND2_X1 inst_443 ( .A2(net_280), .ZN(net_226), .A1(n294) );
INV_X1 inst_633 ( .ZN(net_54), .A(net_53) );
XNOR2_X1 inst_34 ( .ZN(net_615), .B(net_612), .A(net_609) );
XNOR2_X1 inst_12 ( .ZN(net_91), .A(n97), .B(n107) );
NAND2_X1 inst_529 ( .A1(net_410), .ZN(net_404), .A2(net_403) );
NAND2_X1 inst_524 ( .ZN(net_390), .A2(net_389), .A1(n97) );
OR3_X2 inst_56 ( .ZN(net_426), .A1(net_368), .A3(net_341), .A2(n33) );
OR2_X4 inst_71 ( .A2(net_443), .ZN(net_380), .A1(n179) );
INV_X1 inst_655 ( .A(net_588), .ZN(net_580) );
NAND2_X1 inst_308 ( .ZN(net_26), .A2(n68), .A1(n238) );
NOR3_X1 inst_104 ( .ZN(net_470), .A3(net_447), .A1(net_445), .A2(n179) );
NAND2_X1 inst_448 ( .A2(net_231), .ZN(net_230), .A1(n226) );
OR3_X2 inst_60 ( .ZN(net_495), .A2(net_446), .A3(net_425), .A1(net_71) );
NAND2_X1 inst_455 ( .A2(net_265), .ZN(net_239), .A1(n303) );
NOR2_X1 inst_168 ( .ZN(net_523), .A1(net_504), .A2(net_474) );
AND3_X4 inst_675 ( .ZN(net_503), .A2(net_486), .A3(net_433), .A1(net_400) );
NAND2_X1 inst_384 ( .A2(net_168), .ZN(net_147), .A1(n107) );
NAND2_X1 inst_321 ( .A2(net_205), .ZN(net_43), .A1(n20) );
NAND2_X1 inst_496 ( .ZN(net_307), .A2(net_305), .A1(n143) );
INV_X1 inst_653 ( .ZN(net_545), .A(net_531) );
MUX2_X2 inst_608 ( .S(net_444), .Z(net_439), .B(n200), .A(n190) );
NAND2_X1 inst_336 ( .ZN(net_110), .A2(net_64), .A1(n200) );
NAND2_X1 inst_563 ( .ZN(net_515), .A1(net_513), .A2(net_495) );
NAND2_X1 inst_583 ( .ZN(net_598), .A1(net_597), .A2(net_596) );
NAND2_X1 inst_580 ( .A1(net_626), .A2(net_602), .ZN(net_592) );
NOR2_X1 inst_170 ( .ZN(net_518), .A1(net_507), .A2(net_480) );
NAND3_X1 inst_258 ( .ZN(net_479), .A1(net_386), .A3(net_329), .A2(net_123) );
NAND2_X1 inst_376 ( .ZN(net_134), .A2(net_133), .A1(n87) );
NAND4_X1 inst_199 ( .ZN(net_370), .A2(net_307), .A1(net_267), .A4(net_221), .A3(net_169) );
XNOR2_X1 inst_41 ( .ZN(net_644), .B(net_628), .A(net_584) );
NAND2_X1 inst_511 ( .A1(net_333), .ZN(net_329), .A2(net_180) );
NOR2_X1 inst_143 ( .A1(net_535), .A2(net_513), .ZN(net_455) );
NOR2_X1 inst_152 ( .A2(net_295), .ZN(net_292), .A1(net_201) );
NAND3_X1 inst_265 ( .ZN(net_450), .A1(net_416), .A3(net_226), .A2(net_210) );
NAND2_X1 inst_482 ( .ZN(net_281), .A2(net_280), .A1(n58) );
NAND2_X1 inst_468 ( .A2(net_254), .ZN(net_253), .A1(n143) );
AND2_X4 inst_682 ( .A2(net_265), .ZN(net_259), .A1(n143) );
NAND2_X1 inst_544 ( .A2(net_468), .ZN(net_466), .A1(net_465) );
NAND3_X1 inst_238 ( .ZN(net_273), .A1(net_128), .A3(net_102), .A2(net_72) );
NAND2_X1 inst_540 ( .A2(net_479), .A1(net_465), .ZN(net_461) );
NAND2_X1 inst_539 ( .A2(net_477), .A1(net_465), .ZN(net_460) );
NAND2_X1 inst_429 ( .A2(net_220), .ZN(net_208), .A1(n283) );
NAND2_X1 inst_404 ( .ZN(net_340), .A2(net_168), .A1(n77) );
NOR2_X1 inst_178 ( .A2(net_587), .ZN(net_584), .A1(net_576) );
OR2_X4 inst_89 ( .ZN(net_645), .A2(net_644), .A1(net_633) );
NOR2_X1 inst_111 ( .ZN(net_17), .A2(n264), .A1(n257) );
OR2_X4 inst_66 ( .ZN(net_112), .A1(net_84), .A2(net_75) );
NAND2_X1 inst_388 ( .A2(net_168), .ZN(net_151), .A1(n294) );
XOR2_X1 inst_7 ( .Z(net_663), .A(n384), .B(n381) );
NOR2_X1 inst_182 ( .ZN(net_622), .A2(net_614), .A1(net_537) );
NAND2_X1 inst_392 ( .A2(net_165), .ZN(net_155), .A1(n322) );
NOR2_X1 inst_120 ( .A1(net_363), .ZN(net_38), .A2(n1) );
NAND3_X1 inst_273 ( .ZN(net_529), .A3(net_526), .A1(net_525), .A2(net_500) );
NAND2_X1 inst_294 ( .ZN(net_10), .A2(n41), .A1(n33) );
NAND3_X1 inst_222 ( .ZN(net_374), .A1(net_172), .A3(net_109), .A2(n274) );
NAND3_X1 inst_284 ( .A2(net_652), .ZN(net_642), .A3(net_640), .A1(net_635) );
NAND2_X1 inst_489 ( .A2(net_305), .ZN(net_294), .A1(n116) );
NAND4_X1 inst_192 ( .ZN(net_360), .A3(net_359), .A4(net_339), .A2(net_159), .A1(n33) );
NAND3_X1 inst_280 ( .A3(net_610), .A1(net_592), .A2(net_566), .ZN(n393) );
NAND2_X1 inst_366 ( .A1(net_289), .A2(net_125), .ZN(net_122) );
NAND2_X1 inst_346 ( .ZN(net_214), .A2(net_36), .A1(n50) );
NAND2_X1 inst_491 ( .ZN(net_371), .A2(net_305), .A1(n87) );
NAND2_X1 inst_567 ( .A2(net_556), .ZN(net_536), .A1(net_535) );
NAND4_X1 inst_193 ( .ZN(net_362), .A3(net_361), .A4(net_336), .A2(net_162), .A1(n33) );
NOR2_X1 inst_149 ( .A2(net_295), .ZN(net_286), .A1(net_205) );
NAND2_X1 inst_318 ( .A2(net_296), .ZN(net_37), .A1(n20) );
XNOR2_X1 inst_39 ( .ZN(net_632), .A(net_630), .B(net_605) );
NAND3_X1 inst_230 ( .ZN(net_373), .A1(net_172), .A3(net_107), .A2(n274) );

endmodule
