module c6288 (
n341gat,
n409gat,
n443gat,
n205gat,
n52gat,
n392gat,
n239gat,
n154gat,
n86gat,
n69gat,
n103gat,
n307gat,
n375gat,
n256gat,
n290gat,
n324gat,
n477gat,
n358gat,
n460gat,
n273gat,
n494gat,
n222gat,
n18gat,
n35gat,
n188gat,
n528gat,
n511gat,
n426gat,
n171gat,
n120gat,
n1gat,
n137gat,
n6260gat,
n6270gat,
n3211gat,
n2877gat,
n6190gat,
n3552gat,
n6123gat,
n1901gat,
n3895gat,
n6230gat,
n6170gat,
n2223gat,
n6240gat,
n6200gat,
n5971gat,
n6288gat,
n2548gat,
n6287gat,
n4591gat,
n5672gat,
n4946gat,
n6250gat,
n6160gat,
n6220gat,
n6280gat,
n6150gat,
n4241gat,
n545gat,
n6180gat,
n1581gat,
n5308gat,
n6210gat);

// Start PIs
input n341gat;
input n409gat;
input n443gat;
input n205gat;
input n52gat;
input n392gat;
input n239gat;
input n154gat;
input n86gat;
input n69gat;
input n103gat;
input n307gat;
input n375gat;
input n256gat;
input n290gat;
input n324gat;
input n477gat;
input n358gat;
input n460gat;
input n273gat;
input n494gat;
input n222gat;
input n18gat;
input n35gat;
input n188gat;
input n528gat;
input n511gat;
input n426gat;
input n171gat;
input n120gat;
input n1gat;
input n137gat;

// Start POs
output n6260gat;
output n6270gat;
output n3211gat;
output n2877gat;
output n6190gat;
output n3552gat;
output n6123gat;
output n1901gat;
output n3895gat;
output n6230gat;
output n6170gat;
output n2223gat;
output n6240gat;
output n6200gat;
output n5971gat;
output n6288gat;
output n2548gat;
output n6287gat;
output n4591gat;
output n5672gat;
output n4946gat;
output n6250gat;
output n6160gat;
output n6220gat;
output n6280gat;
output n6150gat;
output n4241gat;
output n545gat;
output n6180gat;
output n1581gat;
output n5308gat;
output n6210gat;

// Start wires
wire net_1354;
wire net_1580;
wire net_1317;
wire net_1406;
wire net_1308;
wire net_796;
wire net_416;
wire net_215;
wire net_933;
wire net_1382;
wire net_1244;
wire net_54;
wire net_1215;
wire net_526;
wire net_943;
wire n6240gat;
wire net_834;
wire net_429;
wire net_694;
wire net_129;
wire net_1389;
wire net_648;
wire net_373;
wire net_98;
wire net_1434;
wire net_739;
wire net_980;
wire net_151;
wire net_356;
wire net_53;
wire net_1377;
wire net_1625;
wire net_452;
wire net_1570;
wire net_974;
wire net_545;
wire net_1483;
wire net_284;
wire net_560;
wire net_774;
wire net_923;
wire net_826;
wire net_439;
wire net_259;
wire net_548;
wire n443gat;
wire n52gat;
wire net_1393;
wire net_501;
wire net_1324;
wire net_1231;
wire net_187;
wire net_111;
wire net_264;
wire net_225;
wire net_636;
wire net_263;
wire net_252;
wire net_124;
wire net_343;
wire n6150gat;
wire net_1138;
wire net_160;
wire net_832;
wire net_322;
wire net_511;
wire net_1064;
wire net_815;
wire net_901;
wire net_420;
wire net_1439;
wire net_665;
wire net_447;
wire n6270gat;
wire net_1260;
wire net_871;
wire net_410;
wire net_1492;
wire net_508;
wire net_390;
wire net_35;
wire net_1185;
wire net_1154;
wire net_1090;
wire net_586;
wire net_1347;
wire net_1091;
wire net_703;
wire net_1072;
wire net_239;
wire net_193;
wire n460gat;
wire net_310;
wire net_120;
wire net_292;
wire net_201;
wire net_109;
wire net_80;
wire net_96;
wire net_167;
wire net_1132;
wire net_1490;
wire net_651;
wire net_682;
wire net_989;
wire net_280;
wire net_1538;
wire net_744;
wire net_495;
wire net_34;
wire net_458;
wire net_108;
wire net_1555;
wire net_598;
wire n6220gat;
wire net_685;
wire net_789;
wire net_971;
wire net_593;
wire net_617;
wire net_672;
wire net_777;
wire net_1007;
wire net_554;
wire net_1579;
wire net_1292;
wire net_490;
wire net_742;
wire net_1014;
wire n2223gat;
wire net_1444;
wire net_46;
wire net_584;
wire net_1441;
wire net_969;
wire net_1232;
wire net_1198;
wire net_1525;
wire net_632;
wire net_538;
wire net_165;
wire net_883;
wire net_1605;
wire net_843;
wire net_821;
wire net_1432;
wire net_464;
wire net_366;
wire net_13;
wire net_1312;
wire net_1614;
wire net_747;
wire net_446;
wire net_1359;
wire net_1516;
wire net_1171;
wire net_1540;
wire net_248;
wire net_384;
wire net_1083;
wire net_1499;
wire net_964;
wire net_1453;
wire net_198;
wire net_209;
wire net_1282;
wire net_3;
wire net_1256;
wire net_634;
wire net_294;
wire n256gat;
wire net_1413;
wire net_802;
wire n6287gat;
wire net_371;
wire net_1114;
wire net_1265;
wire net_1053;
wire net_1571;
wire net_1004;
wire net_848;
wire net_485;
wire net_1080;
wire net_997;
wire net_1619;
wire net_1031;
wire net_503;
wire net_256;
wire net_850;
wire net_1161;
wire net_1140;
wire net_82;
wire net_1464;
wire net_64;
wire net_996;
wire net_726;
wire net_679;
wire net_1168;
wire net_1028;
wire net_308;
wire net_75;
wire net_1529;
wire net_959;
wire net_515;
wire net_1334;
wire net_600;
wire net_1546;
wire net_1395;
wire net_757;
wire net_701;
wire net_206;
wire net_125;
wire net_397;
wire net_808;
wire net_223;
wire net_1009;
wire net_1589;
wire net_715;
wire net_235;
wire net_1046;
wire net_890;
wire net_606;
wire net_623;
wire net_1213;
wire net_663;
wire net_1384;
wire net_1379;
wire net_320;
wire net_1322;
wire net_579;
wire net_250;
wire net_769;
wire net_1301;
wire net_312;
wire net_986;
wire net_130;
wire net_1242;
wire net_572;
wire net_286;
wire net_147;
wire net_787;
wire net_481;
wire net_369;
wire net_1241;
wire net_403;
wire net_1079;
wire net_32;
wire net_1025;
wire net_1596;
wire net_935;
wire net_282;
wire net_1511;
wire net_1518;
wire net_645;
wire net_426;
wire net_1188;
wire net_1089;
wire net_1437;
wire net_1194;
wire net_780;
wire net_1634;
wire net_1446;
wire net_841;
wire net_609;
wire net_541;
wire net_414;
wire net_794;
wire net_1048;
wire net_1251;
wire net_799;
wire net_528;
wire net_1404;
wire net_1012;
wire net_456;
wire net_155;
wire net_705;
wire net_1608;
wire net_335;
wire net_1468;
wire net_907;
wire net_506;
wire net_181;
wire net_1221;
wire net_349;
wire n6160gat;
wire net_39;
wire net_1036;
wire net_245;
wire net_1409;
wire net_395;
wire net_331;
wire net_1130;
wire net_493;
wire net_1196;
wire net_816;
wire net_386;
wire net_1428;
wire net_987;
wire net_641;
wire net_277;
wire net_919;
wire net_89;
wire net_1152;
wire net_1226;
wire net_1217;
wire net_290;
wire net_1508;
wire net_680;
wire net_931;
wire net_1372;
wire net_338;
wire net_1039;
wire n545gat;
wire net_721;
wire net_243;
wire net_400;
wire net_759;
wire net_1018;
wire net_602;
wire net_1575;
wire net_175;
wire net_657;
wire net_823;
wire net_1497;
wire net_106;
wire net_1380;
wire net_140;
wire net_740;
wire net_247;
wire net_329;
wire net_279;
wire net_1523;
wire net_1177;
wire net_1163;
wire net_1259;
wire net_698;
wire net_897;
wire net_25;
wire net_1191;
wire net_70;
wire net_691;
wire net_194;
wire net_1341;
wire net_962;
wire net_730;
wire net_615;
wire net_478;
wire net_1128;
wire net_1559;
wire net_441;
wire net_1620;
wire net_596;
wire net_1127;
wire net_138;
wire net_749;
wire net_1261;
wire net_1019;
wire net_804;
wire net_333;
wire net_1616;
wire net_639;
wire net_1119;
wire net_728;
wire net_1314;
wire net_957;
wire net_1287;
wire net_1276;
wire net_1006;
wire net_719;
wire n494gat;
wire net_1238;
wire net_170;
wire net_531;
wire net_471;
wire net_565;
wire net_499;
wire net_77;
wire net_1055;
wire net_20;
wire net_1531;
wire net_878;
wire net_1340;
wire net_1159;
wire net_1033;
wire net_49;
wire net_518;
wire net_861;
wire net_15;
wire net_57;
wire net_71;
wire net_771;
wire net_929;
wire net_1418;
wire n307gat;
wire net_1;
wire net_708;
wire net_696;
wire net_537;
wire net_180;
wire net_1565;
wire net_1361;
wire net_367;
wire net_169;
wire net_51;
wire net_171;
wire net_432;
wire net_1062;
wire net_1208;
wire net_1475;
wire net_1460;
wire net_1142;
wire net_513;
wire net_204;
wire net_1451;
wire net_232;
wire net_604;
wire net_163;
wire net_967;
wire net_1576;
wire net_1421;
wire net_67;
wire net_1180;
wire net_1527;
wire net_1627;
wire net_268;
wire net_1280;
wire net_459;
wire net_1069;
wire net_483;
wire net_48;
wire net_8;
wire net_1149;
wire net_737;
wire net_1411;
wire net_203;
wire net_505;
wire net_176;
wire net_1602;
wire net_1298;
wire net_1416;
wire net_137;
wire net_296;
wire net_992;
wire net_613;
wire net_237;
wire net_782;
wire net_614;
wire net_532;
wire net_1601;
wire net_1156;
wire net_1123;
wire net_93;
wire net_1095;
wire net_578;
wire net_786;
wire net_302;
wire net_1192;
wire net_1131;
wire net_889;
wire net_127;
wire net_1116;
wire net_1558;
wire net_1339;
wire net_984;
wire net_348;
wire net_753;
wire net_1505;
wire net_626;
wire net_1105;
wire net_101;
wire net_906;
wire net_388;
wire net_1272;
wire net_326;
wire net_707;
wire net_589;
wire net_100;
wire n4946gat;
wire net_655;
wire net_686;
wire net_652;
wire net_536;
wire net_1615;
wire net_455;
wire net_1332;
wire net_1594;
wire net_221;
wire net_115;
wire net_1110;
wire net_689;
wire net_751;
wire n120gat;
wire net_393;
wire net_442;
wire net_830;
wire net_542;
wire net_575;
wire net_1279;
wire net_877;
wire net_595;
wire net_378;
wire net_408;
wire net_1320;
wire net_1047;
wire net_724;
wire net_1026;
wire net_423;
wire net_1466;
wire net_1219;
wire net_328;
wire net_1520;
wire net_157;
wire net_42;
wire net_1228;
wire net_1549;
wire net_1205;
wire net_1474;
wire net_1467;
wire net_1401;
wire net_1061;
wire net_874;
wire net_1588;
wire net_66;
wire net_466;
wire net_1632;
wire net_1495;
wire net_1179;
wire net_868;
wire net_765;
wire net_675;
wire net_1342;
wire net_1236;
wire net_1426;
wire net_818;
wire net_1407;
wire net_938;
wire net_1610;
wire net_443;
wire n477gat;
wire net_922;
wire net_522;
wire net_270;
wire n6280gat;
wire net_183;
wire net_1211;
wire net_668;
wire net_1440;
wire net_1183;
wire n18gat;
wire net_1057;
wire net_150;
wire net_1584;
wire net_1488;
wire net_304;
wire net_1011;
wire net_811;
wire net_352;
wire net_1355;
wire n2877gat;
wire net_800;
wire net_977;
wire net_644;
wire net_30;
wire net_643;
wire net_1070;
wire net_1068;
wire net_1462;
wire net_852;
wire net_436;
wire net_1225;
wire net_24;
wire n6200gat;
wire net_622;
wire net_186;
wire net_812;
wire n273gat;
wire net_1050;
wire net_1042;
wire net_1316;
wire net_1385;
wire net_1107;
wire net_1534;
wire net_1621;
wire net_792;
wire net_1000;
wire net_1338;
wire net_1103;
wire net_1035;
wire net_1016;
wire net_767;
wire net_1607;
wire net_1203;
wire net_825;
wire net_219;
wire net_18;
wire net_309;
wire net_1263;
wire net_659;
wire net_131;
wire net_196;
wire net_913;
wire net_29;
wire net_1366;
wire net_358;
wire net_837;
wire net_899;
wire net_1010;
wire net_516;
wire net_31;
wire net_1479;
wire net_927;
wire net_1151;
wire net_956;
wire n3552gat;
wire net_1285;
wire net_713;
wire net_1519;
wire net_693;
wire net_360;
wire net_1175;
wire net_213;
wire net_729;
wire net_863;
wire net_260;
wire net_947;
wire net_438;
wire net_1513;
wire net_1126;
wire net_732;
wire net_580;
wire net_314;
wire net_1325;
wire net_904;
wire net_341;
wire net_1597;
wire net_1373;
wire net_1352;
wire net_952;
wire net_468;
wire net_58;
wire net_1187;
wire net_970;
wire net_798;
wire net_488;
wire n290gat;
wire net_73;
wire net_807;
wire net_1303;
wire net_86;
wire net_1532;
wire net_1503;
wire net_1160;
wire net_1336;
wire net_945;
wire n6260gat;
wire net_179;
wire net_159;
wire net_61;
wire net_1442;
wire net_449;
wire net_383;
wire net_62;
wire net_6;
wire net_553;
wire net_534;
wire net_217;
wire net_1087;
wire net_733;
wire net_1093;
wire net_887;
wire net_903;
wire net_1551;
wire net_763;
wire net_427;
wire net_486;
wire net_135;
wire net_915;
wire net_1121;
wire net_1560;
wire net_473;
wire n6210gat;
wire net_406;
wire n409gat;
wire net_633;
wire net_324;
wire net_113;
wire net_710;
wire net_1049;
wire net_497;
wire net_454;
wire net_462;
wire net_418;
wire net_40;
wire net_872;
wire net_1296;
wire net_1424;
wire n358gat;
wire net_1414;
wire net_709;
wire net_161;
wire net_300;
wire net_1165;
wire net_1066;
wire net_1545;
wire net_1457;
wire net_1233;
wire net_748;
wire net_677;
wire net_95;
wire net_1486;
wire net_1472;
wire net_173;
wire net_78;
wire net_1113;
wire net_990;
wire net_950;
wire net_1436;
wire net_1344;
wire net_1003;
wire net_514;
wire net_1283;
wire net_1084;
wire net_22;
wire net_376;
wire net_1604;
wire net_1500;
wire net_354;
wire net_524;
wire net_1136;
wire net_1134;
wire net_646;
wire net_363;
wire net_445;
wire net_573;
wire net_1391;
wire net_1319;
wire net_1214;
wire net_776;
wire net_866;
wire net_44;
wire net_784;
wire net_1582;
wire net_520;
wire net_422;
wire net_1345;
wire net_1450;
wire net_1032;
wire net_561;
wire net_567;
wire net_45;
wire net_381;
wire net_591;
wire net_746;
wire net_1368;
wire net_981;
wire net_1592;
wire net_272;
wire net_1248;
wire net_1274;
wire net_1097;
wire net_178;
wire net_845;
wire net_1024;
wire net_1590;
wire net_1566;
wire net_762;
wire net_1305;
wire net_1612;
wire net_695;
wire net_839;
wire net_1387;
wire net_1318;
wire net_1201;
wire net_814;
wire net_1581;
wire net_556;
wire net_941;
wire net_893;
wire net_809;
wire net_629;
wire net_55;
wire net_1557;
wire net_559;
wire net_635;
wire n6288gat;
wire net_255;
wire net_1235;
wire net_266;
wire net_1514;
wire net_1037;
wire net_345;
wire net_859;
wire net_620;
wire net_619;
wire net_350;
wire net_1167;
wire net_398;
wire net_1599;
wire net_306;
wire net_954;
wire net_1044;
wire net_1290;
wire net_500;
wire net_1350;
wire net_1626;
wire net_1258;
wire net_1623;
wire net_631;
wire net_11;
wire n324gat;
wire net_1329;
wire net_123;
wire net_1101;
wire net_994;
wire net_1572;
wire net_527;
wire net_262;
wire net_362;
wire net_68;
wire net_318;
wire net_1052;
wire net_1493;
wire net_976;
wire net_316;
wire net_865;
wire net_84;
wire net_670;
wire net_611;
wire net_231;
wire n2548gat;
wire net_103;
wire net_1124;
wire net_226;
wire net_1021;
wire net_1223;
wire net_228;
wire net_926;
wire n1gat;
wire net_966;
wire net_143;
wire net_190;
wire net_1447;
wire net_391;
wire net_1002;
wire net_533;
wire net_145;
wire net_1108;
wire net_911;
wire net_1617;
wire net_1145;
wire net_37;
wire net_582;
wire net_188;
wire net_1553;
wire net_755;
wire net_509;
wire net_661;
wire net_881;
wire net_211;
wire net_133;
wire net_1397;
wire net_1077;
wire net_568;
wire net_47;
wire net_1141;
wire net_1227;
wire net_1008;
wire net_1543;
wire net_1295;
wire net_1443;
wire net_557;
wire net_1288;
wire net_119;
wire net_1275;
wire net_210;
wire net_1429;
wire net_1321;
wire net_168;
wire net_916;
wire net_741;
wire net_1611;
wire net_477;
wire net_940;
wire net_1173;
wire net_385;
wire net_269;
wire net_851;
wire net_1209;
wire net_1431;
wire net_1099;
wire net_469;
wire n392gat;
wire net_1170;
wire net_727;
wire net_847;
wire net_90;
wire net_1043;
wire net_671;
wire net_283;
wire net_85;
wire net_778;
wire net_404;
wire net_770;
wire net_1455;
wire net_1005;
wire net_240;
wire net_1200;
wire net_4;
wire net_1059;
wire net_1630;
wire net_295;
wire net_895;
wire net_1454;
wire net_1239;
wire net_307;
wire net_1082;
wire net_1463;
wire net_344;
wire net_16;
wire net_1412;
wire net_1550;
wire net_884;
wire net_712;
wire net_1507;
wire net_1422;
wire net_257;
wire net_233;
wire net_1255;
wire n4241gat;
wire net_474;
wire net_1562;
wire net_1106;
wire net_472;
wire net_1628;
wire net_1510;
wire net_65;
wire net_958;
wire net_1394;
wire net_1250;
wire net_1481;
wire net_1268;
wire net_995;
wire net_484;
wire net_896;
wire net_1281;
wire net_1115;
wire net_136;
wire net_207;
wire net_944;
wire net_1524;
wire net_700;
wire net_961;
wire net_1528;
wire n69gat;
wire net_1246;
wire net_126;
wire net_278;
wire net_1547;
wire net_571;
wire net_63;
wire net_1162;
wire net_274;
wire net_601;
wire net_1362;
wire net_1075;
wire n205gat;
wire net_321;
wire net_425;
wire net_1307;
wire net_287;
wire net_189;
wire net_1586;
wire net_829;
wire net_833;
wire net_930;
wire net_720;
wire net_99;
wire net_480;
wire net_216;
wire net_934;
wire net_433;
wire net_836;
wire net_544;
wire net_717;
wire net_900;
wire net_1405;
wire n5308gat;
wire net_368;
wire net_224;
wire net_1399;
wire net_684;
wire net_52;
wire net_608;
wire net_1212;
wire net_370;
wire net_510;
wire net_1353;
wire net_1595;
wire net_413;
wire net_1120;
wire net_1020;
wire net_1491;
wire net_716;
wire net_114;
wire net_1269;
wire net_1169;
wire net_973;
wire net_1300;
wire net_1139;
wire net_1034;
wire net_1245;
wire net_1252;
wire net_36;
wire net_860;
wire net_1392;
wire net_870;
wire net_1574;
wire net_253;
wire net_637;
wire net_276;
wire net_311;
wire net_1449;
wire net_494;
wire net_760;
wire net_547;
wire net_873;
wire net_1098;
wire net_154;
wire net_666;
wire net_507;
wire net_616;
wire net_1220;
wire net_238;
wire net_1509;
wire net_817;
wire net_28;
wire net_529;
wire net_704;
wire net_1478;
wire net_587;
wire net_1262;
wire net_97;
wire net_192;
wire n6190gat;
wire net_649;
wire net_793;
wire net_1356;
wire net_1591;
wire net_460;
wire net_1374;
wire net_1164;
wire net_650;
wire net_291;
wire net_457;
wire net_735;
wire net_772;
wire net_857;
wire net_121;
wire net_867;
wire net_200;
wire net_597;
wire net_1367;
wire net_743;
wire net_1133;
wire net_396;
wire net_195;
wire net_1081;
wire n341gat;
wire net_166;
wire net_107;
wire net_1277;
wire net_1237;
wire net_530;
wire net_1541;
wire net_1420;
wire n3895gat;
wire net_849;
wire net_1371;
wire net_594;
wire net_603;
wire net_23;
wire net_271;
wire net_117;
wire net_74;
wire net_673;
wire net_401;
wire net_642;
wire net_1522;
wire net_205;
wire net_1286;
wire net_1158;
wire net_699;
wire net_242;
wire net_359;
wire net_440;
wire net_1445;
wire net_26;
wire net_470;
wire net_758;
wire net_920;
wire n6170gat;
wire net_334;
wire net_1410;
wire net_1461;
wire net_430;
wire net_1073;
wire net_365;
wire net_718;
wire net_882;
wire net_820;
wire net_380;
wire net_141;
wire net_1190;
wire net_467;
wire net_83;
wire net_879;
wire net_1118;
wire net_1556;
wire net_1311;
wire net_372;
wire net_1207;
wire net_437;
wire net_1270;
wire net_56;
wire net_566;
wire net_1552;
wire net_1063;
wire net_968;
wire net_336;
wire net_803;
wire net_1348;
wire net_624;
wire net_555;
wire net_1578;
wire net_2;
wire net_9;
wire net_1613;
wire net_1476;
wire net_1293;
wire net_298;
wire net_790;
wire net_1504;
wire net_688;
wire net_697;
wire net_998;
wire net_475;
wire net_1577;
wire net_563;
wire net_1417;
wire net_1147;
wire net_1054;
wire n3211gat;
wire net_605;
wire net_199;
wire net_502;
wire net_431;
wire net_1564;
wire net_1568;
wire net_835;
wire net_1181;
wire net_924;
wire net_1526;
wire net_1266;
wire net_898;
wire net_1452;
wire net_1357;
wire net_638;
wire net_1333;
wire net_909;
wire net_222;
wire net_1593;
wire net_152;
wire net_313;
wire net_932;
wire net_489;
wire net_714;
wire net_1309;
wire net_1243;
wire net_1484;
wire net_683;
wire net_258;
wire net_607;
wire n5672gat;
wire net_148;
wire net_1376;
wire net_1517;
wire net_1045;
wire net_419;
wire n171gat;
wire net_1360;
wire net_251;
wire net_972;
wire net_1302;
wire net_244;
wire net_664;
wire net_128;
wire net_585;
wire net_936;
wire net_840;
wire net_819;
wire net_1364;
wire net_1438;
wire net_1078;
wire net_549;
wire net_827;
wire net_374;
wire net_785;
wire net_1143;
wire net_1489;
wire net_411;
wire net_854;
wire net_788;
wire net_214;
wire net_1539;
wire net_1369;
wire net_249;
wire net_1088;
wire net_1349;
wire net_979;
wire net_706;
wire net_156;
wire net_1013;
wire net_1530;
wire net_1548;
wire net_112;
wire net_92;
wire net_394;
wire net_810;
wire net_842;
wire net_1264;
wire net_1189;
wire net_139;
wire net_1040;
wire net_551;
wire net_332;
wire net_409;
wire net_1469;
wire n6180gat;
wire n1581gat;
wire net_1229;
wire net_463;
wire net_492;
wire net_656;
wire net_88;
wire net_1536;
wire net_197;
wire net_766;
wire net_81;
wire net_1609;
wire net_1498;
wire net_1381;
wire net_1153;
wire n86gat;
wire net_402;
wire net_1327;
wire net_1199;
wire net_202;
wire net_110;
wire net_379;
wire net_722;
wire net_1569;
wire net_33;
wire net_1403;
wire net_1383;
wire net_988;
wire net_918;
wire net_1254;
wire net_949;
wire net_289;
wire net_450;
wire net_621;
wire net_435;
wire net_1606;
wire net_1386;
wire net_132;
wire net_105;
wire net_1358;
wire net_12;
wire net_1249;
wire net_978;
wire net_1313;
wire net_1129;
wire net_1071;
wire net_1056;
wire net_1224;
wire net_1430;
wire net_569;
wire net_768;
wire net_1017;
wire net_955;
wire net_1206;
wire net_357;
wire net_327;
wire net_1284;
wire n6123gat;
wire net_960;
wire net_630;
wire net_999;
wire net_76;
wire net_1166;
wire net_1029;
wire net_908;
wire net_353;
wire net_822;
wire net_519;
wire net_801;
wire net_1633;
wire net_412;
wire net_1471;
wire net_838;
wire n426gat;
wire net_1480;
wire net_319;
wire net_17;
wire net_453;
wire net_1598;
wire net_581;
wire net_164;
wire net_377;
wire net_731;
wire net_1146;
wire net_87;
wire net_1544;
wire net_288;
wire net_0;
wire net_1038;
wire net_912;
wire net_658;
wire net_1629;
wire net_1459;
wire net_1204;
wire net_805;
wire net_734;
wire net_540;
wire net_512;
wire net_662;
wire net_779;
wire net_862;
wire net_1174;
wire net_1622;
wire net_891;
wire net_951;
wire net_50;
wire net_1328;
wire net_1109;
wire net_806;
wire net_234;
wire net_38;
wire net_342;
wire n1901gat;
wire net_975;
wire net_612;
wire net_19;
wire net_738;
wire n103gat;
wire net_892;
wire net_946;
wire net_1176;
wire net_1150;
wire net_1102;
wire net_1094;
wire net_504;
wire net_855;
wire net_1253;
wire net_674;
wire net_618;
wire net_1076;
wire net_303;
wire net_1331;
wire net_1537;
wire net_491;
wire net_965;
wire net_681;
wire net_1299;
wire net_1148;
wire net_948;
wire net_783;
wire net_1448;
wire net_392;
wire net_118;
wire net_1487;
wire net_1195;
wire net_754;
wire net_421;
wire net_1561;
wire net_1396;
wire net_146;
wire net_1104;
wire net_921;
wire net_550;
wire net_764;
wire net_417;
wire net_122;
wire net_876;
wire net_7;
wire n528gat;
wire net_172;
wire net_1502;
wire net_1533;
wire net_1117;
wire net_1458;
wire n6230gat;
wire net_1240;
wire net_428;
wire net_246;
wire net_94;
wire net_461;
wire net_1186;
wire net_640;
wire net_482;
wire net_991;
wire net_905;
wire net_1060;
wire net_1512;
wire net_775;
wire net_1378;
wire net_149;
wire net_142;
wire n35gat;
wire net_752;
wire net_387;
wire net_654;
wire net_1600;
wire net_1473;
wire net_330;
wire net_858;
wire net_498;
wire net_535;
wire net_888;
wire net_1330;
wire net_158;
wire net_676;
wire net_41;
wire net_577;
wire net_570;
wire net_444;
wire net_525;
wire net_1023;
wire net_844;
wire net_1496;
wire net_1216;
wire net_1210;
wire net_1067;
wire net_325;
wire net_797;
wire net_301;
wire net_1427;
wire net_1271;
wire net_1086;
wire net_1363;
wire net_299;
wire net_1343;
wire n511gat;
wire net_985;
wire net_182;
wire net_60;
wire net_521;
wire net_1197;
wire net_337;
wire net_590;
wire net_267;
wire net_1585;
wire net_1278;
wire net_273;
wire net_424;
wire net_1567;
wire net_576;
wire net_690;
wire net_1521;
wire net_465;
wire net_177;
wire net_523;
wire net_1435;
wire net_1370;
wire net_407;
wire net_476;
wire net_564;
wire net_382;
wire net_725;
wire net_1315;
wire net_583;
wire net_813;
wire net_1178;
wire n239gat;
wire net_953;
wire net_1306;
wire net_351;
wire net_1027;
wire net_894;
wire net_1074;
wire net_1058;
wire net_1041;
wire net_1423;
wire net_340;
wire net_1408;
wire net_1388;
wire net_265;
wire net_517;
wire net_434;
wire net_628;
wire net_791;
wire net_1257;
wire net_1419;
wire net_939;
wire net_1465;
wire net_220;
wire net_14;
wire net_824;
wire net_1051;
wire net_293;
wire net_942;
wire net_1631;
wire net_1337;
wire net_1202;
wire net_1182;
wire net_69;
wire net_1624;
wire net_543;
wire net_1155;
wire n222gat;
wire net_1515;
wire net_925;
wire net_1218;
wire net_625;
wire net_1573;
wire net_339;
wire net_993;
wire net_1494;
wire net_361;
wire net_864;
wire net_1289;
wire net_27;
wire net_317;
wire net_305;
wire net_856;
wire net_1100;
wire net_880;
wire net_1402;
wire net_261;
wire net_191;
wire net_1398;
wire net_558;
wire net_1125;
wire net_660;
wire net_1618;
wire net_227;
wire net_102;
wire net_144;
wire net_59;
wire net_1144;
wire net_162;
wire net_1001;
wire net_781;
wire net_1291;
wire net_230;
wire net_653;
wire net_910;
wire net_1326;
wire net_134;
wire net_1022;
wire net_678;
wire net_546;
wire net_1415;
wire n375gat;
wire net_185;
wire net_702;
wire net_588;
wire net_1477;
wire net_1222;
wire net_928;
wire net_1230;
wire net_1157;
wire net_667;
wire net_853;
wire net_236;
wire net_208;
wire net_1375;
wire net_1015;
wire net_315;
wire net_212;
wire n137gat;
wire net_487;
wire net_552;
wire net_914;
wire net_1542;
wire net_1433;
wire net_415;
wire net_1172;
wire net_1351;
wire net_116;
wire net_347;
wire net_1535;
wire net_346;
wire net_297;
wire net_91;
wire net_756;
wire net_1193;
wire net_1425;
wire net_1122;
wire net_875;
wire net_104;
wire net_1065;
wire net_448;
wire net_1335;
wire net_72;
wire net_886;
wire net_229;
wire net_1092;
wire net_627;
wire net_241;
wire net_687;
wire net_917;
wire net_5;
wire net_405;
wire net_1111;
wire net_983;
wire net_355;
wire net_184;
wire n5971gat;
wire net_599;
wire net_711;
wire net_610;
wire net_1470;
wire net_1456;
wire net_723;
wire net_389;
wire net_831;
wire net_902;
wire net_451;
wire net_1323;
wire net_323;
wire net_1506;
wire net_963;
wire net_1234;
wire net_750;
wire net_846;
wire net_1583;
wire net_275;
wire net_736;
wire net_399;
wire net_539;
wire net_692;
wire net_1184;
wire net_1563;
wire net_153;
wire net_1390;
wire net_218;
wire net_174;
wire net_1112;
wire net_1273;
wire net_375;
wire net_562;
wire net_1365;
wire net_1135;
wire net_1137;
wire net_364;
wire n6250gat;
wire net_1346;
wire net_43;
wire net_1085;
wire net_10;
wire net_1482;
wire net_592;
wire net_21;
wire n188gat;
wire net_1400;
wire net_79;
wire net_647;
wire net_885;
wire net_1267;
wire net_1030;
wire net_1485;
wire net_773;
wire net_285;
wire net_281;
wire net_828;
wire net_869;
wire net_1603;
wire net_1310;
wire n154gat;
wire net_669;
wire net_254;
wire net_937;
wire n4591gat;
wire net_1501;
wire net_1297;
wire net_496;
wire net_761;
wire net_1554;
wire net_1304;
wire net_479;
wire net_574;
wire net_1096;
wire net_1294;
wire net_795;
wire net_982;
wire net_1247;
wire net_1587;
wire net_745;

// Start cells
INV_X1 inst_1574 ( .ZN(net_1241), .A(net_1240) );
NAND2_X1 inst_696 ( .ZN(net_324), .A2(n341gat), .A1(n239gat) );
NAND2_X1 inst_1175 ( .ZN(net_1131), .A1(net_1130), .A2(net_1102) );
NOR2_X1 inst_481 ( .ZN(net_120), .A2(net_35), .A1(net_2) );
XNOR2_X1 inst_228 ( .ZN(net_903), .B(net_869), .A(net_835) );
XNOR2_X1 inst_125 ( .ZN(net_522), .B(net_474), .A(net_443) );
NOR2_X1 inst_486 ( .ZN(net_56), .A2(net_55), .A1(net_1) );
NAND2_X1 inst_1240 ( .ZN(net_1276), .A1(net_1275), .A2(net_1250) );
NAND2_X1 inst_1025 ( .ZN(net_798), .A2(net_741), .A1(net_712) );
NAND2_X1 inst_707 ( .ZN(net_375), .A2(n341gat), .A1(n205gat) );
NAND2_X1 inst_779 ( .ZN(net_119), .A2(net_118), .A1(net_70) );
XNOR2_X1 inst_395 ( .ZN(net_1506), .B(net_1466), .A(net_1453) );
NAND2_X1 inst_841 ( .ZN(net_359), .A1(net_358), .A2(net_357) );
XNOR2_X1 inst_244 ( .ZN(net_954), .A(net_921), .B(net_886) );
AND2_X4 inst_1636 ( .ZN(net_6), .A2(n273gat), .A1(n188gat) );
OR2_X4 inst_452 ( .ZN(net_173), .A1(net_172), .A2(net_171) );
NAND2_X1 inst_689 ( .ZN(net_24), .A1(n69gat), .A2(n273gat) );
XNOR2_X1 inst_430 ( .ZN(net_1621), .B(net_1575), .A(net_1560) );
INV_X1 inst_1521 ( .ZN(net_889), .A(net_888) );
XNOR2_X1 inst_214 ( .ZN(net_856), .A(net_809), .B(net_780) );
AND2_X4 inst_1629 ( .ZN(net_11), .A2(n290gat), .A1(n103gat) );
INV_X1 inst_1558 ( .ZN(net_1135), .A(net_1134) );
NAND2_X1 inst_548 ( .ZN(net_146), .A2(n307gat), .A1(n18gat) );
NOR2_X1 inst_515 ( .ZN(net_195), .A2(net_129), .A1(net_103) );
INV_X1 inst_1501 ( .ZN(net_771), .A(net_770) );
NAND2_X1 inst_1306 ( .ZN(net_1438), .A2(net_1437), .A1(net_1388) );
NAND2_X1 inst_772 ( .ZN(net_44), .A1(net_27), .A2(net_26) );
NAND2_X1 inst_728 ( .ZN(net_905), .A2(n426gat), .A1(n103gat) );
NAND2_X1 inst_944 ( .ZN(net_593), .A1(net_592), .A2(net_568) );
INV_X1 inst_1407 ( .ZN(net_76), .A(net_75) );
INV_X1 inst_1584 ( .ZN(net_1323), .A(net_1322) );
INV_X1 inst_1615 ( .ZN(net_1518), .A(net_1517) );
NAND2_X1 inst_642 ( .ZN(net_248), .A2(n324gat), .A1(n137gat) );
OR2_X4 inst_459 ( .ZN(net_196), .A1(net_195), .A2(net_194) );
NAND2_X1 inst_1018 ( .ZN(net_759), .A1(net_758), .A2(net_757) );
XNOR2_X1 inst_445 ( .A(net_1624), .B(net_1623), .ZN(n6260gat) );
NAND2_X1 inst_850 ( .ZN(net_394), .A2(net_342), .A1(net_290) );
NAND2_X1 inst_709 ( .ZN(net_1556), .A2(n528gat), .A1(n120gat) );
XNOR2_X1 inst_93 ( .ZN(net_385), .B(net_355), .A(net_354) );
NAND2_X1 inst_700 ( .ZN(net_455), .A1(n86gat), .A2(n358gat) );
NAND2_X1 inst_920 ( .ZN(net_521), .A1(net_520), .A2(net_519) );
NAND2_X1 inst_606 ( .ZN(net_690), .A2(n392gat), .A1(n137gat) );
XNOR2_X1 inst_367 ( .ZN(net_1374), .B(net_1355), .A(net_1343) );
NAND2_X1 inst_957 ( .ZN(net_631), .A1(net_591), .A2(net_524) );
NAND2_X1 inst_1228 ( .ZN(net_1255), .A1(net_1254), .A2(net_1253) );
NAND2_X1 inst_979 ( .ZN(net_702), .A1(net_651), .A2(net_602) );
NAND2_X1 inst_853 ( .ZN(net_402), .A2(net_359), .A1(net_307) );
NAND2_X1 inst_1259 ( .ZN(net_1359), .A1(net_1293), .A2(net_1280) );
NAND2_X1 inst_1008 ( .ZN(net_728), .A1(net_727), .A2(net_726) );
XNOR2_X1 inst_139 ( .ZN(net_567), .A(net_526), .B(net_525) );
NAND2_X1 inst_657 ( .ZN(net_1295), .A1(n69gat), .A2(n494gat) );
NAND2_X1 inst_559 ( .ZN(net_735), .A2(n409gat), .A1(n35gat) );
NAND2_X1 inst_584 ( .ZN(net_813), .A2(n409gat), .A1(n137gat) );
NOR2_X1 inst_521 ( .ZN(net_189), .A2(net_144), .A1(net_121) );
NAND2_X1 inst_1316 ( .ZN(net_1496), .A2(net_1429), .A1(net_1380) );
NOR2_X1 inst_470 ( .ZN(net_31), .A1(net_17), .A2(net_16) );
AND2_X4 inst_1655 ( .ZN(net_135), .A1(net_134), .A2(net_133) );
NAND2_X1 inst_535 ( .ZN(net_369), .A2(n341gat), .A1(n188gat) );
OR2_X4 inst_450 ( .ZN(net_112), .A2(net_90), .A1(net_56) );
NAND2_X1 inst_745 ( .ZN(net_352), .A1(n69gat), .A2(n341gat) );
NOR2_X1 inst_520 ( .ZN(net_175), .A2(net_159), .A1(net_95) );
XNOR2_X1 inst_237 ( .ZN(net_930), .B(net_894), .A(net_867) );
XNOR2_X1 inst_148 ( .ZN(net_611), .B(net_573), .A(net_541) );
NAND2_X1 inst_554 ( .ZN(net_807), .A2(n409gat), .A1(n188gat) );
NAND2_X1 inst_1187 ( .ZN(net_1156), .A1(net_1155), .A2(net_1154) );
XNOR2_X1 inst_191 ( .ZN(net_793), .B(net_724), .A(net_700) );
NAND2_X1 inst_1063 ( .ZN(net_860), .A1(net_859), .A2(net_786) );
NAND2_X1 inst_813 ( .ZN(net_288), .A1(net_287), .A2(net_286) );
XNOR2_X1 inst_51 ( .ZN(net_220), .B(net_204), .A(net_203) );
XNOR2_X1 inst_315 ( .ZN(net_1194), .A(net_1183), .B(net_1149) );
XNOR2_X1 inst_80 ( .ZN(net_357), .A(net_306), .B(net_283) );
NAND2_X1 inst_836 ( .ZN(net_347), .A1(net_346), .A2(net_345) );
NAND2_X1 inst_1066 ( .ZN(net_896), .A2(net_838), .A1(net_790) );
INV_X1 inst_1556 ( .ZN(net_1102), .A(net_1101) );
NAND2_X1 inst_974 ( .ZN(net_656), .A1(net_655), .A2(net_654) );
XNOR2_X1 inst_216 ( .ZN(net_825), .B(net_801), .A(net_800) );
NAND2_X1 inst_1059 ( .ZN(net_877), .A1(net_841), .A2(net_799) );
XNOR2_X1 inst_241 ( .ZN(net_932), .B(net_900), .A(net_899) );
NAND2_X1 inst_1075 ( .ZN(net_898), .A1(net_897), .A2(net_896) );
NAND2_X1 inst_862 ( .ZN(net_424), .A2(net_376), .A1(net_296) );
NAND2_X1 inst_1167 ( .ZN(net_1115), .A1(net_1114), .A2(net_1113) );
INV_X1 inst_1617 ( .ZN(net_1535), .A(net_1534) );
NAND2_X1 inst_1116 ( .ZN(net_1018), .A2(net_961), .A1(net_904) );
XNOR2_X1 inst_151 ( .ZN(net_630), .B(net_588), .A(net_563) );
XNOR2_X1 inst_64 ( .ZN(net_282), .B(net_268), .A(net_222) );
NAND2_X1 inst_1001 ( .ZN(net_748), .A2(net_695), .A1(net_635) );
NAND2_X1 inst_743 ( .ZN(net_724), .A2(n409gat), .A1(n239gat) );
XNOR2_X1 inst_415 ( .ZN(net_1566), .B(net_1524), .A(net_1473) );
NAND2_X1 inst_828 ( .ZN(net_309), .A1(net_308), .A2(net_278) );
NAND2_X1 inst_1303 ( .ZN(net_1432), .A1(net_1431), .A2(net_1430) );
NAND2_X1 inst_1104 ( .ZN(net_959), .A1(net_958), .A2(net_933) );
NAND2_X1 inst_892 ( .ZN(net_475), .A1(net_474), .A2(net_444) );
INV_X1 inst_1623 ( .ZN(net_1563), .A(net_1562) );
XNOR2_X1 inst_223 ( .ZN(net_867), .B(net_833), .A(net_832) );
NAND2_X1 inst_1159 ( .ZN(net_1098), .A1(net_1097), .A2(net_1069) );
NAND2_X1 inst_1132 ( .ZN(net_1033), .A1(net_1032), .A2(net_1031) );
INV_X1 inst_1603 ( .ZN(net_1443), .A(net_1442) );
XNOR2_X1 inst_402 ( .ZN(net_1515), .B(net_1469), .A(net_1468) );
NAND2_X1 inst_968 ( .ZN(net_638), .A1(net_637), .A2(net_636) );
NAND2_X1 inst_819 ( .ZN(net_294), .A2(net_259), .A1(net_190) );
XNOR2_X1 inst_340 ( .ZN(net_1268), .B(net_1245), .A(net_1244) );
INV_X1 inst_1468 ( .ZN(net_542), .A(net_541) );
INV_X1 inst_1516 ( .ZN(net_872), .A(net_871) );
NOR2_X1 inst_494 ( .A2(net_92), .ZN(net_73), .A1(net_54) );
XNOR2_X1 inst_329 ( .ZN(net_1244), .B(net_1229), .A(net_1196) );
INV_X1 inst_1561 ( .ZN(net_1150), .A(net_1149) );
NAND2_X1 inst_938 ( .ZN(net_585), .A1(net_584), .A2(net_583) );
NAND2_X1 inst_574 ( .ZN(net_652), .A2(n392gat), .A1(n222gat) );
XNOR2_X1 inst_386 ( .ZN(net_1451), .B(net_1428), .A(net_1399) );
XNOR2_X1 inst_158 ( .ZN(net_649), .B(net_601), .A(net_575) );
XNOR2_X1 inst_141 ( .A(net_539), .B(net_538), .ZN(n3211gat) );
NAND2_X1 inst_1229 ( .ZN(net_1259), .A1(net_1258), .A2(net_1241) );
NAND2_X1 inst_1322 ( .ZN(net_1500), .A1(net_1448), .A2(net_1398) );
NAND2_X1 inst_936 ( .ZN(net_601), .A1(net_555), .A2(net_505) );
INV_X1 inst_1490 ( .ZN(net_675), .A(net_674) );
NOR2_X1 inst_507 ( .ZN(net_103), .A1(net_102), .A2(net_75) );
NAND2_X1 inst_571 ( .ZN(net_1317), .A2(n494gat), .A1(n171gat) );
NAND2_X1 inst_1288 ( .ZN(net_1409), .A2(net_1373), .A1(net_1303) );
NAND2_X1 inst_884 ( .ZN(net_459), .A1(net_458), .A2(net_457) );
NAND2_X1 inst_1154 ( .ZN(net_1082), .A2(net_1081), .A1(net_1039) );
NAND2_X1 inst_711 ( .ZN(net_1402), .A1(n69gat), .A2(n511gat) );
NAND2_X1 inst_827 ( .ZN(net_307), .A1(net_306), .A2(net_282) );
NAND2_X1 inst_552 ( .ZN(net_1097), .A1(n69gat), .A2(n460gat) );
NAND2_X1 inst_599 ( .ZN(net_1428), .A2(n511gat), .A1(n171gat) );
NAND2_X1 inst_1033 ( .ZN(net_799), .A1(net_798), .A2(net_769) );
NOR2_X1 inst_469 ( .ZN(net_42), .A1(net_13), .A2(net_12) );
INV_X1 inst_1564 ( .ZN(net_1182), .A(net_1181) );
NAND2_X1 inst_1348 ( .ZN(net_1590), .A2(net_1514), .A1(net_1479) );
XNOR2_X1 inst_18 ( .ZN(net_160), .A(net_92), .B(net_89) );
NAND2_X1 inst_915 ( .ZN(net_507), .A1(net_506), .A2(net_483) );
NAND2_X1 inst_811 ( .ZN(net_299), .A2(net_267), .A1(net_199) );
NAND2_X1 inst_541 ( .ZN(net_152), .A2(n307gat), .A1(n154gat) );
XNOR2_X1 inst_208 ( .ZN(net_815), .A(net_789), .B(net_788) );
XOR2_X1 inst_9 ( .Z(net_1633), .A(net_1522), .B(net_1521) );
XNOR2_X1 inst_113 ( .ZN(net_482), .B(net_461), .A(net_460) );
NOR2_X1 inst_505 ( .ZN(net_99), .A1(net_98), .A2(net_77) );
NAND2_X1 inst_1365 ( .ZN(net_1574), .A1(net_1573), .A2(net_1547) );
XNOR2_X1 inst_356 ( .ZN(net_1338), .A(net_1302), .B(net_1301) );
NAND2_X1 inst_1058 ( .ZN(net_880), .A1(net_831), .A2(net_797) );
NAND2_X1 inst_1216 ( .ZN(net_1233), .A1(net_1232), .A2(net_1231) );
XNOR2_X1 inst_198 ( .ZN(net_772), .B(net_758), .A(net_757) );
NAND2_X1 inst_1371 ( .ZN(net_1591), .A1(net_1590), .A2(net_1586) );
NAND2_X1 inst_952 ( .ZN(net_606), .A2(net_605), .A1(net_544) );
NAND2_X1 inst_897 ( .ZN(net_498), .A2(net_462), .A1(net_399) );
NAND2_X1 inst_1201 ( .ZN(net_1189), .A1(net_1188), .A2(net_1187) );
AND2_X4 inst_1644 ( .ZN(net_45), .A2(net_44), .A1(net_27) );
INV_X1 inst_1473 ( .ZN(net_566), .A(net_565) );
INV_X1 inst_1594 ( .ZN(net_1368), .A(net_1367) );
NAND2_X1 inst_784 ( .ZN(net_186), .A2(net_124), .A1(net_113) );
NAND2_X1 inst_721 ( .ZN(net_1247), .A2(n477gat), .A1(n137gat) );
NAND2_X1 inst_902 ( .ZN(net_504), .A2(net_467), .A1(net_408) );
NAND2_X1 inst_1272 ( .ZN(net_1360), .A2(net_1359), .A1(net_1353) );
XNOR2_X1 inst_293 ( .ZN(net_1101), .A(net_1079), .B(net_1078) );
NAND2_X1 inst_778 ( .ZN(net_113), .A2(net_112), .A1(net_65) );
NAND2_X1 inst_636 ( .ZN(net_472), .A2(n358gat), .A1(n188gat) );
NAND2_X1 inst_632 ( .ZN(net_1021), .A2(n443gat), .A1(n188gat) );
NAND2_X1 inst_1264 ( .ZN(net_1342), .A1(net_1341), .A2(net_1340) );
NAND2_X1 inst_1366 ( .ZN(net_1576), .A2(net_1575), .A1(net_1561) );
XOR2_X1 inst_0 ( .Z(net_116), .A(net_87), .B(net_63) );
INV_X1 inst_1544 ( .ZN(net_1040), .A(net_1039) );
XNOR2_X1 inst_184 ( .ZN(net_754), .A(net_691), .B(net_674) );
NAND2_X1 inst_690 ( .ZN(net_571), .A1(n86gat), .A2(n375gat) );
XNOR2_X1 inst_433 ( .ZN(net_1609), .B(net_1588), .A(net_1580) );
NAND2_X1 inst_1254 ( .ZN(net_1315), .A1(net_1314), .A2(net_1313) );
NAND2_X1 inst_781 ( .ZN(net_126), .A1(net_125), .A2(net_117) );
NAND2_X1 inst_732 ( .ZN(net_155), .A2(n307gat), .A1(n171gat) );
XNOR2_X1 inst_98 ( .ZN(net_465), .B(net_407), .A(net_377) );
XNOR2_X1 inst_263 ( .ZN(net_995), .B(net_970), .A(net_969) );
XNOR2_X1 inst_185 ( .ZN(net_726), .B(net_705), .A(net_682) );
NAND2_X1 inst_959 ( .ZN(net_636), .A1(net_595), .A2(net_530) );
INV_X1 inst_1442 ( .ZN(net_335), .A(net_334) );
XNOR2_X1 inst_75 ( .ZN(net_362), .A(net_297), .B(net_277) );
XNOR2_X1 inst_332 ( .ZN(net_1277), .B(net_1236), .A(net_1203) );
XNOR2_X1 inst_166 ( .ZN(net_666), .B(net_631), .A(net_630) );
NAND2_X1 inst_868 ( .ZN(net_399), .A1(net_398), .A2(net_388) );
XNOR2_X1 inst_163 ( .A(net_625), .B(net_624), .ZN(n3552gat) );
XNOR2_X1 inst_394 ( .ZN(net_1473), .B(net_1445), .A(net_1444) );
XNOR2_X1 inst_79 ( .ZN(net_338), .B(net_314), .A(net_313) );
NAND2_X1 inst_1289 ( .ZN(net_1394), .A1(net_1393), .A2(net_1381) );
XNOR2_X1 inst_106 ( .ZN(net_439), .B(net_416), .A(net_415) );
INV_X1 inst_1559 ( .ZN(net_1143), .A(net_1142) );
XNOR2_X1 inst_422 ( .ZN(net_1603), .B(net_1564), .A(net_1549) );
XNOR2_X1 inst_201 ( .ZN(net_778), .A(net_746), .B(net_745) );
NAND2_X1 inst_927 ( .ZN(net_550), .A1(net_549), .A2(net_548) );
NAND2_X1 inst_605 ( .ZN(net_784), .A1(n86gat), .A2(n409gat) );
NAND2_X1 inst_1084 ( .ZN(net_920), .A1(net_919), .A2(net_918) );
XNOR2_X1 inst_304 ( .ZN(net_1142), .B(net_1114), .A(net_1113) );
INV_X1 inst_1475 ( .ZN(net_570), .A(net_569) );
INV_X1 inst_1426 ( .ZN(net_231), .A(net_230) );
NAND2_X1 inst_752 ( .ZN(net_1002), .A2(n443gat), .A1(n256gat) );
AND2_X4 inst_1637 ( .ZN(net_17), .A2(n290gat), .A1(n120gat) );
INV_X1 inst_1488 ( .ZN(net_671), .A(net_670) );
NAND2_X1 inst_1027 ( .ZN(net_790), .A1(net_789), .A2(net_788) );
XNOR2_X1 inst_73 ( .ZN(net_332), .B(net_292), .A(net_291) );
NAND2_X1 inst_1143 ( .ZN(net_1054), .A1(net_1053), .A2(net_1030) );
NAND2_X1 inst_1352 ( .ZN(net_1553), .A1(net_1552), .A2(net_1535) );
NAND2_X1 inst_1345 ( .ZN(net_1527), .A1(net_1526), .A2(net_1505) );
XNOR2_X1 inst_378 ( .ZN(net_1430), .A(net_1385), .B(net_1358) );
NAND2_X1 inst_1384 ( .ZN(net_1612), .A1(net_1610), .A2(net_1589) );
INV_X1 inst_1605 ( .ZN(net_1452), .A(net_1451) );
NAND2_X1 inst_890 ( .ZN(net_471), .A1(net_470), .A2(net_442) );
XNOR2_X1 inst_361 ( .ZN(net_1353), .B(net_1326), .A(net_1289) );
NAND2_X1 inst_1024 ( .ZN(net_794), .A2(net_738), .A1(net_708) );
NAND2_X1 inst_1168 ( .ZN(net_1117), .A1(net_1116), .A2(net_1092) );
NAND2_X1 inst_1016 ( .ZN(net_753), .A1(net_752), .A2(net_751) );
INV_X1 inst_1538 ( .ZN(net_994), .A(net_993) );
AND2_X4 inst_1658 ( .ZN(net_147), .A1(net_146), .A2(net_145) );
NAND2_X1 inst_659 ( .ZN(net_16), .A2(n273gat), .A1(n137gat) );
XNOR2_X1 inst_250 ( .ZN(net_945), .A(net_909), .B(net_889) );
NAND2_X1 inst_848 ( .ZN(net_374), .A1(net_373), .A2(net_329) );
INV_X1 inst_1410 ( .ZN(net_82), .A(net_81) );
NAND2_X1 inst_786 ( .ZN(net_170), .A1(net_169), .A2(net_168) );
NAND2_X1 inst_1161 ( .ZN(net_1128), .A2(net_1073), .A1(net_1020) );
INV_X1 inst_1448 ( .ZN(net_382), .A(net_381) );
XNOR2_X1 inst_397 ( .ZN(net_1480), .B(net_1460), .A(net_1459) );
NOR2_X1 inst_504 ( .ZN(net_95), .A1(net_94), .A2(net_85) );
INV_X1 inst_1523 ( .ZN(net_893), .A(net_892) );
INV_X1 inst_1554 ( .ZN(net_1096), .A(net_1095) );
INV_X1 inst_1542 ( .ZN(net_1030), .A(net_1029) );
NAND2_X1 inst_1048 ( .ZN(net_859), .A1(net_806), .A2(net_750) );
XNOR2_X1 inst_440 ( .A(net_1609), .B(net_1608), .ZN(n6210gat) );
NAND2_X1 inst_1297 ( .ZN(net_1419), .A1(net_1418), .A2(net_1417) );
XOR2_X1 inst_2 ( .Z(net_323), .A(net_287), .B(net_286) );
NAND2_X1 inst_644 ( .ZN(net_435), .A2(n358gat), .A1(n1gat) );
NAND2_X1 inst_918 ( .ZN(net_515), .A1(net_514), .A2(net_513) );
INV_X1 inst_1581 ( .ZN(net_1300), .A(net_1299) );
NAND2_X1 inst_1173 ( .ZN(net_1127), .A1(net_1126), .A2(net_1125) );
NAND2_X1 inst_1380 ( .ZN(net_1605), .A2(net_1604), .A1(net_1565) );
NAND2_X1 inst_1091 ( .ZN(net_931), .A1(net_930), .A2(net_929) );
NAND2_X1 inst_1331 ( .ZN(net_1499), .A1(net_1498), .A2(net_1451) );
NAND2_X1 inst_578 ( .ZN(net_907), .A2(n426gat), .A1(n205gat) );
NAND2_X1 inst_888 ( .ZN(net_469), .A1(net_468), .A2(net_431) );
XNOR2_X1 inst_52 ( .ZN(net_236), .A(net_201), .B(net_200) );
NAND2_X1 inst_1393 ( .ZN(net_1625), .A1(net_1624), .A2(net_1623) );
NAND2_X1 inst_668 ( .ZN(net_143), .A2(n307gat), .A1(n205gat) );
NAND2_X1 inst_1236 ( .ZN(net_1301), .A1(net_1246), .A2(net_1230) );
XNOR2_X1 inst_221 ( .ZN(net_845), .B(net_823), .A(net_822) );
NAND2_X1 inst_556 ( .ZN(net_1431), .A2(n511gat), .A1(n103gat) );
NAND2_X1 inst_650 ( .ZN(net_1447), .A2(n511gat), .A1(n120gat) );
XNOR2_X1 inst_289 ( .ZN(net_1093), .A(net_1061), .B(net_1060) );
NAND2_X1 inst_987 ( .ZN(net_693), .A1(net_689), .A2(net_667) );
INV_X1 inst_1498 ( .ZN(net_761), .A(net_760) );
XNOR2_X1 inst_432 ( .ZN(net_1611), .B(net_1594), .A(net_1584) );
NAND2_X1 inst_679 ( .ZN(net_1258), .A2(n494gat), .A1(n239gat) );
XNOR2_X1 inst_420 ( .ZN(net_1630), .B(net_1538), .A(net_1480) );
XNOR2_X1 inst_282 ( .ZN(net_1126), .B(net_1053), .A(net_1029) );
NAND2_X1 inst_1358 ( .ZN(net_1575), .A1(net_1533), .A2(net_1497) );
NOR2_X1 inst_513 ( .ZN(net_121), .A1(net_120), .A2(net_97) );
NAND2_X1 inst_1351 ( .ZN(net_1546), .A1(net_1542), .A2(net_1520) );
NAND2_X1 inst_754 ( .ZN(net_919), .A2(n443gat), .A1(n1gat) );
XNOR2_X1 inst_44 ( .ZN(net_222), .A(net_207), .B(net_206) );
AND2_X4 inst_1630 ( .ZN(net_26), .A2(n273gat), .A1(n103gat) );
NAND2_X1 inst_1305 ( .ZN(net_1455), .A2(net_1406), .A1(net_1364) );
XNOR2_X1 inst_371 ( .ZN(net_1387), .B(net_1370), .A(net_1369) );
INV_X1 inst_1586 ( .ZN(net_1331), .A(net_1330) );
XNOR2_X1 inst_314 ( .ZN(net_1190), .B(net_1158), .A(net_1157) );
XNOR2_X1 inst_435 ( .ZN(net_1606), .A(net_1590), .B(net_1587) );
INV_X1 inst_1572 ( .ZN(net_1215), .A(net_1214) );
NAND2_X1 inst_597 ( .ZN(net_805), .A2(n409gat), .A1(n205gat) );
NAND2_X1 inst_687 ( .ZN(net_476), .A2(n358gat), .A1(n120gat) );
NAND2_X1 inst_774 ( .ZN(net_41), .A2(net_30), .A1(net_15) );
NAND2_X1 inst_621 ( .ZN(net_373), .A2(n341gat), .A1(n120gat) );
INV_X1 inst_1587 ( .ZN(net_1339), .A(net_1338) );
NAND2_X1 inst_1185 ( .ZN(net_1148), .A1(net_1147), .A2(net_1146) );
NAND2_X1 inst_838 ( .ZN(net_350), .A1(net_349), .A2(net_348) );
NAND2_X1 inst_985 ( .ZN(net_714), .A1(net_663), .A2(net_600) );
NAND2_X1 inst_628 ( .ZN(net_596), .A2(n375gat), .A1(n171gat) );
NAND2_X1 inst_815 ( .ZN(net_292), .A2(net_247), .A1(net_182) );
NOR2_X1 inst_472 ( .ZN(net_51), .A1(net_25), .A2(net_24) );
XNOR2_X1 inst_447 ( .A(net_1630), .B(net_1629), .ZN(n6280gat) );
OR2_X4 inst_457 ( .ZN(net_190), .A1(net_189), .A2(net_188) );
INV_X1 inst_1508 ( .ZN(net_787), .A(net_786) );
NAND2_X1 inst_1257 ( .ZN(net_1325), .A1(net_1324), .A2(net_1310) );
NAND2_X1 inst_875 ( .ZN(net_417), .A1(net_416), .A2(net_415) );
NAND2_X1 inst_1391 ( .ZN(net_1622), .A1(net_1621), .A2(net_1620) );
NAND2_X1 inst_1222 ( .ZN(net_1246), .A1(net_1245), .A2(net_1244) );
NAND2_X1 inst_665 ( .ZN(net_262), .A2(n324gat), .A1(n154gat) );
NAND2_X1 inst_1387 ( .ZN(net_1616), .A1(net_1615), .A2(net_1614) );
INV_X1 inst_1405 ( .ZN(net_72), .A(net_71) );
NAND2_X1 inst_1073 ( .ZN(net_881), .A2(net_880), .A1(net_872) );
NAND2_X1 inst_1117 ( .ZN(net_1000), .A1(net_999), .A2(net_976) );
NAND2_X1 inst_1130 ( .ZN(net_1026), .A1(net_1025), .A2(net_998) );
INV_X1 inst_1449 ( .ZN(net_384), .A(net_383) );
XNOR2_X1 inst_127 ( .ZN(net_556), .B(net_508), .A(net_486) );
NAND2_X1 inst_855 ( .ZN(net_391), .A1(net_390), .A2(net_389) );
XNOR2_X1 inst_413 ( .ZN(net_1547), .B(net_1526), .A(net_1504) );
XNOR2_X1 inst_146 ( .ZN(net_581), .B(net_554), .A(net_553) );
INV_X1 inst_1610 ( .ZN(net_1481), .A(net_1480) );
XNOR2_X1 inst_334 ( .ZN(net_1256), .B(net_1227), .A(net_1226) );
NAND2_X1 inst_859 ( .ZN(net_410), .A2(net_368), .A1(net_320) );
XNOR2_X1 inst_187 ( .ZN(net_722), .B(net_707), .A(net_647) );
XNOR2_X1 inst_206 ( .ZN(net_822), .B(net_784), .A(net_760) );
NAND2_X1 inst_1268 ( .ZN(net_1378), .A1(net_1318), .A2(net_1276) );
NAND2_X1 inst_805 ( .ZN(net_289), .A2(net_243), .A1(net_187) );
XNOR2_X1 inst_122 ( .ZN(net_516), .B(net_470), .A(net_441) );
NAND2_X1 inst_1196 ( .ZN(net_1176), .A1(net_1175), .A2(net_1174) );
XNOR2_X1 inst_25 ( .A(net_123), .B(net_122), .ZN(n1901gat) );
XNOR2_X1 inst_354 ( .ZN(net_1328), .B(net_1292), .A(net_1291) );
XNOR2_X1 inst_405 ( .ZN(net_1517), .B(net_1483), .A(net_1482) );
NAND2_X1 inst_1145 ( .ZN(net_1089), .A2(net_1038), .A1(net_982) );
NOR2_X1 inst_492 ( .A2(net_94), .ZN(net_71), .A1(net_40) );
NAND2_X1 inst_1042 ( .ZN(net_819), .A1(net_818), .A2(net_817) );
NAND2_X1 inst_817 ( .ZN(net_314), .A2(net_249), .A1(net_196) );
XNOR2_X1 inst_326 ( .ZN(net_1273), .A(net_1216), .B(net_1190) );
NAND2_X1 inst_1363 ( .ZN(net_1588), .A2(net_1559), .A1(net_1503) );
NOR2_X1 inst_518 ( .ZN(net_184), .A2(net_150), .A1(net_105) );
XNOR2_X1 inst_69 ( .ZN(net_351), .A(net_321), .B(net_281) );
XNOR2_X1 inst_373 ( .ZN(net_1399), .A(net_1379), .B(net_1378) );
XNOR2_X1 inst_82 ( .ZN(net_343), .B(net_324), .A(net_323) );
AND2_X4 inst_1646 ( .ZN(net_47), .A2(net_46), .A1(net_7) );
XNOR2_X1 inst_108 ( .ZN(net_443), .B(net_413), .A(net_412) );
NAND2_X1 inst_844 ( .ZN(net_366), .A1(net_365), .A2(net_331) );
NAND2_X1 inst_595 ( .ZN(net_689), .A2(n392gat), .A1(n120gat) );
XNOR2_X1 inst_22 ( .ZN(net_157), .A(net_94), .B(net_86) );
NAND2_X1 inst_1121 ( .ZN(net_1008), .A1(net_1007), .A2(net_988) );
NAND2_X1 inst_1102 ( .ZN(net_952), .A1(net_951), .A2(net_950) );
OR2_X4 inst_460 ( .ZN(net_199), .A1(net_198), .A2(net_197) );
INV_X1 inst_1455 ( .ZN(net_440), .A(net_439) );
NAND2_X1 inst_1354 ( .ZN(net_1557), .A1(net_1556), .A2(net_1555) );
INV_X1 inst_1429 ( .ZN(net_237), .A(net_236) );
NAND2_X1 inst_970 ( .ZN(net_644), .A1(net_643), .A2(net_642) );
XNOR2_X1 inst_307 ( .ZN(net_1164), .A(net_1128), .B(net_1100) );
NAND2_X1 inst_1278 ( .ZN(net_1395), .A1(net_1346), .A2(net_1285) );
NAND2_X1 inst_767 ( .ZN(net_37), .A1(net_5), .A2(net_4) );
NAND2_X1 inst_638 ( .ZN(net_23), .A2(n290gat), .A1(n239gat) );
XNOR2_X1 inst_161 ( .ZN(net_645), .B(net_612), .A(net_611) );
NAND2_X1 inst_560 ( .ZN(net_1370), .A2(n511gat), .A1(n239gat) );
NAND2_X1 inst_749 ( .ZN(net_1264), .A2(n494gat), .A1(n222gat) );
NAND2_X1 inst_586 ( .ZN(net_1529), .A2(n528gat), .A1(n188gat) );
NAND2_X1 inst_702 ( .ZN(net_474), .A2(n358gat), .A1(n137gat) );
XNOR2_X1 inst_16 ( .ZN(net_136), .B(net_118), .A(net_61) );
INV_X1 inst_1505 ( .ZN(net_779), .A(net_778) );
NAND2_X1 inst_717 ( .ZN(net_1165), .A2(n477gat), .A1(n35gat) );
XNOR2_X1 inst_276 ( .ZN(net_1044), .A(net_1016), .B(net_1015) );
NAND2_X1 inst_1030 ( .ZN(net_823), .A2(net_767), .A1(net_716) );
NAND2_X1 inst_718 ( .ZN(net_1232), .A2(n494gat), .A1(n1gat) );
NAND2_X1 inst_1029 ( .ZN(net_792), .A1(net_791), .A2(net_765) );
XNOR2_X1 inst_156 ( .ZN(net_657), .B(net_609), .A(net_577) );
INV_X1 inst_1466 ( .ZN(net_535), .A(net_534) );
NAND2_X1 inst_950 ( .ZN(net_602), .A1(net_601), .A2(net_576) );
NAND2_X1 inst_1373 ( .ZN(net_1593), .A1(net_1592), .A2(net_1570) );
NAND2_X1 inst_1068 ( .ZN(net_902), .A1(net_850), .A2(net_802) );
NAND2_X1 inst_886 ( .ZN(net_464), .A1(net_463), .A2(net_432) );
NAND2_X1 inst_1203 ( .ZN(net_1227), .A2(net_1166), .A1(net_1129) );
NAND2_X1 inst_802 ( .ZN(net_269), .A1(net_268), .A2(net_223) );
XNOR2_X1 inst_296 ( .ZN(net_1146), .B(net_1106), .A(net_1083) );
XNOR2_X1 inst_91 ( .ZN(net_415), .A(net_369), .B(net_332) );
NAND2_X1 inst_1218 ( .ZN(net_1237), .A1(net_1236), .A2(net_1204) );
NAND2_X1 inst_1324 ( .ZN(net_1492), .A2(net_1441), .A1(net_1394) );
NAND2_X1 inst_905 ( .ZN(net_520), .A2(net_471), .A1(net_411) );
XNOR2_X1 inst_132 ( .ZN(net_553), .B(net_504), .A(net_490) );
XNOR2_X1 inst_342 ( .ZN(net_1291), .B(net_1262), .A(net_1251) );
NOR2_X1 inst_526 ( .ZN(net_1516), .A2(net_1515), .A1(net_1493) );
NAND2_X1 inst_1006 ( .ZN(net_719), .A1(net_718), .A2(net_717) );
NAND2_X1 inst_1178 ( .ZN(net_1138), .A1(net_1137), .A2(net_1136) );
OR2_X4 inst_463 ( .ZN(net_211), .A1(net_210), .A2(net_209) );
INV_X1 inst_1534 ( .ZN(net_984), .A(net_983) );
XNOR2_X1 inst_96 ( .ZN(net_425), .A(net_360), .B(net_327) );
INV_X1 inst_1549 ( .ZN(net_1075), .A(net_1074) );
XNOR2_X1 inst_101 ( .ZN(net_430), .B(net_405), .A(net_404) );
XNOR2_X1 inst_319 ( .ZN(net_1201), .B(net_1172), .A(net_1171) );
INV_X1 inst_1450 ( .ZN(net_386), .A(net_385) );
XNOR2_X1 inst_400 ( .ZN(net_1504), .A(net_1476), .B(net_1475) );
NAND2_X1 inst_614 ( .ZN(net_169), .A2(n307gat), .A1(n256gat) );
NAND2_X1 inst_649 ( .ZN(net_1037), .A2(n460gat), .A1(n1gat) );
NAND2_X1 inst_821 ( .ZN(net_293), .A1(net_292), .A2(net_291) );
XNOR2_X1 inst_261 ( .ZN(net_991), .A(net_965), .B(net_964) );
INV_X1 inst_1464 ( .ZN(net_489), .A(net_488) );
NAND2_X1 inst_1247 ( .ZN(net_1296), .A1(net_1295), .A2(net_1294) );
NAND2_X1 inst_1031 ( .ZN(net_795), .A1(net_794), .A2(net_793) );
NAND2_X1 inst_980 ( .ZN(net_709), .A1(net_656), .A2(net_608) );
NOR2_X1 inst_500 ( .A2(net_98), .ZN(net_88), .A1(net_32) );
INV_X1 inst_1592 ( .ZN(net_1358), .A(net_1357) );
NAND2_X1 inst_945 ( .ZN(net_595), .A1(net_594), .A2(net_570) );
NOR2_X1 inst_510 ( .ZN(net_109), .A1(net_108), .A2(net_79) );
XNOR2_X1 inst_268 ( .ZN(net_1049), .B(net_1013), .A(net_983) );
INV_X1 inst_1518 ( .ZN(net_883), .A(net_882) );
XNOR2_X1 inst_369 ( .ZN(net_1401), .B(net_1361), .A(net_1328) );
INV_X1 inst_1575 ( .ZN(net_1250), .A(net_1249) );
NAND2_X1 inst_995 ( .ZN(net_710), .A2(net_709), .A1(net_679) );
NAND2_X1 inst_550 ( .ZN(net_1292), .A1(n86gat), .A2(n494gat) );
INV_X1 inst_1493 ( .ZN(net_683), .A(net_682) );
NAND2_X1 inst_1258 ( .ZN(net_1327), .A1(net_1326), .A2(net_1290) );
NAND2_X1 inst_830 ( .ZN(net_315), .A1(net_314), .A2(net_313) );
NAND2_X1 inst_603 ( .ZN(net_468), .A2(n358gat), .A1(n103gat) );
XNOR2_X1 inst_327 ( .ZN(net_1238), .B(net_1206), .A(net_1205) );
NAND2_X1 inst_1308 ( .ZN(net_1446), .A1(net_1445), .A2(net_1444) );
XNOR2_X1 inst_85 ( .ZN(net_377), .B(net_352), .A(net_351) );
XNOR2_X1 inst_291 ( .ZN(net_1099), .B(net_1085), .A(net_1051) );
NAND2_X1 inst_1286 ( .ZN(net_1390), .A1(net_1389), .A2(net_1368) );
NAND2_X1 inst_1060 ( .ZN(net_853), .A1(net_852), .A2(net_851) );
XNOR2_X1 inst_266 ( .ZN(net_1042), .B(net_999), .A(net_975) );
NAND2_X1 inst_776 ( .ZN(net_64), .A1(net_63), .A2(net_60) );
INV_X1 inst_1419 ( .ZN(net_217), .A(net_216) );
NAND2_X1 inst_900 ( .ZN(net_502), .A2(net_459), .A1(net_401) );
NAND2_X1 inst_866 ( .ZN(net_395), .A1(net_394), .A2(net_384) );
NAND2_X1 inst_1198 ( .ZN(net_1210), .A2(net_1153), .A1(net_1110) );
XNOR2_X1 inst_77 ( .ZN(net_336), .B(net_319), .A(net_318) );
XNOR2_X1 inst_171 ( .ZN(net_703), .B(net_662), .A(net_620) );
INV_X1 inst_1439 ( .ZN(net_329), .A(net_328) );
NAND2_X1 inst_1362 ( .ZN(net_1594), .A1(net_1557), .A2(net_1501) );
NAND2_X1 inst_558 ( .ZN(net_363), .A2(n341gat), .A1(n103gat) );
NAND2_X1 inst_594 ( .ZN(net_1389), .A2(n511gat), .A1(n222gat) );
XNOR2_X1 inst_145 ( .ZN(net_579), .B(net_549), .A(net_548) );
XNOR2_X1 inst_290 ( .ZN(net_1095), .A(net_1064), .B(net_1063) );
XNOR2_X1 inst_374 ( .ZN(net_1417), .A(net_1359), .B(net_1354) );
XNOR2_X1 inst_272 ( .ZN(net_1034), .A(net_1005), .B(net_1004) );
NOR2_X1 inst_502 ( .ZN(net_91), .A1(net_90), .A2(net_71) );
XNOR2_X1 inst_103 ( .ZN(net_457), .B(net_400), .A(net_385) );
NAND2_X1 inst_814 ( .ZN(net_321), .A2(net_271), .A1(net_185) );
AND2_X4 inst_1632 ( .ZN(net_21), .A1(n35gat), .A2(n290gat) );
XNOR2_X1 inst_248 ( .A(net_919), .B(net_918), .ZN(n4591gat) );
INV_X1 inst_1613 ( .ZN(net_1493), .A(net_1492) );
XNOR2_X1 inst_389 ( .ZN(net_1462), .B(net_1426), .A(net_1425) );
INV_X1 inst_1458 ( .ZN(net_446), .A(net_445) );
NAND2_X1 inst_925 ( .ZN(net_540), .A1(net_539), .A2(net_538) );
NAND2_X1 inst_789 ( .ZN(net_240), .A1(net_239), .A2(net_238) );
INV_X1 inst_1598 ( .ZN(net_1400), .A(net_1399) );
XNOR2_X1 inst_357 ( .ZN(net_1343), .A(net_1307), .B(net_1306) );
NAND2_X1 inst_1120 ( .ZN(net_1006), .A1(net_1005), .A2(net_1004) );
INV_X1 inst_1437 ( .ZN(net_285), .A(net_284) );
NAND2_X1 inst_1382 ( .ZN(net_1608), .A2(net_1607), .A1(net_1591) );
NAND2_X1 inst_1141 ( .ZN(net_1081), .A1(net_1026), .A2(net_974) );
NAND2_X1 inst_809 ( .ZN(net_308), .A2(net_269), .A1(net_208) );
INV_X1 inst_1536 ( .ZN(net_988), .A(net_987) );
NAND2_X1 inst_881 ( .ZN(net_453), .A1(net_452), .A2(net_451) );
NAND2_X1 inst_932 ( .ZN(net_572), .A1(net_571), .A2(net_535) );
NAND2_X1 inst_822 ( .ZN(net_296), .A1(net_295), .A2(net_294) );
NAND2_X1 inst_913 ( .ZN(net_503), .A1(net_502), .A2(net_485) );
XNOR2_X1 inst_180 ( .ZN(net_743), .B(net_690), .A(net_668) );
NAND2_X1 inst_1125 ( .ZN(net_1041), .A2(net_990), .A1(net_931) );
NAND2_X1 inst_1234 ( .ZN(net_1265), .A1(net_1264), .A2(net_1263) );
NAND2_X1 inst_1225 ( .ZN(net_1272), .A2(net_1220), .A1(net_1168) );
NAND2_X1 inst_947 ( .ZN(net_612), .A1(net_572), .A2(net_497) );
NAND2_X1 inst_912 ( .ZN(net_501), .A2(net_500), .A1(net_450) );
NAND2_X1 inst_731 ( .ZN(net_1192), .A1(n52gat), .A2(n477gat) );
NAND2_X1 inst_609 ( .ZN(net_128), .A2(n307gat), .A1(n137gat) );
NAND2_X1 inst_1022 ( .ZN(net_767), .A1(net_766), .A2(net_733) );
NAND2_X1 inst_795 ( .ZN(net_255), .A1(net_254), .A2(net_235) );
XNOR2_X1 inst_301 ( .ZN(net_1134), .B(net_1123), .A(net_1095) );
XNOR2_X1 inst_363 ( .ZN(net_1357), .B(net_1347), .A(net_1311) );
XNOR2_X1 inst_27 ( .ZN(net_203), .A(net_134), .B(net_133) );
XNOR2_X1 inst_247 ( .ZN(net_939), .A(net_914), .B(net_913) );
XNOR2_X1 inst_403 ( .ZN(net_1528), .B(net_1494), .A(net_1449) );
XNOR2_X1 inst_302 ( .ZN(net_1154), .A(net_1111), .B(net_1088) );
AND2_X4 inst_1639 ( .ZN(net_9), .A2(n290gat), .A1(n154gat) );
XNOR2_X1 inst_322 ( .ZN(net_1226), .B(net_1192), .A(net_1162) );
NAND2_X1 inst_673 ( .ZN(net_691), .A2(n392gat), .A1(n171gat) );
NAND2_X1 inst_1223 ( .ZN(net_1248), .A1(net_1247), .A2(net_1215) );
XNOR2_X1 inst_211 ( .ZN(net_842), .B(net_803), .A(net_774) );
NAND2_X1 inst_619 ( .ZN(net_256), .A2(n324gat), .A1(n120gat) );
INV_X1 inst_1588 ( .ZN(net_1344), .A(net_1343) );
NAND2_X1 inst_1151 ( .ZN(net_1073), .A1(net_1072), .A2(net_1047) );
NAND2_X1 inst_681 ( .ZN(net_1072), .A2(n460gat), .A1(n35gat) );
INV_X1 inst_1414 ( .ZN(net_97), .A(net_96) );
NAND2_X1 inst_561 ( .ZN(net_1116), .A2(n460gat), .A1(n171gat) );
XNOR2_X1 inst_412 ( .B(net_1515), .A(net_1492), .ZN(n6150gat) );
OR2_X4 inst_449 ( .ZN(net_58), .A2(net_42), .A1(net_13) );
AND2_X4 inst_1654 ( .ZN(net_132), .A1(net_131), .A2(net_130) );
NAND2_X1 inst_1355 ( .ZN(net_1559), .A1(net_1558), .A2(net_1540) );
NAND2_X1 inst_639 ( .ZN(net_699), .A2(n392gat), .A1(n154gat) );
NAND2_X1 inst_877 ( .ZN(net_423), .A1(net_422), .A2(net_421) );
AND2_X4 inst_1641 ( .ZN(net_4), .A2(n273gat), .A1(n154gat) );
INV_X1 inst_1506 ( .ZN(net_781), .A(net_780) );
XNOR2_X1 inst_155 ( .ZN(net_624), .B(net_603), .A(net_579) );
OR2_X4 inst_464 ( .ZN(net_1577), .A1(net_1516), .A2(n6150gat) );
NAND2_X1 inst_871 ( .ZN(net_406), .A1(net_405), .A2(net_404) );
XNOR2_X1 inst_341 ( .ZN(net_1281), .B(net_1254), .A(net_1253) );
NAND2_X1 inst_962 ( .ZN(net_616), .A1(net_615), .A2(net_614) );
XNOR2_X1 inst_196 ( .ZN(net_768), .B(net_735), .A(net_734) );
INV_X1 inst_1567 ( .ZN(net_1195), .A(net_1194) );
NAND2_X1 inst_532 ( .ZN(net_1011), .A2(n443gat), .A1(n205gat) );
XNOR2_X1 inst_55 ( .ZN(net_291), .A(net_258), .B(net_232) );
NAND2_X1 inst_1171 ( .ZN(net_1124), .A1(net_1123), .A2(net_1096) );
NAND2_X1 inst_641 ( .ZN(net_1009), .A2(n443gat), .A1(n154gat) );
NOR2_X1 inst_498 ( .A2(net_102), .ZN(net_77), .A1(net_38) );
NAND2_X1 inst_684 ( .ZN(net_1486), .A2(n528gat), .A1(n35gat) );
AND2_X4 inst_1651 ( .ZN(net_59), .A2(net_48), .A1(net_23) );
INV_X1 inst_1403 ( .ZN(net_67), .A(net_66) );
NAND2_X1 inst_1361 ( .ZN(net_1568), .A1(net_1567), .A2(net_1566) );
XNOR2_X1 inst_298 ( .ZN(net_1132), .B(net_1104), .A(net_1103) );
NAND2_X1 inst_1327 ( .ZN(net_1484), .A1(net_1483), .A2(net_1482) );
NAND2_X1 inst_1137 ( .ZN(net_1063), .A2(net_1014), .A1(net_949) );
XNOR2_X1 inst_42 ( .ZN(net_216), .A(net_178), .B(net_177) );
XNOR2_X1 inst_323 ( .ZN(net_1231), .B(net_1198), .A(net_1185) );
NAND2_X1 inst_1162 ( .ZN(net_1105), .A1(net_1104), .A2(net_1103) );
NAND2_X1 inst_1389 ( .ZN(net_1619), .A1(net_1618), .A2(net_1617) );
NAND2_X1 inst_588 ( .ZN(net_12), .A2(n273gat), .A1(n239gat) );
INV_X1 inst_1479 ( .ZN(net_582), .A(net_581) );
XNOR2_X1 inst_350 ( .ZN(net_1333), .B(net_1297), .A(net_1281) );
XNOR2_X1 inst_231 ( .ZN(net_886), .B(net_852), .A(net_851) );
NAND2_X1 inst_1138 ( .ZN(net_1043), .A1(net_1042), .A2(net_1041) );
NAND2_X1 inst_1241 ( .ZN(net_1279), .A1(net_1278), .A2(net_1277) );
NAND2_X1 inst_1119 ( .ZN(net_1003), .A1(net_1002), .A2(net_1001) );
INV_X1 inst_1494 ( .ZN(net_701), .A(net_700) );
INV_X1 inst_1433 ( .ZN(net_277), .A(net_276) );
NAND2_X1 inst_1038 ( .ZN(net_810), .A1(net_809), .A2(net_781) );
NAND2_X1 inst_793 ( .ZN(net_251), .A1(net_250), .A2(net_225) );
NAND2_X1 inst_715 ( .ZN(net_894), .A1(n86gat), .A2(n426gat) );
XNOR2_X1 inst_437 ( .A(net_1600), .B(net_1599), .ZN(n6180gat) );
NAND2_X1 inst_1255 ( .ZN(net_1318), .A1(net_1317), .A2(net_1316) );
NAND2_X1 inst_940 ( .ZN(net_605), .A2(net_552), .A1(net_501) );
NAND2_X1 inst_1004 ( .ZN(net_751), .A1(net_692), .A2(net_641) );
INV_X1 inst_1481 ( .ZN(net_623), .A(net_622) );
NAND2_X1 inst_1340 ( .ZN(net_1523), .A1(net_1522), .A2(net_1521) );
XNOR2_X1 inst_189 ( .ZN(net_739), .B(net_711), .A(net_680) );
INV_X1 inst_1452 ( .ZN(net_431), .A(net_430) );
NAND2_X1 inst_1356 ( .ZN(net_1571), .A2(net_1527), .A1(net_1477) );
XNOR2_X1 inst_14 ( .ZN(net_130), .A(net_108), .B(net_80) );
NOR2_X1 inst_475 ( .ZN(net_34), .A2(net_33), .A1(net_29) );
XNOR2_X1 inst_31 ( .ZN(net_180), .A(net_143), .B(net_142) );
NAND2_X1 inst_1045 ( .ZN(net_831), .A1(net_830), .A2(net_829) );
NAND2_X1 inst_528 ( .ZN(net_1526), .A2(n528gat), .A1(n205gat) );
NAND2_X1 inst_865 ( .ZN(net_393), .A2(net_392), .A1(net_344) );
XNOR2_X1 inst_252 ( .ZN(net_1016), .B(net_941), .A(net_911) );
NAND2_X1 inst_903 ( .ZN(net_511), .A2(net_469), .A1(net_406) );
XNOR2_X1 inst_62 ( .ZN(net_313), .A(net_262), .B(net_228) );
NAND2_X1 inst_956 ( .ZN(net_628), .A1(net_589), .A2(net_518) );
INV_X1 inst_1470 ( .ZN(net_560), .A(net_559) );
XNOR2_X1 inst_251 ( .ZN(net_956), .A(net_930), .B(net_929) );
NAND2_X1 inst_1396 ( .ZN(net_1629), .A1(net_1628), .A2(net_1572) );
XNOR2_X1 inst_352 ( .ZN(net_1322), .A(net_1284), .B(net_1283) );
NAND2_X1 inst_575 ( .ZN(net_590), .A2(n375gat), .A1(n120gat) );
NAND2_X1 inst_1074 ( .ZN(net_895), .A1(net_894), .A2(net_868) );
NAND2_X1 inst_846 ( .ZN(net_370), .A1(net_369), .A2(net_333) );
XNOR2_X1 inst_286 ( .ZN(net_1087), .B(net_1072), .A(net_1046) );
NAND2_X1 inst_879 ( .ZN(net_429), .A1(net_428), .A2(net_427) );
INV_X1 inst_1552 ( .ZN(net_1092), .A(net_1091) );
INV_X1 inst_1524 ( .ZN(net_912), .A(net_911) );
NAND2_X1 inst_1213 ( .ZN(net_1254), .A2(net_1193), .A1(net_1138) );
NOR2_X1 inst_484 ( .ZN(net_52), .A2(net_51), .A1(net_25) );
NAND2_X1 inst_627 ( .ZN(net_1216), .A2(n477gat), .A1(n205gat) );
XNOR2_X1 inst_32 ( .ZN(net_177), .B(net_128), .A(net_127) );
XNOR2_X1 inst_344 ( .ZN(net_1302), .B(net_1266), .A(net_1256) );
XNOR2_X1 inst_428 ( .A(net_1578), .B(net_1577), .ZN(n6160gat) );
INV_X1 inst_1602 ( .ZN(net_1436), .A(net_1435) );
NAND2_X1 inst_969 ( .ZN(net_641), .A1(net_640), .A2(net_639) );
NAND2_X1 inst_629 ( .ZN(net_158), .A1(n35gat), .A2(n307gat) );
NAND2_X1 inst_1100 ( .ZN(net_964), .A2(net_922), .A1(net_853) );
XNOR2_X1 inst_407 ( .ZN(net_1543), .A(net_1498), .B(net_1452) );
NAND2_X1 inst_791 ( .ZN(net_247), .A1(net_246), .A2(net_219) );
NAND2_X1 inst_623 ( .ZN(net_1421), .A2(n511gat), .A1(n256gat) );
NAND2_X1 inst_1208 ( .ZN(net_1213), .A1(net_1198), .A2(net_1186) );
NAND2_X1 inst_1072 ( .ZN(net_879), .A1(net_878), .A2(net_877) );
NAND2_X1 inst_1044 ( .ZN(net_824), .A1(net_823), .A2(net_822) );
XNOR2_X1 inst_97 ( .ZN(net_434), .B(net_394), .A(net_383) );
INV_X1 inst_1621 ( .ZN(net_1550), .A(net_1549) );
NAND2_X1 inst_616 ( .ZN(net_1297), .A1(n52gat), .A2(n494gat) );
NAND2_X1 inst_1338 ( .ZN(net_1551), .A2(net_1487), .A1(net_1458) );
NAND2_X1 inst_898 ( .ZN(net_496), .A2(net_456), .A1(net_397) );
NAND2_X1 inst_1191 ( .ZN(net_1166), .A1(net_1165), .A2(net_1164) );
NAND2_X1 inst_775 ( .ZN(net_60), .A2(net_48), .A1(net_22) );
NAND2_X1 inst_533 ( .ZN(net_551), .A2(n375gat), .A1(n222gat) );
NAND2_X1 inst_620 ( .ZN(net_355), .A1(n86gat), .A2(n341gat) );
NAND2_X1 inst_1107 ( .ZN(net_968), .A1(net_967), .A2(net_945) );
NAND2_X1 inst_652 ( .ZN(net_588), .A2(n375gat), .A1(n137gat) );
NAND2_X1 inst_1377 ( .ZN(net_1601), .A1(net_1600), .A2(net_1599) );
XNOR2_X1 inst_137 ( .ZN(net_563), .B(net_517), .A(net_516) );
NAND2_X1 inst_677 ( .ZN(net_921), .A2(n426gat), .A1(n188gat) );
XNOR2_X1 inst_425 ( .ZN(net_1584), .B(net_1567), .A(net_1566) );
INV_X1 inst_1427 ( .ZN(net_233), .A(net_232) );
XNOR2_X1 inst_130 ( .ZN(net_536), .B(net_500), .A(net_449) );
INV_X1 inst_1566 ( .ZN(net_1191), .A(net_1190) );
INV_X1 inst_1532 ( .ZN(net_976), .A(net_975) );
INV_X1 inst_1409 ( .ZN(net_80), .A(net_79) );
NAND2_X1 inst_722 ( .ZN(net_1109), .A2(n460gat), .A1(n256gat) );
XNOR2_X1 inst_227 ( .ZN(net_873), .B(net_843), .A(net_842) );
NAND2_X1 inst_1095 ( .ZN(net_972), .A2(net_928), .A1(net_866) );
NAND2_X1 inst_760 ( .ZN(net_1513), .A1(n86gat), .A2(n528gat) );
NAND2_X1 inst_746 ( .ZN(net_258), .A2(n324gat), .A1(n205gat) );
XNOR2_X1 inst_176 ( .ZN(net_715), .B(net_676), .A(net_645) );
XNOR2_X1 inst_58 ( .ZN(net_274), .A(net_260), .B(net_220) );
XNOR2_X1 inst_87 ( .ZN(net_379), .B(net_349), .A(net_348) );
NAND2_X1 inst_1054 ( .ZN(net_841), .A1(net_840), .A2(net_839) );
NAND2_X1 inst_1336 ( .ZN(net_1511), .A1(net_1510), .A2(net_1509) );
NAND2_X1 inst_1332 ( .ZN(net_1501), .A2(net_1500), .A1(net_1488) );
AND2_X2 inst_1665 ( .ZN(n545gat), .A2(n273gat), .A1(n1gat) );
INV_X1 inst_1469 ( .ZN(net_544), .A(net_543) );
NAND2_X1 inst_972 ( .ZN(net_684), .A2(net_616), .A1(net_585) );
NAND2_X1 inst_983 ( .ZN(net_711), .A1(net_659), .A2(net_610) );
NAND2_X1 inst_800 ( .ZN(net_265), .A1(net_264), .A2(net_227) );
NAND2_X1 inst_780 ( .ZN(net_124), .A1(net_123), .A2(net_122) );
XNOR2_X1 inst_10 ( .ZN(net_122), .B(net_112), .A(net_62) );
XOR2_X1 inst_4 ( .Z(net_513), .A(net_493), .B(net_492) );
INV_X1 inst_1577 ( .ZN(net_1257), .A(net_1256) );
NAND2_X1 inst_1110 ( .ZN(net_1001), .A2(net_942), .A1(net_898) );
NAND2_X1 inst_581 ( .ZN(net_131), .A2(n307gat), .A1(n188gat) );
NAND2_X1 inst_600 ( .ZN(net_15), .A2(n290gat), .A1(n1gat) );
XNOR2_X1 inst_28 ( .ZN(net_166), .A(net_146), .B(net_145) );
NAND2_X1 inst_1194 ( .ZN(net_1170), .A1(net_1169), .A2(net_1143) );
INV_X1 inst_1569 ( .ZN(net_1200), .A(net_1199) );
NAND2_X1 inst_1089 ( .ZN(net_953), .A2(net_910), .A1(net_855) );
XNOR2_X1 inst_49 ( .ZN(net_232), .A(net_189), .B(net_188) );
XNOR2_X1 inst_204 ( .ZN(net_786), .A(net_737), .B(net_723) );
INV_X1 inst_1550 ( .ZN(net_1084), .A(net_1083) );
NAND2_X1 inst_592 ( .ZN(net_470), .A2(n358gat), .A1(n154gat) );
NAND2_X1 inst_1284 ( .ZN(net_1386), .A2(net_1385), .A1(net_1357) );
NAND2_X1 inst_546 ( .ZN(net_925), .A2(n426gat), .A1(n137gat) );
NAND2_X1 inst_993 ( .ZN(net_706), .A2(net_705), .A1(net_683) );
NAND2_X1 inst_1290 ( .ZN(net_1396), .A2(net_1395), .A1(net_1352) );
NAND2_X1 inst_910 ( .ZN(net_497), .A1(net_496), .A2(net_495) );
NAND2_X1 inst_704 ( .ZN(net_989), .A1(n69gat), .A2(n443gat) );
INV_X1 inst_1446 ( .ZN(net_378), .A(net_377) );
NAND2_X1 inst_1291 ( .ZN(net_1398), .A1(net_1397), .A2(net_1374) );
NAND2_X1 inst_693 ( .ZN(net_341), .A2(n341gat), .A1(n1gat) );
XNOR2_X1 inst_390 ( .ZN(net_1464), .B(net_1431), .A(net_1430) );
NAND2_X1 inst_1062 ( .ZN(net_858), .A1(net_857), .A2(net_856) );
XNOR2_X1 inst_359 ( .ZN(net_1379), .B(net_1324), .A(net_1309) );
NAND2_X1 inst_1055 ( .ZN(net_844), .A1(net_843), .A2(net_842) );
NAND2_X1 inst_1276 ( .ZN(net_1373), .A1(net_1372), .A2(net_1339) );
NAND2_X1 inst_765 ( .ZN(net_478), .A2(n358gat), .A1(n171gat) );
XNOR2_X1 inst_256 ( .ZN(net_1005), .B(net_960), .A(net_934) );
NAND2_X1 inst_694 ( .ZN(net_287), .A2(n324gat), .A1(n256gat) );
NAND2_X1 inst_630 ( .ZN(net_1405), .A1(n52gat), .A2(n511gat) );
NAND2_X1 inst_937 ( .ZN(net_609), .A1(net_550), .A2(net_499) );
XNOR2_X1 inst_401 ( .ZN(net_1512), .B(net_1478), .A(net_1464) );
NAND2_X1 inst_1273 ( .ZN(net_1362), .A2(net_1361), .A1(net_1329) );
NAND2_X1 inst_923 ( .ZN(net_530), .A1(net_529), .A2(net_528) );
NOR2_X1 inst_512 ( .ZN(net_115), .A1(net_114), .A2(net_66) );
NAND2_X1 inst_908 ( .ZN(net_523), .A2(net_477), .A1(net_420) );
XNOR2_X1 inst_355 ( .ZN(net_1330), .B(net_1295), .A(net_1294) );
NAND2_X1 inst_1301 ( .ZN(net_1427), .A1(net_1426), .A2(net_1425) );
NAND2_X1 inst_782 ( .ZN(net_138), .A1(net_137), .A2(net_136) );
XNOR2_X1 inst_218 ( .ZN(net_839), .B(net_798), .A(net_768) );
NAND2_X1 inst_647 ( .ZN(net_1391), .A2(n511gat), .A1(n35gat) );
NAND2_X1 inst_1342 ( .ZN(net_1525), .A1(net_1524), .A2(net_1474) );
XOR2_X1 inst_6 ( .Z(net_1151), .A(net_1109), .B(net_1108) );
XNOR2_X1 inst_194 ( .ZN(net_764), .A(net_730), .B(net_729) );
NAND2_X1 inst_1014 ( .ZN(net_747), .A1(net_746), .A2(net_745) );
NAND2_X1 inst_787 ( .ZN(net_187), .A1(net_186), .A2(net_167) );
NAND2_X1 inst_1347 ( .ZN(net_1533), .A1(net_1532), .A2(net_1531) );
NAND2_X1 inst_825 ( .ZN(net_303), .A1(net_302), .A2(net_301) );
AND2_X4 inst_1656 ( .ZN(net_141), .A1(net_140), .A2(net_139) );
NAND2_X1 inst_833 ( .ZN(net_322), .A1(net_321), .A2(net_280) );
XNOR2_X1 inst_123 ( .ZN(net_529), .A(net_480), .B(net_445) );
NOR2_X1 inst_509 ( .ZN(net_107), .A1(net_106), .A2(net_83) );
NAND2_X1 inst_930 ( .ZN(net_555), .A1(net_554), .A2(net_553) );
NAND2_X1 inst_699 ( .ZN(net_1053), .A2(n460gat), .A1(n239gat) );
NAND2_X1 inst_960 ( .ZN(net_639), .A1(net_597), .A2(net_533) );
INV_X1 inst_1462 ( .ZN(net_485), .A(net_484) );
XNOR2_X1 inst_118 ( .ZN(net_490), .B(net_458), .A(net_457) );
INV_X1 inst_1626 ( .ZN(net_1585), .A(net_1584) );
NAND2_X1 inst_935 ( .ZN(net_599), .A1(net_547), .A2(net_503) );
XNOR2_X1 inst_153 ( .ZN(net_637), .A(net_592), .B(net_567) );
XNOR2_X1 inst_442 ( .A(net_1615), .B(net_1614), .ZN(n6230gat) );
XNOR2_X1 inst_38 ( .ZN(net_197), .A(net_161), .B(net_160) );
XNOR2_X1 inst_381 ( .ZN(net_1423), .A(net_1397), .B(net_1375) );
INV_X1 inst_1459 ( .ZN(net_448), .A(net_447) );
NAND2_X1 inst_726 ( .ZN(net_809), .A2(n409gat), .A1(n171gat) );
XNOR2_X1 inst_295 ( .ZN(net_1136), .B(net_1097), .A(net_1068) );
NAND2_X1 inst_883 ( .ZN(net_492), .A2(net_429), .A1(net_391) );
XNOR2_X1 inst_209 ( .ZN(net_829), .B(net_796), .A(net_770) );
NAND2_X1 inst_964 ( .ZN(net_626), .A1(net_625), .A2(net_624) );
NAND2_X1 inst_1087 ( .ZN(net_926), .A1(net_925), .A2(net_893) );
XNOR2_X1 inst_40 ( .ZN(net_212), .A(net_184), .B(net_183) );
XNOR2_X1 inst_320 ( .ZN(net_1203), .B(net_1175), .A(net_1174) );
NAND2_X1 inst_1249 ( .ZN(net_1335), .A2(net_1265), .A1(net_1243) );
XNOR2_X1 inst_167 ( .ZN(net_668), .B(net_628), .A(net_627) );
NAND2_X1 inst_607 ( .ZN(net_960), .A2(n443gat), .A1(n35gat) );
NAND2_X1 inst_1320 ( .ZN(net_1472), .A1(net_1471), .A2(net_1443) );
NAND2_X1 inst_1026 ( .ZN(net_785), .A1(net_784), .A2(net_761) );
NAND2_X1 inst_756 ( .ZN(net_840), .A2(n426gat), .A1(n18gat) );
NAND2_X1 inst_1245 ( .ZN(net_1288), .A1(net_1287), .A2(net_1286) );
NAND2_X1 inst_1375 ( .ZN(net_1598), .A1(net_1597), .A2(net_1596) );
NAND2_X1 inst_1251 ( .ZN(net_1303), .A1(net_1302), .A2(net_1301) );
INV_X1 inst_1416 ( .ZN(net_167), .A(net_166) );
XNOR2_X1 inst_95 ( .ZN(net_387), .B(net_358), .A(net_357) );
NAND2_X1 inst_1318 ( .ZN(net_1467), .A1(net_1466), .A2(net_1454) );
XOR2_X1 inst_1 ( .Z(net_238), .A(net_169), .B(net_168) );
XNOR2_X1 inst_439 ( .B(net_1606), .A(net_1605), .ZN(n6200gat) );
INV_X1 inst_1485 ( .ZN(net_665), .A(net_664) );
NAND2_X1 inst_1188 ( .ZN(net_1187), .A1(net_1131), .A2(net_1080) );
NAND2_X1 inst_1165 ( .ZN(net_1137), .A2(net_1086), .A1(net_1033) );
XNOR2_X1 inst_331 ( .ZN(net_1307), .A(net_1234), .B(net_1201) );
NAND2_X1 inst_1070 ( .ZN(net_900), .A1(net_848), .A2(net_795) );
XNOR2_X1 inst_235 ( .ZN(net_914), .B(net_875), .A(net_845) );
NAND2_X1 inst_750 ( .ZN(net_977), .A1(n52gat), .A2(n443gat) );
XNOR2_X1 inst_317 ( .ZN(net_1218), .B(net_1167), .A(net_1132) );
NAND2_X1 inst_1123 ( .ZN(net_1012), .A1(net_1011), .A2(net_986) );
NAND2_X1 inst_1082 ( .ZN(net_936), .A1(net_895), .A2(net_834) );
NAND2_X1 inst_667 ( .ZN(net_8), .A2(n273gat), .A1(n171gat) );
XNOR2_X1 inst_278 ( .ZN(net_1079), .A(net_1009), .B(net_994) );
NOR2_X1 inst_467 ( .ZN(net_43), .A1(net_9), .A2(net_8) );
NAND2_X1 inst_992 ( .ZN(net_704), .A1(net_703), .A2(net_702) );
XNOR2_X1 inst_105 ( .ZN(net_437), .B(net_422), .A(net_421) );
NOR2_X1 inst_488 ( .ZN(net_92), .A2(net_53), .A1(net_10) );
XNOR2_X1 inst_387 ( .ZN(net_1453), .B(net_1418), .A(net_1417) );
AND2_X4 inst_1628 ( .ZN(net_13), .A2(n290gat), .A1(n222gat) );
NAND2_X1 inst_997 ( .ZN(net_713), .A1(net_699), .A2(net_665) );
NAND2_X1 inst_1329 ( .ZN(net_1495), .A1(net_1494), .A2(net_1450) );
NAND2_X1 inst_857 ( .ZN(net_400), .A2(net_353), .A1(net_322) );
NAND2_X1 inst_1204 ( .ZN(net_1207), .A1(net_1206), .A2(net_1205) );
XNOR2_X1 inst_254 ( .ZN(net_975), .A(net_937), .B(net_936) );
NAND2_X1 inst_654 ( .ZN(net_554), .A1(n52gat), .A2(n375gat) );
NAND2_X1 inst_625 ( .ZN(net_1206), .A1(n86gat), .A2(n477gat) );
XNOR2_X1 inst_225 ( .ZN(net_950), .A(net_847), .B(net_827) );
INV_X1 inst_1511 ( .ZN(net_826), .A(net_825) );
NOR2_X1 inst_508 ( .ZN(net_105), .A1(net_104), .A2(net_81) );
NAND2_X1 inst_568 ( .ZN(net_1211), .A2(n477gat), .A1(n256gat) );
INV_X1 inst_1483 ( .ZN(net_648), .A(net_647) );
INV_X1 inst_1412 ( .ZN(net_86), .A(net_85) );
NOR2_X1 inst_523 ( .ZN(net_198), .A2(net_165), .A1(net_101) );
XNOR2_X1 inst_365 ( .ZN(net_1367), .A(net_1336), .B(net_1335) );
INV_X1 inst_1492 ( .ZN(net_681), .A(net_680) );
NAND2_X1 inst_1181 ( .ZN(net_1169), .A1(net_1117), .A2(net_1059) );
XNOR2_X1 inst_67 ( .ZN(net_318), .A(net_254), .B(net_234) );
NAND2_X1 inst_954 ( .ZN(net_610), .A1(net_609), .A2(net_578) );
XNOR2_X1 inst_181 ( .ZN(net_757), .A(net_699), .B(net_664) );
NAND2_X1 inst_1153 ( .ZN(net_1080), .A1(net_1079), .A2(net_1078) );
NAND2_X1 inst_1135 ( .ZN(net_1057), .A2(net_1008), .A1(net_955) );
INV_X1 inst_1504 ( .ZN(net_777), .A(net_776) );
XNOR2_X1 inst_391 ( .ZN(net_1482), .B(net_1437), .A(net_1387) );
NAND2_X1 inst_661 ( .ZN(net_2), .A2(n273gat), .A1(n222gat) );
NAND2_X1 inst_590 ( .ZN(net_346), .A2(n341gat), .A1(n18gat) );
INV_X1 inst_1548 ( .ZN(net_1069), .A(net_1068) );
NAND2_X1 inst_713 ( .ZN(net_252), .A2(n324gat), .A1(n222gat) );
NAND2_X1 inst_1310 ( .ZN(net_1475), .A1(net_1416), .A2(net_1377) );
XNOR2_X1 inst_202 ( .ZN(net_780), .A(net_752), .B(net_751) );
INV_X1 inst_1401 ( .ZN(net_70), .A(net_61) );
NAND2_X1 inst_634 ( .ZN(net_260), .A2(n324gat), .A1(n103gat) );
XNOR2_X1 inst_419 ( .ZN(net_1597), .B(net_1551), .A(net_1536) );
NAND2_X1 inst_1105 ( .ZN(net_961), .A1(net_960), .A2(net_935) );
NAND2_X1 inst_981 ( .ZN(net_686), .A1(net_685), .A2(net_684) );
NOR2_X1 inst_477 ( .ZN(net_98), .A2(net_31), .A1(net_16) );
NAND2_X1 inst_1368 ( .ZN(net_1592), .A1(net_1568), .A2(net_1525) );
NAND2_X1 inst_1266 ( .ZN(net_1348), .A1(net_1347), .A2(net_1312) );
XNOR2_X1 inst_423 ( .ZN(net_1600), .B(net_1552), .A(net_1534) );
NAND2_X1 inst_1069 ( .ZN(net_876), .A1(net_875), .A2(net_846) );
NAND2_X1 inst_835 ( .ZN(net_342), .A1(net_341), .A2(net_340) );
XNOR2_X1 inst_136 ( .ZN(net_561), .B(net_520), .A(net_519) );
XNOR2_X1 inst_30 ( .ZN(net_209), .A(net_131), .B(net_130) );
XNOR2_X1 inst_330 ( .ZN(net_1249), .B(net_1219), .A(net_1218) );
NAND2_X1 inst_610 ( .ZN(net_830), .A2(n426gat), .A1(n1gat) );
NAND2_X1 inst_1112 ( .ZN(net_1004), .A2(net_944), .A1(net_879) );
NAND2_X1 inst_1036 ( .ZN(net_806), .A1(net_805), .A2(net_777) );
XNOR2_X1 inst_233 ( .ZN(net_890), .B(net_857), .A(net_856) );
NAND2_X1 inst_710 ( .ZN(net_557), .A2(n375gat), .A1(n35gat) );
XNOR2_X1 inst_165 ( .ZN(net_664), .B(net_643), .A(net_642) );
INV_X1 inst_1526 ( .ZN(net_933), .A(net_932) );
INV_X1 inst_1477 ( .ZN(net_578), .A(net_577) );
NAND2_X1 inst_1379 ( .ZN(net_1604), .A1(net_1603), .A2(net_1602) );
NAND2_X1 inst_941 ( .ZN(net_587), .A1(net_586), .A2(net_562) );
XNOR2_X1 inst_271 ( .ZN(net_1029), .A(net_1002), .B(net_1001) );
XNOR2_X1 inst_34 ( .ZN(net_191), .B(net_155), .A(net_154) );
NAND2_X1 inst_1176 ( .ZN(net_1158), .A2(net_1105), .A1(net_1067) );
XNOR2_X1 inst_12 ( .ZN(net_127), .A(net_102), .B(net_76) );
NAND2_X1 inst_1047 ( .ZN(net_857), .A2(net_812), .A1(net_756) );
NAND2_X1 inst_529 ( .ZN(net_1347), .A2(n494gat), .A1(n120gat) );
XNOR2_X1 inst_56 ( .ZN(net_301), .A(net_246), .B(net_218) );
XNOR2_X1 inst_71 ( .ZN(net_328), .B(net_311), .A(net_310) );
XNOR2_X1 inst_308 ( .A(net_1140), .B(net_1139), .ZN(n5308gat) );
INV_X1 inst_1546 ( .ZN(net_1047), .A(net_1046) );
INV_X1 inst_1528 ( .ZN(net_940), .A(net_939) );
NAND2_X1 inst_1230 ( .ZN(net_1304), .A1(net_1233), .A2(net_1213) );
INV_X1 inst_1454 ( .ZN(net_438), .A(net_437) );
XNOR2_X1 inst_60 ( .ZN(net_295), .B(net_252), .A(net_236) );
OR2_X4 inst_455 ( .ZN(net_182), .A1(net_181), .A2(net_180) );
NAND2_X1 inst_1232 ( .ZN(net_1286), .A1(net_1237), .A2(net_1176) );
INV_X1 inst_1424 ( .ZN(net_227), .A(net_226) );
NAND2_X1 inst_1064 ( .ZN(net_863), .A1(net_862), .A2(net_861) );
NAND2_X1 inst_1313 ( .ZN(net_1458), .A1(net_1457), .A2(net_1436) );
INV_X1 inst_1425 ( .ZN(net_229), .A(net_228) );
NAND2_X1 inst_1334 ( .ZN(net_1542), .A2(net_1470), .A1(net_1410) );
NAND2_X1 inst_675 ( .ZN(net_791), .A2(n409gat), .A1(n103gat) );
NAND2_X1 inst_758 ( .ZN(net_694), .A2(n392gat), .A1(n205gat) );
NOR2_X1 inst_496 ( .A2(net_110), .ZN(net_66), .A1(net_47) );
NAND2_X1 inst_860 ( .ZN(net_422), .A2(net_370), .A1(net_293) );
XNOR2_X1 inst_336 ( .ZN(net_1284), .A(net_1221), .B(net_1200) );
NAND2_X1 inst_563 ( .ZN(net_941), .A2(n443gat), .A1(n239gat) );
NAND2_X1 inst_583 ( .ZN(net_1055), .A2(n460gat), .A1(n18gat) );
NAND2_X1 inst_943 ( .ZN(net_591), .A1(net_590), .A2(net_566) );
XNOR2_X1 inst_258 ( .ZN(net_985), .B(net_951), .A(net_950) );
XNOR2_X1 inst_376 ( .ZN(net_1476), .B(net_1389), .A(net_1367) );
XNOR2_X1 inst_143 ( .ZN(net_575), .B(net_546), .A(net_545) );
AND2_X4 inst_1633 ( .ZN(net_14), .A2(n273gat), .A1(n18gat) );
NAND2_X1 inst_1262 ( .ZN(net_1334), .A1(net_1333), .A2(net_1332) );
NAND2_X1 inst_1243 ( .ZN(net_1319), .A2(net_1259), .A1(net_1212) );
XNOR2_X1 inst_265 ( .ZN(net_1032), .B(net_989), .A(net_956) );
NAND2_X1 inst_1211 ( .ZN(net_1222), .A1(net_1221), .A2(net_1199) );
NOR2_X1 inst_482 ( .ZN(net_50), .A2(net_43), .A1(net_9) );
NAND2_X1 inst_1192 ( .ZN(net_1198), .A2(net_1141), .A1(net_1090) );
INV_X1 inst_1593 ( .ZN(net_1366), .A(net_1365) );
NAND2_X1 inst_1040 ( .ZN(net_814), .A1(net_813), .A2(net_773) );
NAND2_X1 inst_682 ( .ZN(net_658), .A2(n392gat), .A1(n18gat) );
NAND2_X1 inst_736 ( .ZN(net_849), .A2(n426gat), .A1(n35gat) );
NAND2_X1 inst_544 ( .ZN(net_927), .A2(n426gat), .A1(n120gat) );
XNOR2_X1 inst_238 ( .ZN(net_911), .A(net_897), .B(net_896) );
NAND2_X1 inst_1093 ( .ZN(net_967), .A2(net_924), .A1(net_858) );
NAND2_X1 inst_539 ( .ZN(net_1221), .A2(n477gat), .A1(n171gat) );
NAND2_X1 inst_724 ( .ZN(net_123), .A2(n307gat), .A1(n1gat) );
NAND2_X1 inst_895 ( .ZN(net_481), .A1(net_480), .A2(net_446) );
XNOR2_X1 inst_178 ( .ZN(net_700), .A(net_685), .B(net_684) );
INV_X1 inst_1596 ( .ZN(net_1382), .A(net_1381) );
XNOR2_X1 inst_111 ( .ZN(net_449), .B(net_428), .A(net_427) );
NAND2_X1 inst_975 ( .ZN(net_659), .A1(net_658), .A2(net_657) );
INV_X1 inst_1430 ( .ZN(net_245), .A(net_244) );
NAND2_X1 inst_734 ( .ZN(net_1440), .A2(n528gat), .A1(n1gat) );
NAND2_X1 inst_1282 ( .ZN(net_1411), .A1(net_1356), .A2(net_1308) );
NAND2_X1 inst_1077 ( .ZN(net_904), .A1(net_903), .A2(net_902) );
NAND2_X1 inst_1210 ( .ZN(net_1220), .A1(net_1219), .A2(net_1218) );
NAND2_X1 inst_1148 ( .ZN(net_1065), .A1(net_1064), .A2(net_1063) );
INV_X1 inst_1435 ( .ZN(net_281), .A(net_280) );
INV_X1 inst_1431 ( .ZN(net_273), .A(net_272) );
NAND2_X1 inst_1398 ( .ZN(net_1632), .A2(net_1631), .A1(net_1539) );
XNOR2_X1 inst_222 ( .ZN(net_899), .B(net_837), .A(net_815) );
XNOR2_X1 inst_284 ( .ZN(net_1083), .A(net_1049), .B(net_1048) );
INV_X1 inst_1555 ( .ZN(net_1100), .A(net_1099) );
NAND2_X1 inst_806 ( .ZN(net_311), .A2(net_257), .A1(net_179) );
NAND2_X1 inst_1293 ( .ZN(net_1406), .A1(net_1405), .A2(net_1404) );
XNOR2_X1 inst_280 ( .A(net_1037), .B(net_1036), .ZN(n4946gat) );
NAND2_X1 inst_763 ( .ZN(net_685), .A2(n392gat), .A1(n256gat) );
XNOR2_X1 inst_346 ( .ZN(net_1299), .B(net_1264), .A(net_1263) );
NOR2_X1 inst_491 ( .A2(net_104), .ZN(net_83), .A1(net_57) );
INV_X1 inst_1467 ( .ZN(net_537), .A(net_536) );
NAND2_X1 inst_1302 ( .ZN(net_1429), .A1(net_1428), .A2(net_1400) );
NAND2_X1 inst_1280 ( .ZN(net_1377), .A1(net_1376), .A2(net_1300) );
NAND2_X1 inst_1052 ( .ZN(net_834), .A1(net_833), .A2(net_832) );
NAND2_X1 inst_978 ( .ZN(net_677), .A1(net_676), .A2(net_646) );
AND2_X4 inst_1648 ( .ZN(net_104), .A2(net_49), .A1(net_18) );
NAND2_X1 inst_1079 ( .ZN(net_908), .A1(net_907), .A2(net_884) );
NAND2_X1 inst_842 ( .ZN(net_361), .A1(net_360), .A2(net_326) );
NAND2_X1 inst_537 ( .ZN(net_789), .A2(n409gat), .A1(n256gat) );
NAND2_X1 inst_826 ( .ZN(net_305), .A2(net_304), .A1(net_245) );
NAND2_X1 inst_551 ( .ZN(net_452), .A1(n35gat), .A2(n358gat) );
INV_X1 inst_1513 ( .ZN(net_836), .A(net_835) );
NAND2_X1 inst_1155 ( .ZN(net_1108), .A2(net_1054), .A1(net_1003) );
NAND2_X1 inst_1051 ( .ZN(net_862), .A2(net_814), .A1(net_759) );
XNOR2_X1 inst_207 ( .ZN(net_832), .B(net_791), .A(net_764) );
XNOR2_X1 inst_353 ( .ZN(net_1311), .A(net_1287), .B(net_1286) );
NOR2_X1 inst_495 ( .A2(net_120), .ZN(net_79), .A1(net_36) );
NOR2_X1 inst_506 ( .ZN(net_101), .A1(net_100), .A2(net_73) );
XNOR2_X1 inst_159 ( .ZN(net_654), .B(net_607), .A(net_581) );
NAND2_X1 inst_872 ( .ZN(net_408), .A1(net_407), .A2(net_378) );
NAND2_X1 inst_951 ( .ZN(net_604), .A1(net_603), .A2(net_580) );
XNOR2_X1 inst_134 ( .ZN(net_543), .B(net_514), .A(net_513) );
INV_X1 inst_1545 ( .ZN(net_1045), .A(net_1044) );
NAND2_X1 inst_1323 ( .ZN(net_1477), .A1(net_1476), .A2(net_1475) );
NAND2_X1 inst_1085 ( .ZN(net_922), .A1(net_921), .A2(net_887) );
XNOR2_X1 inst_333 ( .ZN(net_1251), .B(net_1224), .A(net_1223) );
NAND2_X1 inst_712 ( .ZN(net_573), .A2(n375gat), .A1(n103gat) );
NAND2_X1 inst_1215 ( .ZN(net_1230), .A1(net_1229), .A2(net_1197) );
NAND2_X1 inst_1349 ( .ZN(net_1539), .A2(net_1538), .A1(net_1481) );
XNOR2_X1 inst_131 ( .ZN(net_548), .B(net_498), .A(net_488) );
XNOR2_X1 inst_406 ( .ZN(net_1519), .B(net_1486), .A(net_1485) );
XNOR2_X1 inst_160 ( .ZN(net_622), .B(net_605), .A(net_543) );
OR2_X4 inst_462 ( .ZN(net_208), .A1(net_207), .A2(net_206) );
XNOR2_X1 inst_328 ( .ZN(net_1240), .A(net_1211), .B(net_1210) );
NAND2_X1 inst_869 ( .ZN(net_401), .A1(net_400), .A2(net_386) );
NAND2_X1 inst_1359 ( .ZN(net_1582), .A1(net_1545), .A2(net_1499) );
XNOR2_X1 inst_19 ( .ZN(net_133), .A(net_98), .B(net_78) );
XNOR2_X1 inst_47 ( .ZN(net_228), .A(net_192), .B(net_191) );
XOR2_X1 inst_8 ( .Z(net_1459), .A(net_1421), .B(net_1420) );
NAND2_X1 inst_818 ( .ZN(net_306), .A2(net_251), .A1(net_176) );
XNOR2_X1 inst_370 ( .ZN(net_1404), .B(net_1363), .A(net_1330) );
NAND2_X1 inst_762 ( .ZN(net_1469), .A2(n528gat), .A1(n18gat) );
NAND2_X1 inst_573 ( .ZN(net_958), .A2(n443gat), .A1(n222gat) );
NAND2_X1 inst_1265 ( .ZN(net_1346), .A1(net_1345), .A2(net_1323) );
XNOR2_X1 inst_100 ( .ZN(net_451), .B(net_402), .A(net_379) );
NAND2_X1 inst_965 ( .ZN(net_629), .A1(net_628), .A2(net_627) );
INV_X1 inst_1453 ( .ZN(net_433), .A(net_432) );
NAND2_X1 inst_921 ( .ZN(net_524), .A1(net_523), .A2(net_522) );
XNOR2_X1 inst_279 ( .ZN(net_1051), .A(net_1032), .B(net_1031) );
XNOR2_X1 inst_81 ( .ZN(net_348), .A(net_308), .B(net_279) );
NAND2_X1 inst_612 ( .ZN(net_546), .A1(n69gat), .A2(n375gat) );
NAND2_X1 inst_1321 ( .ZN(net_1498), .A2(net_1446), .A1(net_1396) );
NOR2_X1 inst_525 ( .ZN(net_204), .A2(net_162), .A1(net_93) );
NAND2_X1 inst_1012 ( .ZN(net_741), .A1(net_740), .A2(net_739) );
NAND2_X1 inst_901 ( .ZN(net_500), .A2(net_464), .A1(net_393) );
XNOR2_X1 inst_434 ( .ZN(net_1614), .B(net_1592), .A(net_1569) );
NAND2_X1 inst_790 ( .ZN(net_243), .A1(net_242), .A2(net_241) );
NAND2_X1 inst_1032 ( .ZN(net_797), .A1(net_796), .A2(net_771) );
NAND2_X1 inst_1009 ( .ZN(net_731), .A1(net_730), .A2(net_729) );
NAND2_X1 inst_1206 ( .ZN(net_1212), .A1(net_1211), .A2(net_1210) );
NAND2_X1 inst_751 ( .ZN(net_1130), .A2(n460gat), .A1(n137gat) );
NAND2_X1 inst_906 ( .ZN(net_517), .A2(net_475), .A1(net_414) );
NAND2_X1 inst_845 ( .ZN(net_368), .A1(net_367), .A2(net_337) );
NAND2_X1 inst_1248 ( .ZN(net_1298), .A1(net_1297), .A2(net_1282) );
NAND2_X1 inst_1367 ( .ZN(net_1579), .A1(net_1578), .A2(net_1577) );
NAND2_X1 inst_1392 ( .ZN(net_1624), .A2(net_1622), .A1(net_1576) );
NAND2_X1 inst_733 ( .ZN(net_727), .A2(n409gat), .A1(n1gat) );
XNOR2_X1 inst_377 ( .ZN(net_1425), .B(net_1383), .A(net_1349) );
INV_X1 inst_1476 ( .ZN(net_576), .A(net_575) );
XNOR2_X1 inst_142 ( .ZN(net_598), .B(net_571), .A(net_534) );
XNOR2_X1 inst_78 ( .ZN(net_354), .A(net_299), .B(net_275) );
INV_X1 inst_1487 ( .ZN(net_669), .A(net_668) );
INV_X1 inst_1460 ( .ZN(net_450), .A(net_449) );
NAND2_X1 inst_1344 ( .ZN(net_1552), .A2(net_1511), .A1(net_1456) );
XNOR2_X1 inst_177 ( .ZN(net_718), .B(net_687), .A(net_660) );
NAND2_X1 inst_783 ( .ZN(net_168), .A2(net_126), .A1(net_64) );
NAND2_X1 inst_885 ( .ZN(net_462), .A1(net_461), .A2(net_460) );
INV_X1 inst_1436 ( .ZN(net_283), .A(net_282) );
XNOR2_X1 inst_183 ( .ZN(net_752), .A(net_696), .B(net_672) );
INV_X1 inst_1443 ( .ZN(net_337), .A(net_336) );
NAND2_X1 inst_852 ( .ZN(net_405), .A2(net_364), .A1(net_298) );
NAND2_X1 inst_1142 ( .ZN(net_1050), .A1(net_1049), .A2(net_1048) );
NAND2_X1 inst_928 ( .ZN(net_583), .A2(net_515), .A1(net_494) );
NAND2_X1 inst_1028 ( .ZN(net_818), .A2(net_763), .A1(net_704) );
XNOR2_X1 inst_107 ( .ZN(net_441), .B(net_410), .A(net_409) );
XNOR2_X1 inst_393 ( .A(net_1440), .B(net_1439), .ZN(n6123gat) );
NAND2_X1 inst_615 ( .ZN(net_10), .A2(n273gat), .A1(n120gat) );
INV_X1 inst_1474 ( .ZN(net_568), .A(net_567) );
NAND2_X1 inst_990 ( .ZN(net_698), .A1(net_690), .A2(net_669) );
INV_X1 inst_1539 ( .ZN(net_996), .A(net_995) );
XNOR2_X1 inst_92 ( .ZN(net_418), .A(net_371), .B(net_338) );
XNOR2_X1 inst_345 ( .ZN(net_1289), .B(net_1278), .A(net_1277) );
NAND2_X1 inst_1271 ( .ZN(net_1385), .A1(net_1327), .A2(net_1279) );
NAND2_X1 inst_1050 ( .ZN(net_854), .A2(net_810), .A1(net_753) );
NAND2_X1 inst_1381 ( .ZN(net_1607), .A1(net_1606), .A2(net_1605) );
NAND2_X1 inst_643 ( .ZN(net_687), .A2(n392gat), .A1(n103gat) );
NAND2_X1 inst_1311 ( .ZN(net_1478), .A2(net_1419), .A1(net_1360) );
NAND2_X1 inst_697 ( .ZN(net_254), .A2(n324gat), .A1(n171gat) );
NOR2_X1 inst_487 ( .ZN(net_108), .A2(net_33), .A1(net_28) );
NAND2_X1 inst_1296 ( .ZN(net_1416), .A1(net_1415), .A2(net_1414) );
AND2_X4 inst_1640 ( .ZN(net_25), .A1(n52gat), .A2(n290gat) );
XNOR2_X1 inst_200 ( .ZN(net_776), .A(net_749), .B(net_748) );
XNOR2_X1 inst_57 ( .ZN(net_272), .A(net_250), .B(net_224) );
XNOR2_X1 inst_338 ( .ZN(net_1263), .B(net_1242), .A(net_1181) );
INV_X1 inst_1557 ( .ZN(net_1133), .A(net_1132) );
INV_X1 inst_1553 ( .ZN(net_1094), .A(net_1093) );
NAND2_X1 inst_1237 ( .ZN(net_1306), .A1(net_1248), .A2(net_1189) );
XNOR2_X1 inst_417 ( .ZN(net_1560), .B(net_1529), .A(net_1528) );
NAND2_X1 inst_671 ( .ZN(net_1483), .A2(n528gat), .A1(n222gat) );
AND2_X4 inst_1635 ( .ZN(net_18), .A1(n86gat), .A2(n273gat) );
INV_X1 inst_1616 ( .ZN(net_1520), .A(net_1519) );
NAND2_X1 inst_1307 ( .ZN(net_1441), .A1(net_1440), .A2(net_1439) );
NAND2_X1 inst_1017 ( .ZN(net_756), .A1(net_755), .A2(net_754) );
XNOR2_X1 inst_21 ( .ZN(net_148), .A(net_104), .B(net_82) );
NAND2_X1 inst_579 ( .ZN(net_7), .A2(n290gat), .A1(n171gat) );
INV_X1 inst_1500 ( .ZN(net_769), .A(net_768) );
XNOR2_X1 inst_281 ( .ZN(net_1068), .A(net_1042), .B(net_1041) );
NAND2_X1 inst_1094 ( .ZN(net_970), .A2(net_926), .A1(net_863) );
INV_X1 inst_1606 ( .ZN(net_1454), .A(net_1453) );
NAND2_X1 inst_585 ( .ZN(net_1345), .A2(n494gat), .A1(n154gat) );
NAND2_X1 inst_698 ( .ZN(net_28), .A2(n273gat), .A1(n205gat) );
NAND2_X1 inst_893 ( .ZN(net_477), .A1(net_476), .A2(net_448) );
XNOR2_X1 inst_88 ( .ZN(net_381), .B(net_363), .A(net_362) );
XNOR2_X1 inst_410 ( .ZN(net_1555), .A(net_1500), .B(net_1489) );
XNOR2_X1 inst_316 ( .ZN(net_1196), .B(net_1165), .A(net_1164) );
XNOR2_X1 inst_220 ( .A(net_830), .B(net_829), .ZN(n4241gat) );
INV_X1 inst_1585 ( .ZN(net_1329), .A(net_1328) );
NAND2_X1 inst_1317 ( .ZN(net_1502), .A2(net_1432), .A1(net_1386) );
NAND2_X1 inst_851 ( .ZN(net_407), .A2(net_350), .A1(net_309) );
NAND2_X1 inst_831 ( .ZN(net_317), .A1(net_316), .A2(net_272) );
NAND2_X1 inst_1174 ( .ZN(net_1129), .A1(net_1128), .A2(net_1099) );
XNOR2_X1 inst_360 ( .ZN(net_1351), .B(net_1317), .A(net_1316) );
XNOR2_X1 inst_383 ( .ZN(net_1435), .B(net_1405), .A(net_1404) );
NAND2_X1 inst_1023 ( .ZN(net_801), .A2(net_736), .A1(net_710) );
XNOR2_X1 inst_50 ( .ZN(net_234), .B(net_210), .A(net_209) );
NAND2_X1 inst_773 ( .ZN(net_65), .A2(net_30), .A1(net_14) );
XNOR2_X1 inst_245 ( .ZN(net_969), .A(net_923), .B(net_890) );
NAND2_X1 inst_569 ( .ZN(net_1085), .A1(n52gat), .A2(n460gat) );
NAND2_X1 inst_1080 ( .ZN(net_910), .A1(net_909), .A2(net_888) );
NAND2_X1 inst_1124 ( .ZN(net_1014), .A1(net_1013), .A2(net_984) );
NAND2_X1 inst_678 ( .ZN(net_1471), .A2(n511gat), .A1(n137gat) );
NAND2_X1 inst_624 ( .ZN(net_655), .A2(n392gat), .A1(n35gat) );
NAND2_X1 inst_1103 ( .ZN(net_955), .A1(net_954), .A2(net_953) );
XNOR2_X1 inst_260 ( .ZN(net_1019), .B(net_977), .A(net_939) );
NAND2_X1 inst_1129 ( .ZN(net_1024), .A1(net_1023), .A2(net_996) );
NAND2_X1 inst_854 ( .ZN(net_396), .A2(net_356), .A1(net_300) );
XNOR2_X1 inst_147 ( .ZN(net_634), .A(net_551), .B(net_537) );
NAND2_X1 inst_837 ( .ZN(net_389), .A2(net_325), .A1(net_288) );
XNOR2_X1 inst_313 ( .ZN(net_1205), .A(net_1160), .B(net_1135) );
NAND2_X1 inst_744 ( .ZN(net_1266), .A2(n494gat), .A1(n35gat) );
AND2_X4 inst_1650 ( .ZN(net_57), .A2(net_49), .A1(net_19) );
NAND2_X1 inst_549 ( .ZN(net_740), .A2(n409gat), .A1(n18gat) );
NAND2_X1 inst_1041 ( .ZN(net_833), .A2(net_785), .A1(net_719) );
XNOR2_X1 inst_234 ( .ZN(net_892), .B(net_862), .A(net_861) );
INV_X1 inst_1497 ( .ZN(net_733), .A(net_732) );
NOR2_X1 inst_522 ( .ZN(net_207), .A2(net_141), .A1(net_107) );
XNOR2_X1 inst_236 ( .ZN(net_918), .B(net_880), .A(net_871) );
NAND2_X1 inst_1002 ( .ZN(net_742), .A1(net_693), .A2(net_632) );
NOR2_X1 inst_478 ( .ZN(net_40), .A2(net_39), .A1(net_21) );
NAND2_X1 inst_553 ( .ZN(net_1341), .A2(n511gat), .A1(n1gat) );
XNOR2_X1 inst_65 ( .ZN(net_284), .A(net_264), .B(net_226) );
NAND2_X1 inst_1304 ( .ZN(net_1466), .A2(net_1403), .A1(net_1362) );
NAND2_X1 inst_536 ( .ZN(net_514), .A2(n375gat), .A1(n239gat) );
NAND2_X1 inst_1328 ( .ZN(net_1487), .A1(net_1486), .A2(net_1485) );
XNOR2_X1 inst_242 ( .ZN(net_934), .A(net_903), .B(net_902) );
NAND2_X1 inst_986 ( .ZN(net_692), .A1(net_691), .A2(net_675) );
INV_X1 inst_1618 ( .ZN(net_1537), .A(net_1536) );
INV_X1 inst_1422 ( .ZN(net_223), .A(net_222) );
NAND2_X1 inst_688 ( .ZN(net_149), .A1(n69gat), .A2(n307gat) );
NOR2_X1 inst_516 ( .ZN(net_172), .A2(net_147), .A1(net_91) );
NAND2_X1 inst_804 ( .ZN(net_271), .A1(net_270), .A2(net_213) );
NAND2_X1 inst_1186 ( .ZN(net_1153), .A1(net_1152), .A2(net_1151) );
XNOR2_X1 inst_190 ( .ZN(net_732), .A(net_715), .B(net_714) );
NAND2_X1 inst_1267 ( .ZN(net_1376), .A2(net_1315), .A1(net_1271) );
INV_X1 inst_1507 ( .ZN(net_783), .A(net_782) );
XNOR2_X1 inst_13 ( .ZN(net_163), .A(net_100), .B(net_74) );
NAND2_X1 inst_919 ( .ZN(net_518), .A1(net_517), .A2(net_516) );
NAND2_X1 inst_1221 ( .ZN(net_1243), .A2(net_1242), .A1(net_1182) );
NAND2_X1 inst_1166 ( .ZN(net_1112), .A1(net_1111), .A2(net_1087) );
XNOR2_X1 inst_116 ( .ZN(net_488), .B(net_452), .A(net_451) );
XNOR2_X1 inst_416 ( .ZN(net_1578), .B(net_1542), .A(net_1519) );
NAND2_X1 inst_598 ( .ZN(net_264), .A2(n324gat), .A1(n18gat) );
NAND2_X1 inst_1158 ( .ZN(net_1090), .A1(net_1089), .A2(net_1074) );
NAND2_X1 inst_1133 ( .ZN(net_1038), .A1(net_1037), .A2(net_1036) );
NOR2_X1 inst_471 ( .ZN(net_39), .A1(net_21), .A2(net_20) );
NAND2_X1 inst_799 ( .ZN(net_263), .A1(net_262), .A2(net_229) );
XNOR2_X1 inst_219 ( .ZN(net_835), .B(net_818), .A(net_817) );
NAND2_X1 inst_738 ( .ZN(net_1314), .A2(n494gat), .A1(n205gat) );
INV_X1 inst_1624 ( .ZN(net_1570), .A(net_1569) );
NAND2_X1 inst_719 ( .ZN(net_1326), .A2(n494gat), .A1(n103gat) );
NAND2_X1 inst_840 ( .ZN(net_356), .A1(net_355), .A2(net_354) );
NAND2_X1 inst_1220 ( .ZN(net_1260), .A2(net_1209), .A1(net_1148) );
INV_X1 inst_1406 ( .ZN(net_74), .A(net_73) );
INV_X1 inst_1456 ( .ZN(net_442), .A(net_441) );
XNOR2_X1 inst_255 ( .ZN(net_979), .B(net_958), .A(net_932) );
NAND2_X1 inst_542 ( .ZN(net_1104), .A2(n460gat), .A1(n205gat) );
XNOR2_X1 inst_128 ( .ZN(net_534), .B(net_496), .A(net_495) );
OR2_X4 inst_453 ( .ZN(net_176), .A1(net_175), .A2(net_174) );
NAND2_X1 inst_1134 ( .ZN(net_1066), .A2(net_1012), .A1(net_952) );
NOR2_X1 inst_493 ( .A2(net_100), .ZN(net_81), .A1(net_45) );
XNOR2_X1 inst_23 ( .ZN(net_145), .A(net_90), .B(net_72) );
NAND2_X1 inst_896 ( .ZN(net_508), .A2(net_453), .A1(net_403) );
XNOR2_X1 inst_339 ( .ZN(net_1336), .B(net_1258), .A(net_1240) );
NAND2_X1 inst_1113 ( .ZN(net_982), .A2(net_981), .A1(net_962) );
XNOR2_X1 inst_351 ( .ZN(net_1340), .B(net_1304), .A(net_1268) );
INV_X1 inst_1609 ( .ZN(net_1474), .A(net_1473) );
XNOR2_X1 inst_408 ( .ZN(net_1534), .B(net_1507), .A(net_1506) );
NAND2_X1 inst_973 ( .ZN(net_653), .A1(net_652), .A2(net_622) );
NAND2_X1 inst_1144 ( .ZN(net_1056), .A1(net_1055), .A2(net_1035) );
XNOR2_X1 inst_325 ( .ZN(net_1253), .B(net_1208), .A(net_1179) );
OR2_X4 inst_461 ( .ZN(net_205), .A1(net_204), .A2(net_203) );
XNOR2_X1 inst_385 ( .ZN(net_1449), .B(net_1415), .A(net_1414) );
NAND2_X1 inst_829 ( .ZN(net_312), .A1(net_311), .A2(net_310) );
NAND2_X1 inst_812 ( .ZN(net_319), .A2(net_263), .A1(net_193) );
NAND2_X1 inst_1197 ( .ZN(net_1178), .A1(net_1177), .A2(net_1145) );
XNOR2_X1 inst_197 ( .ZN(net_770), .B(net_740), .A(net_739) );
XNOR2_X1 inst_179 ( .ZN(net_730), .B(net_689), .A(net_666) );
XNOR2_X1 inst_24 ( .ZN(net_201), .B(net_125), .A(net_116) );
NAND2_X1 inst_955 ( .ZN(net_643), .A1(net_587), .A2(net_521) );
XNOR2_X1 inst_114 ( .ZN(net_484), .B(net_455), .A(net_454) );
NAND2_X1 inst_1122 ( .ZN(net_1010), .A1(net_1009), .A2(net_993) );
NAND2_X1 inst_1209 ( .ZN(net_1217), .A1(net_1216), .A2(net_1191) );
XNOR2_X1 inst_76 ( .ZN(net_334), .A(net_295), .B(net_294) );
NAND2_X1 inst_617 ( .ZN(net_239), .A2(n324gat), .A1(n239gat) );
INV_X1 inst_1560 ( .ZN(net_1145), .A(net_1144) );
INV_X1 inst_1611 ( .ZN(net_1489), .A(net_1488) );
NAND2_X1 inst_1127 ( .ZN(net_1020), .A1(net_1019), .A2(net_1018) );
XNOR2_X1 inst_150 ( .ZN(net_627), .A(net_586), .B(net_561) );
XNOR2_X1 inst_172 ( .ZN(net_678), .B(net_650), .A(net_649) );
XNOR2_X1 inst_362 ( .ZN(net_1412), .A(net_1345), .B(net_1322) );
INV_X1 inst_1530 ( .ZN(net_957), .A(net_956) );
XNOR2_X1 inst_277 ( .ZN(net_1046), .A(net_1019), .B(net_1018) );
INV_X1 inst_1510 ( .ZN(net_821), .A(net_820) );
XNOR2_X1 inst_83 ( .A(net_341), .B(net_340), .ZN(n2548gat) );
XNOR2_X1 inst_121 ( .ZN(net_526), .A(net_463), .B(net_433) );
NAND2_X1 inst_887 ( .ZN(net_467), .A1(net_466), .A2(net_465) );
XNOR2_X1 inst_306 ( .ZN(net_1144), .B(net_1121), .A(net_1120) );
NAND2_X1 inst_534 ( .ZN(net_615), .A2(n392gat), .A1(n239gat) );
NAND2_X1 inst_1065 ( .ZN(net_866), .A1(net_865), .A2(net_864) );
NAND2_X1 inst_1057 ( .ZN(net_850), .A1(net_849), .A2(net_826) );
NAND2_X1 inst_596 ( .ZN(net_539), .A2(n375gat), .A1(n1gat) );
AND2_X4 inst_1663 ( .ZN(net_162), .A1(net_161), .A2(net_160) );
XNOR2_X1 inst_90 ( .ZN(net_383), .B(net_346), .A(net_345) );
XNOR2_X1 inst_140 ( .ZN(net_569), .A(net_529), .B(net_528) );
XNOR2_X1 inst_267 ( .ZN(net_1036), .A(net_981), .B(net_963) );
NAND2_X1 inst_847 ( .ZN(net_372), .A1(net_371), .A2(net_339) );
NAND2_X1 inst_748 ( .ZN(net_676), .A1(n86gat), .A2(n392gat) );
NAND2_X1 inst_1146 ( .ZN(net_1059), .A1(net_1058), .A2(net_1057) );
NAND2_X1 inst_716 ( .ZN(net_480), .A2(n358gat), .A1(n205gat) );
NAND2_X1 inst_637 ( .ZN(net_0), .A1(n35gat), .A2(n273gat) );
NAND2_X1 inst_530 ( .ZN(net_270), .A1(n69gat), .A2(n324gat) );
NAND2_X1 inst_547 ( .ZN(net_549), .A2(n375gat), .A1(n18gat) );
NAND2_X1 inst_792 ( .ZN(net_249), .A1(net_248), .A2(net_215) );
NAND2_X1 inst_720 ( .ZN(net_909), .A2(n426gat), .A1(n171gat) );
NAND2_X1 inst_958 ( .ZN(net_633), .A2(net_593), .A1(net_527) );
NAND2_X1 inst_1217 ( .ZN(net_1235), .A1(net_1234), .A2(net_1202) );
NAND2_X1 inst_1353 ( .ZN(net_1554), .A1(net_1551), .A2(net_1537) );
XNOR2_X1 inst_368 ( .ZN(net_1381), .B(net_1372), .A(net_1338) );
NAND2_X1 inst_1010 ( .ZN(net_736), .A1(net_735), .A2(net_734) );
NAND2_X1 inst_803 ( .ZN(net_286), .A2(net_240), .A1(net_170) );
NAND2_X1 inst_769 ( .ZN(net_30), .A1(net_15), .A2(net_14) );
XNOR2_X1 inst_174 ( .ZN(net_682), .B(net_658), .A(net_657) );
XNOR2_X1 inst_274 ( .ZN(net_1039), .B(net_1023), .A(net_995) );
INV_X1 inst_1607 ( .ZN(net_1463), .A(net_1462) );
NAND2_X1 inst_1277 ( .ZN(net_1393), .A2(net_1342), .A1(net_1305) );
NAND2_X1 inst_1200 ( .ZN(net_1229), .A2(net_1156), .A1(net_1112) );
NAND2_X1 inst_662 ( .ZN(net_1183), .A2(n477gat), .A1(n222gat) );
NAND2_X1 inst_701 ( .ZN(net_1013), .A2(n443gat), .A1(n103gat) );
XNOR2_X1 inst_164 ( .ZN(net_660), .B(net_618), .A(net_617) );
NAND2_X1 inst_867 ( .ZN(net_397), .A1(net_396), .A2(net_382) );
INV_X1 inst_1533 ( .ZN(net_980), .A(net_979) );
NAND2_X1 inst_820 ( .ZN(net_290), .A1(net_289), .A2(net_284) );
NAND2_X1 inst_1199 ( .ZN(net_1184), .A1(net_1183), .A2(net_1150) );
XOR2_X1 inst_5 ( .Z(net_614), .A(net_584), .B(net_583) );
INV_X1 inst_1441 ( .ZN(net_333), .A(net_332) );
XNOR2_X1 inst_157 ( .ZN(net_620), .B(net_599), .A(net_598) );
NAND2_X1 inst_729 ( .ZN(net_1415), .A2(n511gat), .A1(n205gat) );
AND2_X4 inst_1662 ( .ZN(net_159), .A1(net_158), .A2(net_157) );
INV_X1 inst_1440 ( .ZN(net_331), .A(net_330) );
XNOR2_X1 inst_213 ( .ZN(net_851), .B(net_805), .A(net_776) );
XNOR2_X1 inst_68 ( .ZN(net_340), .A(net_289), .B(net_285) );
INV_X1 inst_1465 ( .ZN(net_491), .A(net_490) );
NAND2_X1 inst_604 ( .ZN(net_349), .A1(n52gat), .A2(n341gat) );
XNOR2_X1 inst_53 ( .A(net_242), .B(net_241), .ZN(n2223gat) );
NAND2_X1 inst_1253 ( .ZN(net_1308), .A1(net_1307), .A2(net_1306) );
NAND2_X1 inst_1007 ( .ZN(net_725), .A1(net_724), .A2(net_701) );
XNOR2_X1 inst_205 ( .ZN(net_817), .B(net_766), .A(net_732) );
NAND2_X1 inst_753 ( .ZN(net_1522), .A2(n528gat), .A1(n256gat) );
AND2_X4 inst_1645 ( .ZN(net_102), .A2(net_37), .A1(net_4) );
NAND2_X1 inst_1285 ( .ZN(net_1420), .A2(net_1371), .A1(net_1321) );
XNOR2_X1 inst_380 ( .ZN(net_1444), .B(net_1395), .A(net_1351) );
NAND2_X1 inst_1179 ( .ZN(net_1141), .A1(net_1140), .A2(net_1139) );
NAND2_X1 inst_946 ( .ZN(net_597), .A1(net_596), .A2(net_560) );
NAND2_X1 inst_651 ( .ZN(net_1155), .A2(n477gat), .A1(n18gat) );
XNOR2_X1 inst_292 ( .ZN(net_1113), .A(net_1076), .B(net_1028) );
NAND2_X1 inst_999 ( .ZN(net_716), .A1(net_715), .A2(net_714) );
AND2_X4 inst_1643 ( .ZN(net_38), .A2(net_37), .A1(net_5) );
INV_X1 inst_1591 ( .ZN(net_1354), .A(net_1353) );
NAND2_X1 inst_1157 ( .ZN(net_1111), .A2(net_1056), .A1(net_1006) );
INV_X1 inst_1515 ( .ZN(net_868), .A(net_867) );
XNOR2_X1 inst_379 ( .ZN(net_1439), .A(net_1393), .B(net_1382) );
NAND2_X1 inst_926 ( .ZN(net_547), .A1(net_546), .A2(net_545) );
INV_X1 inst_1463 ( .ZN(net_487), .A(net_486) );
XNOR2_X1 inst_186 ( .ZN(net_720), .A(net_703), .B(net_702) );
XNOR2_X1 inst_17 ( .ZN(net_154), .A(net_110), .B(net_69) );
NAND2_X1 inst_1325 ( .ZN(net_1479), .A1(net_1478), .A2(net_1465) );
NAND2_X1 inst_706 ( .ZN(net_1544), .A2(n528gat), .A1(n154gat) );
NAND2_X1 inst_759 ( .ZN(net_811), .A2(n409gat), .A1(n154gat) );
NAND2_X1 inst_1287 ( .ZN(net_1392), .A1(net_1391), .A2(net_1366) );
XNOR2_X1 inst_249 ( .ZN(net_965), .A(net_907), .B(net_885) );
NAND2_X1 inst_863 ( .ZN(net_413), .A2(net_372), .A1(net_315) );
NAND2_X1 inst_839 ( .ZN(net_353), .A1(net_352), .A2(net_351) );
NAND2_X1 inst_1015 ( .ZN(net_750), .A1(net_749), .A2(net_748) );
INV_X1 inst_1472 ( .ZN(net_564), .A(net_563) );
XNOR2_X1 inst_240 ( .ZN(net_937), .B(net_905), .A(net_873) );
AND2_X4 inst_1649 ( .ZN(net_100), .A2(net_44), .A1(net_26) );
NAND2_X1 inst_1385 ( .ZN(net_1613), .A1(net_1612), .A2(net_1611) );
NAND2_X1 inst_1169 ( .ZN(net_1119), .A1(net_1118), .A2(net_1094) );
XNOR2_X1 inst_110 ( .ZN(net_447), .B(net_419), .A(net_418) );
INV_X1 inst_1573 ( .ZN(net_1239), .A(net_1238) );
INV_X1 inst_1480 ( .ZN(net_621), .A(net_620) );
NAND2_X1 inst_891 ( .ZN(net_473), .A1(net_472), .A2(net_438) );
NAND2_X1 inst_1183 ( .ZN(net_1175), .A1(net_1122), .A2(net_1082) );
NAND2_X1 inst_1390 ( .ZN(net_1620), .A1(net_1619), .A2(net_1583) );
XNOR2_X1 inst_74 ( .ZN(net_345), .A(net_316), .B(net_273) );
NAND2_X1 inst_1235 ( .ZN(net_1267), .A1(net_1266), .A2(net_1257) );
XNOR2_X1 inst_288 ( .ZN(net_1091), .A(net_1058), .B(net_1057) );
XNOR2_X1 inst_229 ( .ZN(net_882), .B(net_865), .A(net_864) );
XNOR2_X1 inst_396 ( .ZN(net_1509), .B(net_1455), .A(net_1433) );
XNOR2_X1 inst_99 ( .ZN(net_454), .B(net_396), .A(net_381) );
INV_X1 inst_1489 ( .ZN(net_673), .A(net_672) );
AND2_X4 inst_1661 ( .ZN(net_156), .A1(net_155), .A2(net_154) );
NAND2_X1 inst_669 ( .ZN(net_367), .A2(n341gat), .A1(n154gat) );
NAND2_X1 inst_1298 ( .ZN(net_1422), .A1(net_1421), .A2(net_1420) );
NAND2_X1 inst_664 ( .ZN(net_246), .A2(n324gat), .A1(n188gat) );
NAND2_X1 inst_1394 ( .ZN(net_1627), .A2(net_1625), .A1(net_1574) );
NAND2_X1 inst_1160 ( .ZN(net_1125), .A2(net_1071), .A1(net_1017) );
XNOR2_X1 inst_283 ( .ZN(net_1074), .B(net_1055), .A(net_1034) );
XNOR2_X1 inst_311 ( .ZN(net_1181), .B(net_1152), .A(net_1151) );
NAND2_X1 inst_917 ( .ZN(net_512), .A1(net_511), .A2(net_510) );
INV_X1 inst_1597 ( .ZN(net_1388), .A(net_1387) );
XNOR2_X1 inst_372 ( .ZN(net_1414), .B(net_1376), .A(net_1299) );
INV_X1 inst_1600 ( .ZN(net_1424), .A(net_1423) );
NAND2_X1 inst_988 ( .ZN(net_695), .A1(net_694), .A2(net_671) );
XNOR2_X1 inst_215 ( .ZN(net_861), .B(net_811), .A(net_782) );
XNOR2_X1 inst_169 ( .ZN(net_672), .A(net_637), .B(net_636) );
INV_X1 inst_1418 ( .ZN(net_215), .A(net_214) );
XNOR2_X1 inst_421 ( .ZN(net_1569), .B(net_1544), .A(net_1543) );
NAND2_X1 inst_1315 ( .ZN(net_1494), .A2(net_1427), .A1(net_1384) );
NAND2_X1 inst_1092 ( .ZN(net_951), .A1(net_908), .A2(net_860) );
NAND2_X1 inst_555 ( .ZN(net_766), .A1(n69gat), .A2(n409gat) );
NAND2_X1 inst_849 ( .ZN(net_376), .A1(net_375), .A2(net_335) );
NAND2_X1 inst_816 ( .ZN(net_316), .A2(net_265), .A1(net_173) );
XNOR2_X1 inst_431 ( .ZN(net_1618), .B(net_1582), .A(net_1562) );
XOR2_X1 inst_3 ( .Z(net_427), .A(net_390), .B(net_389) );
XNOR2_X1 inst_348 ( .ZN(net_1309), .A(net_1273), .B(net_1272) );
NAND2_X1 inst_1172 ( .ZN(net_1147), .A2(net_1098), .A1(net_1043) );
NAND2_X1 inst_1184 ( .ZN(net_1177), .A2(net_1124), .A1(net_1065) );
NAND2_X1 inst_1090 ( .ZN(net_947), .A1(net_906), .A2(net_844) );
NAND2_X1 inst_889 ( .ZN(net_506), .A2(net_436), .A1(net_395) );
NAND2_X1 inst_577 ( .ZN(net_1372), .A2(n511gat), .A1(n18gat) );
AND2_X4 inst_1657 ( .ZN(net_144), .A1(net_143), .A2(net_142) );
NAND2_X1 inst_566 ( .ZN(net_140), .A1(n52gat), .A2(n307gat) );
NAND2_X1 inst_1399 ( .ZN(net_1634), .A1(net_1633), .A2(net_1632) );
NAND2_X1 inst_1239 ( .ZN(net_1274), .A1(net_1273), .A2(net_1272) );
NAND2_X1 inst_1364 ( .ZN(net_1572), .A1(net_1571), .A2(net_1518) );
XNOR2_X1 inst_36 ( .ZN(net_174), .A(net_140), .B(net_139) );
NAND2_X1 inst_656 ( .ZN(net_1123), .A2(n460gat), .A1(n103gat) );
NAND2_X1 inst_1370 ( .ZN(net_1589), .A1(net_1588), .A2(net_1581) );
NAND2_X1 inst_645 ( .ZN(net_458), .A1(n69gat), .A2(n358gat) );
XNOR2_X1 inst_45 ( .ZN(net_224), .B(net_175), .A(net_174) );
NOR2_X1 inst_503 ( .ZN(net_93), .A1(net_92), .A2(net_88) );
OR2_X4 inst_451 ( .ZN(net_118), .A2(net_87), .A1(net_59) );
NAND2_X1 inst_1108 ( .ZN(net_971), .A1(net_970), .A2(net_969) );
XNOR2_X1 inst_269 ( .ZN(net_1027), .B(net_1011), .A(net_985) );
NAND2_X1 inst_1190 ( .ZN(net_1161), .A1(net_1160), .A2(net_1134) );
OR2_X4 inst_458 ( .ZN(net_193), .A1(net_192), .A2(net_191) );
XNOR2_X1 inst_444 ( .A(net_1621), .B(net_1620), .ZN(n6250gat) );
INV_X1 inst_1562 ( .ZN(net_1163), .A(net_1162) );
INV_X1 inst_1495 ( .ZN(net_721), .A(net_720) );
NAND2_X1 inst_797 ( .ZN(net_259), .A1(net_258), .A2(net_233) );
NAND2_X1 inst_1097 ( .ZN(net_942), .A1(net_941), .A2(net_912) );
NAND2_X1 inst_686 ( .ZN(net_1324), .A2(n494gat), .A1(n188gat) );
NAND2_X1 inst_741 ( .ZN(net_897), .A2(n426gat), .A1(n256gat) );
NOR2_X1 inst_514 ( .ZN(net_181), .A2(net_132), .A1(net_109) );
INV_X1 inst_1541 ( .ZN(net_1028), .A(net_1027) );
NAND2_X1 inst_967 ( .ZN(net_635), .A1(net_634), .A2(net_633) );
NAND2_X1 inst_685 ( .ZN(net_923), .A2(n426gat), .A1(n154gat) );
NAND2_X1 inst_1350 ( .ZN(net_1545), .A1(net_1544), .A2(net_1543) );
XNOR2_X1 inst_63 ( .ZN(net_280), .A(net_266), .B(net_230) );
INV_X1 inst_1522 ( .ZN(net_891), .A(net_890) );
XNOR2_X1 inst_119 ( .ZN(net_531), .A(net_472), .B(net_437) );
NAND2_X1 inst_939 ( .ZN(net_607), .A1(net_558), .A2(net_509) );
INV_X1 inst_1543 ( .ZN(net_1035), .A(net_1034) );
NAND2_X1 inst_676 ( .ZN(net_1224), .A2(n477gat), .A1(n103gat) );
NAND2_X1 inst_1118 ( .ZN(net_1031), .A2(net_978), .A1(net_915) );
NAND2_X1 inst_1115 ( .ZN(net_1015), .A2(net_959), .A1(net_901) );
NAND2_X1 inst_1233 ( .ZN(net_1261), .A1(net_1260), .A2(net_1239) );
NAND2_X1 inst_1227 ( .ZN(net_1278), .A2(net_1225), .A1(net_1178) );
NAND2_X1 inst_874 ( .ZN(net_414), .A1(net_413), .A2(net_412) );
NAND2_X1 inst_1019 ( .ZN(net_788), .A2(net_725), .A1(net_686) );
NAND2_X1 inst_1021 ( .ZN(net_796), .A2(net_728), .A1(net_706) );
NAND2_X1 inst_1386 ( .ZN(net_1615), .A1(net_1613), .A2(net_1595) );
NOR2_X1 inst_473 ( .ZN(net_33), .A1(net_29), .A2(net_28) );
AND2_X4 inst_1652 ( .A2(net_65), .A1(net_41), .ZN(n1581gat) );
NAND2_X1 inst_1131 ( .ZN(net_1048), .A2(net_1000), .A1(net_938) );
NAND2_X1 inst_1076 ( .ZN(net_901), .A1(net_900), .A2(net_899) );
XNOR2_X1 inst_217 ( .ZN(net_827), .B(net_794), .A(net_793) );
INV_X1 inst_1622 ( .ZN(net_1561), .A(net_1560) );
NAND2_X1 inst_572 ( .ZN(net_662), .A1(n69gat), .A2(n392gat) );
NAND2_X1 inst_1357 ( .ZN(net_1573), .A2(net_1530), .A1(net_1495) );
NAND2_X1 inst_742 ( .ZN(net_1070), .A2(n460gat), .A1(n222gat) );
NAND2_X1 inst_691 ( .ZN(net_360), .A2(n341gat), .A1(n222gat) );
NAND2_X1 inst_1101 ( .ZN(net_949), .A1(net_948), .A2(net_947) );
XNOR2_X1 inst_427 ( .ZN(net_1626), .B(net_1571), .A(net_1517) );
XNOR2_X1 inst_257 ( .ZN(net_983), .A(net_948), .B(net_947) );
NOR2_X1 inst_485 ( .ZN(net_54), .A2(net_53), .A1(net_11) );
NAND2_X1 inst_770 ( .ZN(net_49), .A1(net_19), .A2(net_18) );
NAND2_X1 inst_565 ( .ZN(net_1558), .A2(n528gat), .A1(n103gat) );
NAND2_X1 inst_1195 ( .ZN(net_1173), .A1(net_1172), .A2(net_1171) );
NAND2_X1 inst_861 ( .ZN(net_416), .A2(net_366), .A1(net_303) );
NAND2_X1 inst_672 ( .ZN(net_250), .A1(n35gat), .A2(n324gat) );
INV_X1 inst_1471 ( .ZN(net_562), .A(net_561) );
XNOR2_X1 inst_138 ( .ZN(net_565), .B(net_523), .A(net_522) );
NAND2_X1 inst_622 ( .ZN(net_1007), .A2(n443gat), .A1(n171gat) );
INV_X1 inst_1404 ( .ZN(net_69), .A(net_68) );
NAND2_X1 inst_1205 ( .ZN(net_1209), .A1(net_1208), .A2(net_1180) );
NAND2_X1 inst_1189 ( .ZN(net_1159), .A1(net_1158), .A2(net_1157) );
NAND2_X1 inst_1283 ( .ZN(net_1384), .A2(net_1383), .A1(net_1350) );
XNOR2_X1 inst_409 ( .ZN(net_1536), .B(net_1510), .A(net_1509) );
NAND2_X1 inst_1269 ( .ZN(net_1356), .A1(net_1355), .A2(net_1344) );
INV_X1 inst_1525 ( .ZN(net_917), .A(net_916) );
NAND2_X1 inst_1339 ( .ZN(net_1514), .A1(net_1513), .A2(net_1512) );
NAND2_X1 inst_1202 ( .ZN(net_1193), .A1(net_1192), .A2(net_1163) );
NAND2_X1 inst_899 ( .ZN(net_494), .A1(net_493), .A2(net_492) );
NAND2_X1 inst_1312 ( .ZN(net_1456), .A1(net_1455), .A2(net_1434) );
INV_X1 inst_1540 ( .ZN(net_998), .A(net_997) );
XNOR2_X1 inst_33 ( .ZN(net_171), .A(net_158), .B(net_157) );
NAND2_X1 inst_703 ( .ZN(net_137), .A2(n307gat), .A1(n222gat) );
AND2_X4 inst_1660 ( .ZN(net_153), .A1(net_152), .A2(net_151) );
XNOR2_X1 inst_312 ( .ZN(net_1185), .B(net_1155), .A(net_1154) );
NAND2_X1 inst_660 ( .ZN(net_493), .A2(n358gat), .A1(n256gat) );
NAND2_X1 inst_977 ( .ZN(net_705), .A1(net_626), .A2(net_604) );
NOR2_X1 inst_517 ( .ZN(net_178), .A2(net_135), .A1(net_99) );
INV_X1 inst_1620 ( .ZN(net_1548), .A(net_1547) );
INV_X1 inst_1576 ( .ZN(net_1252), .A(net_1251) );
XNOR2_X1 inst_309 ( .ZN(net_1162), .B(net_1137), .A(net_1136) );
NAND2_X1 inst_1261 ( .ZN(net_1363), .A1(net_1298), .A2(net_1255) );
XNOR2_X1 inst_232 ( .ZN(net_888), .A(net_854), .B(net_821) );
XNOR2_X1 inst_347 ( .ZN(net_1313), .A(net_1270), .B(net_1195) );
NAND2_X1 inst_768 ( .ZN(net_46), .A1(net_7), .A2(net_6) );
NAND2_X1 inst_663 ( .ZN(net_584), .A2(n375gat), .A1(n256gat) );
XNOR2_X1 inst_297 ( .ZN(net_1139), .A(net_1089), .B(net_1075) );
NAND2_X1 inst_755 ( .ZN(net_1355), .A2(n494gat), .A1(n137gat) );
NAND2_X1 inst_1067 ( .ZN(net_870), .A1(net_869), .A2(net_836) );
NAND2_X1 inst_1395 ( .ZN(net_1628), .A1(net_1627), .A2(net_1626) );
XNOR2_X1 inst_310 ( .ZN(net_1179), .B(net_1147), .A(net_1146) );
NAND2_X1 inst_1214 ( .ZN(net_1228), .A1(net_1227), .A2(net_1226) );
NAND2_X1 inst_1043 ( .ZN(net_843), .A2(net_792), .A1(net_731) );
XNOR2_X1 inst_253 ( .ZN(net_962), .B(net_943), .A(net_916) );
NAND2_X1 inst_971 ( .ZN(net_651), .A1(net_650), .A2(net_649) );
INV_X1 inst_1417 ( .ZN(net_213), .A(net_212) );
NAND2_X1 inst_1219 ( .ZN(net_1262), .A2(net_1207), .A1(net_1161) );
XNOR2_X1 inst_162 ( .ZN(net_647), .B(net_615), .A(net_614) );
NAND2_X1 inst_589 ( .ZN(net_594), .A2(n375gat), .A1(n188gat) );
NAND2_X1 inst_794 ( .ZN(net_253), .A1(net_252), .A2(net_237) );
NAND2_X1 inst_1005 ( .ZN(net_755), .A1(net_713), .A2(net_644) );
NAND2_X1 inst_1330 ( .ZN(net_1497), .A1(net_1496), .A2(net_1463) );
NAND2_X1 inst_1147 ( .ZN(net_1062), .A1(net_1061), .A2(net_1060) );
INV_X1 inst_1580 ( .ZN(net_1290), .A(net_1289) );
NAND2_X1 inst_602 ( .ZN(net_134), .A2(n307gat), .A1(n120gat) );
XNOR2_X1 inst_59 ( .ZN(net_276), .B(net_256), .A(net_216) );
XNOR2_X1 inst_135 ( .ZN(net_559), .B(net_532), .A(net_531) );
INV_X1 inst_1408 ( .ZN(net_78), .A(net_77) );
NAND2_X1 inst_996 ( .ZN(net_712), .A2(net_711), .A1(net_681) );
XNOR2_X1 inst_37 ( .ZN(net_188), .B(net_137), .A(net_136) );
INV_X1 inst_1527 ( .ZN(net_935), .A(net_934) );
NAND2_X1 inst_1098 ( .ZN(net_944), .A1(net_943), .A2(net_917) );
AND2_X4 inst_1664 ( .ZN(net_165), .A1(net_164), .A2(net_163) );
NAND2_X1 inst_740 ( .ZN(net_390), .A2(n341gat), .A1(n256gat) );
INV_X1 inst_1447 ( .ZN(net_380), .A(net_379) );
XNOR2_X1 inst_264 ( .ZN(net_997), .A(net_973), .B(net_972) );
INV_X1 inst_1496 ( .ZN(net_723), .A(net_722) );
XNOR2_X1 inst_84 ( .ZN(net_421), .A(net_375), .B(net_334) );
INV_X1 inst_1565 ( .ZN(net_1186), .A(net_1185) );
NAND2_X1 inst_924 ( .ZN(net_533), .A1(net_532), .A2(net_531) );
NAND2_X1 inst_1333 ( .ZN(net_1503), .A1(net_1502), .A2(net_1490) );
XNOR2_X1 inst_303 ( .ZN(net_1149), .A(net_1126), .B(net_1125) );
XNOR2_X1 inst_173 ( .ZN(net_680), .B(net_655), .A(net_654) );
NAND2_X1 inst_723 ( .ZN(net_1219), .A2(n477gat), .A1(n188gat) );
XNOR2_X1 inst_224 ( .ZN(net_878), .B(net_849), .A(net_825) );
NAND2_X1 inst_611 ( .ZN(net_63), .A2(n290gat), .A1(n256gat) );
XNOR2_X1 inst_287 ( .ZN(net_1103), .A(net_1066), .B(net_980) );
XNOR2_X1 inst_426 ( .ZN(net_1586), .A(net_1558), .B(net_1541) );
NAND2_X1 inst_618 ( .ZN(net_1023), .A2(n443gat), .A1(n137gat) );
INV_X1 inst_1551 ( .ZN(net_1088), .A(net_1087) );
AND2_X4 inst_1647 ( .ZN(net_110), .A2(net_46), .A1(net_6) );
NAND2_X1 inst_648 ( .ZN(net_1460), .A2(n528gat), .A1(n239gat) );
NAND2_X1 inst_1260 ( .ZN(net_1361), .A1(net_1296), .A2(net_1261) );
NAND2_X1 inst_1275 ( .ZN(net_1371), .A1(net_1370), .A2(net_1369) );
NAND2_X1 inst_1088 ( .ZN(net_928), .A1(net_927), .A2(net_883) );
XNOR2_X1 inst_270 ( .ZN(net_1061), .A(net_1007), .B(net_987) );
NOR2_X1 inst_474 ( .ZN(net_32), .A2(net_31), .A1(net_17) );
XNOR2_X1 inst_26 ( .ZN(net_194), .A(net_152), .B(net_151) );
NAND2_X1 inst_766 ( .ZN(net_1510), .A1(n52gat), .A2(n528gat) );
NOR2_X1 inst_490 ( .ZN(net_106), .A2(net_51), .A1(net_24) );
NAND2_X1 inst_984 ( .ZN(net_688), .A1(net_687), .A2(net_661) );
NAND2_X1 inst_801 ( .ZN(net_267), .A1(net_266), .A2(net_231) );
NAND2_X1 inst_626 ( .ZN(net_650), .A1(n52gat), .A2(n392gat) );
NAND2_X1 inst_1376 ( .ZN(net_1599), .A2(net_1598), .A1(net_1554) );
NAND2_X1 inst_692 ( .ZN(net_737), .A2(n409gat), .A1(n222gat) );
INV_X1 inst_1517 ( .ZN(net_874), .A(net_873) );
NAND2_X1 inst_1292 ( .ZN(net_1403), .A1(net_1402), .A2(net_1401) );
XNOR2_X1 inst_70 ( .ZN(net_326), .B(net_304), .A(net_244) );
XNOR2_X1 inst_129 ( .ZN(net_545), .B(net_502), .A(net_484) );
NAND2_X1 inst_870 ( .ZN(net_403), .A1(net_402), .A2(net_380) );
NAND2_X1 inst_1309 ( .ZN(net_1448), .A1(net_1447), .A2(net_1423) );
INV_X1 inst_1531 ( .ZN(net_963), .A(net_962) );
XNOR2_X1 inst_11 ( .ZN(net_142), .A(net_120), .B(net_96) );
NAND2_X1 inst_631 ( .ZN(net_1234), .A2(n477gat), .A1(n154gat) );
NAND2_X1 inst_1056 ( .ZN(net_848), .A1(net_847), .A2(net_828) );
XNOR2_X1 inst_188 ( .ZN(net_734), .B(net_709), .A(net_678) );
INV_X1 inst_1619 ( .ZN(net_1541), .A(net_1540) );
XNOR2_X1 inst_441 ( .A(net_1612), .B(net_1611), .ZN(n6220gat) );
AND2_X4 inst_1659 ( .ZN(net_150), .A1(net_149), .A2(net_148) );
INV_X1 inst_1503 ( .ZN(net_775), .A(net_774) );
NAND2_X1 inst_798 ( .ZN(net_261), .A1(net_260), .A2(net_221) );
NAND2_X1 inst_808 ( .ZN(net_297), .A2(net_261), .A1(net_205) );
INV_X1 inst_1537 ( .ZN(net_992), .A(net_991) );
NAND2_X1 inst_557 ( .ZN(net_592), .A2(n375gat), .A1(n205gat) );
NAND2_X1 inst_777 ( .ZN(net_96), .A2(net_70), .A1(net_58) );
XNOR2_X1 inst_398 ( .ZN(net_1488), .B(net_1471), .A(net_1442) );
NAND2_X1 inst_1128 ( .ZN(net_1022), .A1(net_1021), .A2(net_992) );
XNOR2_X1 inst_436 ( .A(net_1597), .B(net_1596), .ZN(n6170gat) );
INV_X1 inst_1434 ( .ZN(net_279), .A(net_278) );
NAND2_X1 inst_1383 ( .ZN(net_1610), .A1(net_1609), .A2(net_1608) );
NAND2_X1 inst_1037 ( .ZN(net_808), .A1(net_807), .A2(net_779) );
INV_X1 inst_1461 ( .ZN(net_483), .A(net_482) );
NAND2_X1 inst_823 ( .ZN(net_298), .A1(net_297), .A2(net_276) );
NAND2_X1 inst_933 ( .ZN(net_603), .A1(net_540), .A2(net_507) );
XNOR2_X1 inst_300 ( .ZN(net_1188), .A(net_1118), .B(net_1093) );
NAND2_X1 inst_1250 ( .ZN(net_1332), .A1(net_1267), .A2(net_1228) );
XNOR2_X1 inst_102 ( .ZN(net_432), .B(net_392), .A(net_343) );
NAND2_X1 inst_1226 ( .ZN(net_1275), .A1(net_1222), .A2(net_1170) );
NAND2_X1 inst_1013 ( .ZN(net_744), .A1(net_743), .A2(net_742) );
XNOR2_X1 inst_446 ( .A(net_1627), .B(net_1626), .ZN(n6270gat) );
XNOR2_X1 inst_364 ( .ZN(net_1365), .A(net_1333), .B(net_1332) );
INV_X1 inst_1457 ( .ZN(net_444), .A(net_443) );
XNOR2_X1 inst_144 ( .ZN(net_577), .B(net_557), .A(net_556) );
XNOR2_X1 inst_195 ( .ZN(net_800), .B(net_762), .A(net_720) );
INV_X1 inst_1438 ( .ZN(net_327), .A(net_326) );
NAND2_X1 inst_824 ( .ZN(net_300), .A1(net_299), .A2(net_274) );
XNOR2_X1 inst_411 ( .ZN(net_1540), .A(net_1502), .B(net_1491) );
NAND2_X1 inst_1224 ( .ZN(net_1270), .A1(net_1217), .A2(net_1159) );
NAND2_X1 inst_1170 ( .ZN(net_1122), .A1(net_1121), .A2(net_1120) );
NAND2_X1 inst_1150 ( .ZN(net_1071), .A1(net_1070), .A2(net_1045) );
XNOR2_X1 inst_124 ( .ZN(net_510), .B(net_476), .A(net_447) );
NAND2_X1 inst_880 ( .ZN(net_436), .A1(net_435), .A2(net_434) );
INV_X1 inst_1413 ( .ZN(net_89), .A(net_88) );
NAND2_X1 inst_680 ( .ZN(net_1025), .A2(n443gat), .A1(n120gat) );
NAND2_X1 inst_785 ( .ZN(net_200), .A2(net_138), .A1(net_119) );
NAND2_X1 inst_737 ( .ZN(net_1114), .A2(n460gat), .A1(n188gat) );
NAND2_X1 inst_961 ( .ZN(net_613), .A1(net_612), .A2(net_611) );
NAND2_X1 inst_876 ( .ZN(net_420), .A1(net_419), .A2(net_418) );
INV_X1 inst_1590 ( .ZN(net_1352), .A(net_1351) );
NAND2_X1 inst_545 ( .ZN(net_266), .A1(n86gat), .A2(n324gat) );
INV_X1 inst_1589 ( .ZN(net_1350), .A(net_1349) );
NAND2_X1 inst_1270 ( .ZN(net_1383), .A1(net_1325), .A2(net_1274) );
XNOR2_X1 inst_399 ( .ZN(net_1490), .A(net_1447), .B(net_1424) );
NAND2_X1 inst_1388 ( .ZN(net_1617), .A1(net_1616), .A2(net_1593) );
NAND2_X1 inst_527 ( .ZN(net_625), .A2(n392gat), .A1(n1gat) );
NAND2_X1 inst_1326 ( .ZN(net_1521), .A2(net_1461), .A1(net_1422) );
XNOR2_X1 inst_226 ( .ZN(net_871), .B(net_840), .A(net_839) );
NAND2_X1 inst_1180 ( .ZN(net_1167), .A1(net_1115), .A2(net_1077) );
XNOR2_X1 inst_414 ( .ZN(net_1549), .B(net_1513), .A(net_1512) );
XNOR2_X1 inst_61 ( .ZN(net_278), .B(net_270), .A(net_212) );
XNOR2_X1 inst_203 ( .ZN(net_782), .B(net_755), .A(net_754) );
NAND2_X1 inst_531 ( .ZN(net_803), .A2(n409gat), .A1(n120gat) );
NAND2_X1 inst_562 ( .ZN(net_1121), .A2(n460gat), .A1(n120gat) );
XNOR2_X1 inst_212 ( .ZN(net_820), .B(net_807), .A(net_778) );
NAND2_X1 inst_1299 ( .ZN(net_1437), .A2(net_1390), .A1(net_1337) );
NAND2_X1 inst_1139 ( .ZN(net_1076), .A2(net_1022), .A1(net_966) );
NOR2_X1 inst_499 ( .A2(net_106), .ZN(net_85), .A1(net_52) );
INV_X1 inst_1519 ( .ZN(net_885), .A(net_884) );
NAND2_X1 inst_1372 ( .ZN(net_1596), .A2(net_1579), .A1(net_1546) );
XNOR2_X1 inst_335 ( .A(net_1232), .B(net_1231), .ZN(n5672gat) );
NAND2_X1 inst_1360 ( .ZN(net_1565), .A1(net_1564), .A2(net_1550) );
NAND2_X1 inst_674 ( .ZN(net_999), .A1(n86gat), .A2(n443gat) );
INV_X1 inst_1571 ( .ZN(net_1204), .A(net_1203) );
INV_X1 inst_1451 ( .ZN(net_388), .A(net_387) );
NOR2_X1 inst_466 ( .ZN(net_35), .A1(net_3), .A2(net_2) );
NAND2_X1 inst_658 ( .ZN(net_19), .A1(n69gat), .A2(n290gat) );
NAND2_X1 inst_989 ( .ZN(net_697), .A1(net_696), .A2(net_673) );
OR2_X4 inst_456 ( .ZN(net_185), .A1(net_184), .A2(net_183) );
NAND2_X1 inst_832 ( .ZN(net_320), .A1(net_319), .A2(net_318) );
INV_X1 inst_1491 ( .ZN(net_679), .A(net_678) );
INV_X1 inst_1402 ( .A(net_65), .ZN(net_62) );
XNOR2_X1 inst_275 ( .ZN(net_1064), .A(net_1025), .B(net_997) );
XNOR2_X1 inst_117 ( .ZN(net_495), .B(net_468), .A(net_430) );
NAND2_X1 inst_858 ( .ZN(net_398), .A2(net_347), .A1(net_317) );
XNOR2_X1 inst_438 ( .A(net_1603), .B(net_1602), .ZN(n6190gat) );
NAND2_X1 inst_1109 ( .ZN(net_974), .A1(net_973), .A2(net_972) );
NOR2_X1 inst_501 ( .A2(net_108), .ZN(net_68), .A1(net_34) );
NAND2_X1 inst_1341 ( .ZN(net_1538), .A2(net_1484), .A1(net_1438) );
NAND2_X1 inst_587 ( .ZN(net_869), .A1(n52gat), .A2(n426gat) );
NAND2_X1 inst_1081 ( .ZN(net_929), .A1(net_876), .A2(net_824) );
XNOR2_X1 inst_154 ( .ZN(net_640), .A(net_594), .B(net_569) );
NAND2_X1 inst_666 ( .ZN(net_1532), .A2(n528gat), .A1(n171gat) );
XNOR2_X1 inst_324 ( .ZN(net_1214), .A(net_1188), .B(net_1187) );
NOR2_X1 inst_465 ( .ZN(net_55), .A1(net_1), .A2(net_0) );
NAND2_X1 inst_1182 ( .ZN(net_1172), .A2(net_1119), .A1(net_1062) );
XNOR2_X1 inst_54 ( .ZN(net_244), .B(net_239), .A(net_238) );
XNOR2_X1 inst_109 ( .ZN(net_445), .A(net_425), .B(net_424) );
NAND2_X1 inst_570 ( .ZN(net_1445), .A2(n511gat), .A1(n154gat) );
INV_X1 inst_1570 ( .ZN(net_1202), .A(net_1201) );
NAND2_X1 inst_640 ( .ZN(net_586), .A2(n375gat), .A1(n154gat) );
INV_X1 inst_1482 ( .ZN(net_646), .A(net_645) );
INV_X1 inst_1420 ( .ZN(net_219), .A(net_218) );
NAND2_X1 inst_1314 ( .ZN(net_1461), .A1(net_1460), .A2(net_1459) );
XNOR2_X1 inst_43 ( .ZN(net_218), .B(net_181), .A(net_180) );
INV_X1 inst_1612 ( .ZN(net_1491), .A(net_1490) );
INV_X1 inst_1478 ( .ZN(net_580), .A(net_579) );
NAND2_X1 inst_1156 ( .ZN(net_1086), .A1(net_1085), .A2(net_1052) );
INV_X1 inst_1444 ( .ZN(net_339), .A(net_338) );
NAND2_X1 inst_1231 ( .ZN(net_1283), .A1(net_1235), .A2(net_1173) );
XNOR2_X1 inst_94 ( .ZN(net_412), .B(net_367), .A(net_336) );
NAND2_X1 inst_1114 ( .ZN(net_990), .A1(net_989), .A2(net_957) );
OR2_X4 inst_454 ( .ZN(net_179), .A1(net_178), .A2(net_177) );
XNOR2_X1 inst_375 ( .ZN(net_1407), .B(net_1391), .A(net_1365) );
NAND2_X1 inst_942 ( .ZN(net_589), .A1(net_588), .A2(net_564) );
NAND2_X1 inst_1295 ( .ZN(net_1413), .A1(net_1412), .A2(net_1411) );
NAND2_X1 inst_904 ( .ZN(net_532), .A2(net_479), .A1(net_417) );
XNOR2_X1 inst_262 ( .ZN(net_993), .A(net_967), .B(net_946) );
NAND2_X1 inst_1378 ( .ZN(net_1602), .A2(net_1601), .A1(net_1553) );
XNOR2_X1 inst_243 ( .ZN(net_948), .A(net_927), .B(net_882) );
XNOR2_X1 inst_285 ( .ZN(net_1157), .A(net_1070), .B(net_1044) );
XNOR2_X1 inst_424 ( .ZN(net_1580), .B(net_1556), .A(net_1555) );
NAND2_X1 inst_591 ( .ZN(net_943), .A2(n443gat), .A1(n18gat) );
NOR2_X1 inst_497 ( .A2(net_114), .ZN(net_75), .A1(net_50) );
XNOR2_X1 inst_15 ( .ZN(net_139), .A(net_106), .B(net_84) );
NAND2_X1 inst_757 ( .ZN(net_1245), .A2(n494gat), .A1(n18gat) );
INV_X1 inst_1627 ( .ZN(net_1587), .A(net_1586) );
XNOR2_X1 inst_343 ( .ZN(net_1294), .B(net_1260), .A(net_1238) );
NAND2_X1 inst_1035 ( .ZN(net_804), .A1(net_803), .A2(net_775) );
NAND2_X1 inst_1335 ( .ZN(net_1508), .A1(net_1507), .A2(net_1506) );
INV_X1 inst_1563 ( .ZN(net_1180), .A(net_1179) );
NAND2_X1 inst_1106 ( .ZN(net_966), .A1(net_965), .A2(net_964) );
XNOR2_X1 inst_337 ( .ZN(net_1287), .B(net_1247), .A(net_1214) );
NAND2_X1 inst_543 ( .ZN(net_1418), .A1(n86gat), .A2(n511gat) );
NAND2_X1 inst_929 ( .ZN(net_552), .A1(net_551), .A2(net_536) );
NAND2_X1 inst_982 ( .ZN(net_707), .A2(net_653), .A1(net_606) );
NAND2_X1 inst_1212 ( .ZN(net_1225), .A1(net_1224), .A2(net_1223) );
NAND2_X1 inst_1397 ( .ZN(net_1631), .A1(net_1630), .A2(net_1629) );
NAND2_X1 inst_1256 ( .ZN(net_1321), .A1(net_1320), .A2(net_1319) );
NAND2_X1 inst_1078 ( .ZN(net_906), .A1(net_905), .A2(net_874) );
NAND2_X1 inst_670 ( .ZN(net_875), .A1(n69gat), .A2(n426gat) );
XNOR2_X1 inst_299 ( .ZN(net_1171), .A(net_1116), .B(net_1091) );
INV_X1 inst_1423 ( .ZN(net_225), .A(net_224) );
NAND2_X1 inst_1034 ( .ZN(net_802), .A1(net_801), .A2(net_800) );
NOR2_X1 inst_476 ( .ZN(net_36), .A2(net_35), .A1(net_3) );
XNOR2_X1 inst_418 ( .ZN(net_1562), .B(net_1532), .A(net_1531) );
NAND2_X1 inst_864 ( .ZN(net_419), .A2(net_374), .A1(net_312) );
NAND2_X1 inst_1207 ( .ZN(net_1242), .A2(net_1184), .A1(net_1127) );
XNOR2_X1 inst_86 ( .ZN(net_404), .B(net_373), .A(net_328) );
NAND2_X1 inst_949 ( .ZN(net_600), .A1(net_599), .A2(net_598) );
XNOR2_X1 inst_20 ( .ZN(net_151), .A(net_114), .B(net_67) );
NAND2_X1 inst_1369 ( .ZN(net_1583), .A2(net_1582), .A1(net_1563) );
NAND2_X1 inst_613 ( .ZN(net_371), .A2(n341gat), .A1(n137gat) );
NAND2_X1 inst_1039 ( .ZN(net_812), .A1(net_811), .A2(net_783) );
NAND2_X1 inst_714 ( .ZN(net_466), .A1(n52gat), .A2(n358gat) );
XNOR2_X1 inst_349 ( .ZN(net_1316), .B(net_1275), .A(net_1249) );
INV_X1 inst_1428 ( .ZN(net_235), .A(net_234) );
NOR2_X1 inst_483 ( .ZN(net_94), .A2(net_39), .A1(net_20) );
NAND2_X1 inst_576 ( .ZN(net_358), .A1(n35gat), .A2(n341gat) );
XNOR2_X1 inst_259 ( .ZN(net_987), .A(net_954), .B(net_953) );
NAND2_X1 inst_1046 ( .ZN(net_865), .A2(net_804), .A1(net_744) );
XNOR2_X1 inst_246 ( .ZN(net_973), .A(net_925), .B(net_892) );
NAND2_X1 inst_1020 ( .ZN(net_763), .A1(net_762), .A2(net_721) );
NAND2_X1 inst_1061 ( .ZN(net_855), .A1(net_854), .A2(net_820) );
NAND2_X1 inst_635 ( .ZN(net_1118), .A2(n460gat), .A1(n154gat) );
NAND2_X1 inst_1177 ( .ZN(net_1160), .A2(net_1107), .A1(net_1050) );
NAND2_X1 inst_807 ( .ZN(net_302), .A2(net_255), .A1(net_211) );
NAND2_X1 inst_705 ( .ZN(net_242), .A2(n324gat), .A1(n1gat) );
NAND2_X1 inst_1244 ( .ZN(net_1285), .A1(net_1284), .A2(net_1283) );
XNOR2_X1 inst_72 ( .ZN(net_330), .B(net_302), .A(net_301) );
NAND2_X1 inst_911 ( .ZN(net_499), .A1(net_498), .A2(net_489) );
NAND2_X1 inst_976 ( .ZN(net_663), .A1(net_662), .A2(net_621) );
INV_X1 inst_1578 ( .ZN(net_1269), .A(net_1268) );
NOR2_X1 inst_519 ( .ZN(net_210), .A2(net_156), .A1(net_111) );
NAND2_X1 inst_1279 ( .ZN(net_1397), .A2(net_1348), .A1(net_1288) );
AND2_X2 inst_1666 ( .A1(net_1634), .A2(net_1523), .ZN(n6287gat) );
AND2_X4 inst_1634 ( .ZN(net_1), .A2(n290gat), .A1(n18gat) );
NAND2_X1 inst_909 ( .ZN(net_528), .A2(net_473), .A1(net_423) );
NAND2_X1 inst_1003 ( .ZN(net_745), .A1(net_697), .A2(net_638) );
NAND2_X1 inst_582 ( .ZN(net_461), .A2(n358gat), .A1(n18gat) );
NAND2_X1 inst_1096 ( .ZN(net_938), .A1(net_937), .A2(net_936) );
NAND2_X1 inst_683 ( .ZN(net_837), .A2(n426gat), .A1(n239gat) );
NAND2_X1 inst_735 ( .ZN(net_696), .A2(n392gat), .A1(n188gat) );
INV_X1 inst_1529 ( .ZN(net_946), .A(net_945) );
NAND2_X1 inst_1053 ( .ZN(net_838), .A1(net_837), .A2(net_816) );
XNOR2_X1 inst_115 ( .ZN(net_486), .B(net_466), .A(net_465) );
AND2_X4 inst_1653 ( .ZN(net_129), .A1(net_128), .A2(net_127) );
XNOR2_X1 inst_210 ( .ZN(net_864), .A(net_813), .B(net_772) );
NAND2_X1 inst_894 ( .ZN(net_479), .A1(net_478), .A2(net_440) );
NAND2_X1 inst_994 ( .ZN(net_708), .A2(net_707), .A1(net_648) );
NAND2_X1 inst_761 ( .ZN(net_1426), .A2(n511gat), .A1(n188gat) );
XNOR2_X1 inst_239 ( .ZN(net_916), .A(net_878), .B(net_877) );
INV_X1 inst_1582 ( .ZN(net_1310), .A(net_1309) );
NAND2_X1 inst_1294 ( .ZN(net_1410), .A1(net_1409), .A2(net_1407) );
NAND2_X1 inst_1193 ( .ZN(net_1168), .A2(net_1167), .A1(net_1133) );
INV_X1 inst_1625 ( .ZN(net_1581), .A(net_1580) );
INV_X1 inst_1432 ( .ZN(net_275), .A(net_274) );
XNOR2_X1 inst_175 ( .ZN(net_749), .A(net_652), .B(net_623) );
NAND2_X1 inst_593 ( .ZN(net_1140), .A2(n477gat), .A1(n1gat) );
NAND2_X1 inst_725 ( .ZN(net_762), .A1(n52gat), .A2(n409gat) );
NAND2_X1 inst_747 ( .ZN(net_1208), .A1(n69gat), .A2(n477gat) );
NAND2_X1 inst_843 ( .ZN(net_364), .A1(net_363), .A2(net_362) );
NAND2_X1 inst_601 ( .ZN(net_20), .A1(n52gat), .A2(n273gat) );
NAND2_X1 inst_1337 ( .ZN(net_1524), .A2(net_1472), .A1(net_1413) );
XNOR2_X1 inst_133 ( .ZN(net_541), .B(net_511), .A(net_510) );
NAND2_X1 inst_1263 ( .ZN(net_1337), .A1(net_1336), .A2(net_1335) );
XNOR2_X1 inst_112 ( .A(net_435), .B(net_434), .ZN(n2877gat) );
NAND2_X1 inst_916 ( .ZN(net_509), .A1(net_508), .A2(net_487) );
NAND2_X1 inst_764 ( .ZN(net_463), .A2(n358gat), .A1(n222gat) );
AND2_X4 inst_1638 ( .ZN(net_22), .A2(n273gat), .A1(n256gat) );
NOR2_X1 inst_479 ( .ZN(net_61), .A2(net_42), .A1(net_12) );
XNOR2_X1 inst_305 ( .ZN(net_1174), .A(net_1130), .B(net_1101) );
INV_X1 inst_1595 ( .ZN(net_1375), .A(net_1374) );
INV_X1 inst_1547 ( .ZN(net_1052), .A(net_1051) );
NAND2_X1 inst_1111 ( .ZN(net_978), .A1(net_977), .A2(net_940) );
XNOR2_X1 inst_29 ( .ZN(net_183), .B(net_164), .A(net_163) );
INV_X1 inst_1583 ( .ZN(net_1312), .A(net_1311) );
NAND2_X1 inst_1149 ( .ZN(net_1067), .A2(net_1066), .A1(net_979) );
NAND2_X1 inst_771 ( .ZN(net_48), .A1(net_23), .A2(net_22) );
INV_X1 inst_1445 ( .ZN(net_344), .A(net_343) );
NAND2_X1 inst_1281 ( .ZN(net_1380), .A1(net_1379), .A2(net_1378) );
INV_X1 inst_1509 ( .ZN(net_816), .A(net_815) );
NAND2_X1 inst_878 ( .ZN(net_426), .A1(net_425), .A2(net_424) );
NAND2_X1 inst_1274 ( .ZN(net_1364), .A2(net_1363), .A1(net_1331) );
XNOR2_X1 inst_126 ( .ZN(net_538), .B(net_506), .A(net_482) );
NOR2_X1 inst_480 ( .ZN(net_114), .A2(net_43), .A1(net_8) );
INV_X1 inst_1512 ( .ZN(net_828), .A(net_827) );
AND2_X4 inst_1631 ( .ZN(net_3), .A2(n290gat), .A1(n205gat) );
NAND2_X1 inst_538 ( .ZN(net_847), .A2(n426gat), .A1(n222gat) );
NAND2_X1 inst_564 ( .ZN(net_1320), .A2(n494gat), .A1(n256gat) );
NAND2_X1 inst_646 ( .ZN(net_5), .A2(n290gat), .A1(n137gat) );
NAND2_X1 inst_1319 ( .ZN(net_1470), .A1(net_1469), .A2(net_1468) );
NAND2_X1 inst_1300 ( .ZN(net_1457), .A2(net_1392), .A1(net_1334) );
NAND2_X1 inst_963 ( .ZN(net_619), .A1(net_618), .A2(net_617) );
NAND2_X1 inst_1140 ( .ZN(net_1078), .A1(net_1024), .A2(net_971) );
XNOR2_X1 inst_382 ( .ZN(net_1433), .B(net_1402), .A(net_1401) );
XNOR2_X1 inst_35 ( .ZN(net_206), .B(net_149), .A(net_148) );
NAND2_X1 inst_739 ( .ZN(net_164), .A1(n86gat), .A2(n307gat) );
NAND2_X1 inst_948 ( .ZN(net_618), .A1(net_574), .A2(net_512) );
NAND2_X1 inst_1086 ( .ZN(net_924), .A1(net_923), .A2(net_891) );
XNOR2_X1 inst_358 ( .ZN(net_1349), .B(net_1314), .A(net_1313) );
XNOR2_X1 inst_48 ( .ZN(net_230), .B(net_198), .A(net_197) );
NAND2_X1 inst_907 ( .ZN(net_525), .A2(net_481), .A1(net_426) );
XNOR2_X1 inst_46 ( .ZN(net_226), .B(net_172), .A(net_171) );
NAND2_X1 inst_934 ( .ZN(net_574), .A1(net_573), .A2(net_542) );
NAND2_X1 inst_922 ( .ZN(net_527), .A1(net_526), .A2(net_525) );
INV_X1 inst_1614 ( .ZN(net_1505), .A(net_1504) );
NAND2_X1 inst_1000 ( .ZN(net_758), .A1(net_698), .A2(net_629) );
NAND2_X1 inst_1126 ( .ZN(net_1017), .A1(net_1016), .A2(net_1015) );
INV_X1 inst_1502 ( .ZN(net_773), .A(net_772) );
XNOR2_X1 inst_443 ( .A(net_1618), .B(net_1617), .ZN(n6240gat) );
NAND2_X1 inst_796 ( .ZN(net_257), .A1(net_256), .A2(net_217) );
NAND2_X1 inst_633 ( .ZN(net_365), .A2(n341gat), .A1(n171gat) );
NOR2_X1 inst_524 ( .ZN(net_192), .A2(net_153), .A1(net_115) );
NAND2_X1 inst_655 ( .ZN(net_268), .A1(n52gat), .A2(n324gat) );
XNOR2_X1 inst_104 ( .ZN(net_460), .B(net_398), .A(net_387) );
XNOR2_X1 inst_448 ( .B(net_1633), .A(net_1632), .ZN(n6288gat) );
NAND2_X1 inst_1049 ( .ZN(net_852), .A2(net_808), .A1(net_747) );
XNOR2_X1 inst_168 ( .ZN(net_670), .A(net_634), .B(net_633) );
INV_X1 inst_1568 ( .ZN(net_1197), .A(net_1196) );
INV_X1 inst_1499 ( .ZN(net_765), .A(net_764) );
NAND2_X1 inst_914 ( .ZN(net_505), .A1(net_504), .A2(net_491) );
NAND2_X1 inst_695 ( .ZN(net_1236), .A2(n477gat), .A1(n120gat) );
NAND2_X1 inst_730 ( .ZN(net_1507), .A1(n69gat), .A2(n528gat) );
AND2_X4 inst_1642 ( .ZN(net_29), .A2(n290gat), .A1(n188gat) );
XNOR2_X1 inst_384 ( .ZN(net_1442), .A(net_1412), .B(net_1411) );
NAND2_X1 inst_727 ( .ZN(net_428), .A2(n358gat), .A1(n239gat) );
NAND2_X1 inst_873 ( .ZN(net_411), .A1(net_410), .A2(net_409) );
NAND2_X1 inst_1252 ( .ZN(net_1305), .A2(net_1304), .A1(net_1269) );
XNOR2_X1 inst_321 ( .ZN(net_1223), .B(net_1177), .A(net_1144) );
NAND2_X1 inst_653 ( .ZN(net_161), .A2(n307gat), .A1(n103gat) );
NAND2_X1 inst_991 ( .ZN(net_717), .A1(net_677), .A2(net_613) );
NAND2_X1 inst_1343 ( .ZN(net_1564), .A2(net_1508), .A1(net_1467) );
NAND2_X1 inst_608 ( .ZN(net_27), .A1(n86gat), .A2(n290gat) );
NAND2_X1 inst_834 ( .ZN(net_325), .A1(net_324), .A2(net_323) );
NAND2_X1 inst_882 ( .ZN(net_456), .A1(net_455), .A2(net_454) );
XNOR2_X1 inst_170 ( .ZN(net_674), .A(net_640), .B(net_639) );
NAND2_X1 inst_580 ( .ZN(net_1152), .A2(n477gat), .A1(n239gat) );
NAND2_X1 inst_966 ( .ZN(net_632), .A1(net_631), .A2(net_630) );
NAND2_X1 inst_1246 ( .ZN(net_1293), .A1(net_1292), .A2(net_1291) );
NOR2_X1 inst_511 ( .ZN(net_111), .A1(net_110), .A2(net_68) );
XNOR2_X1 inst_41 ( .ZN(net_214), .B(net_195), .A(net_194) );
XNOR2_X1 inst_199 ( .ZN(net_774), .A(net_743), .B(net_742) );
NAND2_X1 inst_1164 ( .ZN(net_1110), .A1(net_1109), .A2(net_1108) );
NAND2_X1 inst_1346 ( .ZN(net_1530), .A1(net_1529), .A2(net_1528) );
NAND2_X1 inst_708 ( .ZN(net_125), .A2(n307gat), .A1(n239gat) );
NAND2_X1 inst_1374 ( .ZN(net_1595), .A2(net_1594), .A1(net_1585) );
XNOR2_X1 inst_152 ( .ZN(net_617), .B(net_590), .A(net_565) );
NAND2_X1 inst_1238 ( .ZN(net_1271), .A1(net_1270), .A2(net_1194) );
NAND2_X1 inst_953 ( .ZN(net_608), .A1(net_607), .A2(net_582) );
NAND2_X1 inst_1071 ( .ZN(net_913), .A1(net_870), .A2(net_819) );
NAND2_X1 inst_1163 ( .ZN(net_1107), .A1(net_1106), .A2(net_1084) );
INV_X1 inst_1421 ( .ZN(net_221), .A(net_220) );
NAND2_X1 inst_1099 ( .ZN(net_981), .A2(net_920), .A1(net_881) );
NOR2_X1 inst_468 ( .ZN(net_53), .A1(net_11), .A2(net_10) );
NAND2_X1 inst_1152 ( .ZN(net_1077), .A2(net_1076), .A1(net_1027) );
NAND2_X1 inst_1242 ( .ZN(net_1280), .A1(net_1262), .A2(net_1252) );
INV_X1 inst_1604 ( .ZN(net_1450), .A(net_1449) );
INV_X1 inst_1400 ( .ZN(net_87), .A(net_60) );
NAND2_X1 inst_1011 ( .ZN(net_738), .A1(net_737), .A2(net_722) );
XNOR2_X1 inst_429 ( .ZN(net_1623), .A(net_1573), .B(net_1548) );
NAND2_X1 inst_540 ( .ZN(net_1567), .A2(n528gat), .A1(n137gat) );
XNOR2_X1 inst_404 ( .ZN(net_1531), .B(net_1496), .A(net_1462) );
INV_X1 inst_1599 ( .ZN(net_1408), .A(net_1407) );
NAND2_X1 inst_998 ( .ZN(net_729), .A1(net_688), .A2(net_619) );
XNOR2_X1 inst_89 ( .ZN(net_409), .B(net_365), .A(net_330) );
INV_X1 inst_1520 ( .ZN(net_887), .A(net_886) );
XNOR2_X1 inst_388 ( .ZN(net_1468), .A(net_1409), .B(net_1408) );
XNOR2_X1 inst_66 ( .ZN(net_310), .A(net_248), .B(net_214) );
INV_X1 inst_1535 ( .ZN(net_986), .A(net_985) );
XOR2_X1 inst_7 ( .Z(net_1369), .A(net_1320), .B(net_1319) );
XNOR2_X1 inst_392 ( .ZN(net_1485), .B(net_1457), .A(net_1435) );
XNOR2_X1 inst_182 ( .ZN(net_746), .A(net_694), .B(net_670) );
XNOR2_X1 inst_273 ( .ZN(net_1058), .B(net_1021), .A(net_991) );
XNOR2_X1 inst_120 ( .ZN(net_519), .A(net_478), .B(net_439) );
XNOR2_X1 inst_294 ( .ZN(net_1120), .A(net_1081), .B(net_1040) );
NAND2_X1 inst_788 ( .ZN(net_202), .A1(net_201), .A2(net_200) );
NOR2_X1 inst_489 ( .ZN(net_90), .A2(net_55), .A1(net_0) );
NAND2_X1 inst_931 ( .ZN(net_558), .A1(net_557), .A2(net_556) );
XNOR2_X1 inst_192 ( .A(net_727), .B(net_726), .ZN(n3895gat) );
INV_X1 inst_1514 ( .ZN(net_846), .A(net_845) );
XNOR2_X1 inst_366 ( .A(net_1341), .B(net_1340), .ZN(n5971gat) );
INV_X1 inst_1579 ( .ZN(net_1282), .A(net_1281) );
NAND2_X1 inst_1083 ( .ZN(net_915), .A1(net_914), .A2(net_913) );
INV_X1 inst_1608 ( .ZN(net_1465), .A(net_1464) );
NAND2_X1 inst_567 ( .ZN(net_1106), .A1(n86gat), .A2(n460gat) );
INV_X1 inst_1411 ( .ZN(net_84), .A(net_83) );
XNOR2_X1 inst_149 ( .ZN(net_642), .A(net_596), .B(net_559) );
XNOR2_X1 inst_193 ( .ZN(net_760), .A(net_718), .B(net_717) );
XNOR2_X1 inst_318 ( .ZN(net_1199), .B(net_1169), .A(net_1142) );
NAND2_X1 inst_810 ( .ZN(net_304), .A2(net_253), .A1(net_202) );
NAND2_X1 inst_1136 ( .ZN(net_1060), .A2(net_1010), .A1(net_968) );
XNOR2_X1 inst_39 ( .ZN(net_241), .B(net_186), .A(net_166) );
XNOR2_X1 inst_230 ( .ZN(net_884), .A(net_859), .B(net_787) );
INV_X1 inst_1601 ( .ZN(net_1434), .A(net_1433) );
INV_X1 inst_1484 ( .ZN(net_661), .A(net_660) );
INV_X1 inst_1415 ( .ZN(net_117), .A(net_116) );
NAND2_X1 inst_856 ( .ZN(net_392), .A2(net_361), .A1(net_305) );
INV_X1 inst_1486 ( .ZN(net_667), .A(net_666) );

endmodule
