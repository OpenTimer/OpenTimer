module aes_core (
x7198,
x3951,
x3290,
x1373,
x3332,
x5505,
x5409,
x5926,
x2945,
x2197,
x6246,
x3376,
x2835,
x2978,
x3346,
x4481,
x2103,
x2531,
x1413,
x2077,
x5244,
x4496,
x1701,
x3791,
x5825,
x4285,
x1580,
x4384,
x2481,
x2382,
x2344,
x6655,
x2547,
x6631,
x3279,
x1731,
x2035,
x7607,
x1497,
x4215,
x4706,
x5188,
x2618,
x1808,
x7296,
x7443,
x1963,
x1932,
x5328,
x1362,
x6680,
x3463,
x1674,
x2260,
x2401,
x6089,
x6544,
x6043,
x3820,
x1781,
x6571,
x6145,
x2554,
x2087,
x2139,
x3416,
x2745,
x3608,
x6870,
x2367,
x6710,
x6521,
x5873,
x3021,
x7497,
x6797,
x7698,
x2855,
x7558,
x4848,
x1639,
x3058,
x2160,
x1526,
x2971,
x2881,
x3178,
x3052,
x2659,
x339831,
x7467,
x4345,
x6404,
x4781,
x4980,
x3771,
x2333,
x6071,
x1457,
x7235,
x1845,
x3989,
x2230,
x7042,
x4261,
x1354,
x3106,
x3220,
x5669,
x3268,
x1765,
x3491,
x6461,
x4668,
x3311,
x1446,
x1401,
x4815,
x2508,
x2468,
x6280,
x4099,
x3199,
x2357,
x4139,
x2280,
x4545,
x2784,
x5053,
x5464,
x1869,
x3863,
x4172,
x6832,
x2802,
x6494,
x6764,
x1471,
x4416,
x7135,
x2767,
x1651,
x2249,
x5637,
x5099,
x6966,
x6300,
x7268,
x6012,
x7413,
x2149,
x2957,
x3322,
x6600,
x4734,
x3117,
x4642,
x4319,
x6430,
x2042,
x3732,
x5568,
x6320,
x2420,
x1662,
x4041,
x2219,
x2650,
x3635,
x3163,
x3007,
x2571,
x5903,
x2115,
x2666,
x6110,
x3136,
x2985,
x3910,
x1747,
x3354,
x2457,
x1483,
x5145,
x1623,
x3339,
x2027,
x6585,
x5360,
x4916,
x1718,
x3001,
x5957,
x4603,
x3147,
x6740,
x2914,
x6912,
x6936,
x1948,
x6381,
x6697,
x5754,
x2011,
x1551,
x4444,
x1510,
x2428,
x2240,
x3701,
x3242,
x7527,
x2713,
x3667,
x1425,
x5723,
x2272,
x1987,
x3090,
x5537,
x2127,
x1912,
x1878,
x3153,
x6178,
x5290,
x7336,
x2174,
x2809,
x2688,
x5992,
x5853,
x5685,
x2639,
x6203,
x2298,
x3014,
x1891,
x7366,
x3553,
x7584,
x7088,
x5787,
x6224,
x2019,
x3079,
x4888,
x7000,
x6350,
x1975,
x3209,
x7642,
x1603,
x5605,
x5015,
x1686,
x2186,
x3521,
x7654,
x7158,
x643,
x492,
x346,
x140,
x1159,
x804,
x556,
x1283,
x1299,
x315,
x473,
x329,
x815,
x1247,
x1087,
x936,
x1032,
x912,
x55,
x532,
x733,
x1215,
x277,
x8,
x659,
x1134,
x876,
x71,
x161,
x256,
x957,
x90,
x1275,
x697,
x184,
x779,
x503,
x246,
x452,
x132,
x122,
x585,
x151,
x1330,
x424,
x598,
x1204,
x887,
x23,
x222,
x797,
x610,
x233,
x311,
x1259,
x839,
x0,
x107,
x629,
x1306,
x323,
x368,
x771,
x392,
x675,
x353,
x511,
x763,
x570,
x546,
x683,
x462,
x266,
x603,
x445,
x1192,
x1322,
x480,
x215,
x288,
x615,
x899,
x866,
x790,
x1121,
x648,
x745,
x990,
x33,
x636,
x622,
x756,
x1103,
x975,
x1291,
x205,
x1005,
x848,
x1044,
x361,
x173,
x668,
x719,
x522,
x304,
x592,
x339,
x687,
x1068,
x563,
x708,
x1021,
x1176,
x402,
x1314,
x16,
x923,
x539,
x1238,
x833,
x413,
x1146,
x844,
x577,
x856,
x726,
x296,
x826,
x1227);

// Start PIs
input x7198;
input x3951;
input x3290;
input x1373;
input x3332;
input x5505;
input x5409;
input x5926;
input x2945;
input x2197;
input x6246;
input x3376;
input x2835;
input x2978;
input x3346;
input x4481;
input x2103;
input x2531;
input x1413;
input x2077;
input x5244;
input x4496;
input x1701;
input x3791;
input x5825;
input x4285;
input x1580;
input x4384;
input x2481;
input x2382;
input x2344;
input x6655;
input x2547;
input x6631;
input x3279;
input x1731;
input x2035;
input x7607;
input x1497;
input x4215;
input x4706;
input x5188;
input x2618;
input x1808;
input x7296;
input x7443;
input x1963;
input x1932;
input x5328;
input x1362;
input x6680;
input x3463;
input x1674;
input x2260;
input x2401;
input x6089;
input x6544;
input x6043;
input x3820;
input x1781;
input x6571;
input x6145;
input x2554;
input x2087;
input x2139;
input x3416;
input x2745;
input x3608;
input x6870;
input x2367;
input x6710;
input x6521;
input x5873;
input x3021;
input x7497;
input x6797;
input x7698;
input x2855;
input x7558;
input x4848;
input x1639;
input x3058;
input x2160;
input x1526;
input x2971;
input x2881;
input x3178;
input x3052;
input x2659;
input x339831;
input x7467;
input x4345;
input x6404;
input x4781;
input x4980;
input x3771;
input x2333;
input x6071;
input x1457;
input x7235;
input x1845;
input x3989;
input x2230;
input x7042;
input x4261;
input x1354;
input x3106;
input x3220;
input x5669;
input x3268;
input x1765;
input x3491;
input x6461;
input x4668;
input x3311;
input x1446;
input x1401;
input x4815;
input x2508;
input x2468;
input x6280;
input x4099;
input x3199;
input x2357;
input x4139;
input x2280;
input x4545;
input x2784;
input x5053;
input x5464;
input x1869;
input x3863;
input x4172;
input x6832;
input x2802;
input x6494;
input x6764;
input x1471;
input x4416;
input x7135;
input x2767;
input x1651;
input x2249;
input x5637;
input x5099;
input x6966;
input x6300;
input x7268;
input x6012;
input x7413;
input x2149;
input x2957;
input x3322;
input x6600;
input x4734;
input x3117;
input x4642;
input x4319;
input x6430;
input x2042;
input x3732;
input x5568;
input x6320;
input x2420;
input x1662;
input x4041;
input x2219;
input x2650;
input x3635;
input x3163;
input x3007;
input x2571;
input x5903;
input x2115;
input x2666;
input x6110;
input x3136;
input x2985;
input x3910;
input x1747;
input x3354;
input x2457;
input x1483;
input x5145;
input x1623;
input x3339;
input x2027;
input x6585;
input x5360;
input x4916;
input x1718;
input x3001;
input x5957;
input x4603;
input x3147;
input x6740;
input x2914;
input x6912;
input x6936;
input x1948;
input x6381;
input x6697;
input x5754;
input x2011;
input x1551;
input x4444;
input x1510;
input x2428;
input x2240;
input x3701;
input x3242;
input x7527;
input x2713;
input x3667;
input x1425;
input x5723;
input x2272;
input x1987;
input x3090;
input x5537;
input x2127;
input x1912;
input x1878;
input x3153;
input x6178;
input x5290;
input x7336;
input x2174;
input x2809;
input x2688;
input x5992;
input x5853;
input x5685;
input x2639;
input x6203;
input x2298;
input x3014;
input x1891;
input x7366;
input x3553;
input x7584;
input x7088;
input x5787;
input x6224;
input x2019;
input x3079;
input x4888;
input x7000;
input x6350;
input x1975;
input x3209;
input x7642;
input x1603;
input x5605;
input x5015;
input x1686;
input x2186;
input x3521;
input x7654;
input x7158;

// Start POs
output x643;
output x492;
output x346;
output x140;
output x1159;
output x804;
output x556;
output x1283;
output x1299;
output x315;
output x473;
output x329;
output x815;
output x1247;
output x1087;
output x936;
output x1032;
output x912;
output x55;
output x532;
output x733;
output x1215;
output x277;
output x8;
output x659;
output x1134;
output x876;
output x71;
output x161;
output x256;
output x957;
output x90;
output x1275;
output x697;
output x184;
output x779;
output x503;
output x246;
output x452;
output x132;
output x122;
output x585;
output x151;
output x1330;
output x424;
output x598;
output x1204;
output x887;
output x23;
output x222;
output x797;
output x610;
output x233;
output x311;
output x1259;
output x839;
output x0;
output x107;
output x629;
output x1306;
output x323;
output x368;
output x771;
output x392;
output x675;
output x353;
output x511;
output x763;
output x570;
output x546;
output x683;
output x462;
output x266;
output x603;
output x445;
output x1192;
output x1322;
output x480;
output x215;
output x288;
output x615;
output x899;
output x866;
output x790;
output x1121;
output x648;
output x745;
output x990;
output x33;
output x636;
output x622;
output x756;
output x1103;
output x975;
output x1291;
output x205;
output x1005;
output x848;
output x1044;
output x361;
output x173;
output x668;
output x719;
output x522;
output x304;
output x592;
output x339;
output x687;
output x1068;
output x563;
output x708;
output x1021;
output x1176;
output x402;
output x1314;
output x16;
output x923;
output x539;
output x1238;
output x833;
output x413;
output x1146;
output x844;
output x577;
output x856;
output x726;
output x296;
output x826;
output x1227;

// Start wires
wire net_15987;
wire net_19401;
wire net_8631;
wire net_4065;
wire x3332;
wire x492;
wire net_11968;
wire net_4854;
wire net_2418;
wire net_16075;
wire net_7279;
wire net_11788;
wire net_4598;
wire net_21710;
wire net_12833;
wire net_1897;
wire net_980;
wire net_5499;
wire net_53;
wire net_9803;
wire net_12029;
wire net_7081;
wire net_10629;
wire net_11370;
wire net_5515;
wire net_3996;
wire net_22259;
wire net_18920;
wire net_17083;
wire net_15044;
wire net_6241;
wire net_7298;
wire net_4382;
wire net_13988;
wire net_13226;
wire net_12501;
wire net_21509;
wire net_8105;
wire net_4306;
wire net_21875;
wire net_264;
wire net_12959;
wire net_11178;
wire net_18857;
wire net_3904;
wire net_17256;
wire net_8914;
wire net_20731;
wire net_17057;
wire net_21295;
wire net_11757;
wire net_9072;
wire net_2769;
wire net_22546;
wire net_3707;
wire net_14405;
wire net_2082;
wire net_5035;
wire net_22713;
wire net_20115;
wire net_22580;
wire net_22232;
wire net_4832;
wire net_4464;
wire net_8577;
wire net_22602;
wire net_16142;
wire net_17675;
wire net_15913;
wire net_18014;
wire net_21560;
wire net_703;
wire net_22200;
wire net_5330;
wire net_193;
wire net_11377;
wire net_9989;
wire net_12447;
wire net_14381;
wire net_6773;
wire net_5273;
wire net_12413;
wire net_16843;
wire net_2942;
wire net_22364;
wire net_18119;
wire net_13993;
wire net_19378;
wire net_18314;
wire net_22812;
wire net_17574;
wire net_13916;
wire net_4442;
wire net_3134;
wire net_13458;
wire net_5523;
wire net_1720;
wire net_14164;
wire net_16825;
wire net_13885;
wire net_8191;
wire net_15098;
wire net_6104;
wire net_2060;
wire net_2051;
wire net_6087;
wire net_4535;
wire net_16807;
wire net_6426;
wire net_593;
wire net_21589;
wire net_19877;
wire net_5563;
wire net_10156;
wire net_18422;
wire net_16544;
wire net_6238;
wire net_20893;
wire net_17216;
wire net_2765;
wire net_15665;
wire net_15085;
wire net_22321;
wire x4848;
wire net_8341;
wire net_21500;
wire net_18353;
wire net_11044;
wire net_18683;
wire x266;
wire net_16383;
wire net_9597;
wire net_10343;
wire net_15449;
wire net_10320;
wire net_1198;
wire net_3975;
wire net_2862;
wire net_8100;
wire net_2457;
wire net_22504;
wire net_18237;
wire net_8260;
wire x790;
wire net_21923;
wire net_5533;
wire net_19340;
wire net_1516;
wire net_22578;
wire net_20576;
wire net_6782;
wire net_6473;
wire net_18777;
wire net_17317;
wire net_1083;
wire net_21976;
wire net_3423;
wire net_964;
wire net_2913;
wire x3268;
wire net_17245;
wire net_16018;
wire net_18257;
wire net_13729;
wire net_6402;
wire net_11003;
wire net_2268;
wire net_17930;
wire net_14352;
wire net_17384;
wire net_17044;
wire net_2846;
wire net_13331;
wire net_11685;
wire net_9479;
wire x3311;
wire net_4369;
wire net_18283;
wire net_16364;
wire net_21121;
wire net_20092;
wire net_6401;
wire net_10007;
wire net_4929;
wire net_3959;
wire net_4309;
wire net_8873;
wire net_12393;
wire net_11226;
wire net_6573;
wire net_1140;
wire net_18060;
wire net_2764;
wire net_1464;
wire net_16423;
wire net_22212;
wire net_11985;
wire net_4973;
wire net_3196;
wire net_14740;
wire net_5962;
wire net_515;
wire net_21883;
wire net_10620;
wire net_6806;
wire net_5121;
wire net_223;
wire net_15725;
wire net_7146;
wire net_2077;
wire net_20250;
wire net_15028;
wire net_19237;
wire net_7496;
wire net_16933;
wire net_2745;
wire net_19306;
wire net_16856;
wire net_13973;
wire net_5084;
wire net_3965;
wire net_19454;
wire net_13827;
wire net_15008;
wire net_6706;
wire net_7212;
wire net_572;
wire net_5289;
wire net_10955;
wire net_9614;
wire net_7850;
wire net_1662;
wire net_10396;
wire net_14615;
wire net_1079;
wire net_10148;
wire net_6760;
wire net_5198;
wire net_14318;
wire net_3235;
wire net_4938;
wire net_7099;
wire net_20367;
wire net_13261;
wire net_2391;
wire net_2802;
wire net_7965;
wire net_4614;
wire net_2906;
wire net_456;
wire x2115;
wire net_18332;
wire net_11299;
wire net_7238;
wire net_16750;
wire net_8533;
wire net_19279;
wire net_3428;
wire net_15781;
wire net_14528;
wire net_22117;
wire net_493;
wire net_16378;
wire net_6374;
wire net_6080;
wire net_14306;
wire net_6506;
wire net_987;
wire x797;
wire net_15963;
wire net_19098;
wire net_6167;
wire net_3620;
wire net_7781;
wire net_13824;
wire net_20703;
wire net_8475;
wire net_3271;
wire net_13183;
wire net_11197;
wire net_10675;
wire net_13098;
wire net_12568;
wire net_12276;
wire net_12418;
wire net_18816;
wire net_721;
wire net_9033;
wire net_7779;
wire x6697;
wire net_8164;
wire net_15590;
wire net_12127;
wire x392;
wire net_21369;
wire net_20142;
wire net_13634;
wire net_1018;
wire net_11085;
wire net_20181;
wire net_11701;
wire net_13289;
wire net_18519;
wire net_6591;
wire net_823;
wire net_9067;
wire net_9269;
wire net_7271;
wire net_4788;
wire x2713;
wire net_19844;
wire net_11774;
wire net_9541;
wire net_7892;
wire net_11028;
wire net_17367;
wire net_5428;
wire net_1191;
wire net_13688;
wire net_16311;
wire net_2255;
wire net_4754;
wire net_17485;
wire net_17596;
wire net_8970;
wire net_16236;
wire net_7471;
wire net_12918;
wire net_21303;
wire net_16257;
wire net_1019;
wire net_1616;
wire net_17389;
wire net_6180;
wire net_10348;
wire net_16064;
wire net_19182;
wire net_16625;
wire net_15902;
wire net_9415;
wire net_14181;
wire net_4342;
wire net_12863;
wire net_2969;
wire net_7518;
wire net_21126;
wire net_12522;
wire net_12351;
wire net_5490;
wire net_12960;
wire net_18734;
wire net_13167;
wire net_15078;
wire net_11406;
wire net_8886;
wire net_2985;
wire net_19272;
wire net_19766;
wire net_11551;
wire net_537;
wire net_18750;
wire net_12943;
wire net_11310;
wire net_10893;
wire net_12477;
wire net_22761;
wire net_19904;
wire net_13446;
wire net_5501;
wire net_19784;
wire net_18880;
wire net_12294;
wire net_3252;
wire net_17130;
wire net_18753;
wire net_16184;
wire net_5790;
wire net_5891;
wire net_513;
wire net_22780;
wire net_12020;
wire net_22487;
wire net_7950;
wire net_1576;
wire net_1421;
wire net_14282;
wire net_12462;
wire net_17742;
wire net_8737;
wire net_2736;
wire net_1280;
wire net_459;
wire net_12616;
wire net_9239;
wire x7654;
wire net_6590;
wire net_18510;
wire net_3412;
wire net_2113;
wire net_13305;
wire net_9397;
wire net_4793;
wire net_21314;
wire net_19253;
wire net_20567;
wire net_22319;
wire net_4760;
wire net_3915;
wire net_12737;
wire net_19772;
wire net_14424;
wire x5926;
wire net_21569;
wire net_18938;
wire net_5606;
wire net_19241;
wire net_8063;
wire net_19652;
wire net_8353;
wire net_22021;
wire net_5150;
wire net_22686;
wire net_9212;
wire net_12713;
wire net_8176;
wire net_21240;
wire net_11493;
wire net_7709;
wire net_12672;
wire net_18275;
wire net_1659;
wire net_19252;
wire net_589;
wire net_21441;
wire net_20728;
wire net_18329;
wire net_1814;
wire net_17851;
wire net_11610;
wire net_5981;
wire net_22100;
wire net_16703;
wire net_20304;
wire net_21722;
wire net_10186;
wire net_7319;
wire net_8698;
wire net_724;
wire net_9826;
wire net_9123;
wire net_8058;
wire net_2384;
wire net_16784;
wire net_16229;
wire net_7760;
wire net_5889;
wire net_2480;
wire net_9943;
wire net_12181;
wire net_9868;
wire net_874;
wire net_13706;
wire net_15909;
wire net_22180;
wire net_15264;
wire net_11399;
wire net_4277;
wire net_7907;
wire net_12107;
wire net_3674;
wire net_22642;
wire net_7555;
wire net_22028;
wire net_21236;
wire net_6187;
wire net_4966;
wire net_17749;
wire net_15522;
wire net_14973;
wire net_5244;
wire net_10178;
wire net_20917;
wire net_11182;
wire net_12857;
wire net_436;
wire net_18713;
wire net_2837;
wire net_7963;
wire net_7181;
wire net_5641;
wire net_21004;
wire net_11157;
wire net_2824;
wire net_1777;
wire net_12983;
wire net_8263;
wire net_18602;
wire net_15706;
wire net_13647;
wire net_20161;
wire net_12325;
wire net_7246;
wire net_12153;
wire net_12134;
wire net_5556;
wire net_17534;
wire net_1702;
wire net_21791;
wire net_4403;
wire net_7974;
wire net_6358;
wire net_16728;
wire net_1838;
wire net_11365;
wire net_10857;
wire net_358;
wire net_1973;
wire net_8748;
wire net_2934;
wire net_11427;
wire net_18026;
wire net_1285;
wire net_10364;
wire net_5912;
wire net_20498;
wire net_3112;
wire net_15320;
wire net_1175;
wire net_13207;
wire net_13118;
wire net_22559;
wire net_9453;
wire net_18361;
wire net_19964;
wire net_15970;
wire net_9934;
wire net_5722;
wire net_20547;
wire net_9312;
wire net_9191;
wire net_2922;
wire net_1742;
wire net_11884;
wire net_18003;
wire net_22681;
wire net_21208;
wire net_7641;
wire net_19914;
wire net_17427;
wire net_21155;
wire net_11823;
wire net_6890;
wire net_20691;
wire net_22632;
wire net_22575;
wire net_8011;
wire net_17988;
wire net_15368;
wire net_19898;
wire net_13734;
wire net_3370;
wire net_7025;
wire x7135;
wire net_13040;
wire net_15830;
wire net_9497;
wire net_3947;
wire net_3441;
wire net_18213;
wire net_4947;
wire net_16915;
wire net_4015;
wire net_3662;
wire net_12730;
wire net_16586;
wire net_8729;
wire net_9187;
wire net_22228;
wire net_13441;
wire net_16688;
wire net_6349;
wire net_16451;
wire net_16086;
wire net_10756;
wire net_17879;
wire net_18549;
wire net_3539;
wire net_2031;
wire net_1560;
wire net_4414;
wire net_12451;
wire net_4409;
wire net_17831;
wire net_12160;
wire net_10453;
wire net_6754;
wire net_17870;
wire net_13690;
wire net_8538;
wire net_9684;
wire net_20571;
wire net_8715;
wire net_14227;
wire net_13111;
wire net_21201;
wire net_7724;
wire net_6489;
wire net_1545;
wire net_20349;
wire x503;
wire net_4662;
wire net_18627;
wire net_8204;
wire net_10798;
wire net_18254;
wire net_13838;
wire net_2332;
wire net_20439;
wire net_12491;
wire net_2715;
wire net_1941;
wire net_14915;
wire net_13074;
wire net_13968;
wire net_14276;
wire net_3899;
wire net_17052;
wire net_1319;
wire net_8757;
wire net_3080;
wire net_11075;
wire net_15091;
wire net_1582;
wire net_4016;
wire net_22245;
wire net_6028;
wire net_13747;
wire net_2333;
wire net_6544;
wire net_6464;
wire net_17210;
wire net_1368;
wire net_1248;
wire x3147;
wire net_2238;
wire net_845;
wire net_10745;
wire net_8003;
wire net_22799;
wire net_10973;
wire net_9081;
wire net_695;
wire net_18987;
wire net_7692;
wire net_14086;
wire net_2671;
wire net_20933;
wire net_6787;
wire net_6569;
wire net_19407;
wire net_12761;
wire net_18542;
wire net_5896;
wire net_12788;
wire net_15169;
wire net_12610;
wire net_19697;
wire net_14605;
wire net_2198;
wire net_9043;
wire net_16341;
wire net_19148;
wire net_5250;
wire net_6435;
wire net_6661;
wire net_20470;
wire net_2940;
wire net_8672;
wire net_16346;
wire net_5583;
wire net_2095;
wire net_20332;
wire net_19988;
wire net_4681;
wire net_6955;
wire net_5231;
wire net_9726;
wire net_2314;
wire net_9905;
wire net_5454;
wire net_2613;
wire net_18958;
wire net_15311;
wire net_9995;
wire net_9010;
wire net_8849;
wire net_11479;
wire net_231;
wire net_10197;
wire net_16122;
wire net_17519;
wire x5787;
wire net_3024;
wire net_18860;
wire net_4691;
wire net_18520;
wire x7000;
wire net_22013;
wire net_20291;
wire net_19205;
wire net_17445;
wire net_12381;
wire net_17110;
wire net_4223;
wire net_11321;
wire net_2297;
wire net_13052;
wire net_9439;
wire net_3325;
wire net_6171;
wire net_582;
wire net_12485;
wire net_16671;
wire net_15331;
wire net_17187;
wire net_7419;
wire net_2341;
wire net_661;
wire net_3360;
wire net_13537;
wire net_15648;
wire net_11854;
wire net_17289;
wire net_9086;
wire net_18461;
wire net_10006;
wire net_22421;
wire net_9460;
wire net_17165;
wire net_18639;
wire net_21336;
wire net_210;
wire net_916;
wire net_3395;
wire net_22425;
wire net_21458;
wire net_11641;
wire net_4335;
wire net_851;
wire net_9924;
wire net_14865;
wire net_13247;
wire net_2426;
wire net_18196;
wire net_7405;
wire net_12237;
wire net_3310;
wire net_671;
wire net_8817;
wire net_8846;
wire net_14425;
wire net_12431;
wire net_6830;
wire net_6965;
wire net_20475;
wire net_8734;
wire net_18436;
wire net_16545;
wire net_12978;
wire net_9054;
wire net_17999;
wire net_15473;
wire net_307;
wire net_20101;
wire net_13938;
wire net_3547;
wire net_14497;
wire net_3543;
wire net_11470;
wire net_15298;
wire net_5104;
wire net_15248;
wire net_14774;
wire net_6069;
wire net_17935;
wire net_2656;
wire net_22388;
wire net_6326;
wire net_19883;
wire net_3922;
wire net_3212;
wire net_6530;
wire net_9632;
wire net_1764;
wire net_17684;
wire net_14067;
wire net_3513;
wire net_9968;
wire net_13290;
wire net_4042;
wire net_19713;
wire net_9691;
wire net_3335;
wire net_5377;
wire net_3682;
wire net_6456;
wire net_22266;
wire net_18198;
wire net_12245;
wire net_5655;
wire net_18168;
wire net_16839;
wire net_7856;
wire net_2667;
wire net_12818;
wire net_17238;
wire net_22569;
wire net_5431;
wire net_8443;
wire net_480;
wire net_7662;
wire net_4507;
wire net_4986;
wire net_2897;
wire net_18611;
wire net_5810;
wire net_19423;
wire net_836;
wire net_22623;
wire net_13817;
wire net_18382;
wire net_2161;
wire net_18551;
wire net_12075;
wire net_10671;
wire net_6568;
wire net_8408;
wire net_6059;
wire net_20501;
wire net_370;
wire net_22101;
wire net_16470;
wire net_16026;
wire net_20241;
wire net_21197;
wire net_13429;
wire net_6443;
wire net_1169;
wire net_13416;
wire net_7057;
wire net_7013;
wire net_13677;
wire net_9238;
wire net_7389;
wire net_2206;
wire net_21733;
wire net_11206;
wire net_1392;
wire net_14575;
wire net_6121;
wire net_311;
wire net_2479;
wire net_22529;
wire net_10132;
wire net_15453;
wire net_11119;
wire net_4469;
wire net_11452;
wire net_17726;
wire net_14598;
wire x402;
wire net_16280;
wire net_12527;
wire net_21660;
wire net_17899;
wire net_9986;
wire net_13210;
wire net_2520;
wire net_10166;
wire net_10768;
wire net_19851;
wire net_10704;
wire x2280;
wire net_6676;
wire net_2197;
wire net_15943;
wire net_19274;
wire net_10521;
wire net_5399;
wire net_10220;
wire net_12089;
wire net_9473;
wire net_14658;
wire net_2905;
wire net_10372;
wire net_200;
wire net_4435;
wire net_16489;
wire net_22089;
wire net_16032;
wire net_8612;
wire net_5220;
wire net_16463;
wire net_5995;
wire net_16208;
wire net_14706;
wire net_1853;
wire net_9741;
wire net_10119;
wire net_10240;
wire net_2170;
wire net_6851;
wire net_15304;
wire net_15026;
wire net_2678;
wire net_17605;
wire net_11036;
wire net_8346;
wire net_9119;
wire net_16965;
wire net_10256;
wire net_8906;
wire net_6698;
wire net_18228;
wire net_11267;
wire net_18301;
wire net_21502;
wire net_10381;
wire net_20508;
wire net_19354;
wire net_15609;
wire net_7717;
wire net_6988;
wire net_20129;
wire net_6281;
wire net_6209;
wire net_2864;
wire net_1998;
wire net_9341;
wire net_13621;
wire net_11656;
wire net_19525;
wire net_2795;
wire net_20748;
wire net_13587;
wire net_5540;
wire net_16214;
wire net_16166;
wire net_21046;
wire net_1918;
wire net_12790;
wire net_21250;
wire net_19050;
wire net_18421;
wire net_15388;
wire net_19716;
wire net_5870;
wire net_7894;
wire net_3236;
wire net_17964;
wire net_5837;
wire net_3201;
wire net_11812;
wire net_11169;
wire net_8147;
wire net_8096;
wire net_5613;
wire net_17510;
wire net_9560;
wire net_8966;
wire net_7163;
wire net_17889;
wire net_8024;
wire net_6897;
wire net_12912;
wire net_5300;
wire net_12359;
wire net_8926;
wire net_22584;
wire net_19313;
wire net_19411;
wire net_18677;
wire net_19543;
wire x0;
wire net_20839;
wire net_5803;
wire net_5410;
wire net_22405;
wire net_14838;
wire net_3650;
wire net_22009;
wire net_2465;
wire net_15544;
wire net_5078;
wire net_5447;
wire net_12043;
wire net_15230;
wire net_14465;
wire net_8485;
wire net_20402;
wire net_10388;
wire net_7462;
wire net_9900;
wire net_6023;
wire net_13862;
wire net_898;
wire net_14855;
wire net_6136;
wire net_10416;
wire net_16288;
wire net_15548;
wire net_13023;
wire net_8364;
wire net_7229;
wire net_7045;
wire net_22589;
wire net_8640;
wire x1551;
wire x1510;
wire net_20441;
wire net_1376;
wire net_5005;
wire net_13409;
wire net_8810;
wire net_6885;
wire net_22697;
wire net_6701;
wire net_18792;
wire net_1980;
wire net_13793;
wire net_20832;
wire net_9303;
wire net_1302;
wire net_244;
wire net_7341;
wire net_8687;
wire net_2395;
wire net_6012;
wire net_5347;
wire net_5439;
wire net_4002;
wire net_1989;
wire net_18642;
wire net_2855;
wire net_1795;
wire net_13310;
wire net_9247;
wire net_18878;
wire net_12186;
wire net_17597;
wire net_1539;
wire net_9626;
wire net_16538;
wire net_17193;
wire net_4261;
wire net_18871;
wire x3553;
wire net_10123;
wire net_3490;
wire net_3035;
wire net_7646;
wire net_14417;
wire net_22136;
wire net_15191;
wire x522;
wire net_11483;
wire net_13434;
wire net_16100;
wire net_6359;
wire net_12082;
wire net_11131;
wire net_7430;
wire net_20532;
wire net_20007;
wire net_7437;
wire net_1469;
wire net_15749;
wire net_11626;
wire net_18927;
wire net_4081;
wire net_15694;
wire net_2436;
wire net_81;
wire net_19136;
wire net_18427;
wire net_16811;
wire net_16403;
wire net_20741;
wire net_16454;
wire net_10793;
wire net_22735;
wire net_14176;
wire net_19168;
wire net_22439;
wire net_11878;
wire net_621;
wire net_10018;
wire net_5153;
wire net_13316;
wire net_10375;
wire net_105;
wire net_22726;
wire net_12586;
wire net_18246;
wire net_7729;
wire net_5598;
wire net_12591;
wire net_19473;
wire net_11276;
wire net_3985;
wire net_14492;
wire net_18648;
wire net_14801;
wire net_12390;
wire net_9792;
wire net_18770;
wire net_21755;
wire net_9552;
wire net_10229;
wire net_9689;
wire net_18101;
wire net_12663;
wire net_13032;
wire net_999;
wire net_15783;
wire net_8549;
wire net_21416;
wire net_10888;
wire net_8838;
wire net_20028;
wire net_13924;
wire net_22777;
wire net_9752;
wire net_4994;
wire net_19937;
wire net_3588;
wire net_9151;
wire net_1480;
wire net_18912;
wire net_22128;
wire net_14759;
wire net_15839;
wire net_7700;
wire net_4952;
wire net_21037;
wire net_377;
wire net_20277;
wire net_8836;
wire net_288;
wire net_16640;
wire net_2649;
wire net_1459;
wire net_12252;
wire net_7290;
wire net_5265;
wire net_11650;
wire net_22164;
wire net_7749;
wire net_3741;
wire net_13257;
wire net_4470;
wire net_9168;
wire net_540;
wire net_20785;
wire net_20280;
wire net_2642;
wire net_6650;
wire net_891;
wire net_19616;
wire net_12899;
wire net_9388;
wire net_5224;
wire net_3065;
wire net_21546;
wire net_5821;
wire net_4167;
wire net_15011;
wire net_7796;
wire net_6746;
wire net_4711;
wire net_10236;
wire net_5868;
wire net_18059;
wire net_10358;
wire net_18336;
wire net_16437;
wire net_4802;
wire net_22140;
wire net_16635;
wire net_618;
wire net_18786;
wire net_21515;
wire net_9075;
wire net_3688;
wire net_5759;
wire net_21768;
wire net_12001;
wire net_12399;
wire net_22721;
wire net_20387;
wire net_8256;
wire net_6970;
wire net_19921;
wire net_14907;
wire net_21084;
wire net_19107;
wire net_14255;
wire net_5945;
wire net_6148;
wire net_754;
wire net_10785;
wire net_7193;
wire net_921;
wire net_9113;
wire net_21801;
wire net_7989;
wire net_17569;
wire net_20499;
wire net_11581;
wire net_4957;
wire net_14900;
wire net_3308;
wire net_12607;
wire net_10274;
wire net_16772;
wire net_2192;
wire net_1533;
wire net_20203;
wire net_16440;
wire net_16336;
wire net_8565;
wire net_7999;
wire net_7681;
wire net_21007;
wire net_9138;
wire net_15525;
wire net_11158;
wire net_9884;
wire net_3502;
wire net_14014;
wire net_22535;
wire net_21686;
wire net_4827;
wire net_654;
wire net_17248;
wire net_330;
wire net_3506;
wire net_19750;
wire net_22137;
wire net_20609;
wire net_16953;
wire net_8082;
wire net_19317;
wire net_14538;
wire net_9116;
wire net_570;
wire net_444;
wire net_525;
wire net_3829;
wire net_3646;
wire net_1210;
wire net_1067;
wire net_15575;
wire net_6624;
wire net_5058;
wire net_18746;
wire net_16882;
wire net_14920;
wire net_5998;
wire net_7820;
wire net_16971;
wire net_14681;
wire net_16569;
wire net_6200;
wire net_6259;
wire net_15206;
wire net_3933;
wire net_19218;
wire net_20461;
wire net_18584;
wire net_21669;
wire net_11629;
wire net_22296;
wire net_16300;
wire net_20066;
wire net_19793;
wire net_22111;
wire net_9325;
wire net_4820;
wire net_21988;
wire net_13486;
wire net_10055;
wire net_7577;
wire net_16579;
wire net_15828;
wire net_22169;
wire net_9409;
wire net_9404;
wire net_1178;
wire net_20844;
wire net_9722;
wire net_5573;
wire net_17372;
wire net_7098;
wire net_19369;
wire net_3825;
wire net_11142;
wire net_6218;
wire net_17177;
wire net_16097;
wire net_12380;
wire net_340;
wire net_6039;
wire net_16057;
wire net_15885;
wire net_15435;
wire net_2634;
wire net_434;
wire net_6915;
wire net_8434;
wire net_7024;
wire net_6936;
wire net_14200;
wire net_1797;
wire net_20671;
wire net_21224;
wire net_9443;
wire net_19674;
wire net_11086;
wire net_69;
wire net_19817;
wire net_14732;
wire net_4906;
wire net_4524;
wire net_339;
wire net_7686;
wire net_17848;
wire net_13105;
wire net_3468;
wire net_10443;
wire net_11775;
wire net_18918;
wire net_12753;
wire net_20266;
wire net_2710;
wire net_19492;
wire net_15722;
wire net_2660;
wire net_14486;
wire net_8624;
wire net_10083;
wire net_8087;
wire net_5389;
wire net_3671;
wire net_8236;
wire net_8651;
wire net_20630;
wire net_21804;
wire net_3691;
wire net_21662;
wire net_17562;
wire net_678;
wire net_15771;
wire net_21361;
wire net_16503;
wire net_11631;
wire net_8979;
wire net_928;
wire net_15251;
wire net_5459;
wire net_13363;
wire net_208;
wire net_9225;
wire net_20296;
wire net_7878;
wire net_8215;
wire net_2744;
wire net_2377;
wire net_415;
wire net_116;
wire net_3251;
wire net_2786;
wire net_347;
wire net_14784;
wire net_13526;
wire net_11059;
wire net_19977;
wire net_3794;
wire net_22756;
wire net_12664;
wire net_15997;
wire net_20011;
wire net_20229;
wire net_7306;
wire net_22147;
wire net_20708;
wire net_20992;
wire net_16551;
wire net_1335;
wire net_19854;
wire net_18874;
wire net_21973;
wire net_15716;
wire net_19994;
wire net_21918;
wire net_15519;
wire net_12210;
wire net_5477;
wire net_18154;
wire net_16932;
wire net_2212;
wire net_22538;
wire net_19518;
wire net_5453;
wire net_20341;
wire net_11535;
wire net_7730;
wire net_16725;
wire x1912;
wire net_16499;
wire net_3571;
wire x7336;
wire net_22031;
wire net_4642;
wire net_610;
wire net_8130;
wire net_16889;
wire net_21115;
wire net_7870;
wire net_19812;
wire net_19049;
wire net_15187;
wire net_2344;
wire net_10588;
wire net_1323;
wire net_21216;
wire net_14130;
wire net_1506;
wire net_10470;
wire net_17836;
wire net_13386;
wire net_6496;
wire net_13193;
wire net_22416;
wire net_539;
wire net_16617;
wire net_13068;
wire net_692;
wire net_22284;
wire net_16094;
wire net_18971;
wire net_4568;
wire net_10807;
wire net_17551;
wire net_4377;
wire net_16660;
wire net_15130;
wire net_14261;
wire net_7704;
wire net_13125;
wire net_15104;
wire net_10311;
wire net_1400;
wire net_885;
wire net_9202;
wire net_11698;
wire x1975;
wire net_14320;
wire net_9918;
wire net_18276;
wire net_21391;
wire net_10770;
wire net_6822;
wire net_11607;
wire net_6594;
wire net_3517;
wire net_761;
wire net_496;
wire net_20639;
wire net_11396;
wire net_1554;
wire net_22156;
wire net_7101;
wire net_16779;
wire net_22562;
wire net_22192;
wire net_21326;
wire net_10638;
wire net_4370;
wire net_18980;
wire net_4979;
wire net_14613;
wire net_12578;
wire net_2249;
wire net_19459;
wire net_16106;
wire x1299;
wire net_5686;
wire net_15129;
wire net_739;
wire net_22305;
wire net_21033;
wire net_8760;
wire net_20095;
wire net_19956;
wire net_20057;
wire net_17529;
wire net_17472;
wire x2978;
wire net_826;
wire net_15069;
wire net_1738;
wire net_10384;
wire net_10504;
wire net_14887;
wire net_19154;
wire net_16178;
wire net_11644;
wire net_6716;
wire net_20313;
wire net_2624;
wire net_11761;
wire net_343;
wire net_20947;
wire net_19336;
wire net_19655;
wire net_17038;
wire net_20114;
wire net_7313;
wire net_9672;
wire net_8456;
wire x246;
wire net_5236;
wire net_4424;
wire net_19416;
wire net_7541;
wire net_9615;
wire net_7451;
wire net_2487;
wire net_7803;
wire net_19487;
wire net_19067;
wire net_8227;
wire net_17649;
wire net_13132;
wire net_15674;
wire net_2975;
wire net_17201;
wire net_4625;
wire net_5257;
wire net_8220;
wire net_2779;
wire net_14187;
wire net_11552;
wire net_17494;
wire net_16225;
wire net_6392;
wire net_18990;
wire net_15158;
wire net_9346;
wire net_11352;
wire net_8169;
wire net_1490;
wire net_9274;
wire net_4282;
wire net_15216;
wire net_17066;
wire net_11806;
wire net_12774;
wire net_18923;
wire net_17926;
wire net_22824;
wire net_19520;
wire net_15565;
wire net_14765;
wire net_14342;
wire net_5742;
wire net_19624;
wire net_4356;
wire net_21788;
wire net_685;
wire net_8466;
wire net_20684;
wire net_18808;
wire net_16307;
wire net_12349;
wire net_19196;
wire net_17711;
wire net_11843;
wire net_4052;
wire net_8513;
wire net_21942;
wire net_18224;
wire net_8681;
wire net_15953;
wire x1639;
wire net_16897;
wire net_22133;
wire net_17049;
wire net_13469;
wire net_10652;
wire net_7160;
wire net_20962;
wire net_17633;
wire net_12876;
wire net_4686;
wire net_1946;
wire net_2733;
wire net_17204;
wire net_14280;
wire net_18697;
wire net_6764;
wire net_13252;
wire net_6769;
wire net_3612;
wire net_11634;
wire net_1605;
wire net_12795;
wire net_18726;
wire net_21571;
wire net_22772;
wire net_18702;
wire net_5118;
wire x745;
wire net_747;
wire net_20206;
wire net_15597;
wire net_2305;
wire net_1653;
wire net_14125;
wire net_5842;
wire net_9817;
wire net_7377;
wire net_16023;
wire net_22617;
wire net_21934;
wire net_2258;
wire net_22571;
wire net_11168;
wire net_12510;
wire net_14327;
wire net_17397;
wire net_19178;
wire net_6500;
wire net_17276;
wire net_2367;
wire net_21991;
wire net_15977;
wire net_14697;
wire net_4573;
wire net_4127;
wire net_16900;
wire net_2810;
wire net_13546;
wire net_1053;
wire net_11292;
wire net_1004;
wire net_21627;
wire net_4921;
wire net_17939;
wire net_11716;
wire net_11359;
wire net_21751;
wire net_3232;
wire net_13356;
wire net_4498;
wire net_21837;
wire net_19865;
wire net_3228;
wire net_19870;
wire net_2282;
wire net_10029;
wire net_20192;
wire net_1546;
wire net_11367;
wire net_8542;
wire net_15695;
wire net_6042;
wire net_13654;
wire net_20174;
wire net_18849;
wire net_16390;
wire net_1046;
wire net_19573;
wire net_19016;
wire net_11502;
wire net_10332;
wire net_4960;
wire net_1213;
wire net_22768;
wire net_2265;
wire net_8118;
wire net_16948;
wire net_10163;
wire net_22370;
wire net_16479;
wire net_5795;
wire net_12812;
wire net_769;
wire net_1780;
wire net_13668;
wire net_19761;
wire net_16132;
wire net_19600;
wire net_1025;
wire net_3758;
wire net_15062;
wire net_13157;
wire net_10403;
wire net_7502;
wire net_15807;
wire net_1089;
wire net_12169;
wire net_16359;
wire net_11998;
wire net_16386;
wire net_4528;
wire net_6233;
wire net_5625;
wire net_16695;
wire net_4141;
wire net_19482;
wire net_18292;
wire net_14094;
wire net_12535;
wire net_10669;
wire net_5146;
wire net_16713;
wire net_8701;
wire net_22498;
wire net_5326;
wire net_12921;
wire net_17923;
wire net_4394;
wire net_18082;
wire net_15421;
wire net_5953;
wire net_12442;
wire net_11047;
wire net_12702;
wire net_9433;
wire net_10816;
wire net_14124;
wire net_13248;
wire net_3626;
wire net_15924;
wire net_12095;
wire net_5779;
wire net_14798;
wire net_21844;
wire net_6417;
wire net_4726;
wire net_20590;
wire net_15475;
wire net_14377;
wire net_13086;
wire net_9588;
wire net_18033;
wire net_17220;
wire net_14572;
wire net_5344;
wire net_20584;
wire net_7492;
wire net_12468;
wire net_5364;
wire net_18945;
wire net_8743;
wire net_6388;
wire net_13478;
wire net_740;
wire net_4072;
wire net_11090;
wire net_21700;
wire net_5825;
wire net_3183;
wire net_19687;
wire net_17863;
wire net_3908;
wire net_4837;
wire net_730;
wire net_4150;
wire net_8049;
wire net_7094;
wire net_5405;
wire net_22494;
wire net_22448;
wire net_11931;
wire net_2105;
wire net_20704;
wire net_16371;
wire net_7226;
wire net_1127;
wire net_6381;
wire net_17226;
wire net_9458;
wire net_11243;
wire net_6420;
wire net_13831;
wire net_18176;
wire net_7465;
wire net_9297;
wire net_15732;
wire net_4143;
wire net_12900;
wire net_18768;
wire net_8679;
wire net_7285;
wire net_5140;
wire net_3123;
wire net_2955;
wire net_19232;
wire net_20951;
wire net_22390;
wire net_771;
wire net_2301;
wire net_2978;
wire net_19226;
wire net_15033;
wire net_5185;
wire net_13139;
wire net_21816;
wire net_19297;
wire net_3950;
wire x6224;
wire net_22179;
wire net_22214;
wire net_1062;
wire net_14395;
wire net_4936;
wire net_3293;
wire net_22208;
wire net_4120;
wire net_9246;
wire net_7733;
wire net_16263;
wire net_14987;
wire net_6050;
wire net_21016;
wire net_13214;
wire net_5188;
wire net_4590;
wire net_18343;
wire net_18096;
wire net_6116;
wire net_16512;
wire net_1411;
wire net_12549;
wire net_505;
wire net_4088;
wire net_16862;
wire net_10471;
wire net_3723;
wire net_14724;
wire net_10493;
wire net_10426;
wire net_7152;
wire net_6527;
wire net_992;
wire net_21243;
wire net_7485;
wire net_15933;
wire net_9781;
wire net_6727;
wire net_782;
wire net_22565;
wire net_22054;
wire net_10527;
wire net_13576;
wire net_11106;
wire net_18347;
wire net_22399;
wire net_6291;
wire net_4186;
wire net_13328;
wire net_4738;
wire net_3314;
wire net_7422;
wire net_2971;
wire net_22359;
wire net_5776;
wire net_17102;
wire net_13322;
wire net_10339;
wire net_20481;
wire net_8072;
wire net_8244;
wire net_2836;
wire net_10615;
wire net_5689;
wire net_7429;
wire net_1805;
wire net_4667;
wire net_11536;
wire x3791;
wire net_10660;
wire net_3635;
wire net_17838;
wire net_13559;
wire net_7120;
wire net_1110;
wire net_17423;
wire net_15356;
wire net_442;
wire net_14999;
wire net_22084;
wire net_13789;
wire net_22393;
wire net_21597;
wire net_16594;
wire net_7202;
wire net_20238;
wire net_21696;
wire net_3087;
wire net_17402;
wire net_14627;
wire net_13900;
wire net_1821;
wire net_19539;
wire net_42;
wire net_11675;
wire net_7480;
wire net_3865;
wire net_1588;
wire net_9029;
wire net_4037;
wire net_3937;
wire net_1495;
wire net_17080;
wire net_18800;
wire net_2992;
wire net_12974;
wire net_17227;
wire net_16329;
wire net_3522;
wire net_668;
wire net_7601;
wire net_18142;
wire net_15758;
wire net_3079;
wire net_14203;
wire net_17733;
wire net_8040;
wire net_5814;
wire net_20657;
wire net_12707;
wire net_1070;
wire net_20723;
wire net_21913;
wire net_8878;
wire net_1225;
wire net_812;
wire net_22079;
wire x3052;
wire net_19709;
wire net_14993;
wire net_13805;
wire net_18830;
wire net_6314;
wire net_6972;
wire net_1107;
wire net_16563;
wire net_22807;
wire net_15850;
wire net_11053;
wire net_18581;
wire net_15621;
wire net_3384;
wire net_1203;
wire net_13347;
wire net_22658;
wire net_15055;
wire net_9011;
wire net_12402;
wire net_12176;
wire net_10867;
wire net_10715;
wire net_5321;
wire net_11434;
wire net_12789;
wire net_21863;
wire net_22377;
wire net_20674;
wire net_17440;
wire x687;
wire net_17652;
wire net_5884;
wire net_863;
wire net_7131;
wire net_6468;
wire net_3164;
wire net_22709;
wire net_16527;
wire net_16998;
wire net_14058;
wire net_13150;
wire net_904;
wire net_19292;
wire net_21102;
wire net_15580;
wire net_12850;
wire net_14226;
wire net_13552;
wire net_58;
wire net_16244;
wire net_6777;
wire net_12286;
wire net_6633;
wire net_8126;
wire net_22349;
wire net_6092;
wire net_16813;
wire net_6559;
wire net_15553;
wire net_11360;
wire net_9183;
wire net_15688;
wire net_4845;
wire net_1160;
wire net_18630;
wire net_15917;
wire net_159;
wire net_11147;
wire net_9379;
wire net_3268;
wire net_18939;
wire net_5863;
wire net_11615;
wire net_9523;
wire net_10181;
wire x936;
wire net_19171;
wire net_9354;
wire net_14834;
wire net_2875;
wire x6300;
wire net_12952;
wire net_20967;
wire net_10213;
wire x2149;
wire net_324;
wire net_20982;
wire net_6848;
wire net_11724;
wire net_10284;
wire net_10074;
wire net_13397;
wire net_5480;
wire net_14675;
wire net_10309;
wire net_18761;
wire net_16354;
wire net_7257;
wire net_17776;
wire net_13047;
wire net_9706;
wire net_14248;
wire net_14103;
wire net_17616;
wire net_12647;
wire net_10964;
wire net_5046;
wire net_3066;
wire net_19054;
wire net_20698;
wire net_6270;
wire net_15385;
wire net_20451;
wire net_6275;
wire net_17805;
wire net_4181;
wire net_376;
wire net_20199;
wire net_21895;
wire net_19131;
wire net_17909;
wire net_2133;
wire net_17703;
wire net_13643;
wire net_16978;
wire net_4817;
wire net_13374;
wire net_2515;
wire net_19020;
wire net_3173;
wire net_8038;
wire net_3738;
wire net_17393;
wire net_7994;
wire net_15529;
wire net_5298;
wire net_5119;
wire net_422;
wire net_4290;
wire net_21056;
wire net_18048;
wire net_14739;
wire net_1345;
wire net_1450;
wire net_561;
wire net_12694;
wire net_4899;
wire net_20216;
wire net_5955;
wire net_8501;
wire net_4299;
wire net_2290;
wire net_12741;
wire net_2851;
wire net_17140;
wire net_8427;
wire net_14640;
wire net_21536;
wire net_14019;
wire net_21434;
wire net_3772;
wire net_7901;
wire net_20226;
wire net_4868;
wire net_2698;
wire net_6552;
wire net_18653;
wire net_8453;
wire net_3450;
wire net_14412;
wire net_14813;
wire net_3528;
wire net_8559;
wire net_18005;
wire net_8956;
wire net_350;
wire net_4270;
wire net_8332;
wire net_13178;
wire net_7606;
wire net_13275;
wire net_18075;
wire net_3117;
wire net_20745;
wire net_16753;
wire net_14245;
wire net_19325;
wire net_11816;
wire net_3482;
wire net_6648;
wire net_7375;
wire x2688;
wire net_15712;
wire net_19923;
wire net_21194;
wire net_3369;
wire net_9020;
wire net_1101;
wire net_994;
wire net_21425;
wire net_12828;
wire net_12268;
wire net_18919;
wire net_19333;
wire net_21554;
wire net_6685;
wire net_11837;
wire net_4166;
wire net_4608;
wire net_21615;
wire net_15122;
wire net_3340;
wire net_21284;
wire net_4545;
wire net_3844;
wire net_1849;
wire net_10045;
wire net_5486;
wire net_16647;
wire net_13516;
wire net_14994;
wire net_14637;
wire net_11122;
wire net_1108;
wire net_22791;
wire net_8583;
wire net_9756;
wire net_1878;
wire net_16598;
wire net_16820;
wire net_16231;
wire net_17314;
wire net_13070;
wire net_16678;
wire net_9255;
wire net_16435;
wire net_11446;
wire net_20883;
wire net_3890;
wire net_5975;
wire net_133;
wire net_20105;
wire net_7528;
wire net_4025;
wire net_16112;
wire net_9194;
wire net_15459;
wire net_7078;
wire net_7008;
wire net_11957;
wire net_3882;
wire net_557;
wire net_3043;
wire net_15288;
wire net_7860;
wire net_6611;
wire net_19134;
wire net_13891;
wire net_11386;
wire net_12316;
wire net_1991;
wire net_1611;
wire net_18201;
wire net_20257;
wire net_22523;
wire net_14046;
wire net_1431;
wire net_1714;
wire net_21939;
wire net_18135;
wire net_19214;
wire net_13014;
wire net_11970;
wire net_16945;
wire net_18827;
wire net_8868;
wire net_240;
wire net_15115;
wire net_20435;
wire net_15872;
wire net_18147;
wire net_17261;
wire net_17588;
wire net_295;
wire net_22132;
wire net_8411;
wire net_18558;
wire net_13425;
wire net_9241;
wire net_20871;
wire net_5935;
wire net_17326;
wire net_22265;
wire net_13490;
wire net_7753;
wire net_15236;
wire net_14879;
wire net_12115;
wire net_7720;
wire net_16462;
wire net_22453;
wire net_11239;
wire net_12619;
wire net_6691;
wire net_12967;
wire net_278;
wire net_20775;
wire net_18208;
wire net_6864;
wire net_21479;
wire net_19029;
wire net_9063;
wire net_4874;
wire net_10090;
wire net_16794;
wire net_13309;
wire x7497;
wire net_17952;
wire net_2443;
wire net_22064;
wire x7698;
wire net_10736;
wire net_1307;
wire net_4514;
wire net_21370;
wire x570;
wire net_15857;
wire net_17499;
wire net_19880;
wire net_15753;
wire net_6940;
wire net_5591;
wire net_4810;
wire net_15413;
wire net_4418;
wire net_17959;
wire net_5385;
wire net_14145;
wire net_22597;
wire net_6099;
wire net_9786;
wire net_12679;
wire net_7630;
wire net_19445;
wire net_21310;
wire net_13854;
wire net_13712;
wire net_3776;
wire net_17954;
wire net_1252;
wire net_9173;
wire net_7739;
wire net_19643;
wire net_9095;
wire net_7784;
wire net_16700;
wire net_10731;
wire net_507;
wire net_10097;
wire net_8981;
wire net_1902;
wire net_17115;
wire net_7111;
wire net_2600;
wire net_5734;
wire net_22749;
wire net_20724;
wire net_3563;
wire net_12224;
wire net_8726;
wire net_6585;
wire net_9565;
wire net_19868;
wire net_11936;
wire net_4491;
wire net_11543;
wire net_8282;
wire net_7538;
wire net_16737;
wire net_1962;
wire net_291;
wire net_9502;
wire net_7351;
wire net_1964;
wire net_857;
wire net_867;
wire net_21452;
wire net_5964;
wire net_15618;
wire net_396;
wire net_22515;
wire net_21741;
wire net_14845;
wire net_10602;
wire net_17468;
wire net_8851;
wire net_10535;
wire net_20539;
wire net_1541;
wire net_14966;
wire net_14216;
wire net_9748;
wire net_15683;
wire net_5177;
wire net_271;
wire net_3329;
wire net_10067;
wire net_6111;
wire net_12208;
wire net_14693;
wire net_3611;
wire net_2064;
wire net_15274;
wire net_5333;
wire net_1925;
wire net_1909;
wire net_16664;
wire net_1410;
wire net_365;
wire net_21992;
wire net_13412;
wire net_19350;
wire net_18043;
wire net_3344;
wire net_12060;
wire net_8374;
wire net_10729;
wire net_4413;
wire net_13849;
wire net_8719;
wire net_4313;
wire net_21813;
wire net_16483;
wire net_16830;
wire net_11000;
wire net_22463;
wire net_16448;
wire net_8313;
wire net_16630;
wire net_9339;
wire net_19287;
wire net_7128;
wire net_7915;
wire net_22592;
wire net_13723;
wire net_13730;
wire net_4892;
wire net_803;
wire net_19706;
wire net_10884;
wire net_14713;
wire net_14111;
wire net_7764;
wire net_6375;
wire net_17501;
wire net_1476;
wire net_1293;
wire net_14939;
wire net_11098;
wire net_2883;
wire net_8665;
wire net_11742;
wire net_2681;
wire net_12159;
wire net_9629;
wire net_18181;
wire net_17791;
wire net_5136;
wire net_22247;
wire net_22067;
wire net_18598;
wire net_4855;
wire net_14668;
wire net_22419;
wire net_19320;
wire net_1266;
wire net_1452;
wire net_2773;
wire net_17995;
wire net_909;
wire net_4529;
wire net_4898;
wire net_152;
wire x5754;
wire net_11575;
wire net_3105;
wire net_2138;
wire net_16153;
wire net_258;
wire net_11192;
wire net_10761;
wire net_16196;
wire net_12935;
wire net_12054;
wire net_19033;
wire net_19017;
wire net_13983;
wire net_20850;
wire net_5083;
wire net_2446;
wire net_18576;
wire net_7171;
wire net_20370;
wire net_11999;
wire net_15644;
wire x3090;
wire net_7605;
wire net_585;
wire net_7611;
wire net_17754;
wire net_7809;
wire net_14823;
wire net_11913;
wire net_11347;
wire net_12061;
wire net_10593;
wire net_14514;
wire net_20715;
wire net_10293;
wire net_20780;
wire net_12632;
wire net_788;
wire net_19567;
wire net_9090;
wire net_214;
wire net_22033;
wire net_20543;
wire net_8113;
wire net_13028;
wire net_8144;
wire net_3578;
wire net_12455;
wire net_13903;
wire net_8804;
wire net_21064;
wire net_20042;
wire net_6310;
wire x173;
wire net_5097;
wire net_7329;
wire net_18409;
wire net_4259;
wire net_2565;
wire net_17890;
wire net_8018;
wire net_21259;
wire net_19777;
wire net_13229;
wire net_22272;
wire net_6783;
wire net_5908;
wire net_2118;
wire net_463;
wire net_15281;
wire net_17946;
wire net_9487;
wire net_197;
wire net_18867;
wire net_2560;
wire net_9331;
wire net_5017;
wire net_3709;
wire net_21027;
wire net_13085;
wire net_12803;
wire net_7588;
wire net_11468;
wire net_5352;
wire net_2595;
wire net_22314;
wire net_1383;
wire net_7302;
wire net_2751;
wire net_9663;
wire net_9165;
wire net_20798;
wire net_18462;
wire net_4446;
wire net_14160;
wire net_10484;
wire net_6269;
wire net_6176;
wire net_14170;
wire net_13672;
wire net_21520;
wire net_11116;
wire net_13497;
wire net_1683;
wire net_22092;
wire net_17178;
wire net_17027;
wire net_12515;
wire net_978;
wire net_15510;
wire net_1313;
wire net_7618;
wire net_3331;
wire net_15855;
wire net_16891;
wire net_11994;
wire net_13286;
wire net_5712;
wire net_14446;
wire net_10877;
wire net_8383;
wire net_9954;
wire net_6360;
wire net_17351;
wire net_17298;
wire net_1789;
wire net_14035;
wire net_13142;
wire net_13940;
wire net_19722;
wire net_3219;
wire net_20412;
wire net_7520;
wire net_4587;
wire net_20124;
wire net_18286;
wire net_2576;
wire net_2352;
wire net_1038;
wire net_19729;
wire net_6931;
wire net_4241;
wire net_9920;
wire net_8168;
wire net_22070;
wire net_5710;
wire net_5369;
wire net_3763;
wire net_15445;
wire net_6333;
wire net_19730;
wire net_11338;
wire net_14662;
wire net_7697;
wire net_22016;
wire net_2277;
wire net_17162;
wire net_6078;
wire net_975;
wire net_21098;
wire net_5421;
wire net_21605;
wire net_15538;
wire net_4650;
wire net_19374;
wire net_15805;
wire net_13061;
wire net_15735;
wire net_6160;
wire net_5874;
wire net_18489;
wire net_2006;
wire net_13570;
wire net_1331;
wire net_20562;
wire net_18474;
wire net_19193;
wire net_12307;
wire net_20556;
wire net_15071;
wire net_5826;
wire net_18908;
wire net_13912;
wire net_18065;
wire net_16071;
wire net_8604;
wire net_2728;
wire net_17070;
wire net_18109;
wire net_4636;
wire net_122;
wire net_20287;
wire net_6264;
wire net_19129;
wire net_17991;
wire net_13619;
wire net_12847;
wire net_11514;
wire net_10026;
wire x1322;
wire net_16550;
wire net_9262;
wire net_18456;
wire net_14752;
wire net_4092;
wire net_17406;
wire net_12300;
wire net_8595;
wire net_94;
wire net_21483;
wire net_19676;
wire net_11760;
wire net_10751;
wire net_15361;
wire net_4486;
wire net_9427;
wire net_19383;
wire net_18054;
wire net_9131;
wire net_15905;
wire net_17197;
wire net_10983;
wire net_7262;
wire net_387;
wire net_22275;
wire net_15327;
wire net_3275;
wire net_7447;
wire net_6297;
wire net_18524;
wire net_17660;
wire net_10828;
wire net_5291;
wire net_1893;
wire net_20373;
wire net_16509;
wire net_15355;
wire net_1932;
wire net_9639;
wire net_8896;
wire net_11620;
wire net_8268;
wire net_21161;
wire net_19692;
wire net_3836;
wire net_15777;
wire net_14554;
wire net_1957;
wire net_10102;
wire net_13743;
wire net_13231;
wire net_9368;
wire net_15377;
wire net_7581;
wire net_2572;
wire net_60;
wire net_2414;
wire net_20636;
wire net_19003;
wire net_1846;
wire net_21074;
wire net_20826;
wire net_20423;
wire net_13381;
wire net_5667;
wire net_20152;
wire net_11222;
wire net_9662;
wire x2802;
wire net_7888;
wire net_12475;
wire net_11066;
wire net_13984;
wire net_4254;
wire net_13760;
wire net_3815;
wire net_3555;
wire net_17810;
wire net_18538;
wire net_5739;
wire net_2371;
wire net_21437;
wire net_6794;
wire net_14077;
wire net_21948;
wire net_21785;
wire net_19060;
wire net_13368;
wire net_11014;
wire net_16622;
wire net_8396;
wire net_12546;
wire net_9640;
wire net_7843;
wire net_7392;
wire net_3982;
wire net_1388;
wire net_4709;
wire net_14409;
wire net_14959;
wire net_20818;
wire net_19546;
wire net_9858;
wire net_3391;
wire net_15018;
wire net_2730;
wire x6430;
wire net_6835;
wire net_13553;
wire net_4655;
wire net_1624;
wire net_6618;
wire net_12332;
wire net_20324;
wire net_1638;
wire net_21340;
wire net_20640;
wire net_7455;
wire net_3875;
wire net_12146;
wire net_9319;
wire net_14436;
wire net_10135;
wire net_5268;
wire net_11389;
wire net_20923;
wire net_22353;
wire net_21856;
wire net_14980;
wire net_6335;
wire net_2153;
wire net_17692;
wire net_1939;
wire net_9582;
wire net_8781;
wire net_3098;
wire net_7242;
wire net_20136;
wire net_14190;
wire net_6288;
wire net_4673;
wire net_5762;
wire net_9061;
wire net_10249;
wire net_16852;
wire net_20088;
wire net_7828;
wire net_162;
wire net_21348;
wire net_15751;
wire net_14952;
wire net_8301;
wire net_7776;
wire net_653;
wire net_14301;
wire net_13160;
wire net_22531;
wire net_16909;
wire net_5066;
wire net_13919;
wire net_14718;
wire net_11735;
wire net_12030;
wire net_21941;
wire net_3145;
wire net_9558;
wire net_15879;
wire net_13694;
wire net_3694;
wire net_16001;
wire net_18661;
wire net_14880;
wire net_10262;
wire net_11592;
wire net_3855;
wire net_236;
wire net_12324;
wire net_9286;
wire net_552;
wire net_10823;
wire net_8206;
wire net_1787;
wire net_19942;
wire net_17897;
wire net_3551;
wire net_6654;
wire net_7440;
wire net_14791;
wire net_13390;
wire net_22625;
wire net_9518;
wire net_7067;
wire net_17300;
wire net_16980;
wire net_15143;
wire net_16910;
wire net_8329;
wire net_104;
wire x3667;
wire net_19496;
wire net_14402;
wire net_21233;
wire net_3416;
wire net_7198;
wire net_18686;
wire net_5166;
wire net_17609;
wire net_15992;
wire net_21371;
wire net_14595;
wire net_4886;
wire net_9878;
wire net_17479;
wire net_15655;
wire net_10914;
wire net_14070;
wire net_12039;
wire net_8522;
wire net_6659;
wire net_12192;
wire net_6877;
wire net_711;
wire net_17882;
wire net_19435;
wire net_20857;
wire net_20270;
wire net_15635;
wire net_18952;
wire net_17309;
wire net_8618;
wire net_4700;
wire net_846;
wire net_17152;
wire net_3017;
wire net_11864;
wire net_4677;
wire net_16880;
wire net_20073;
wire net_8033;
wire net_21317;
wire net_20232;
wire net_16515;
wire net_10996;
wire net_10038;
wire net_5768;
wire net_18021;
wire net_2607;
wire net_7799;
wire net_15210;
wire net_7957;
wire net_10971;
wire net_14755;
wire net_19940;
wire net_21020;
wire net_8769;
wire net_13870;
wire net_5023;
wire net_79;
wire net_2168;
wire net_18072;
wire net_17091;
wire net_1885;
wire net_1030;
wire net_14357;
wire net_10406;
wire net_6929;
wire net_16272;
wire net_10682;
wire net_19949;
wire net_15498;
wire net_11498;
wire net_10031;
wire net_4773;
wire net_4201;
wire net_4273;
wire net_1969;
wire net_22782;
wire net_7991;
wire net_15514;
wire net_12306;
wire net_8009;
wire net_7064;
wire net_17007;
wire net_933;
wire net_22682;
wire net_12532;
wire net_12036;
wire net_10860;
wire net_3377;
wire net_373;
wire net_16573;
wire net_21254;
wire net_16357;
wire net_452;
wire net_16046;
wire net_3683;
wire net_20937;
wire net_1483;
wire net_8067;
wire net_3031;
wire net_17707;
wire net_20212;
wire net_2645;
wire net_20652;
wire net_10433;
wire net_5356;
wire net_14386;
wire net_8078;
wire net_7674;
wire net_7386;
wire net_6684;
wire net_4278;
wire net_2674;
wire net_16847;
wire net_13801;
wire net_10193;
wire net_8934;
wire net_22815;
wire net_7059;
wire net_14428;
wire net_19295;
wire net_1671;
wire net_4764;
wire x4285;
wire net_665;
wire net_1746;
wire net_2222;
wire net_21173;
wire net_2825;
wire net_17343;
wire net_7209;
wire net_18478;
wire net_3670;
wire net_14647;
wire net_5940;
wire x4215;
wire net_5985;
wire net_7925;
wire net_16565;
wire net_6606;
wire net_10182;
wire net_20104;
wire net_10376;
wire net_4861;
wire net_11666;
wire x1963;
wire net_109;
wire net_1706;
wire net_16691;
wire net_3574;
wire net_22701;
wire net_18796;
wire net_5994;
wire net_10852;
wire net_2921;
wire net_3289;
wire net_8829;
wire net_10225;
wire net_3114;
wire net_3415;
wire net_10019;
wire net_744;
wire net_16430;
wire net_8276;
wire net_15620;
wire net_18430;
wire net_17530;
wire net_7985;
wire net_4136;
wire net_2011;
wire net_19756;
wire net_15023;
wire net_22348;
wire net_777;
wire net_4806;
wire net_13203;
wire net_7185;
wire net_3157;
wire net_7532;
wire net_490;
wire net_18297;
wire net_17746;
wire net_14805;
wire net_11497;
wire net_19529;
wire net_12677;
wire net_18782;
wire net_12130;
wire net_13930;
wire net_6009;
wire net_22184;
wire net_3462;
wire net_20494;
wire net_21151;
wire net_5670;
wire net_4439;
wire net_5602;
wire net_7638;
wire net_2841;
wire net_20274;
wire net_10106;
wire net_19749;
wire net_11889;
wire net_7255;
wire net_5813;
wire net_1977;
wire net_2938;
wire net_14009;
wire net_14568;
wire net_22153;
wire net_1171;
wire net_10691;
wire net_9680;
wire net_248;
wire net_3594;
wire net_20307;
wire net_17989;
wire net_6548;
wire net_5341;
wire net_16995;
wire x5669;
wire net_16562;
wire net_14064;
wire net_13583;
wire net_15268;
wire net_18616;
wire net_18580;
wire net_1767;
wire net_4010;
wire net_21445;
wire net_21148;
wire net_7333;
wire net_11827;
wire net_22441;
wire net_1640;
wire net_12956;
wire net_13788;
wire net_2724;
wire net_11916;
wire net_12090;
wire net_20283;
wire net_15762;
wire net_1741;
wire net_16708;
wire net_10141;
wire net_16163;
wire net_4227;
wire net_20955;
wire net_7550;
wire net_959;
wire net_5381;
wire net_11476;
wire net_7911;
wire net_3051;
wire net_2345;
wire net_6981;
wire net_16643;
wire net_6460;
wire x1651;
wire net_6660;
wire net_2164;
wire net_11079;
wire net_5659;
wire net_11797;
wire net_3751;
wire net_21095;
wire net_19517;
wire net_22024;
wire net_20912;
wire net_5311;
wire net_4564;
wire net_2338;
wire net_15685;
wire net_2616;
wire net_8200;
wire net_282;
wire net_1596;
wire net_17039;
wire net_10804;
wire net_4296;
wire net_11857;
wire net_10908;
wire net_11693;
wire net_2370;
wire net_2047;
wire net_22676;
wire net_8320;
wire net_9647;
wire net_12733;
wire net_2693;
wire net_13115;
wire net_11212;
wire net_16711;
wire net_12765;
wire net_12185;
wire net_9621;
wire net_907;
wire net_18909;
wire net_14473;
wire net_3076;
wire net_16103;
wire net_21908;
wire net_2719;
wire net_6343;
wire net_9688;
wire net_21026;
wire net_16126;
wire net_641;
wire net_2798;
wire net_5071;
wire net_10977;
wire net_3869;
wire net_22650;
wire net_14335;
wire net_1152;
wire net_21799;
wire net_1226;
wire net_14212;
wire net_10525;
wire net_5315;
wire net_15533;
wire net_14976;
wire net_10257;
wire net_3805;
wire x6936;
wire net_19740;
wire net_15865;
wire net_16764;
wire net_3942;
wire net_15823;
wire net_15352;
wire net_7836;
wire net_13199;
wire net_1818;
wire net_12783;
wire net_11850;
wire net_13335;
wire net_8646;
wire net_19426;
wire net_9371;
wire net_17013;
wire net_1523;
wire net_1656;
wire net_17095;
wire net_6522;
wire net_20353;
wire net_16315;
wire net_17558;
wire net_15179;
wire net_691;
wire net_6951;
wire net_5551;
wire net_3178;
wire net_2701;
wire net_17356;
wire net_10422;
wire net_20380;
wire net_1863;
wire net_20479;
wire net_15108;
wire net_19653;
wire net_10774;
wire net_8399;
wire net_2519;
wire net_471;
wire net_18210;
wire net_18000;
wire net_1055;
wire net_3894;
wire net_878;
wire net_518;
wire net_57;
wire net_11136;
wire net_10172;
wire net_14523;
wire net_13533;
wire net_929;
wire net_18853;
wire net_17045;
wire net_2523;
wire net_21489;
wire net_11779;
wire net_4210;
wire net_3954;
wire net_12939;
wire net_11811;
wire net_5726;
wire net_1565;
wire net_5262;
wire net_21109;
wire net_14487;
wire net_169;
wire net_17738;
wire net_15347;
wire net_9948;
wire net_21527;
wire net_16869;
wire net_12986;
wire net_2234;
wire net_16318;
wire net_12120;
wire net_17000;
wire net_15629;
wire net_17727;
wire net_6828;
wire net_10481;
wire net_967;
wire net_19396;
wire net_13056;
wire net_4420;
wire net_21778;
wire net_19633;
wire net_8007;
wire net_13861;
wire net_4318;
wire net_22542;
wire net_12358;
wire net_11475;
wire net_22752;
wire net_4910;
wire net_17172;
wire net_1645;
wire net_2962;
wire net_21292;
wire net_16428;
wire net_4365;
wire net_176;
wire net_19571;
wire net_12410;
wire net_15036;
wire net_614;
wire net_17570;
wire net_21499;
wire net_19343;
wire net_12505;
wire net_22645;
wire net_8293;
wire net_3194;
wire net_3572;
wire net_22832;
wire net_5537;
wire net_4740;
wire net_8338;
wire net_1192;
wire net_10697;
wire net_6857;
wire net_14368;
wire net_4542;
wire net_11753;
wire net_11705;
wire net_15093;
wire net_8730;
wire net_4061;
wire net_12201;
wire net_3156;
wire net_20663;
wire net_12109;
wire net_2482;
wire net_21677;
wire net_13043;
wire net_7275;
wire net_707;
wire net_19362;
wire net_6534;
wire net_21838;
wire net_5039;
wire net_11174;
wire net_6867;
wire net_18038;
wire net_18175;
wire net_4850;
wire net_13828;
wire net_4531;
wire net_14778;
wire net_575;
wire net_5833;
wire net_18184;
wire net_4715;
wire net_7169;
wire net_3697;
wire net_18993;
wire net_20679;
wire net_11374;
wire net_14810;
wire net_12582;
wire net_6193;
wire net_16188;
wire net_15962;
wire net_6431;
wire net_3618;
wire net_19057;
wire net_9156;
wire net_7562;
wire net_15893;
wire net_14012;
wire net_10842;
wire net_16829;
wire net_5512;
wire net_765;
wire net_1342;
wire net_2633;
wire net_1666;
wire net_20036;
wire net_4193;
wire net_15661;
wire net_8573;
wire net_19200;
wire net_8253;
wire net_17249;
wire net_21300;
wire net_2099;
wire net_15390;
wire net_5745;
wire net_6750;
wire net_5182;
wire net_7612;
wire net_18757;
wire net_13454;
wire net_18088;
wire net_16659;
wire net_9809;
wire net_10302;
wire net_22256;
wire net_17679;
wire net_16308;
wire net_16137;
wire net_8195;
wire net_5850;
wire net_5646;
wire net_2021;
wire net_11248;
wire net_1068;
wire net_22508;
wire x3058;
wire net_186;
wire net_2495;
wire net_15229;
wire net_12823;
wire net_6672;
wire net_16803;
wire net_1050;
wire net_17670;
wire net_2760;
wire net_5914;
wire net_21901;
wire net_4751;
wire net_15910;
wire net_2271;
wire net_5327;
wire net_19472;
wire net_21125;
wire net_16036;
wire net_14083;
wire net_18902;
wire net_12164;
wire net_6125;
wire net_7143;
wire net_16014;
wire net_7983;
wire net_10324;
wire net_3130;
wire net_8572;
wire net_15157;
wire net_20688;
wire net_16478;
wire net_17340;
wire net_5704;
wire net_4289;
wire net_9775;
wire net_9510;
wire net_13806;
wire net_4712;
wire net_11340;
wire net_20997;
wire net_260;
wire net_2947;
wire net_15729;
wire net_12552;
wire net_11784;
wire net_3137;
wire net_8649;
wire net_12423;
wire net_20835;
wire net_1597;
wire net_16911;
wire net_7946;
wire net_8785;
wire net_7593;
wire net_3988;
wire net_17056;
wire net_2761;
wire net_19901;
wire net_6396;
wire net_3788;
wire net_22236;
wire net_15605;
wire net_4355;
wire net_21268;
wire net_16007;
wire net_10623;
wire net_1503;
wire net_3961;
wire net_8430;
wire net_4639;
wire net_19302;
wire net_8628;
wire net_11089;
wire net_5494;
wire net_9299;
wire net_17885;
wire net_20788;
wire net_11928;
wire net_9574;
wire net_12638;
wire net_9606;
wire net_12362;
wire net_11409;
wire net_6595;
wire net_13663;
wire net_11653;
wire net_21653;
wire net_13866;
wire net_17362;
wire net_5443;
wire net_5211;
wire net_4731;
wire net_2989;
wire net_497;
wire net_22631;
wire net_6720;
wire net_19281;
wire net_12494;
wire net_7658;
wire net_15291;
wire net_8160;
wire net_1414;
wire net_4153;
wire net_19468;
wire net_11307;
wire net_10927;
wire net_9864;
wire net_300;
wire net_2652;
wire net_5526;
wire net_10149;
wire net_21368;
wire net_20336;
wire net_1233;
wire net_2720;
wire net_6351;
wire net_15058;
wire net_12917;
wire net_1834;
wire net_6027;
wire net_4925;
wire net_17285;
wire net_13213;
wire net_15258;
wire net_13024;
wire net_13313;
wire net_19908;
wire net_15690;
wire net_11355;
wire net_5474;
wire net_14363;
wire net_9745;
wire net_21764;
wire net_8984;
wire net_12565;
wire net_15888;
wire net_13405;
wire net_10203;
wire net_11946;
wire net_21796;
wire net_13603;
wire net_5194;
wire net_12025;
wire net_22725;
wire net_3150;
wire net_9596;
wire net_21116;
wire net_15967;
wire net_20758;
wire net_3979;
wire net_8822;
wire net_21657;
wire net_15927;
wire net_12712;
wire net_839;
wire net_13542;
wire net_11778;
wire net_7095;
wire net_20764;
wire net_18754;
wire net_19094;
wire net_4660;
wire net_21307;
wire net_13013;
wire net_17719;
wire net_18504;
wire net_11294;
wire net_7805;
wire net_19099;
wire net_11313;
wire net_954;
wire net_19848;
wire net_18415;
wire net_22262;
wire net_13094;
wire net_4565;
wire net_9051;
wire net_9037;
wire net_15048;
wire net_8796;
wire net_11271;
wire net_8962;
wire net_10897;
wire net_16957;
wire net_16412;
wire net_10152;
wire net_20606;
wire net_15671;
wire x2298;
wire net_16253;
wire net_19233;
wire net_13359;
wire net_13265;
wire net_14456;
wire net_9545;
wire net_10411;
wire net_18730;
wire net_12445;
wire net_21959;
wire net_11989;
wire net_4790;
wire net_12048;
wire net_17383;
wire net_5363;
wire net_21227;
wire net_7529;
wire net_22124;
wire net_8888;
wire net_6665;
wire net_16921;
wire net_4900;
wire net_9807;
wire net_13222;
wire net_22292;
wire net_6502;
wire net_14888;
wire net_14783;
wire net_7305;
wire net_6163;
wire net_3011;
wire net_17577;
wire net_13079;
wire net_10643;
wire net_18229;
wire net_13187;
wire net_10021;
wire net_19509;
wire net_12946;
wire net_6817;
wire net_6000;
wire net_22605;
wire net_9079;
wire net_8863;
wire net_20188;
wire net_14859;
wire net_11930;
wire net_13628;
wire net_12466;
wire net_9536;
wire net_17592;
wire net_12887;
wire net_3010;
wire net_881;
wire net_12657;
wire net_17877;
wire x296;
wire net_21602;
wire net_10544;
wire net_2805;
wire net_1397;
wire net_14619;
wire net_14231;
wire net_15182;
wire net_4474;
wire net_18373;
wire net_14623;
wire net_17566;
wire net_21549;
wire net_16290;
wire x473;
wire net_1954;
wire net_21395;
wire net_13036;
wire net_7615;
wire x2197;
wire net_22692;
wire net_21633;
wire net_17272;
wire net_14294;
wire net_14924;
wire net_2041;
wire net_17933;
wire net_13090;
wire net_16628;
wire net_11830;
wire net_10354;
wire net_20971;
wire net_21829;
wire net_21803;
wire net_7937;
wire net_18056;
wire net_7930;
wire net_7196;
wire net_16613;
wire net_12197;
wire net_14143;
wire net_2423;
wire net_7535;
wire net_6723;
wire net_20486;
wire net_13875;
wire net_12379;
wire net_11283;
wire net_895;
wire net_10781;
wire net_6412;
wire net_18475;
wire net_14469;
wire net_11603;
wire net_5990;
wire x2035;
wire net_22789;
wire net_14358;
wire net_15202;
wire net_12006;
wire net_8240;
wire net_7048;
wire net_9715;
wire net_7767;
wire net_17683;
wire net_8831;
wire net_12394;
wire net_10683;
wire net_1255;
wire net_12603;
wire net_1250;
wire net_22472;
wire net_8247;
wire net_13928;
wire net_16395;
wire net_15176;
wire net_16937;
wire net_207;
wire net_21542;
wire net_3643;
wire net_18743;
wire net_19045;
wire net_15149;
wire x6571;
wire net_16775;
wire net_13639;
wire net_17782;
wire net_12102;
wire net_13382;
wire net_11874;
wire net_1689;
wire net_10345;
wire net_10271;
wire net_20023;
wire net_6186;
wire net_17783;
wire net_15466;
wire net_8569;
wire net_5698;
wire net_274;
wire net_13987;
wire net_22664;
wire net_1075;
wire net_9387;
wire net_13360;
wire net_6204;
wire net_930;
wire net_2387;
wire net_12599;
wire net_9316;
wire net_8358;
wire net_4723;
wire net_2267;
wire net_21354;
wire net_20736;
wire net_7323;
wire net_4769;
wire net_19382;
wire net_20399;
wire net_18217;
wire net_16740;
wire net_13590;
wire net_10016;
wire net_4888;
wire net_9539;
wire net_18013;
wire net_14636;
wire net_17528;
wire net_21871;
wire net_19008;
wire net_3304;
wire net_15382;
wire net_2549;
wire net_20383;
wire net_11024;
wire net_8654;
wire net_14390;
wire net_3465;
wire net_18658;
wire net_6217;
wire net_637;
wire net_15787;
wire net_13062;
wire net_2390;
wire net_5436;
wire net_2686;
wire net_5577;
wire net_1509;
wire net_529;
wire net_18493;
wire net_9447;
wire net_3495;
wire net_9887;
wire net_2553;
wire net_17548;
wire net_4881;
wire net_19787;
wire net_18113;
wire net_8506;
wire net_6477;
wire net_11303;
wire x844;
wire net_16076;
wire net_121;
wire net_19682;
wire net_5228;
wire net_7475;
wire net_15324;
wire net_16305;
wire net_19613;
wire net_16908;
wire net_9762;
wire net_15579;
wire net_3820;
wire net_3799;
wire net_4175;
wire net_22500;
wire net_19825;
wire net_10938;
wire net_2664;
wire net_18403;
wire net_14206;
wire net_21808;
wire net_11202;
wire net_849;
wire net_14161;
wire net_17563;
wire net_10577;
wire net_7470;
wire net_5294;
wire net_11681;
wire net_14545;
wire net_5751;
wire net_401;
wire net_8165;
wire net_17376;
wire net_10720;
wire net_3798;
wire net_14906;
wire net_2714;
wire net_2183;
wire net_2557;
wire net_14903;
wire net_14265;
wire net_9229;
wire net_11361;
wire net_26;
wire net_758;
wire net_14955;
wire net_13754;
wire net_6874;
wire net_22520;
wire net_14482;
wire net_10846;
wire net_13563;
wire net_7682;
wire x6320;
wire net_21426;
wire net_5504;
wire net_18233;
wire net_15133;
wire net_22152;
wire net_4998;
wire net_19903;
wire net_3255;
wire net_22224;
wire net_12303;
wire net_9848;
wire net_6564;
wire x5903;
wire net_16052;
wire net_15835;
wire net_20751;
wire net_9797;
wire net_12973;
wire net_10946;
wire net_22336;
wire net_20262;
wire net_16098;
wire net_5306;
wire net_9577;
wire net_9938;
wire net_11539;
wire net_16893;
wire net_2917;
wire net_8404;
wire net_15630;
wire net_6711;
wire net_3221;
wire net_16936;
wire net_21212;
wire net_7708;
wire net_605;
wire net_3411;
wire net_4987;
wire net_22280;
wire net_10447;
wire net_17291;
wire net_9233;
wire net_9527;
wire net_924;
wire net_8883;
wire net_12255;
wire net_17323;
wire net_5469;
wire net_9205;
wire net_10980;
wire net_16444;
wire net_7829;
wire net_2348;
wire net_489;
wire net_21525;
wire net_14911;
wire net_21366;
wire net_17476;
wire net_5457;
wire net_21930;
wire net_6143;
wire net_4646;
wire net_18774;
wire net_2748;
wire net_9991;
wire net_18150;
wire net_11561;
wire net_9611;
wire net_19645;
wire net_9135;
wire net_8060;
wire net_251;
wire net_15772;
wire net_21666;
wire net_840;
wire net_9206;
wire net_10632;
wire net_8086;
wire net_17845;
wire net_6933;
wire net_20466;
wire net_15429;
wire net_5789;
wire net_20269;
wire net_13281;
wire net_12928;
wire net_11229;
wire net_9914;
wire net_411;
wire net_2137;
wire net_20346;
wire net_22289;
wire net_11689;
wire net_15075;
wire net_12220;
wire net_11256;
wire net_12688;
wire net_20061;
wire net_7874;
wire net_7293;
wire net_22144;
wire net_8975;
wire net_1862;
wire net_13889;
wire net_10052;
wire net_2317;
wire net_6248;
wire net_16118;
wire net_8135;
wire net_16885;
wire net_10584;
wire net_6035;
wire net_6492;
wire net_3583;
wire net_112;
wire net_21088;
wire net_8183;
wire net_19030;
wire net_10536;
wire net_8219;
wire net_15802;
wire net_2373;
wire net_11694;
wire net_14109;
wire net_19598;
wire net_20902;
wire net_17310;
wire net_19813;
wire net_16332;
wire net_10943;
wire net_7746;
wire net_9282;
wire net_15137;
wire net_1609;
wire net_402;
wire net_7847;
wire net_4047;
wire net_3448;
wire net_22534;
wire net_21761;
wire net_7108;
wire net_33;
wire net_3248;
wire net_12450;
wire net_2274;
wire net_11597;
wire net_22283;
wire net_12681;
wire net_17602;
wire net_11488;
wire net_13859;
wire net_10950;
wire net_19984;
wire net_18842;
wire net_12345;
wire net_2359;
wire net_16835;
wire net_21887;
wire net_20649;
wire net_15038;
wire net_16701;
wire net_13101;
wire net_12574;
wire net_15432;
wire net_11585;
wire net_16473;
wire net_10127;
wire net_4102;
wire net_6908;
wire net_1430;
wire net_22737;
wire net_9964;
wire net_6892;
wire net_21465;
wire net_2478;
wire net_6429;
wire net_2563;
wire net_18040;
wire net_12435;
wire net_9484;
wire net_9243;
wire net_8051;
wire net_5679;
wire net_16729;
wire net_3408;
wire net_4870;
wire net_630;
wire net_76;
wire net_12514;
wire net_2202;
wire x71;
wire net_2490;
wire net_8841;
wire net_14861;
wire net_4428;
wire net_1791;
wire net_4339;
wire net_1471;
wire net_9975;
wire net_8997;
wire net_7667;
wire net_3608;
wire net_18079;
wire net_17088;
wire net_16602;
wire net_14892;
wire net_912;
wire net_17034;
wire net_20907;
wire net_19112;
wire net_13562;
wire net_7018;
wire net_4517;
wire net_15315;
wire x5188;
wire net_3841;
wire net_1928;
wire net_1328;
wire net_22435;
wire net_9871;
wire net_16458;
wire net_2859;
wire net_3848;
wire net_2884;
wire net_20719;
wire net_5372;
wire net_4942;
wire net_13616;
wire x2554;
wire net_3205;
wire net_22429;
wire net_1094;
wire net_3487;
wire net_2749;
wire net_855;
wire net_674;
wire net_18935;
wire net_19926;
wire net_11032;
wire net_9506;
wire net_303;
wire net_10041;
wire net_21332;
wire net_15821;
wire net_18647;
wire net_9982;
wire net_2475;
wire net_9925;
wire net_18328;
wire net_2937;
wire net_7792;
wire net_7657;
wire net_7400;
wire net_6191;
wire net_21442;
wire net_17168;
wire net_14744;
wire net_12249;
wire net_16746;
wire net_12993;
wire net_7865;
wire net_4743;
wire net_20003;
wire net_13767;
wire net_17960;
wire net_9478;
wire net_2439;
wire net_13297;
wire net_19504;
wire net_11048;
wire net_172;
wire net_4341;
wire net_13460;
wire net_15300;
wire x4781;
wire net_4048;
wire net_17234;
wire net_16962;
wire net_10749;
wire net_4570;
wire net_17832;
wire net_16284;
wire net_10244;
wire net_18449;
wire net_6689;
wire net_22384;
wire net_12233;
wire net_13934;
wire net_7034;
wire net_6446;
wire net_8029;
wire net_11939;
wire net_9050;
wire net_6198;
wire net_3733;
wire net_19365;
wire net_3881;
wire net_12263;
wire net_8598;
wire net_11944;
wire net_10519;
wire net_20512;
wire net_14136;
wire net_15481;
wire net_8091;
wire net_8057;
wire net_6258;
wire net_8361;
wire net_19512;
wire net_1758;
wire net_13840;
wire net_8813;
wire net_18571;
wire net_16549;
wire net_14868;
wire net_11802;
wire net_1769;
wire net_9115;
wire net_6694;
wire net_15504;
wire net_1567;
wire net_17940;
wire net_8020;
wire net_6322;
wire net_12087;
wire net_15286;
wire net_11186;
wire net_8152;
wire net_18193;
wire net_9520;
wire net_19286;
wire net_22479;
wire net_14930;
wire net_476;
wire net_2783;
wire net_17513;
wire net_14461;
wire net_6055;
wire net_7079;
wire net_382;
wire net_11412;
wire net_11259;
wire net_5301;
wire net_583;
wire net_7041;
wire net_16987;
wire net_15947;
wire net_9408;
wire net_17996;
wire net_14173;
wire net_16734;
wire net_17967;
wire net_13055;
wire net_9695;
wire net_4719;
wire net_17071;
wire net_10379;
wire net_19712;
wire net_17827;
wire net_15234;
wire net_9005;
wire net_4460;
wire net_220;
wire net_1465;
wire net_11153;
wire net_13599;
wire net_4982;
wire net_16407;
wire net_543;
wire net_625;
wire net_22401;
wire net_3760;
wire net_17469;
wire net_16944;
wire net_11411;
wire net_10708;
wire net_21219;
wire net_17796;
wire net_20445;
wire net_15543;
wire net_17506;
wire net_11637;
wire net_21386;
wire net_14509;
wire net_13790;
wire net_4331;
wire net_2909;
wire net_4953;
wire net_15464;
wire net_9607;
wire net_21486;
wire net_20519;
wire net_4697;
wire net_5638;
wire net_7899;
wire net_19278;
wire net_15594;
wire net_12157;
wire net_10562;
wire net_20406;
wire net_1694;
wire net_12844;
wire net_4991;
wire net_910;
wire net_15940;
wire net_12356;
wire net_15332;
wire net_18514;
wire net_5394;
wire net_21744;
wire net_7944;
wire net_2412;
wire net_16247;
wire net_12070;
wire net_4265;
wire net_18717;
wire net_14563;
wire net_4158;
wire net_13442;
wire net_17078;
wire net_13527;
wire net_315;
wire net_1375;
wire net_18411;
wire net_4006;
wire net_16969;
wire net_8212;
wire net_1351;
wire net_17455;
wire net_18673;
wire net_1535;
wire net_16859;
wire net_2400;
wire net_5543;
wire net_18261;
wire net_8661;
wire net_10959;
wire net_2034;
wire net_15189;
wire net_14963;
wire net_8921;
wire net_1808;
wire net_3256;
wire net_22402;
wire net_13122;
wire net_18164;
wire net_20768;
wire net_15003;
wire net_14916;
wire net_13438;
wire net_10567;
wire x5853;
wire net_3322;
wire net_2533;
wire net_10267;
wire net_1913;
wire net_12297;
wire net_16024;
wire net_13243;
wire net_11526;
wire net_7830;
wire net_20394;
wire net_16413;
wire net_9673;
wire net_9016;
wire net_7642;
wire net_20791;
wire net_11904;
wire net_9732;
wire net_9264;
wire net_15244;
wire net_6615;
wire net_12279;
wire net_7409;
wire net_7671;
wire net_1760;
wire net_7714;
wire net_3926;
wire net_4849;
wire net_5758;
wire net_3403;
wire net_10002;
wire net_21265;
wire net_6977;
wire net_10718;
wire net_3093;
wire net_7935;
wire net_12820;
wire net_6886;
wire net_647;
wire net_3247;
wire net_20978;
wire net_15745;
wire x6350;
wire net_19820;
wire net_17975;
wire net_18962;
wire net_6452;
wire net_8684;
wire net_2464;
wire net_12272;
wire net_9492;
wire net_3839;
wire net_6513;
wire net_17722;
wire net_17349;
wire net_2732;
wire net_21420;
wire net_13483;
wire net_11809;
wire net_8368;
wire net_7345;
wire net_19719;
wire net_1096;
wire net_21405;
wire net_795;
wire net_8153;
wire net_18425;
wire net_11403;
wire net_1406;
wire net_9093;
wire net_22037;
wire net_15754;
wire net_19535;
wire net_18965;
wire net_8490;
wire net_18986;
wire net_10463;
wire net_1434;
wire net_22803;
wire net_6996;
wire net_3668;
wire net_19601;
wire net_14728;
wire net_6096;
wire net_21648;
wire net_9823;
wire net_10012;
wire net_5130;
wire net_11870;
wire net_5617;
wire net_21593;
wire net_4946;
wire net_20727;
wire net_774;
wire net_15101;
wire net_18804;
wire net_10071;
wire net_6958;
wire net_20807;
wire net_8892;
wire net_13235;
wire net_7221;
wire net_501;
wire net_21239;
wire x2077;
wire net_3679;
wire net_4489;
wire net_12344;
wire net_5818;
wire net_20052;
wire net_21019;
wire net_20806;
wire net_6213;
wire net_4692;
wire net_9769;
wire net_6644;
wire net_20357;
wire net_7481;
wire net_9170;
wire net_13327;
wire net_447;
wire net_19893;
wire net_9180;
wire net_19830;
wire net_15126;
wire net_13279;
wire net_5772;
wire net_6318;
wire net_11219;
wire net_19391;
wire net_14031;
wire net_10755;
wire net_16590;
wire net_13371;
wire net_9703;
wire net_22072;
wire net_12368;
wire net_8952;
wire net_20438;
wire net_13944;
wire net_10923;
wire net_19582;
wire net_7900;
wire net_18563;
wire net_14038;
wire net_4106;
wire net_2951;
wire net_8621;
wire net_3631;
wire net_12854;
wire net_18707;
wire net_2293;
wire net_20177;
wire net_16681;
wire net_10105;
wire net_1802;
wire x107;
wire net_15100;
wire net_7694;
wire net_5482;
wire net_22655;
wire net_19147;
wire net_10456;
wire net_7637;
wire net_11318;
wire net_18045;
wire net_20610;
wire net_2755;
wire net_12172;
wire net_21694;
wire x683;
wire net_13850;
wire net_1678;
wire net_21067;
wire net_46;
wire net_14997;
wire net_6638;
wire net_3366;
wire net_10210;
wire net_15338;
wire net_19587;
wire net_18628;
wire net_21277;
wire net_8271;
wire net_7737;
wire net_7206;
wire net_22614;
wire net_6757;
wire net_17656;
wire net_8511;
wire net_7757;
wire net_11726;
wire net_15442;
wire net_21532;
wire net_10934;
wire net_3436;
wire net_18069;
wire net_18136;
wire net_14159;
wire net_15500;
wire net_21261;
wire net_10812;
wire net_8708;
wire net_19638;
wire net_7725;
wire net_3911;
wire net_17441;
wire net_13913;
wire net_12866;
wire net_5337;
wire net_22596;
wire net_15557;
wire net_8638;
wire net_17929;
wire net_3365;
wire net_10711;
wire net_18390;
wire net_14372;
wire net_14099;
wire net_12698;
wire net_8587;
wire net_1114;
wire net_10619;
wire net_13431;
wire net_7090;
wire net_3388;
wire net_10664;
wire net_4116;
wire net_3218;
wire net_18386;
wire net_13005;
wire net_21773;
wire net_4632;
wire net_20516;
wire net_12283;
wire net_18525;
wire net_8171;
wire net_7266;
wire net_6738;
wire net_18700;
wire net_6690;
wire net_6565;
wire net_18559;
wire net_3811;
wire net_19839;
wire net_1028;
wire net_14287;
wire net_1529;
wire net_600;
wire net_14021;
wire net_397;
wire net_11126;
wire net_7602;
wire net_5595;
wire net_19876;
wire net_10968;
wire net_9894;
wire net_12373;
wire net_1384;
wire net_17518;
wire net_17181;
wire net_8712;
wire net_3918;
wire net_9107;
wire net_5280;
wire net_320;
wire net_6844;
wire net_16240;
wire net_4916;
wire net_6902;
wire net_15211;
wire net_9251;
wire net_9103;
wire net_12530;
wire net_7063;
wire net_21220;
wire net_19379;
wire net_986;
wire net_1242;
wire net_15980;
wire net_6556;
wire net_4346;
wire net_1241;
wire net_15571;
wire net_13153;
wire net_11953;
wire net_3690;
wire net_15584;
wire net_20974;
wire net_7524;
wire net_11833;
wire net_11019;
wire net_21399;
wire net_13998;
wire net_13197;
wire net_19104;
wire net_17581;
wire net_3001;
wire net_3121;
wire net_10368;
wire net_4841;
wire net_4621;
wire net_10289;
wire net_10217;
wire net_1634;
wire net_10305;
wire net_6271;
wire net_609;
wire net_12034;
wire net_13343;
wire net_19869;
wire net_19175;
wire net_22639;
wire net_6155;
wire net_3083;
wire net_5693;
wire net_17612;
wire net_9782;
wire net_1221;
wire net_15419;
wire net_7158;
wire net_6911;
wire net_4895;
wire net_20130;
wire net_9851;
wire x887;
wire net_14943;
wire net_816;
wire net_16005;
wire net_16082;
wire net_9100;
wire net_3264;
wire net_7363;
wire net_2092;
wire net_16872;
wire net_13209;
wire net_7134;
wire net_12745;
wire net_8669;
wire net_18230;
wire net_21867;
wire net_1217;
wire net_13879;
wire net_7028;
wire net_22795;
wire net_9719;
wire net_2933;
wire net_8141;
wire net_3381;
wire net_10818;
wire net_16344;
wire net_14156;
wire net_8848;
wire net_18895;
wire net_4118;
wire net_4577;
wire net_22326;
wire net_17913;
wire net_4970;
wire net_20572;
wire net_1575;
wire net_17821;
wire net_3279;
wire net_657;
wire net_8495;
wire net_5042;
wire net_1727;
wire net_17644;
wire net_16367;
wire net_329;
wire net_16757;
wire net_5809;
wire net_4600;
wire net_21611;
wire net_14633;
wire net_12848;
wire net_1924;
wire net_4287;
wire net_1825;
wire net_3168;
wire x445;
wire net_16674;
wire net_10078;
wire net_14714;
wire net_10558;
wire net_962;
wire net_7914;
wire net_8695;
wire net_13731;
wire net_7817;
wire net_596;
wire net_11840;
wire net_1261;
wire net_22125;
wire net_20887;
wire net_2120;
wire net_15081;
wire net_4705;
wire net_10430;
wire net_14167;
wire net_7566;
wire net_14735;
wire net_13512;
wire net_18657;
wire net_20666;
wire net_12893;
wire net_565;
wire net_2569;
wire net_21281;
wire net_2832;
wire net_21339;
wire net_4478;
wire net_2149;
wire net_18904;
wire net_13174;
wire net_9736;
wire net_22332;
wire net_15654;
wire net_10611;
wire net_17304;
wire net_10363;
wire net_16785;
wire net_5062;
wire net_6518;
wire net_4236;
wire net_19243;
wire net_11618;
wire net_19593;
wire net_17772;
wire net_22197;
wire net_18372;
wire net_4813;
wire net_21205;
wire net_14679;
wire net_10986;
wire net_232;
wire net_21643;
wire net_16260;
wire net_6538;
wire net_14273;
wire net_18787;
wire net_21438;
wire net_21052;
wire net_12778;
wire net_2167;
wire net_2880;
wire net_20317;
wire net_16350;
wire net_15408;
wire net_7923;
wire net_11062;
wire net_2996;
wire x3290;
wire net_20080;
wire net_6386;
wire net_15147;
wire net_4465;
wire net_532;
wire net_2501;
wire net_3530;
wire net_13179;
wire net_21623;
wire net_20695;
wire net_19483;
wire net_14751;
wire net_14817;
wire net_18516;
wire net_8223;
wire net_889;
wire net_12609;
wire net_1116;
wire net_20170;
wire net_21288;
wire net_13018;
wire net_16879;
wire net_5253;
wire net_17542;
wire net_4373;
wire net_13135;
wire net_9289;
wire net_17498;
wire net_18832;
wire net_11521;
wire net_2814;
wire net_689;
wire net_751;
wire net_16294;
wire net_15172;
wire net_15222;
wire net_22159;
wire net_14670;
wire net_2363;
wire x2547;
wire net_22820;
wire net_14346;
wire net_15882;
wire net_3659;
wire net_6578;
wire net_5232;
wire net_13708;
wire net_10512;
wire net_20588;
wire net_3724;
wire net_13129;
wire net_16556;
wire net_16174;
wire net_4593;
wire net_20891;
wire net_15615;
wire net_15561;
wire net_20943;
wire net_1426;
wire net_20821;
wire net_12649;
wire net_11111;
wire net_9813;
wire net_1407;
wire net_3147;
wire net_4903;
wire net_15343;
wire net_5409;
wire net_12949;
wire net_16043;
wire net_3263;
wire net_20196;
wire net_10093;
wire net_21575;
wire net_14610;
wire net_20877;
wire net_16941;
wire net_14129;
wire net_19862;
wire net_17137;
wire net_4931;
wire net_16548;
wire net_17715;
wire net_22369;
wire net_10509;
wire net_7261;
wire net_8613;
wire net_8233;
wire net_6189;
wire net_22176;
wire net_5114;
wire net_15920;
wire net_4398;
wire net_1042;
wire net_4783;
wire net_4076;
wire net_15703;
wire net_7788;
wire net_17409;
wire net_19458;
wire net_1000;
wire net_21323;
wire net_1995;
wire net_17208;
wire net_2545;
wire net_20767;
wire net_18979;
wire net_5158;
wire net_17751;
wire net_2870;
wire net_14769;
wire net_18358;
wire net_22671;
wire net_6182;
wire net_20526;
wire net_22097;
wire net_4320;
wire net_11847;
wire net_2596;
wire net_10835;
wire net_2970;
wire net_14388;
wire net_12369;
wire net_18117;
wire net_14001;
wire net_9001;
wire net_2584;
wire net_16279;
wire net_14052;
wire net_20310;
wire net_17764;
wire net_18099;
wire net_22374;
wire net_20156;
wire net_18451;
wire net_7546;
wire net_11963;
wire net_952;
wire net_14305;
wire net_4097;
wire net_11743;
wire net_5170;
wire net_3185;
wire net_19025;
wire net_17433;
wire net_13821;
wire net_14290;
wire net_9048;
wire net_3300;
wire net_19952;
wire net_86;
wire net_21945;
wire net_6438;
wire net_2245;
wire net_20755;
wire net_22115;
wire net_7268;
wire net_21629;
wire net_12963;
wire net_8187;
wire net_7570;
wire net_13773;
wire net_4231;
wire net_383;
wire net_4068;
wire net_20098;
wire net_14055;
wire net_3140;
wire net_15625;
wire net_6765;
wire net_18500;
wire net_16203;
wire net_427;
wire net_7823;
wire net_135;
wire net_22030;
wire net_1121;
wire x7413;
wire net_21187;
wire net_18123;
wire net_22046;
wire net_19222;
wire net_13687;
wire net_7288;
wire net_13897;
wire net_7559;
wire net_18809;
wire net_7381;
wire net_21094;
wire net_4329;
wire net_16904;
wire net_11094;
wire net_6409;
wire net_2777;
wire net_17464;
wire net_1049;
wire net_13531;
wire net_9440;
wire net_3901;
wire net_17867;
wire net_21927;
wire net_10674;
wire net_18693;
wire net_14674;
wire net_9364;
wire net_6707;
wire net_8437;
wire net_9278;
wire net_7582;
wire net_6229;
wire net_8608;
wire net_5199;
wire net_21460;
wire net_12905;
wire net_19577;
wire net_19544;
wire net_12388;
wire net_9293;
wire net_18739;
wire net_2591;
wire net_14534;
wire net_10552;
wire net_8985;
wire net_22762;
wire net_10880;
wire net_17789;
wire net_5189;
wire net_11896;
wire net_5791;
wire net_3968;
wire net_1283;
wire net_16652;
wire net_22550;
wire net_12875;
wire net_4554;
wire net_18885;
wire net_354;
wire net_19663;
wire net_14607;
wire net_17067;
wire net_12428;
wire net_21670;
wire net_15001;
wire net_16267;
wire net_21584;
wire net_15973;
wire net_18017;
wire net_12099;
wire net_3356;
wire net_11423;
wire net_7175;
wire net_5465;
wire net_12640;
wire net_21469;
wire net_3886;
wire net_7281;
wire net_22172;
wire net_1592;
wire net_21848;
wire net_13650;
wire net_2085;
wire net_4406;
wire net_17416;
wire net_16668;
wire net_12557;
wire net_5621;
wire net_15425;
wire net_8764;
wire net_10297;
wire net_1637;
wire net_3702;
wire net_9374;
wire net_6480;
wire net_6425;
wire net_5971;
wire net_19620;
wire net_6220;
wire net_16639;
wire net_8915;
wire net_7629;
wire net_18315;
wire net_11324;
wire net_5854;
wire net_14519;
wire net_4555;
wire net_2070;
wire net_11661;
wire net_16389;
wire net_10605;
wire net_4124;
wire net_16191;
wire net_18934;
wire net_16698;
wire net_12372;
wire net_3981;
wire net_13659;
wire net_3161;
wire net_6107;
wire net_4303;
wire net_1290;
wire net_12924;
wire net_4147;
wire net_22309;
wire net_21833;
wire net_21413;
wire net_4056;
wire net_21736;
wire net_17337;
wire net_12589;
wire net_3297;
wire net_14028;
wire net_11766;
wire net_5249;
wire net_13474;
wire net_12205;
wire net_3424;
wire net_18941;
wire net_15371;
wire net_6364;
wire net_22238;
wire net_21859;
wire net_10169;
wire net_5087;
wire net_13218;
wire net_11983;
wire net_15397;
wire net_3104;
wire net_5508;
wire net_15066;
wire net_2278;
wire net_3072;
wire net_15409;
wire net_7286;
wire net_1021;
wire net_18680;
wire net_19477;
wire net_10498;
wire net_5269;
wire net_10488;
wire net_1737;
wire net_9979;
wire net_16375;
wire net_10657;
wire net_6801;
wire net_21012;
wire net_3607;
wire net_4654;
wire net_8541;
wire net_20781;
wire net_4917;
wire net_1145;
wire net_8424;
wire net_9306;
wire net_2261;
wire net_9411;
wire net_18949;
wire net_3061;
wire net_19063;
wire net_7414;
wire net_21023;
wire net_2958;
wire net_21890;
wire net_11328;
wire net_20222;
wire net_14131;
wire net_5918;
wire net_18105;
wire net_10827;
wire net_19999;
wire net_119;
wire net_22005;
wire net_15869;
wire net_22080;
wire net_16069;
wire net_6853;
wire net_13961;
wire net_13624;
wire net_21780;
wire net_6307;
wire net_4192;
wire net_21704;
wire net_11977;
wire net_14586;
wire net_17330;
wire net_11733;
wire net_11141;
wire net_11568;
wire net_90;
wire net_4583;
wire net_20377;
wire net_22518;
wire net_18488;
wire net_18222;
wire net_12290;
wire net_4663;
wire net_21166;
wire net_14330;
wire net_19552;
wire net_5822;
wire net_4084;
wire net_4500;
wire net_8045;
wire net_20128;
wire net_15351;
wire net_8591;
wire net_5879;
wire net_14250;
wire net_15812;
wire net_8562;
wire net_2056;
wire net_5716;
wire net_17293;
wire net_7884;
wire net_12217;
wire net_10800;
wire net_9147;
wire net_1628;
wire net_3476;
wire net_15162;
wire net_13957;
wire net_7347;
wire net_4823;
wire net_12519;
wire net_2512;
wire net_12997;
wire net_1936;
wire net_3802;
wire net_14749;
wire net_21390;
wire net_18219;
wire net_10035;
wire net_14339;
wire net_126;
wire net_2708;
wire net_8773;
wire net_8705;
wire net_18996;
wire net_17523;
wire net_10873;
wire net_9958;
wire net_2211;
wire net_19725;
wire net_18279;
wire net_7425;
wire net_21609;
wire net_5479;
wire net_16050;
wire net_13001;
wire net_20540;
wire net_14090;
wire net_8388;
wire net_8777;
wire net_19387;
wire net_9998;
wire net_1732;
wire net_5926;
wire net_7866;
wire net_6348;
wire net_21905;
wire net_18485;
wire net_9390;
wire net_12149;
wire net_20814;
wire net_900;
wire net_19734;
wire net_7597;
wire net_19125;
wire net_21273;
wire net_5528;
wire net_2001;
wire net_1491;
wire net_10879;
wire net_14442;
wire net_8306;
wire net_10918;
wire net_5390;
wire net_20552;
wire net_18527;
wire net_1034;
wire net_11559;
wire x205;
wire net_16218;
wire net_15634;
wire net_11510;
wire net_17758;
wire net_21774;
wire net_17437;
wire net_3439;
wire net_20327;
wire net_18323;
wire net_13332;
wire x304;
wire net_18159;
wire net_11398;
wire net_1959;
wire net_21344;
wire net_20081;
wire net_18212;
wire net_15372;
wire net_11506;
wire net_12320;
wire net_14884;
wire net_21223;
wire net_17667;
wire net_19156;
wire net_460;
wire net_7356;
wire net_6797;
wire net_6074;
wire net_4206;
wire net_16983;
wire net_15566;
wire net_15365;
wire net_20417;
wire net_1133;
wire net_15797;
wire net_14788;
wire net_14222;
wire net_6131;
wire net_17062;
wire net_11712;
wire net_10724;
wire net_166;
wire net_14429;
wire net_11027;
wire net_21143;
wire net_13954;
wire net_5489;
wire net_13164;
wire net_3871;
wire net_18915;
wire net_4455;
wire net_10995;
wire net_8788;
wire net_3352;
wire net_18634;
wire net_7507;
wire net_3832;
wire net_17119;
wire net_5663;
wire net_6017;
wire net_10062;
wire net_20627;
wire net_17688;
wire net_6925;
wire net_334;
wire net_10930;
wire net_2453;
wire net_3062;
wire net_19640;
wire net_9586;
wire net_5738;
wire net_12629;
wire net_22193;
wire net_10952;
wire net_13797;
wire net_16539;
wire net_18364;
wire net_12626;
wire net_14042;
wire net_6790;
wire net_3768;
wire net_2286;
wire net_16716;
wire net_1552;
wire net_13785;
wire net_9380;
wire net_14833;
wire net_14015;
wire net_17556;
wire net_20681;
wire net_14539;
wire net_22511;
wire net_5674;
wire net_14532;
wire net_14591;
wire net_7954;
wire net_3215;
wire net_3717;
wire net_298;
wire net_1933;
wire net_20927;
wire net_998;
wire net_12620;
wire net_4657;
wire net_2157;
wire net_8945;
wire net_15491;
wire net_10317;
wire net_11154;
wire net_13148;
wire net_12457;
wire net_9328;
wire net_19946;
wire net_13763;
wire x5360;
wire net_14194;
wire net_2405;
wire net_14929;
wire net_835;
wire net_21822;
wire net_7459;
wire net_15381;
wire net_18592;
wire net_13683;
wire net_9321;
wire net_19227;
wire net_10466;
wire net_20603;
wire net_6459;
wire net_17905;
wire net_14795;
wire net_638;
wire net_20761;
wire x763;
wire net_17916;
wire net_5633;
wire net_18978;
wire net_10028;
wire net_5766;
wire net_11519;
wire net_12801;
wire net_19974;
wire net_1783;
wire net_22460;
wire net_7771;
wire net_1874;
wire net_9554;
wire net_14948;
wire net_19431;
wire net_14308;
wire net_17251;
wire net_22106;
wire net_14447;
wire net_3499;
wire net_5206;
wire net_4777;
wire net_17972;
wire net_13192;
wire net_14108;
wire net_12808;
wire net_785;
wire net_9152;
wire net_16490;
wire net_21376;
wire net_20078;
wire net_5883;
wire x6203;
wire net_4215;
wire net_17920;
wire net_9874;
wire net_6677;
wire net_10902;
wire net_13633;
wire net_10409;
wire net_9657;
wire net_20853;
wire net_7479;
wire net_3746;
wire net_1349;
wire net_19626;
wire net_979;
wire net_19151;
wire net_156;
wire net_13251;
wire net_11820;
wire net_12563;
wire net_2015;
wire net_6658;
wire net_19934;
wire net_9676;
wire net_5202;
wire net_4877;
wire net_4170;
wire net_3101;
wire net_12336;
wire net_6268;
wire net_12723;
wire net_20320;
wire net_21078;
wire net_20432;
wire net_3876;
wire net_16576;
wire net_5982;
wire net_22120;
wire net_1887;
wire net_13146;
wire net_7444;
wire net_5470;
wire net_14851;
wire net_4033;
wire net_4245;
wire net_11868;
wire net_9514;
wire net_5568;
wire net_3047;
wire net_16792;
wire net_8910;
wire net_9532;
wire net_6944;
wire net_22585;
wire net_6883;
wire net_2657;
wire net_15119;
wire x329;
wire net_12259;
wire net_11438;
wire net_20779;
wire net_14696;
wire net_8415;
wire net_20838;
wire net_7742;
wire net_2629;
wire net_2486;
wire net_20456;
wire net_15196;
wire net_7117;
wire x277;
wire net_16235;
wire net_1206;
wire net_8381;
wire net_3653;
wire net_13494;
wire x2531;
wire net_1166;
wire net_22063;
wire net_17958;
wire net_18241;
wire net_10765;
wire net_801;
wire net_2620;
wire net_7450;
wire net_1718;
wire net_2581;
wire net_20111;
wire net_18318;
wire net_5093;
wire net_9417;
wire net_7372;
wire net_11921;
wire net_10391;
wire net_15612;
wire net_8482;
wire net_2129;
wire net_21170;
wire net_19735;
wire net_5968;
wire net_18131;
wire net_6234;
wire net_15112;
wire net_18896;
wire net_9833;
wire net_16156;
wire net_8856;
wire net_11382;
wire net_21408;
wire net_7115;
wire net_5906;
wire net_11391;
wire net_8462;
wire net_16797;
wire net_17412;
wire net_2325;
wire net_8807;
wire net_19560;
wire net_19011;
wire net_22456;
wire net_13715;
wire net_806;
wire x6680;
wire net_11907;
wire net_9901;
wire net_21475;
wire net_16159;
wire net_21516;
wire net_18829;
wire net_18398;
wire net_16814;
wire net_8940;
wire net_4021;
wire net_22490;
wire net_17593;
wire net_10960;
wire net_946;
wire net_17156;
wire net_22406;
wire net_2194;
wire net_21752;
wire net_5010;
wire net_3559;
wire net_8370;
wire net_4682;
wire net_15261;
wire net_10114;
wire net_19551;
wire net_20772;
wire net_10402;
wire net_20400;
wire net_12499;
wire net_10732;
wire net_3564;
wire net_1448;
wire net_21079;
wire net_392;
wire net_20986;
wire net_5683;
wire net_7003;
wire net_2452;
wire net_11463;
wire net_19144;
wire net_10336;
wire net_3523;
wire net_4162;
wire net_17651;
wire net_5549;
wire net_3712;
wire net_21130;
wire net_6680;
wire x3771;
wire net_16299;
wire net_17814;
wire net_1186;
wire net_22083;
wire net_4747;
wire net_14829;
wire net_7074;
wire net_17263;
wire net_10607;
wire net_10437;
wire net_2216;
wire net_10410;
wire net_16522;
wire net_7399;
wire net_3773;
wire net_1773;
wire net_9057;
wire net_21999;
wire net_8731;
wire net_21505;
wire net_18618;
wire net_19329;
wire net_19118;
wire net_19558;
wire net_22834;
wire net_17619;
wire net_5073;
wire net_4452;
wire net_20426;
wire net_2447;
wire net_22744;
wire net_7433;
wire net_14116;
wire net_5417;
wire net_15237;
wire net_8137;
wire net_14643;
wire net_17451;
wire net_182;
wire net_4359;
wire net_19412;
wire net_14506;
wire net_11260;
wire net_21032;
wire net_19079;
wire net_9547;
wire net_18051;
wire net_14872;
wire net_14237;
wire net_16581;
wire net_11442;
wire net_1435;
wire net_1370;
wire net_9462;
wire net_3568;
wire net_4482;
wire net_6470;
wire net_19037;
wire net_8459;
wire net_1970;
wire net_1306;
wire net_1858;
wire net_19563;
wire net_14551;
wire x55;
wire net_14846;
wire net_11332;
wire net_22801;
wire net_20236;
wire net_11196;
wire net_12242;
wire net_791;
wire net_20032;
wire net_14207;
wire net_9422;
wire net_1419;
wire net_3239;
wire net_8554;
wire net_2188;
wire net_17864;
wire net_20930;
wire net_12064;
wire net_13882;
wire net_19324;
wire x2042;
wire net_21673;
wire net_20225;
wire net_17124;
wire net_20849;
wire net_17622;
wire net_14841;
wire net_7410;
wire net_12471;
wire net_7219;
wire net_13272;
wire net_19918;
wire net_6824;
wire net_14651;
wire net_361;
wire net_2890;
wire net_11547;
wire net_20474;
wire net_16991;
wire net_1905;
wire net_19126;
wire net_2540;
wire net_20593;
wire net_2230;
wire x598;
wire net_144;
wire net_227;
wire net_22467;
wire net_13758;
wire net_4183;
wire net_18368;
wire net_10237;
wire net_16788;
wire net_14664;
wire net_3592;
wire net_19072;
wire net_5961;
wire net_13728;
wire net_12543;
wire x233;
wire net_7156;
wire net_14413;
wire net_12636;
wire net_4969;
wire net_18926;
wire net_16817;
wire net_1415;
wire net_7052;
wire net_8859;
wire net_6379;
wire net_3317;
wire net_22790;
wire net_11746;
wire net_8140;
wire net_14934;
wire net_18531;
wire net_18162;
wire net_11638;
wire net_9161;
wire net_10120;
wire net_11910;
wire net_1230;
wire net_18126;
wire net_6047;
wire net_15418;
wire net_20710;
wire net_22096;
wire net_6862;
wire net_6064;
wire net_18204;
wire net_16850;
wire net_15455;
wire net_15317;
wire net_20535;
wire net_20865;
wire net_18577;
wire net_12046;
wire net_7585;
wire net_22002;
wire net_22310;
wire net_10597;
wire net_18138;
wire net_2039;
wire net_11579;
wire net_12067;
wire net_1456;
wire net_9198;
wire net_2227;
wire net_20876;
wire net_16822;
wire net_10280;
wire net_8876;
wire net_20707;
wire net_6968;
wire net_22048;
wire net_11041;
wire net_19780;
wire net_13509;
wire net_13844;
wire net_8752;
wire net_11209;
wire net_218;
wire net_12338;
wire net_16975;
wire net_7110;
wire net_22829;
wire net_9335;
wire net_5173;
wire net_1273;
wire net_3283;
wire net_20046;
wire net_18863;
wire net_9025;
wire net_4433;
wire net_17023;
wire net_13907;
wire net_11995;
wire net_2114;
wire net_2506;
wire net_22528;
wire net_5012;
wire net_9644;
wire net_16183;
wire net_7124;
wire net_18172;
wire net_11235;
wire net_21137;
wire net_11990;
wire net_21682;
wire net_16060;
wire net_14073;
wire net_285;
wire net_18078;
wire x1603;
wire net_2499;
wire net_11567;
wire net_1297;
wire net_18822;
wire net_8901;
wire net_2177;
wire net_6581;
wire x726;
wire net_6916;
wire net_16322;
wire net_18381;
wire net_17840;
wire net_5030;
wire net_19881;
wire net_1317;
wire net_215;
wire net_2394;
wire net_1382;
wire net_11593;
wire net_13408;
wire net_18171;
wire net_15513;
wire net_19852;
wire net_6442;
wire net_15487;
wire net_4508;
wire net_17336;
wire net_20602;
wire net_8093;
wire net_3498;
wire net_12831;
wire net_13580;
wire net_21724;
wire net_9658;
wire net_19422;
wire net_5954;
wire net_14321;
wire net_6119;
wire net_14020;
wire net_9960;
wire net_16190;
wire net_14949;
wire x1701;
wire net_10672;
wire net_16486;
wire net_10476;
wire net_16502;
wire net_2207;
wire net_263;
wire net_16027;
wire net_8509;
wire net_14139;
wire net_3483;
wire net_6838;
wire net_10548;
wire net_17936;
wire net_19867;
wire net_12528;
wire net_4189;
wire net_20043;
wire net_19034;
wire net_16826;
wire net_22313;
wire net_9256;
wire net_1090;
wire net_14850;
wire net_3685;
wire net_7030;
wire net_7012;
wire net_14107;
wire net_9007;
wire net_4285;
wire net_8643;
wire net_15862;
wire net_10726;
wire net_201;
wire net_5077;
wire net_20016;
wire net_17315;
wire net_9496;
wire net_3280;
wire net_17426;
wire net_9666;
wire net_3085;
wire net_4043;
wire net_12631;
wire net_12207;
wire net_20716;
wire net_1852;
wire net_11236;
wire net_11912;
wire net_9515;
wire net_6129;
wire x3416;
wire net_2780;
wire net_18631;
wire net_789;
wire net_15240;
wire net_10769;
wire net_3244;
wire net_12819;
wire net_9041;
wire x5873;
wire net_15282;
wire net_18460;
wire net_12080;
wire net_3833;
wire net_9967;
wire net_8664;
wire net_7256;
wire net_19476;
wire net_19703;
wire net_14870;
wire net_8143;
wire net_22380;
wire net_5137;
wire net_17502;
wire net_11569;
wire net_1860;
wire net_18197;
wire net_14587;
wire net_8025;
wire net_1432;
wire x2333;
wire net_1312;
wire net_9474;
wire net_5463;
wire net_22475;
wire net_16144;
wire net_8843;
wire net_8435;
wire net_4801;
wire net_16546;
wire net_19922;
wire net_5334;
wire net_22420;
wire net_16452;
wire net_5290;
wire net_22561;
wire net_14958;
wire net_17488;
wire net_3546;
wire net_8002;
wire net_1453;
wire net_14328;
wire net_13802;
wire net_13075;
wire net_9603;
wire net_21335;
wire net_3542;
wire net_634;
wire net_5374;
wire net_8516;
wire net_20254;
wire net_14177;
wire net_9630;
wire net_8055;
wire net_14066;
wire x6461;
wire net_371;
wire net_15474;
wire net_13786;
wire net_7752;
wire net_2787;
wire net_22663;
wire net_2466;
wire net_4904;
wire net_8580;
wire net_4699;
wire net_7710;
wire net_7975;
wire net_8872;
wire net_18749;
wire net_7574;
wire net_20029;
wire net_13921;
wire net_22227;
wire net_18199;
wire net_5217;
wire net_17794;
wire net_679;
wire net_19907;
wire net_2680;
wire net_8116;
wire net_8924;
wire net_308;
wire net_12218;
wire net_22389;
wire net_6327;
wire net_22734;
wire net_890;
wire net_21898;
wire x804;
wire net_15693;
wire net_7228;
wire net_9019;
wire net_13401;
wire net_17269;
wire net_9162;
wire net_13646;
wire net_13595;
wire net_2471;
wire net_21112;
wire net_18643;
wire net_17524;
wire net_2404;
wire net_21482;
wire net_481;
wire net_16417;
wire net_5346;
wire net_18879;
wire net_16925;
wire net_6891;
wire net_11482;
wire net_21974;
wire net_1188;
wire net_13855;
wire net_1446;
wire net_541;
wire net_20215;
wire net_20760;
wire net_19605;
wire net_18309;
wire net_13380;
wire net_1251;
wire net_8157;
wire net_20729;
wire net_17725;
wire net_16301;
wire net_8830;
wire net_1697;
wire net_15748;
wire net_15741;
wire net_4222;
wire net_12238;
wire net_1753;
wire net_4163;
wire net_14418;
wire net_20140;
wire net_5548;
wire net_14760;
wire net_14298;
wire net_4264;
wire net_9749;
wire net_18492;
wire net_17806;
wire net_15205;
wire net_9908;
wire x2457;
wire net_11418;
wire net_7525;
wire net_17539;
wire net_3071;
wire net_8611;
wire net_21455;
wire net_14238;
wire net_10925;
wire net_9568;
wire net_7149;
wire net_9994;
wire net_7619;
wire net_16404;
wire net_2998;
wire net_15549;
wire net_243;
wire x6381;
wire net_8905;
wire net_6882;
wire net_2854;
wire net_22051;
wire net_10730;
wire net_17567;
wire net_8867;
wire net_4132;
wire net_8925;
wire net_4990;
wire net_7721;
wire net_9292;
wire net_16831;
wire net_11056;
wire net_13588;
wire net_8326;
wire net_19133;
wire net_1915;
wire net_17094;
wire net_15289;
wire net_13566;
wire net_10992;
wire net_8280;
wire net_18428;
wire net_4334;
wire net_16111;
wire net_14650;
wire net_17541;
wire net_19493;
wire net_15295;
wire net_18662;
wire net_12738;
wire net_18399;
wire net_13779;
wire net_12497;
wire net_21350;
wire net_18304;
wire net_18721;
wire net_14452;
wire x2639;
wire net_18557;
wire net_17893;
wire net_13607;
wire net_21162;
wire net_15131;
wire net_17730;
wire net_9195;
wire net_17103;
wire net_12714;
wire net_7164;
wire net_19715;
wire net_12313;
wire net_19860;
wire net_14645;
wire net_9670;
wire net_21847;
wire net_22071;
wire net_14684;
wire net_7633;
wire net_19314;
wire net_13393;
wire net_18716;
wire net_17873;
wire net_8994;
wire net_3202;
wire net_13422;
wire net_4059;
wire net_6376;
wire net_6736;
wire net_7461;
wire net_15032;
wire net_15389;
wire net_10380;
wire net_5612;
wire net_2668;
wire net_13480;
wire net_19610;
wire net_2677;
wire net_15307;
wire net_14498;
wire net_15545;
wire net_10415;
wire net_20030;
wire net_11540;
wire net_11741;
wire net_3916;
wire net_6852;
wire net_22068;
wire net_8312;
wire net_13937;
wire net_18679;
wire net_21606;
wire net_14466;
wire net_12590;
wire x7158;
wire net_18666;
wire net_5900;
wire net_6206;
wire net_3990;
wire x7198;
wire net_20050;
wire net_10221;
wire net_20732;
wire net_3856;
wire net_9210;
wire net_17111;
wire net_20020;
wire net_17478;
wire net_5345;
wire net_8363;
wire net_4885;
wire net_21983;
wire net_17961;
wire net_14459;
wire net_21528;
wire net_19106;
wire net_22626;
wire net_21006;
wire net_19436;
wire net_3501;
wire net_21769;
wire net_16758;
wire net_7862;
wire net_12775;
wire net_6678;
wire net_15070;
wire net_7916;
wire net_20288;
wire net_13600;
wire net_19318;
wire net_8081;
wire net_15524;
wire net_13982;
wire net_14013;
wire net_8835;
wire net_1272;
wire net_17743;
wire net_10273;
wire net_3505;
wire net_4001;
wire net_5059;
wire net_21217;
wire net_655;
wire net_3536;
wire net_6878;
wire net_16918;
wire net_8534;
wire net_10059;
wire net_17634;
wire net_18350;
wire net_16275;
wire net_12961;
wire net_9110;
wire net_20221;
wire net_14403;
wire net_423;
wire net_3036;
wire net_20390;
wire net_18446;
wire net_328;
wire net_10103;
wire net_10565;
wire net_7934;
wire net_7977;
wire net_9060;
wire net_3294;
wire x1932;
wire net_3016;
wire net_4477;
wire net_12933;
wire net_9117;
wire net_11717;
wire net_3749;
wire net_2746;
wire net_12592;
wire net_9403;
wire net_5024;
wire net_15820;
wire net_18267;
wire net_14574;
wire net_11863;
wire net_2594;
wire net_15574;
wire net_22138;
wire net_17452;
wire net_17151;
wire net_5944;
wire net_15436;
wire net_811;
wire net_1684;
wire net_20973;
wire net_14549;
wire net_30;
wire net_1462;
wire net_15019;
wire net_9150;
wire net_4993;
wire net_21754;
wire net_21521;
wire net_1926;
wire net_3115;
wire net_19843;
wire net_20843;
wire net_16621;
wire net_14158;
wire net_14809;
wire net_3518;
wire net_13069;
wire net_10261;
wire net_22482;
wire net_19929;
wire net_18335;
wire net_3680;
wire net_6926;
wire net_14319;
wire net_3984;
wire net_20507;
wire net_13317;
wire net_3615;
wire net_21540;
wire net_9559;
wire net_13172;
wire net_3055;
wire net_9844;
wire net_17813;
wire net_15782;
wire net_21436;
wire net_17230;
wire net_2845;
wire net_3095;
wire net_6510;
wire net_12585;
wire net_11358;
wire net_4586;
wire net_14986;
wire net_21394;
wire x848;
wire net_13141;
wire net_1763;
wire net_6168;
wire net_7291;
wire net_18338;
wire net_15476;
wire net_11067;
wire net_22127;
wire net_12999;
wire net_3278;
wire net_12277;
wire net_4386;
wire net_20278;
wire net_20786;
wire net_20137;
wire net_8837;
wire net_1513;
wire net_15014;
wire net_16447;
wire net_21492;
wire net_19122;
wire net_10668;
wire net_12701;
wire net_4613;
wire net_7763;
wire net_20500;
wire net_11388;
wire net_10084;
wire net_20592;
wire net_73;
wire net_3135;
wire net_5266;
wire net_5165;
wire net_22668;
wire net_8473;
wire net_21545;
wire net_18518;
wire net_8209;
wire net_1899;
wire net_20702;
wire net_15715;
wire net_19920;
wire net_8890;
wire net_4746;
wire net_16614;
wire net_12198;
wire net_1843;
wire net_6031;
wire net_17196;
wire net_22146;
wire net_12211;
wire net_7019;
wire net_534;
wire net_22333;
wire net_3793;
wire net_21977;
wire net_9261;
wire net_13523;
wire net_8659;
wire net_6823;
wire net_17316;
wire net_1551;
wire net_14951;
wire net_486;
wire net_20360;
wire net_18083;
wire net_14753;
wire net_12898;
wire net_406;
wire net_21805;
wire net_20063;
wire net_22003;
wire net_4190;
wire net_5391;
wire net_12448;
wire net_8967;
wire net_15186;
wire net_3640;
wire net_18455;
wire net_748;
wire net_10587;
wire net_20231;
wire net_6917;
wire net_13124;
wire net_10778;
wire net_3958;
wire net_19938;
wire net_12270;
wire net_5427;
wire net_19433;
wire net_16337;
wire net_15259;
wire net_11621;
wire net_20109;
wire net_11684;
wire net_14902;
wire net_514;
wire net_18766;
wire x122;
wire net_3645;
wire net_1604;
wire net_6499;
wire net_5755;
wire net_20395;
wire net_524;
wire net_13816;
wire net_21706;
wire net_17295;
wire net_21663;
wire net_4368;
wire net_7109;
wire net_20646;
wire net_13002;
wire net_22424;
wire net_18190;
wire net_22727;
wire net_3748;
wire net_15164;
wire net_10786;
wire net_9355;
wire net_14789;
wire net_21446;
wire net_19957;
wire net_12083;
wire net_5067;
wire net_10935;
wire net_1097;
wire net_11756;
wire net_12227;
wire net_14172;
wire net_762;
wire net_17176;
wire net_19785;
wire net_17373;
wire net_3589;
wire net_22297;
wire net_4943;
wire net_17766;
wire net_15827;
wire net_8400;
wire net_6173;
wire net_893;
wire net_3330;
wire net_11163;
wire net_255;
wire net_21579;
wire net_20469;
wire net_9641;
wire net_619;
wire net_13618;
wire net_9085;
wire net_17275;
wire net_19210;
wire net_3932;
wire net_7233;
wire net_11177;
wire net_7689;
wire net_14802;
wire net_21637;
wire net_7104;
wire net_14909;
wire net_19818;
wire net_3444;
wire net_4922;
wire net_3800;
wire net_21860;
wire net_3285;
wire net_20672;
wire net_17990;
wire net_7278;
wire net_22530;
wire net_4425;
wire net_18771;
wire net_68;
wire net_4933;
wire net_5834;
wire net_17623;
wire net_4044;
wire net_14862;
wire net_11300;
wire net_21857;
wire net_13285;
wire net_11699;
wire net_5875;
wire net_4630;
wire net_21225;
wire net_16091;
wire net_15636;
wire net_976;
wire net_6287;
wire net_20361;
wire net_2709;
wire net_5309;
wire net_20265;
wire net_10321;
wire net_20906;
wire net_11630;
wire net_611;
wire net_19859;
wire net_7879;
wire net_17849;
wire net_3514;
wire net_5441;
wire net_19644;
wire net_20249;
wire net_17560;
wire net_6077;
wire net_10849;
wire net_4907;
wire net_6567;
wire net_4107;
wire net_18285;
wire net_2160;
wire net_3692;
wire net_3477;
wire net_391;
wire net_6361;
wire net_9268;
wire net_9723;
wire net_5040;
wire net_20121;
wire net_21360;
wire net_18108;
wire net_5820;
wire net_6692;
wire net_4172;
wire net_16735;
wire x826;
wire net_13892;
wire net_8123;
wire net_12417;
wire net_22757;
wire net_1141;
wire net_6253;
wire net_10621;
wire net_16372;
wire net_3243;
wire net_4867;
wire net_22503;
wire net_7871;
wire net_19199;
wire net_2104;
wire net_5564;
wire net_17040;
wire net_6190;
wire net_19540;
wire net_2766;
wire net_3771;
wire net_20950;
wire net_12469;
wire net_2417;
wire net_16004;
wire net_14406;
wire net_22110;
wire net_741;
wire x2103;
wire net_5509;
wire net_20116;
wire net_17862;
wire net_15092;
wire net_7853;
wire net_6472;
wire net_13765;
wire net_3789;
wire net_15664;
wire net_13288;
wire net_19355;
wire net_18783;
wire net_9598;
wire net_11947;
wire net_12977;
wire net_2850;
wire net_20667;
wire net_770;
wire net_13905;
wire net_12901;
wire net_1005;
wire net_15711;
wire net_11792;
wire net_11198;
wire net_21276;
wire net_1059;
wire net_3891;
wire net_4918;
wire net_16650;
wire net_18903;
wire net_17240;
wire net_1796;
wire net_10328;
wire net_21980;
wire net_5187;
wire net_7501;
wire net_11368;
wire net_11291;
wire net_19260;
wire net_1507;
wire net_2310;
wire net_18354;
wire net_7466;
wire net_474;
wire net_16901;
wire net_16358;
wire net_12518;
wire net_11421;
wire net_11934;
wire net_18076;
wire net_11940;
wire net_7947;
wire net_16310;
wire net_11855;
wire net_12244;
wire net_944;
wire net_16019;
wire net_10008;
wire x1781;
wire net_17385;
wire net_18236;
wire net_21030;
wire net_13477;
wire net_12538;
wire net_21718;
wire net_11002;
wire net_7199;
wire net_22217;
wire net_21834;
wire net_21294;
wire net_12580;
wire net_17003;
wire net_63;
wire net_15709;
wire net_13669;
wire net_19574;
wire net_12028;
wire net_287;
wire net_17492;
wire net_189;
wire net_10414;
wire net_21882;
wire net_20946;
wire net_9893;
wire net_9860;
wire net_15988;
wire net_3755;
wire net_6036;
wire net_433;
wire net_22012;
wire net_11709;
wire net_22813;
wire net_8296;
wire net_4443;
wire net_224;
wire net_15886;
wire net_1898;
wire net_19481;
wire net_9073;
wire net_608;
wire net_1212;
wire net_3604;
wire net_4383;
wire net_5331;
wire net_13194;
wire net_3706;
wire net_21246;
wire net_16387;
wire net_7062;
wire net_12879;
wire net_11997;
wire net_8299;
wire net_12832;
wire net_18066;
wire net_18443;
wire net_22654;
wire net_6416;
wire net_16696;
wire net_15923;
wire net_13227;
wire net_17573;
wire net_873;
wire net_1811;
wire net_13884;
wire net_12374;
wire net_11080;
wire net_20297;
wire net_20189;
wire net_2588;
wire net_20591;
wire net_7802;
wire x1314;
wire net_18921;
wire net_9771;
wire net_704;
wire net_12906;
wire net_3997;
wire net_1356;
wire net_14542;
wire net_8913;
wire net_4393;
wire net_6541;
wire net_3816;
wire net_6101;
wire net_13457;
wire net_5539;
wire net_9056;
wire net_1711;
wire net_14527;
wire net_2084;
wire net_8186;
wire net_11590;
wire x4416;
wire net_9530;
wire net_5085;
wire net_7031;
wire net_7349;
wire net_12653;
wire net_8680;
wire net_20583;
wire net_16506;
wire net_4836;
wire net_9602;
wire net_17366;
wire net_15265;
wire net_11663;
wire x7268;
wire net_7270;
wire net_9283;
wire net_21650;
wire net_12892;
wire net_2526;
wire net_18758;
wire net_16237;
wire net_9414;
wire net_21304;
wire net_18838;
wire net_7338;
wire net_1644;
wire net_12126;
wire net_2800;
wire net_19204;
wire net_14225;
wire net_7940;
wire net_17354;
wire net_17695;
wire net_8255;
wire net_1190;
wire net_3225;
wire x2420;
wire net_19351;
wire net_19163;
wire net_4093;
wire net_6449;
wire net_15535;
wire net_4799;
wire net_16269;
wire net_13812;
wire net_8721;
wire net_12021;
wire net_9829;
wire net_6066;
wire net_17361;
wire net_15140;
wire net_19824;
wire net_2191;
wire net_21933;
wire net_14698;
wire net_13318;
wire net_21382;
wire net_13304;
wire net_22486;
wire net_10690;
wire net_17672;
wire net_15077;
wire net_13168;
wire net_12617;
wire net_15639;
wire net_12416;
wire net_12352;
wire net_14249;
wire net_22670;
wire net_21739;
wire net_1577;
wire net_22760;
wire net_17714;
wire net_1054;
wire net_4595;
wire net_20182;
wire net_22209;
wire net_21127;
wire net_17595;
wire net_19345;
wire net_2727;
wire net_18225;
wire net_16185;
wire net_5605;
wire net_2257;
wire net_10640;
wire net_14741;
wire net_3418;
wire net_18751;
wire net_5491;
wire net_20963;
wire net_13217;
wire net_12044;
wire net_2968;
wire net_7314;
wire net_10649;
wire net_5989;
wire net_19534;
wire net_16105;
wire net_12339;
wire net_2643;
wire net_5845;
wire net_21953;
wire net_19464;
wire net_22302;
wire net_9591;
wire net_3722;
wire net_18034;
wire net_11117;
wire net_17739;
wire net_18331;
wire net_1517;
wire net_19402;
wire net_19307;
wire net_16416;
wire net_11218;
wire net_5980;
wire net_6705;
wire net_9192;
wire net_15217;
wire net_21956;
wire net_1690;
wire net_20464;
wire x1878;
wire x648;
wire net_16606;
wire net_22187;
wire net_19738;
wire net_20312;
wire net_11924;
wire net_2093;
wire net_2997;
wire net_14831;
wire net_15027;
wire net_14186;
wire net_9076;
wire net_7239;
wire net_18776;
wire net_11787;
wire net_19370;
wire net_17138;
wire net_15099;
wire net_18419;
wire net_9549;
wire net_20696;
wire net_4357;
wire net_16878;
wire net_16714;
wire net_2536;
wire net_5890;
wire net_20645;
wire net_7968;
wire net_19455;
wire net_2949;
wire net_3429;
wire net_22251;
wire net_10954;
wire net_9032;
wire net_1708;
wire net_12398;
wire net_5519;
wire net_17215;
wire net_15966;
wire net_13112;
wire net_12575;
wire net_13050;
wire net_722;
wire net_5420;
wire net_17065;
wire net_12094;
wire net_18044;
wire net_20890;
wire net_14612;
wire net_13099;
wire net_5798;
wire net_11351;
wire net_14313;
wire net_5223;
wire net_8216;
wire net_435;
wire net_12077;
wire net_1830;
wire net_21790;
wire net_20910;
wire x140;
wire net_20442;
wire net_22689;
wire net_5156;
wire net_6481;
wire net_1649;
wire net_6603;
wire net_1837;
wire net_6973;
wire net_2427;
wire net_8075;
wire net_1071;
wire net_3378;
wire net_18607;
wire net_5004;
wire net_5817;
wire net_9776;
wire net_18499;
wire net_1701;
wire net_5675;
wire net_11156;
wire net_14007;
wire net_8678;
wire net_12175;
wire net_1633;
wire net_11132;
wire net_12150;
wire net_5251;
wire net_8694;
wire net_15759;
wire net_319;
wire net_18435;
wire net_2670;
wire net_1743;
wire net_2597;
wire net_5913;
wire net_87;
wire net_7640;
wire net_11887;
wire net_4139;
wire net_2923;
wire net_7545;
wire net_512;
wire net_16646;
wire net_19595;
wire net_17878;
wire net_3102;
wire net_18027;
wire net_7510;
wire net_16221;
wire net_13513;
wire net_5780;
wire net_5721;
wire net_7904;
wire net_19762;
wire net_13119;
wire net_16368;
wire net_16243;
wire net_16999;
wire net_3371;
wire net_17898;
wire net_5317;
wire net_13953;
wire net_15874;
wire net_21701;
wire net_6800;
wire net_9375;
wire net_12673;
wire x6521;
wire net_17143;
wire net_21005;
wire net_15212;
wire net_1875;
wire net_5862;
wire net_3420;
wire net_21568;
wire net_3887;
wire net_18009;
wire net_16964;
wire net_7050;
wire net_7484;
wire net_22022;
wire net_13373;
wire net_22260;
wire net_15045;
wire net_12189;
wire net_22510;
wire net_8736;
wire net_16585;
wire net_12953;
wire net_5178;
wire net_17035;
wire net_7678;
wire net_17463;
wire net_2835;
wire net_4543;
wire net_4871;
wire net_6599;
wire net_20454;
wire net_1240;
wire net_9213;
wire net_3000;
wire net_16761;
wire net_12200;
wire net_15002;
wire net_22318;
wire net_15768;
wire net_20985;
wire net_12674;
wire net_17533;
wire net_13048;
wire net_858;
wire net_9338;
wire net_22636;
wire net_15583;
wire net_8986;
wire net_4766;
wire net_6004;
wire net_21723;
wire net_16167;
wire net_8504;
wire net_13549;
wire net_9867;
wire net_7995;
wire net_3735;
wire net_10870;
wire net_11422;
wire net_1427;
wire net_5123;
wire net_17980;
wire net_3921;
wire net_7075;
wire net_19899;
wire net_5899;
wire net_4098;
wire net_5478;
wire net_7251;
wire x3199;
wire net_19794;
wire net_16494;
wire net_12106;
wire net_9827;
wire net_11029;
wire net_18676;
wire net_17702;
wire net_14762;
wire net_20376;
wire net_22444;
wire net_10308;
wire net_6020;
wire net_7172;
wire net_1677;
wire net_20654;
wire net_13260;
wire net_7089;
wire net_2811;
wire net_6788;
wire net_22027;
wire net_21105;
wire net_19698;
wire net_2612;
wire net_8791;
wire net_5230;
wire net_19149;
wire net_2042;
wire net_7189;
wire net_20939;
wire net_13626;
wire net_17218;
wire net_11649;
wire net_18270;
wire net_6649;
wire net_10949;
wire net_3488;
wire x3322;
wire net_3023;
wire net_17010;
wire net_19987;
wire net_5584;
wire net_1202;
wire net_14373;
wire net_19408;
wire net_20934;
wire net_10890;
wire net_925;
wire net_4932;
wire net_19829;
wire net_6776;
wire net_7452;
wire net_21357;
wire net_12827;
wire net_5384;
wire net_17250;
wire net_15680;
wire net_11317;
wire net_10974;
wire net_12074;
wire net_4661;
wire net_2695;
wire net_21904;
wire net_10196;
wire net_11054;
wire net_14337;
wire net_13336;
wire net_12851;
wire net_12611;
wire net_7404;
wire net_8564;
wire net_20490;
wire net_7783;
wire net_14477;
wire net_22613;
wire net_18107;
wire net_6284;
wire net_9436;
wire net_7132;
wire net_2313;
wire net_21043;
wire net_59;
wire net_11655;
wire net_22524;
wire net_9044;
wire net_6172;
wire net_7595;
wire net_230;
wire net_18472;
wire net_4214;
wire net_20754;
wire net_19752;
wire net_18861;
wire net_6985;
wire net_3349;
wire net_4782;
wire net_1222;
wire net_3404;
wire net_19744;
wire net_14080;
wire net_21824;
wire net_20478;
wire net_22572;
wire net_14291;
wire net_19965;
wire net_17734;
wire net_3810;
wire net_14560;
wire net_9172;
wire net_12018;
wire net_19639;
wire net_15689;
wire net_4739;
wire net_4156;
wire net_8823;
wire net_12685;
wire net_13693;
wire net_12459;
wire net_3440;
wire net_6904;
wire net_19223;
wire net_3358;
wire net_1776;
wire net_3368;
wire net_5747;
wire net_15897;
wire net_4014;
wire net_14723;
wire net_19442;
wire net_15626;
wire net_21001;
wire net_18116;
wire net_7204;
wire net_17017;
wire net_2132;
wire net_2292;
wire net_9313;
wire net_12367;
wire net_1880;
wire net_17856;
wire net_3862;
wire net_184;
wire net_5103;
wire net_17901;
wire net_5855;
wire net_10757;
wire net_14087;
wire net_11247;
wire net_10427;
wire net_15359;
wire net_7203;
wire net_18214;
wire net_18967;
wire net_17089;
wire net_1867;
wire net_18626;
wire net_9498;
wire net_8205;
wire net_1949;
wire net_2650;
wire net_13568;
wire net_10455;
wire net_22160;
wire net_1804;
wire net_21926;
wire net_17554;
wire net_2331;
wire net_14520;
wire net_6667;
wire net_16741;
wire net_16042;
wire net_4291;
wire net_12389;
wire net_8637;
wire net_14483;
wire net_1135;
wire net_1365;
wire net_16768;
wire net_11674;
wire net_43;
wire net_1346;
wire net_5047;
wire net_18957;
wire net_17199;
wire net_11478;
wire net_15946;
wire net_13865;
wire net_13835;
wire net_9220;
wire net_9277;
wire net_1801;
wire net_18819;
wire net_15650;
wire net_14364;
wire net_4350;
wire net_6029;
wire net_8955;
wire net_15724;
wire net_669;
wire net_937;
wire net_11252;
wire net_10179;
wire net_21501;
wire net_8452;
wire net_9575;
wire net_8030;
wire net_20096;
wire net_479;
wire net_8740;
wire net_12769;
wire net_6086;
wire net_2030;
wire x1227;
wire net_1587;
wire net_17077;
wire net_13232;
wire net_11025;
wire net_21404;
wire net_796;
wire net_18610;
wire net_22514;
wire net_20790;
wire net_648;
wire net_11901;
wire net_22102;
wire net_16109;
wire net_6884;
wire net_12040;
wire net_8150;
wire net_16888;
wire net_14300;
wire net_14443;
wire net_7054;
wire net_11950;
wire net_7625;
wire net_3658;
wire net_20531;
wire net_12560;
wire net_22598;
wire net_19566;
wire net_14146;
wire net_6964;
wire net_9148;
wire net_15871;
wire net_15414;
wire net_18550;
wire net_17953;
wire net_8237;
wire net_17951;
wire net_17123;
wire net_8556;
wire net_7649;
wire net_16793;
wire net_15804;
wire net_12179;
wire net_10739;
wire net_10232;
wire net_20869;
wire net_15840;
wire net_8725;
wire net_20699;
wire net_4492;
wire net_6700;
wire net_14655;
wire net_1961;
wire net_10831;
wire net_1260;
wire net_10124;
wire net_20568;
wire net_9832;
wire net_15375;
wire net_239;
wire net_18824;
wire net_13396;
wire net_310;
wire net_18899;
wire net_14599;
wire net_10367;
wire net_2437;
wire net_10792;
wire net_14772;
wire net_8982;
wire net_9917;
wire net_13498;
wire net_5886;
wire net_14960;
wire net_17755;
wire net_20070;
wire net_13711;
wire net_682;
wire net_17580;
wire net_1963;
wire net_7122;
wire net_108;
wire net_21071;
wire net_17114;
wire net_13558;
wire net_16033;
wire net_12049;
wire net_17976;
wire net_8989;
wire net_3560;
wire net_5804;
wire net_17908;
wire net_1007;
wire net_15497;
wire net_7000;
wire net_14837;
wire net_4772;
wire net_7007;
wire net_11415;
wire net_1292;
wire net_7197;
wire net_10703;
wire net_7861;
wire net_10771;
wire net_20872;
wire net_12262;
wire net_11039;
wire net_2796;
wire net_18202;
wire net_11400;
wire net_16526;
wire net_15845;
wire net_21938;
wire net_19044;
wire net_5016;
wire net_4024;
wire net_6699;
wire net_9544;
wire net_20631;
wire net_12443;
wire net_6280;
wire net_17086;
wire net_8043;
wire net_1937;
wire net_15114;
wire net_7215;
wire net_21403;
wire net_18308;
wire net_1956;
wire net_11339;
wire net_13433;
wire net_1614;
wire net_13491;
wire net_12911;
wire net_19500;
wire net_11958;
wire net_16597;
wire net_7119;
wire net_10255;
wire net_3209;
wire net_21063;
wire net_19111;
wire net_12791;
wire net_21471;
wire net_4891;
wire net_8688;
wire net_10874;
wire net_8412;
wire net_19326;
wire net_21232;
wire net_7716;
wire net_294;
wire net_17606;
wire net_15305;
wire x563;
wire net_9837;
wire net_10797;
wire net_2429;
wire net_9217;
wire net_1265;
wire net_10822;
wire net_6224;
wire net_14694;
wire net_8697;
wire net_11203;
wire net_12984;
wire net_19089;
wire net_19888;
wire net_8039;
wire net_1619;
wire net_5468;
wire net_12727;
wire net_18742;
wire net_2124;
wire net_5934;
wire net_15247;
wire net_1161;
wire net_7070;
wire net_19140;
wire net_4671;
wire net_17587;
wire net_13606;
wire net_12695;
wire net_7663;
wire net_21132;
wire net_11385;
wire net_10721;
wire net_8500;
wire net_1395;
wire net_8877;
wire net_9360;
wire net_22620;
wire net_21258;
wire net_15005;
wire net_11875;
wire net_17128;
wire net_22452;
wire net_14678;
wire net_5353;
wire net_16195;
wire net_8756;
wire net_5270;
wire net_22462;
wire net_9921;
wire net_12456;
wire net_18218;
wire net_2445;
wire net_3396;
wire net_6640;
wire net_5324;
wire net_15452;
wire net_10592;
wire net_16836;
wire net_20601;
wire net_4511;
wire net_7395;
wire net_13419;
wire net_2894;
wire net_15643;
wire net_13714;
wire net_6999;
wire net_1988;
wire net_7388;
wire net_20544;
wire net_3718;
wire net_4419;
wire net_15619;
wire net_5284;
wire net_16488;
wire net_11125;
wire net_3525;
wire net_10696;
wire net_20240;
wire net_6850;
wire net_20819;
wire net_13508;
wire net_1608;
wire net_506;
wire net_3769;
wire net_12802;
wire net_8019;
wire net_21730;
wire net_9330;
wire net_12836;
wire net_3775;
wire net_8278;
wire x3136;
wire net_5432;
wire net_6586;
wire net_19082;
wire net_5096;
wire net_16020;
wire net_7589;
wire net_12055;
wire net_6909;
wire net_290;
wire net_6476;
wire net_13676;
wire net_6315;
wire net_10913;
wire net_3313;
wire net_9987;
wire net_20608;
wire net_8803;
wire net_5769;
wire net_3591;
wire net_5729;
wire net_16812;
wire net_16207;
wire net_13341;
wire net_15025;
wire net_16464;
wire net_11926;
wire net_12430;
wire net_4436;
wire net_22091;
wire net_15775;
wire net_2329;
wire net_22831;
wire net_16801;
wire net_2150;
wire net_7129;
wire net_2065;
wire net_10003;
wire net_20345;
wire net_13244;
wire net_10030;
wire net_17467;
wire net_8373;
wire net_2927;
wire net_7397;
wire net_16634;
wire net_11831;
wire net_11838;
wire net_194;
wire net_4856;
wire net_13941;
wire net_11264;
wire net_9448;
wire net_21457;
wire net_1128;
wire net_2713;
wire net_13161;
wire net_11582;
wire net_15354;
wire net_12539;
wire net_11320;
wire net_20753;
wire net_1119;
wire net_9637;
wire net_4312;
wire net_19522;
wire net_20886;
wire net_5299;
wire net_8852;
wire net_3345;
wire net_18319;
wire net_10125;
wire net_18582;
wire net_7855;
wire net_11642;
wire net_11006;
wire net_7127;
wire net_7448;
wire net_11900;
wire net_18042;
wire net_19446;
wire net_10742;
wire net_3328;
wire net_14812;
wire net_10174;
wire net_16328;
wire net_2107;
wire net_22742;
wire net_180;
wire net_13462;
wire net_17107;
wire net_6859;
wire net_22246;
wire net_5657;
wire net_4367;
wire net_3290;
wire net_3731;
wire net_1475;
wire net_10241;
wire net_18207;
wire net_14112;
wire net_16459;
wire net_16738;
wire net_10601;
wire net_5446;
wire net_12719;
wire net_21090;
wire net_2173;
wire net_18597;
wire net_9053;
wire net_6865;
wire net_7539;
wire net_20386;
wire net_14785;
wire net_6263;
wire net_5590;
wire net_11673;
wire net_19802;
wire net_14334;
wire x2945;
wire net_5476;
wire net_3744;
wire net_11851;
wire net_21917;
wire net_21379;
wire net_4635;
wire net_14912;
wire net_12193;
wire net_20557;
wire net_18946;
wire net_6570;
wire net_8309;
wire net_15360;
wire net_6939;
wire net_12968;
wire net_4485;
wire net_1558;
wire net_22537;
wire net_8603;
wire x1413;
wire net_4641;
wire net_17405;
wire net_10958;
wire net_10806;
wire net_19597;
wire net_14138;
wire net_455;
wire net_11515;
wire net_16072;
wire net_10294;
wire net_115;
wire net_7498;
wire net_3339;
wire net_6303;
wire net_22459;
wire net_9428;
wire net_7352;
wire net_1832;
wire net_12474;
wire net_20810;
wire net_12622;
wire net_1026;
wire net_16095;
wire net_2215;
wire net_22413;
wire net_15376;
wire net_6453;
wire net_2573;
wire net_22274;
wire net_9369;
wire net_20801;
wire net_10312;
wire net_7378;
wire net_19004;
wire net_21378;
wire net_3993;
wire net_13673;
wire net_21028;
wire net_20825;
wire net_1401;
wire net_20625;
wire net_19995;
wire net_3909;
wire net_11858;
wire net_17800;
wire net_7889;
wire net_14394;
wire net_7248;
wire net_13311;
wire net_17557;
wire net_443;
wire net_6367;
wire net_6495;
wire net_18907;
wire net_8486;
wire net_20491;
wire x6870;
wire net_17661;
wire net_18389;
wire net_20323;
wire net_12364;
wire net_7956;
wire net_14034;
wire net_11346;
wire net_1990;
wire net_7456;
wire net_18155;
wire net_10442;
wire net_17350;
wire net_16391;
wire net_9951;
wire net_18843;
wire net_7880;
wire net_19368;
wire net_11988;
wire net_11601;
wire net_622;
wire net_17028;
wire net_14854;
wire net_11993;
wire net_20251;
wire net_11277;
wire net_5909;
wire net_11225;
wire net_19373;
wire net_1338;
wire net_20168;
wire net_7842;
wire net_19627;
wire net_2053;
wire net_6623;
wire net_2180;
wire x33;
wire net_4242;
wire net_2119;
wire net_3220;
wire net_4720;
wire net_21510;
wire net_18152;
wire net_13108;
wire net_8627;
wire net_7474;
wire net_5920;
wire net_6124;
wire net_22785;
wire net_8384;
wire net_6992;
wire net_13519;
wire net_2007;
wire net_5143;
wire net_5763;
wire net_7703;
wire net_20766;
wire net_16211;
wire net_19386;
wire net_713;
wire net_10653;
wire net_5711;
wire net_17329;
wire net_16898;
wire net_13338;
wire net_8700;
wire net_11104;
wire net_729;
wire net_21876;
wire net_21097;
wire net_19076;
wire net_9222;
wire net_4197;
wire net_17292;
wire net_14893;
wire net_20920;
wire net_13156;
wire net_7093;
wire net_7324;
wire net_13948;
wire net_9169;
wire net_8447;
wire net_5366;
wire net_19257;
wire net_14596;
wire net_8711;
wire net_13571;
wire net_19339;
wire net_341;
wire net_13611;
wire net_14733;
wire net_12992;
wire net_970;
wire net_13362;
wire net_13389;
wire net_8653;
wire net_15539;
wire net_15984;
wire net_13917;
wire net_13184;
wire net_20563;
wire net_3044;
wire net_5929;
wire net_21347;
wire net_17257;
wire net_17457;
wire net_11145;
wire net_14745;
wire net_20650;
wire net_20074;
wire net_13726;
wire net_14071;
wire net_14233;
wire net_12038;
wire net_10100;
wire net_20012;
wire net_2163;
wire net_19943;
wire net_3417;
wire net_3307;
wire net_13301;
wire net_12534;
wire net_553;
wire net_4212;
wire net_6133;
wire net_7797;
wire net_21318;
wire net_20880;
wire net_8300;
wire net_6239;
wire net_15991;
wire net_4701;
wire net_18262;
wire net_20271;
wire net_10889;
wire net_15906;
wire net_462;
wire net_418;
wire net_15415;
wire net_15105;
wire net_161;
wire net_20424;
wire net_7988;
wire net_17615;
wire net_8660;
wire net_1486;
wire net_2606;
wire net_19179;
wire net_18687;
wire net_78;
wire net_1839;
wire net_2320;
wire net_20858;
wire net_1665;
wire net_20079;
wire net_11076;
wire net_14515;
wire net_13744;
wire net_8525;
wire net_8349;
wire net_20860;
wire net_18900;
wire net_16179;
wire net_3550;
wire net_16663;
wire net_20411;
wire net_19219;
wire net_12377;
wire net_11172;
wire net_19941;
wire net_16056;
wire net_21989;
wire net_21819;
wire net_6893;
wire net_9466;
wire net_2224;
wire net_7066;
wire net_21169;
wire net_10037;
wire x1483;
wire net_15404;
wire net_5733;
wire net_15847;
wire net_21786;
wire net_2458;
wire net_9324;
wire net_17164;
wire net_19770;
wire net_3435;
wire net_2635;
wire net_16789;
wire net_3374;
wire net_5207;
wire net_15490;
wire net_13540;
wire net_5572;
wire net_21922;
wire net_15068;
wire net_8283;
wire net_1037;
wire net_21512;
wire net_2019;
wire net_18379;
wire net_4676;
wire net_8395;
wire net_6675;
wire net_13033;
wire net_7549;
wire net_20929;
wire net_19155;
wire net_20641;
wire net_6793;
wire net_15793;
wire net_17668;
wire net_6242;
wire net_14433;
wire net_15012;
wire net_1623;
wire net_2982;
wire net_6948;
wire net_4410;
wire net_21949;
wire net_21419;
wire net_19139;
wire net_7230;
wire net_16849;
wire net_5785;
wire net_14047;
wire net_18245;
wire net_17514;
wire net_18537;
wire net_20085;
wire net_14251;
wire net_13657;
wire net_8650;
wire net_7190;
wire net_10907;
wire net_16000;
wire net_18299;
wire net_8596;
wire net_19978;
wire net_20366;
wire net_10984;
wire net_103;
wire net_12147;
wire net_20924;
wire net_19809;
wire net_12166;
wire net_6651;
wire net_19763;
wire net_16009;
wire net_5485;
wire net_7243;
wire net_18974;
wire net_12004;
wire net_3554;
wire net_20025;
wire net_22497;
wire net_22163;
wire net_12323;
wire net_1920;
wire net_4101;
wire net_21687;
wire net_17628;
wire net_2010;
wire net_18913;
wire net_11665;
wire net_8782;
wire net_6941;
wire net_20344;
wire net_8321;
wire net_9139;
wire net_16853;
wire net_18507;
wire net_4672;
wire net_8862;
wire net_6743;
wire net_1723;
wire net_22322;
wire net_8465;
wire net_2900;
wire net_20004;
wire net_14790;
wire net_17648;
wire net_11015;
wire net_5152;
wire net_5718;
wire net_8190;
wire net_17396;
wire net_21327;
wire net_4376;
wire net_17288;
wire net_14397;
wire net_19588;
wire net_18881;
wire net_19495;
wire net_20150;
wire net_16868;
wire net_2306;
wire net_12382;
wire net_2873;
wire net_3272;
wire net_14618;
wire net_2254;
wire net_2861;
wire net_20141;
wire net_18235;
wire net_11844;
wire net_14343;
wire net_9570;
wire net_4574;
wire net_18701;
wire net_1209;
wire net_15936;
wire net_13076;
wire net_4038;
wire net_847;
wire net_10157;
wire net_4787;
wire net_11740;
wire net_283;
wire net_12864;
wire net_22775;
wire net_13505;
wire net_5117;
wire net_18875;
wire net_4690;
wire net_12796;
wire net_5020;
wire net_14126;
wire net_7316;
wire net_5445;
wire net_18725;
wire net_7428;
wire net_10023;
wire net_10990;
wire net_7958;
wire net_16559;
wire net_344;
wire net_14102;
wire net_4757;
wire net_18735;
wire net_15956;
wire net_2269;
wire net_884;
wire net_14184;
wire net_712;
wire net_1422;
wire net_2281;
wire net_12940;
wire net_17655;
wire net_4497;
wire net_11527;
wire net_18960;
wire net_6670;
wire net_15061;
wire net_1106;
wire net_15817;
wire net_13629;
wire net_8483;
wire net_2972;
wire net_20191;
wire net_5611;
wire net_11311;
wire net_10836;
wire net_15252;
wire net_22204;
wire net_2241;
wire net_13006;
wire net_17430;
wire net_9522;
wire net_8615;
wire net_1547;
wire net_15596;
wire net_13053;
wire net_8768;
wire net_20523;
wire net_5122;
wire net_20207;
wire net_12495;
wire net_11146;
wire net_19335;
wire net_5423;
wire net_13972;
wire net_7971;
wire net_6507;
wire net_9912;
wire net_22685;
wire net_10395;
wire net_21036;
wire net_7344;
wire net_20959;
wire net_16956;
wire net_5055;
wire net_14886;
wire net_7303;
wire net_17392;
wire net_4794;
wire net_2625;
wire net_4149;
wire net_5687;
wire net_19451;
wire net_19469;
wire net_21746;
wire net_6849;
wire net_10292;
wire net_1595;
wire net_5849;
wire net_20873;
wire net_15656;
wire net_114;
wire net_19547;
wire net_12919;
wire net_3432;
wire net_2974;
wire net_20675;
wire net_6519;
wire net_14517;
wire net_3895;
wire net_8339;
wire net_13660;
wire net_20993;
wire net_11736;
wire net_2734;
wire net_12888;
wire net_18603;
wire net_15508;
wire net_13133;
wire net_10637;
wire net_12569;
wire net_6761;
wire net_20407;
wire net_14857;
wire net_7827;
wire net_3146;
wire net_6294;
wire net_18118;
wire net_21183;
wire net_21570;
wire net_6390;
wire net_9347;
wire net_20746;
wire net_10496;
wire net_5237;
wire net_22231;
wire net_19417;
wire net_16601;
wire net_14825;
wire net_17643;
wire net_11553;
wire net_3022;
wire net_8226;
wire net_21695;
wire x2357;
wire net_10989;
wire net_19185;
wire net_16808;
wire net_7495;
wire net_21591;
wire net_9616;
wire net_5741;
wire net_6391;
wire net_21174;
wire net_19521;
wire net_8476;
wire net_6308;
wire net_18513;
wire net_16170;
wire net_17344;
wire net_5700;
wire net_7441;
wire net_22825;
wire net_9671;
wire net_15405;
wire net_9159;
wire net_11899;
wire net_14260;
wire net_18684;
wire net_18473;
wire net_4706;
wire net_21759;
wire net_594;
wire net_5532;
wire net_17203;
wire net_11336;
wire net_9818;
wire net_17225;
wire net_22579;
wire net_14310;
wire net_11892;
wire net_8512;
wire net_22365;
wire net_11690;
wire net_6188;
wire net_4402;
wire net_6328;
wire net_2074;
wire net_16254;
wire net_8428;
wire net_5256;
wire net_16842;
wire net_5274;
wire net_10183;
wire net_2577;
wire net_11091;
wire net_8286;
wire net_2954;
wire net_15890;
wire net_3274;
wire net_17762;
wire net_20484;
wire net_16143;
wire net_2953;
wire net_15731;
wire net_6380;
wire net_467;
wire net_22447;
wire net_2910;
wire x4041;
wire net_19300;
wire net_8728;
wire net_4851;
wire net_2081;
wire net_9245;
wire net_10522;
wire net_21889;
wire net_5195;
wire net_11426;
wire net_18132;
wire net_14555;
wire net_19053;
wire net_3165;
wire net_12644;
wire net_22643;
wire net_22178;
wire net_21083;
wire net_22042;
wire net_18858;
wire net_4965;
wire x23;
wire net_22241;
wire net_12295;
wire net_8648;
wire net_2302;
wire net_21108;
wire net_12523;
wire net_18280;
wire net_14601;
wire net_8545;
wire net_19397;
wire net_19634;
wire net_13649;
wire net_19771;
wire net_22694;
wire net_5502;
wire net_6805;
wire net_6387;
wire net_6403;
wire net_7734;
wire net_18344;
wire net_13873;
wire net_12409;
wire net_15916;
wire net_15294;
wire net_2368;
wire net_18482;
wire net_19667;
wire net_19001;
wire net_12908;
wire net_3966;
wire net_6330;
wire net_607;
wire net_21466;
wire x7527;
wire net_12392;
wire net_8106;
wire net_22601;
wire net_9739;
wire x1425;
wire net_4142;
wire net_1045;
wire net_20173;
wire net_3497;
wire net_22211;
wire net_3905;
wire net_13087;
wire net_21921;
wire net_15392;
wire net_13249;
wire net_4939;
wire net_17246;
wire net_3601;
wire net_9933;
wire x6178;
wire net_22712;
wire net_16133;
wire net_4538;
wire net_19041;
wire net_14648;
wire net_13044;
wire net_12052;
wire net_18073;
wire net_15550;
wire net_20660;
wire net_11167;
wire net_16685;
wire net_12662;
wire net_4527;
wire net_6419;
wire net_18187;
wire net_8548;
wire net_21715;
wire net_4144;
wire net_4716;
wire net_7586;
wire net_2079;
wire net_1731;
wire net_2052;
wire net_16038;
wire net_9089;
wire net_16541;
wire net_9648;
wire net_9463;
wire net_6912;
wire net_12813;
wire net_17419;
wire net_13276;
wire net_17202;
wire net_5952;
wire net_11769;
wire net_15422;
wire net_3636;
wire net_21015;
wire net_7184;
wire net_14095;
wire net_4727;
wire net_17769;
wire net_5032;
wire net_11046;
wire net_1536;
wire net_5852;
wire net_6232;
wire net_12504;
wire net_3478;
wire net_1498;
wire net_8117;
wire net_18089;
wire net_10815;
wire net_20538;
wire net_5561;
wire net_5626;
wire net_949;
wire net_19660;
wire net_14000;
wire net_12401;
wire net_10936;
wire net_7813;
wire net_20851;
wire net_4111;
wire net_9392;
wire net_14267;
wire net_10616;
wire net_12947;
wire net_12287;
wire net_18359;
wire net_18141;
wire net_12722;
wire net_14283;
wire net_20176;
wire net_8262;
wire net_9028;
wire net_2296;
wire x3376;
wire net_9438;
wire net_13994;
wire net_21912;
wire net_3385;
wire net_17798;
wire net_357;
wire net_6954;
wire net_9179;
wire net_12934;
wire net_20331;
wire net_7849;
wire net_3451;
wire net_18769;
wire net_7085;
wire net_8790;
wire net_2694;
wire net_21728;
wire net_17184;
wire net_12280;
wire net_5607;
wire net_2096;
wire net_3118;
wire net_5555;
wire net_18560;
wire net_18521;
wire net_22036;
wire net_22806;
wire net_21864;
wire net_20998;
wire net_15330;
wire net_11501;
wire net_1829;
wire net_16434;
wire net_14240;
wire net_13904;
wire net_9780;
wire x7296;
wire net_662;
wire net_862;
wire net_16121;
wire net_50;
wire net_2307;
wire net_7168;
wire net_14822;
wire net_8127;
wire net_4174;
wire net_5396;
wire net_738;
wire net_4080;
wire net_4325;
wire net_1150;
wire net_504;
wire net_22547;
wire net_18831;
wire net_10333;
wire net_9789;
wire x2367;
wire net_6634;
wire x6710;
wire net_11537;
wire net_7698;
wire net_17839;
wire net_16593;
wire net_21708;
wire net_18348;
wire net_3120;
wire net_14324;
wire net_18274;
wire net_4504;
wire net_1561;
wire net_20517;
wire net_12161;
wire net_3269;
wire net_11455;
wire net_22392;
wire net_17332;
wire net_10472;
wire net_4421;
wire net_18360;
wire net_6666;
wire net_17048;
wire net_19835;
wire net_17775;
wire net_13329;
wire net_9855;
wire net_1940;
wire net_13323;
wire net_11449;
wire net_10452;
wire net_8635;
wire net_11516;
wire net_16670;
wire net_12781;
wire net_14621;
wire net_11528;
wire net_991;
wire net_3912;
wire net_6528;
wire net_13204;
wire net_18253;
wire net_6753;
wire net_3088;
wire net_19531;
wire net_21969;
wire net_19242;
wire net_11107;
wire net_4607;
wire net_12484;
wire net_2979;
wire net_20692;
wire net_20035;
wire net_17925;
wire net_16712;
wire net_10714;
wire net_2772;
wire net_9564;
wire net_21596;
wire net_19398;
wire net_8491;
wire net_5775;
wire net_4180;
wire net_15562;
wire net_13839;
wire net_12116;
wire net_12180;
wire net_2347;
wire net_11710;
wire net_14777;
wire net_2684;
wire net_3806;
wire net_10795;
wire net_10352;
wire net_521;
wire net_3972;
wire net_14275;
wire net_9003;
wire net_14738;
wire net_2754;
wire net_267;
wire net_1585;
wire x2784;
wire net_13748;
wire net_11613;
wire net_20319;
wire net_9143;
wire net_18541;
wire net_11099;
wire net_22398;
wire net_15761;
wire net_6898;
wire net_7421;
wire net_16618;
wire net_3663;
wire net_22430;
wire net_10885;
wire net_3260;
wire net_5110;
wire net_13017;
wire net_9186;
wire net_6465;
wire net_6486;
wire net_6048;
wire net_13177;
wire net_18652;
wire net_2716;
wire x2249;
wire net_11815;
wire net_20954;
wire net_6551;
wire net_4750;
wire net_20614;
wire net_15868;
wire net_13346;
wire net_4558;
wire net_12858;
wire net_21537;
wire net_21209;
wire net_8394;
wire net_15521;
wire net_2828;
wire net_12749;
wire net_824;
wire net_3458;
wire net_1822;
wire net_18801;
wire net_9755;
wire net_19256;
wire net_13038;
wire net_1972;
wire net_15559;
wire net_17945;
wire net_12267;
wire net_3126;
wire net_993;
wire net_10555;
wire net_20106;
wire net_5974;
wire net_21387;
wire net_9456;
wire net_1100;
wire net_7035;
wire net_15121;
wire net_21285;
wire net_14995;
wire net_2817;
wire net_18039;
wire net_22792;
wire net_6686;
wire net_10046;
wire net_17931;
wire net_21618;
wire net_21150;
wire net_15128;
wire net_5996;
wire net_6730;
wire net_13823;
wire net_1326;
wire net_22376;
wire net_7488;
wire net_134;
wire net_546;
wire net_4648;
wire net_14638;
wire net_4546;
wire net_22708;
wire net_19449;
wire net_10065;
wire net_13735;
wire net_13320;
wire net_8062;
wire net_17987;
wire net_12424;
wire net_3701;
wire net_18712;
wire net_17147;
wire net_14296;
wire net_4736;
wire net_7592;
wire net_5592;
wire net_5642;
wire net_8012;
wire net_7906;
wire net_4974;
wire net_3883;
wire net_1542;
wire net_17546;
wire net_1172;
wire net_9124;
wire net_13703;
wire net_8431;
wire net_4230;
wire net_14626;
wire net_16747;
wire net_16228;
wire net_9503;
wire net_4860;
wire net_22341;
wire net_2237;
wire net_21555;
wire net_21311;
wire net_2566;
wire net_8352;
wire net_3953;
wire net_21235;
wire net_917;
wire net_3730;
wire net_21149;
wire net_19739;
wire net_2874;
wire net_10965;
wire net_8942;
wire net_14535;
wire net_9685;
wire net_2993;
wire net_18146;
wire net_10921;
wire net_3067;
wire net_13950;
wire net_10075;
wire net_4288;
wire net_21253;
wire net_323;
wire net_5402;
wire net_963;
wire net_10301;
wire net_20326;
wire net_16534;
wire net_9482;
wire net_7368;
wire net_4689;
wire net_10216;
wire net_153;
wire net_2389;
wire net_19130;
wire net_12328;
wire net_6276;
wire net_7556;
wire net_375;
wire net_562;
wire net_16692;
wire net_364;
wire net_8675;
wire net_14380;
wire net_12770;
wire net_20510;
wire net_17802;
wire net_11723;
wire net_3172;
wire net_10485;
wire net_13772;
wire net_11706;
wire net_4239;
wire net_14011;
wire net_5516;
wire net_7177;
wire net_6313;
wire net_16535;
wire net_6341;
wire net_20211;
wire net_8161;
wire net_6840;
wire net_18111;
wire net_12810;
wire net_18567;
wire net_3171;
wire net_21055;
wire net_7514;
wire net_14217;
wire net_12742;
wire net_17511;
wire net_14472;
wire net_10091;
wire net_8173;
wire net_1247;
wire net_21894;
wire net_3673;
wire net_18793;
wire net_11149;
wire net_2388;
wire net_19617;
wire net_15383;
wire net_14006;
wire net_16396;
wire net_1215;
wire net_5169;
wire net_5248;
wire net_15578;
wire net_129;
wire net_19381;
wire net_21117;
wire net_284;
wire net_6655;
wire net_12743;
wire net_439;
wire net_22379;
wire net_18322;
wire net_259;
wire net_3582;
wire net_3351;
wire net_4094;
wire net_18977;
wire net_18505;
wire net_21496;
wire net_10153;
wire net_3119;
wire net_1231;
wire net_5841;
wire net_19009;
wire net_19664;
wire x957;
wire net_6205;
wire net_815;
wire net_7875;
wire net_18951;
wire net_11304;
wire x4384;
wire net_15049;
wire net_18022;
wire net_6514;
wire net_7897;
wire net_7670;
wire net_5632;
wire net_10279;
wire net_586;
wire net_10845;
wire net_1347;
wire net_1091;
wire net_15926;
wire net_13145;
wire net_16724;
wire net_22722;
wire net_18112;
wire net_3745;
wire net_22568;
wire net_22123;
wire net_11713;
wire net_9879;
wire net_16030;
wire net_3708;
wire net_20596;
wire net_5830;
wire net_5227;
wire net_7536;
wire net_14259;
wire net_7042;
wire net_6073;
wire net_7478;
wire x2087;
wire net_21398;
wire net_22293;
wire net_16302;
wire net_16202;
wire net_2556;
wire net_8599;
wire net_19614;
wire net_16271;
wire net_3519;
wire net_2740;
wire net_14756;
wire net_7294;
wire net_20364;
wire net_672;
wire net_18548;
wire net_15015;
wire net_8834;
wire net_5212;
wire net_16938;
wire net_16914;
wire net_2027;
wire net_13761;
wire net_11680;
wire net_7021;
wire net_3610;
wire net_8963;
wire net_5784;
wire net_1953;
wire net_15177;
wire net_17630;
wire net_21167;
wire net_14295;
wire net_3925;
wire net_21548;
wire net_3847;
wire net_4473;
wire net_8230;
wire net_4582;
wire net_18339;
wire net_4547;
wire net_20460;
wire net_14205;
wire net_7819;
wire net_14455;
wire net_8954;
wire net_15154;
wire net_22143;
wire net_18837;
wire net_10136;
wire net_16776;
wire net_4640;
wire net_17520;
wire net_10926;
wire net_11602;
wire net_21765;
wire net_19432;
wire net_7071;
wire net_7982;
wire net_13264;
wire net_802;
wire net_16610;
wire net_12194;
wire net_19797;
wire net_12930;
wire net_4997;
wire net_14359;
wire net_9230;
wire net_6620;
wire net_20268;
wire net_17817;
wire net_17784;
wire net_4824;
wire x5464;
wire net_15181;
wire net_7049;
wire net_14189;
wire net_13404;
wire net_1636;
wire net_7568;
wire net_9714;
wire net_16293;
wire net_3257;
wire net_4458;
wire net_10899;
wire net_20235;
wire net_75;
wire net_10344;
wire net_10270;
wire net_21159;
wire net_16777;
wire net_1334;
wire net_18374;
wire net_10782;
wire net_20504;
wire net_757;
wire net_206;
wire net_10087;
wire net_10894;
wire net_15430;
wire net_14134;
wire net_235;
wire net_22788;
wire net_13121;
wire net_14970;
wire net_11695;
wire net_12223;
wire net_2961;
wire net_18775;
wire net_5108;
wire net_7652;
wire net_5631;
wire net_3644;
wire net_21365;
wire net_21031;
wire net_16333;
wire net_12273;
wire net_3081;
wire net_12927;
wire net_11279;
wire net_20465;
wire net_10283;
wire net_4879;
wire net_6144;
wire net_17842;
wire net_14570;
wire net_2630;
wire net_1985;
wire net_2340;
wire net_32;
wire net_21042;
wire net_14421;
wire net_14883;
wire net_20977;
wire net_2275;
wire net_10752;
wire net_3976;
wire net_9619;
wire net_10939;
wire net_22168;
wire net_13128;
wire net_841;
wire net_20062;
wire net_10803;
wire net_1750;
wire net_6411;
wire net_3346;
wire net_20901;
wire net_8269;
wire net_528;
wire net_335;
wire net_4878;
wire net_15778;
wire net_3464;
wire net_9132;
wire net_181;
wire net_9661;
wire net_6784;
wire net_15796;
wire net_12214;
wire net_3333;
wire net_11556;
wire net_6011;
wire net_10631;
wire net_9014;
wire net_13530;
wire net_6177;
wire net_3649;
wire net_2539;
wire net_18055;
wire net_17555;
wire net_21110;
wire net_6216;
wire net_386;
wire net_12680;
wire net_20797;
wire net_6150;
wire net_10051;
wire net_20642;
wire net_1790;
wire net_8166;
wire net_4103;
wire net_21762;
wire net_20165;
wire net_11221;
wire net_6130;
wire net_15719;
wire net_10583;
wire net_19145;
wire net_12718;
wire net_7573;
wire net_1709;
wire net_19814;
wire net_10981;
wire net_10080;
wire net_17294;
wire net_9698;
wire net_5707;
wire net_18404;
wire net_13622;
wire net_175;
wire net_12650;
wire net_1850;
wire net_4429;
wire net_21301;
wire net_6365;
wire net_1992;
wire net_15606;
wire net_17377;
wire net_12346;
wire net_897;
wire net_21427;
wire net_20017;
wire net_7384;
wire net_11362;
wire net_25;
wire net_2853;
wire net_10578;
wire net_2705;
wire net_21213;
wire net_5164;
wire net_615;
wire net_6712;
wire net_19319;
wire net_18104;
wire net_441;
wire net_16338;
wire net_14224;
wire net_22006;
wire net_17564;
wire net_17279;
wire net_6032;
wire net_17627;
wire net_2663;
wire net_17949;
wire net_728;
wire net_1276;
wire net_5473;
wire net_7774;
wire net_21809;
wire net_14905;
wire net_170;
wire net_17353;
wire net_15138;
wire net_16495;
wire net_5305;
wire net_20245;
wire net_10741;
wire net_22281;
wire net_20391;
wire net_17299;
wire net_17050;
wire net_16986;
wire net_14661;
wire net_21823;
wire net_3321;
wire net_15836;
wire net_15342;
wire net_15631;
wire net_13764;
wire net_708;
wire net_20750;
wire net_7685;
wire net_16667;
wire net_3216;
wire net_20261;
wire net_171;
wire net_20067;
wire net_9796;
wire net_16631;
wire net_15134;
wire net_19358;
wire net_10013;
wire net_6563;
wire net_10528;
wire net_18289;
wire net_604;
wire net_14578;
wire net_17322;
wire net_19209;
wire net_15465;
wire net_16507;
wire net_12385;
wire net_483;
wire net_15439;
wire net_16519;
wire net_1149;
wire net_9937;
wire net_8097;
wire net_15507;
wire net_16283;
wire net_16025;
wire net_15318;
wire net_2131;
wire net_6681;
wire net_16568;
wire net_5651;
wire net_13461;
wire net_12845;
wire net_18484;
wire net_15981;
wire net_19781;
wire net_7153;
wire net_19872;
wire net_13632;
wire net_11369;
wire net_20125;
wire net_2228;
wire net_12357;
wire net_786;
wire net_5141;
wire net_11801;
wire net_11564;
wire net_8998;
wire net_17308;
wire net_9470;
wire net_127;
wire net_17896;
wire net_9892;
wire net_9080;
wire net_8461;
wire net_3577;
wire net_10137;
wire net_1815;
wire net_3840;
wire net_4361;
wire net_22049;
wire net_15458;
wire net_6145;
wire net_3782;
wire net_13250;
wire net_877;
wire net_14680;
wire net_2799;
wire net_6868;
wire net_19215;
wire net_6834;
wire net_8092;
wire x151;
wire net_3734;
wire net_14135;
wire net_14524;
wire net_8021;
wire net_15714;
wire x2618;
wire net_22816;
wire net_9654;
wire net_11570;
wire net_11232;
wire net_4066;
wire net_20864;
wire net_13296;
wire net_6257;
wire net_14869;
wire net_8026;
wire net_3284;
wire net_20047;
wire net_1474;
wire net_4297;
wire net_18675;
wire net_15482;
wire net_12088;
wire net_2784;
wire net_17108;
wire net_15642;
wire x2401;
wire net_13843;
wire net_8753;
wire net_675;
wire net_21192;
wire net_8355;
wire net_2867;
wire net_3472;
wire net_9120;
wire net_10700;
wire net_7578;
wire net_22249;
wire net_1768;
wire net_20711;
wire net_16010;
wire net_19670;
wire net_12950;
wire net_7677;
wire net_20151;
wire net_304;
wire net_17968;
wire net_16427;
wire net_9791;
wire net_7326;
wire net_14967;
wire net_19515;
wire net_4347;
wire net_10551;
wire net_7731;
wire net_15431;
wire net_22471;
wire net_20443;
wire net_18660;
wire net_12731;
wire net_20258;
wire net_20112;
wire net_15517;
wire net_1316;
wire net_6845;
wire net_6545;
wire net_17311;
wire net_792;
wire net_15744;
wire net_13848;
wire net_6223;
wire net_13782;
wire net_8842;
wire net_2203;
wire net_4430;
wire net_13415;
wire net_5373;
wire net_5678;
wire net_18635;
wire x636;
wire net_18242;
wire net_219;
wire net_19127;
wire net_3609;
wire net_18125;
wire net_9976;
wire net_19608;
wire net_2476;
wire net_15791;
wire net_13798;
wire net_913;
wire net_4518;
wire net_5378;
wire net_5338;
wire net_14938;
wire net_13591;
wire net_15423;
wire net_4330;
wire net_7756;
wire net_4019;
wire net_15037;
wire net_4152;
wire net_10832;
wire net_360;
wire net_21798;
wire net_13561;
wire net_7017;
wire net_14832;
wire net_2324;
wire net_18925;
wire net_11688;
wire net_22286;
wire net_20340;
wire net_16961;
wire net_4805;
wire net_21879;
wire x2508;
wire net_13259;
wire net_3316;
wire net_10162;
wire net_3032;
wire net_9507;
wire net_17484;
wire net_1373;
wire net_1352;
wire net_2885;
wire net_16605;
wire net_10735;
wire x1146;
wire net_4696;
wire net_17127;
wire net_8814;
wire net_17087;
wire net_1187;
wire net_17079;
wire net_7408;
wire net_4988;
wire net_3206;
wire net_21745;
wire net_17163;
wire net_2858;
wire net_18696;
wire net_20706;
wire net_15470;
wire net_22731;
wire net_14806;
wire net_14703;
wire net_15004;
wire net_5569;
wire net_12234;
wire net_12047;
wire net_1442;
wire net_18410;
wire net_16400;
wire net_10042;
wire net_11544;
wire net_20224;
wire net_15188;
wire net_16968;
wire net_17411;
wire net_12298;
wire net_1894;
wire net_22428;
wire net_9645;
wire net_10694;
wire net_2431;
wire net_8213;
wire net_633;
wire net_5750;
wire net_10115;
wire net_1914;
wire net_15996;
wire net_14944;
wire net_2408;
wire net_9904;
wire net_6627;
wire net_20446;
wire net_5943;
wire net_6974;
wire net_22186;
wire net_15022;
wire net_14669;
wire net_15540;
wire net_1457;
wire net_2741;
wire net_7010;
wire net_19443;
wire net_18982;
wire net_5414;
wire net_14876;
wire net_4011;
wire net_17721;
wire net_1436;
wire net_9199;
wire net_4338;
wire net_10054;
wire net_10725;
wire net_3392;
wire net_9571;
wire net_2551;
wire net_11572;
wire net_21451;
wire net_21264;
wire net_12547;
wire net_14348;
wire net_6323;
wire net_20970;
wire net_21087;
wire net_2891;
wire net_14314;
wire net_8928;
wire net_11261;
wire net_20637;
wire net_15269;
wire net_22478;
wire net_20938;
wire net_19164;
wire net_18672;
wire net_2401;
wire net_14502;
wire net_22736;
wire net_15530;
wire net_1305;
wire net_17735;
wire net_16482;
wire net_14493;
wire net_1387;
wire net_1581;
wire net_11808;
wire net_4468;
wire net_2413;
wire net_7786;
wire net_14462;
wire net_2792;
wire net_345;
wire net_19711;
wire net_2965;
wire net_2128;
wire net_16722;
wire net_9990;
wire net_17438;
wire net_11891;
wire net_19621;
wire net_5302;
wire net_21080;
wire net_11489;
wire net_9344;
wire net_5080;
wire net_11140;
wire net_17219;
wire net_13584;
wire net_21353;
wire net_21142;
wire net_2461;
wire net_14654;
wire net_1766;
wire net_2582;
wire net_8974;
wire net_7898;
wire net_10419;
wire net_3872;
wire net_4956;
wire net_17098;
wire net_11867;
wire net_22588;
wire net_19027;
wire net_9407;
wire net_4447;
wire net_10357;
wire net_15826;
wire x1891;
wire net_10226;
wire net_13933;
wire net_9235;
wire net_8990;
wire net_14166;
wire net_8794;
wire net_20916;
wire net_9834;
wire net_12667;
wire net_13536;
wire net_13443;
wire net_17155;
wire net_10387;
wire net_1759;
wire net_12996;
wire net_15308;
wire net_12752;
wire net_3764;
wire net_19505;
wire net_12964;
wire net_18395;
wire net_11636;
wire net_2541;
wire net_12310;
wire net_3689;
wire net_12635;
wire net_533;
wire net_7436;
wire net_911;
wire net_7775;
wire net_12017;
wire net_10047;
wire net_9608;
wire net_6637;
wire net_9015;
wire net_7053;
wire net_5570;
wire net_15463;
wire net_22337;
wire net_11745;
wire net_9457;
wire net_13709;
wire net_7962;
wire net_47;
wire net_17981;
wire net_6485;
wire net_22440;
wire net_5312;
wire net_5861;
wire net_20284;
wire net_18182;
wire net_1443;
wire net_20989;
wire net_16699;
wire net_11888;
wire net_8691;
wire net_18815;
wire net_16498;
wire net_2840;
wire net_16929;
wire net_14721;
wire net_3463;
wire net_4005;
wire net_6008;
wire net_17910;
wire net_16763;
wire net_11883;
wire net_20146;
wire net_3199;
wire net_8001;
wire net_3597;
wire net_5671;
wire net_15602;
wire net_16422;
wire net_269;
wire net_5043;
wire net_3193;
wire net_20575;
wire net_3131;
wire net_10107;
wire net_12171;
wire net_20300;
wire net_3179;
wire net_1945;
wire net_10064;
wire net_7207;
wire net_10858;
wire net_19186;
wire net_4073;
wire net_5159;
wire net_1833;
wire net_8496;
wire net_2831;
wire net_3029;
wire net_18296;
wire net_9622;
wire net_7818;
wire net_5725;
wire net_12779;
wire net_19635;
wire net_8252;
wire net_18688;
wire net_6523;
wire net_17182;
wire net_22436;
wire net_5064;
wire net_20330;
wire net_6024;
wire net_17876;
wire net_21488;
wire net_11780;
wire net_12154;
wire net_15755;
wire net_8172;
wire net_19858;
wire net_7912;
wire net_16408;
wire net_5380;
wire net_22409;
wire net_10173;
wire net_8519;
wire net_5648;
wire net_14246;
wire net_18006;
wire net_11152;
wire net_16147;
wire net_11251;
wire net_10644;
wire net_3980;
wire net_10566;
wire net_1481;
wire net_10392;
wire net_7922;
wire net_16875;
wire x6544;
wire net_20513;
wire net_700;
wire net_5000;
wire net_11433;
wire net_9947;
wire net_21315;
wire net_11043;
wire net_6043;
wire net_18300;
wire net_5216;
wire net_21231;
wire net_15195;
wire net_18681;
wire net_11819;
wire net_1673;
wire net_21659;
wire net_11941;
wire net_3480;
wire net_6715;
wire net_8933;
wire net_4135;
wire net_6982;
wire net_2945;
wire net_19392;
wire net_17826;
wire net_16682;
wire net_12855;
wire net_3665;
wire net_717;
wire net_544;
wire net_15587;
wire net_12305;
wire net_10505;
wire net_15328;
wire net_8201;
wire net_9659;
wire net_20564;
wire net_20683;
wire net_18251;
wire net_3402;
wire net_2223;
wire net_6957;
wire net_8008;
wire net_2673;
wire x990;
wire net_19117;
wire net_3500;
wire net_6164;
wire net_20520;
wire net_19231;
wire net_9358;
wire net_5903;
wire net_17706;
wire net_1245;
wire net_3660;
wire net_19066;
wire net_5806;
wire net_18632;
wire net_870;
wire net_7135;
wire net_7176;
wire net_7521;
wire net_10819;
wire net_7941;
wire net_13642;
wire net_12012;
wire net_14581;
wire net_6286;
wire net_17855;
wire net_12874;
wire net_12668;
wire net_20430;
wire net_11645;
wire net_5127;
wire net_17031;
wire net_14155;
wire net_10922;
wire net_7362;
wire net_21171;
wire net_14084;
wire net_16649;
wire net_19015;
wire net_2920;
wire net_1591;
wire net_7695;
wire net_1747;
wire net_650;
wire net_19968;
wire net_20164;
wire net_15080;
wire net_9761;
wire net_19790;
wire net_597;
wire net_17852;
wire net_14065;
wire net_17321;
wire net_15767;
wire net_5984;
wire net_10482;
wire net_8272;
wire net_22082;
wire net_15109;
wire net_14281;
wire net_6336;
wire net_12481;
wire net_8889;
wire net_10853;
wire net_18161;
wire net_19026;
wire net_603;
wire net_4913;
wire net_22433;
wire net_642;
wire net_16314;
wire net_9806;
wire net_2699;
wire net_1158;
wire net_6989;
wire net_11496;
wire net_8006;
wire net_11082;
wire net_10775;
wire net_11530;
wire net_13964;
wire net_19427;
wire net_470;
wire net_2702;
wire net_430;
wire net_2834;
wire net_11659;
wire net_15255;
wire net_17442;
wire net_17346;
wire net_21900;
wire net_15903;
wire net_83;
wire net_3129;
wire net_22818;
wire net_18526;
wire net_21101;
wire net_8568;
wire net_19693;
wire net_12353;
wire net_20359;
wire net_18797;
wire net_11771;
wire net_1063;
wire net_4218;
wire net_14644;
wire net_12571;
wire net_18546;
wire net_9127;
wire net_7297;
wire net_13577;
wire net_15089;
wire net_17763;
wire net_1504;
wire net_475;
wire net_6737;
wire net_21066;
wire net_9432;
wire net_7216;
wire net_21291;
wire net_14272;
wire net_11137;
wire net_14024;
wire net_13768;
wire net_6903;
wire net_2470;
wire net_11474;
wire net_1568;
wire net_14288;
wire net_6756;
wire x629;
wire net_1526;
wire net_13860;
wire net_1884;
wire net_12341;
wire net_3919;
wire net_16920;
wire net_2646;
wire net_20658;
wire net_3936;
wire net_4364;
wire net_13198;
wire net_6645;
wire net_19983;
wire net_17538;
wire net_1360;
wire net_6344;
wire net_22023;
wire net_3364;
wire net_5316;
wire net_21238;
wire net_14420;
wire net_1364;
wire net_6003;
wire net_5050;
wire net_20292;
wire net_19677;
wire net_14727;
wire net_17550;
wire net_827;
wire net_549;
wire net_21221;
wire net_20358;
wire net_10192;
wire net_11050;
wire net_22019;
wire net_21795;
wire net_4563;
wire net_2337;
wire net_14928;
wire net_6945;
wire net_1369;
wire net_6900;
wire net_11068;
wire net_19404;
wire net_4695;
wire net_21331;
wire net_8622;
wire net_1013;
wire net_16865;
wire net_1530;
wire net_16345;
wire net_16809;
wire net_13869;
wire net_3075;
wire net_842;
wire net_11783;
wire net_2336;
wire net_1705;
wire net_14977;
wire net_6571;
wire net_9500;
wire net_11215;
wire net_21911;
wire net_8951;
wire net_21374;
wire net_6560;
wire net_19831;
wire net_10325;
wire net_8199;
wire net_20911;
wire net_3739;
wire net_8455;
wire net_492;
wire net_11392;
wire net_3678;
wire net_7234;
wire net_8797;
wire net_2639;
wire net_21481;
wire net_8071;
wire net_22675;
wire net_16085;
wire net_13370;
wire net_16702;
wire net_3695;
wire net_5450;
wire net_1327;
wire net_17650;
wire net_22549;
wire net_4968;
wire net_21907;
wire net_21563;
wire net_15337;
wire net_12734;
wire net_2248;
wire net_4971;
wire net_11532;
wire net_3866;
wire net_6772;
wire net_13473;
wire net_7787;
wire net_19264;
wire net_13223;
wire net_14548;
wire net_12024;
wire net_12920;
wire net_4300;
wire net_9578;
wire net_22076;
wire net_4776;
wire net_17676;
wire x6246;
wire net_10477;
wire net_15167;
wire net_13820;
wire net_2868;
wire net_6083;
wire net_19842;
wire net_21193;
wire net_16037;
wire net_15074;
wire net_8295;
wire net_2946;
wire net_11373;
wire net_1284;
wire net_4397;
wire net_13977;
wire net_13732;
wire net_13095;
wire net_6671;
wire net_16376;
wire net_3929;
wire net_16321;
wire net_9942;
wire net_13888;
wire net_7567;
wire net_15536;
wire net_18530;
wire net_17422;
wire net_16477;
wire net_2066;
wire net_18439;
wire net_13925;
wire net_9310;
wire net_19167;
wire net_7415;
wire net_8109;
wire net_1146;
wire net_11679;
wire net_4612;
wire net_15815;
wire net_4519;
wire net_17671;
wire net_18097;
wire net_16905;
wire net_8584;
wire net_16739;
wire net_13881;
wire net_17239;
wire net_16015;
wire net_9897;
wire net_18933;
wire net_5495;
wire net_13071;
wire net_9511;
wire net_8284;
wire net_2762;
wire net_21830;
wire net_17525;
wire net_11828;
wire net_20782;
wire net_22753;
wire net_6439;
wire net_6247;
wire net_14569;
wire net_6424;
wire net_4619;
wire net_6377;
wire net_21770;
wire net_10161;
wire net_22507;
wire net_2089;
wire net_6352;
wire net_12429;
wire net_3797;
wire net_15391;
wire net_9718;
wire net_3535;
wire net_22206;
wire net_12248;
wire net_1195;
wire net_18174;
wire net_17884;
wire net_16821;
wire net_2502;
wire net_1396;
wire net_16919;
wire net_4069;
wire net_7225;
wire net_20099;
wire net_2737;
wire net_6397;
wire x215;
wire net_5126;
wire net_18515;
wire net_18408;
wire net_14828;
wire net_12108;
wire net_2481;
wire net_21678;
wire net_4539;
wire net_15698;
wire net_15094;
wire net_19361;
wire net_10624;
wire net_22043;
wire net_8104;
wire net_14210;
wire net_17134;
wire x2230;
wire net_2617;
wire net_1060;
wire net_22717;
wire net_12699;
wire net_4846;
wire net_20968;
wire net_12101;
wire net_1715;
wire net_19341;
wire net_15961;
wire net_9913;
wire net_14842;
wire net_7583;
wire net_9234;
wire net_15221;
wire net_14557;
wire net_6577;
wire net_1216;
wire net_19578;
wire net_4599;
wire net_14583;
wire net_2815;
wire net_15040;
wire net_3785;
wire net_18994;
wire net_11240;
wire net_1271;
wire net_1086;
wire net_19347;
wire net_22648;
wire net_18465;
wire net_9593;
wire net_10978;
wire net_13453;
wire net_1197;
wire net_7613;
wire net_5744;
wire net_5858;
wire net_21585;
wire net_11752;
wire net_21667;
wire net_18018;
wire net_576;
wire net_8932;
wire net_1654;
wire net_8438;
wire net_3005;
wire net_11183;
wire net_12902;
wire net_19344;
wire net_10679;
wire net_21735;
wire net_11272;
wire net_725;
wire net_22181;
wire net_3931;
wire net_17591;
wire net_22555;
wire net_21308;
wire net_18369;
wire net_6183;
wire net_21607;
wire net_14766;
wire net_894;
wire net_16219;
wire net_13914;
wire net_10545;
wire net_17718;
wire net_18496;
wire net_1423;
wire net_13012;
wire net_2902;
wire net_1871;
wire net_517;
wire net_628;
wire net_22114;
wire net_18030;
wire net_3494;
wire net_6600;
wire net_21047;
wire net_12123;
wire net_10377;
wire net_21506;
wire net_19093;
wire net_14018;
wire net_21320;
wire net_10204;
wire net_9555;
wire net_9036;
wire x5568;
wire x1275;
wire net_17482;
wire net_22306;
wire net_17691;
wire net_6406;
wire net_10322;
wire net_1289;
wire net_19275;
wire net_3138;
wire net_14858;
wire x2571;
wire net_11982;
wire net_20527;
wire net_15786;
wire net_13377;
wire net_12867;
wire net_6922;
wire net_17061;
wire net_19460;
wire net_11162;
wire net_5895;
wire net_21411;
wire net_12446;
wire net_5876;
wire net_20185;
wire net_22263;
wire net_2723;
wire net_17365;
wire net_15144;
wire net_5157;
wire net_13504;
wire net_2552;
wire net_3229;
wire net_1001;
wire net_13778;
wire net_781;
wire net_3765;
wire net_8479;
wire net_20836;
wire net_15323;
wire net_13063;
wire net_21242;
wire net_5241;
wire net_7506;
wire net_5967;
wire net_6818;
wire net_16677;
wire net_13188;
wire net_22710;
wire net_16353;
wire net_185;
wire net_7357;
wire net_17195;
wire net_16194;
wire net_22366;
wire net_14687;
wire net_16540;
wire net_4321;
wire net_4631;
wire net_18452;
wire net_1015;
wire net_2980;
wire net_14685;
wire net_16717;
wire net_9863;
wire net_22693;
wire net_19247;
wire x2240;
wire net_20774;
wire net_9772;
wire net_11964;
wire net_5794;
wire net_14748;
wire net_7766;
wire net_17489;
wire net_11759;
wire net_6856;
wire net_20485;
wire net_15660;
wire net_2146;
wire net_405;
wire net_11927;
wire net_19656;
wire net_1111;
wire net_11614;
wire net_2651;
wire net_4281;
wire net_8259;
wire net_3971;
wire net_16841;
wire net_16224;
wire net_3155;
wire net_7969;
wire net_19486;
wire net_20587;
wire net_831;
wire net_4728;
wire net_5442;
wire net_21826;
wire net_451;
wire net_1234;
wire net_750;
wire net_12558;
wire net_20437;
wire net_7835;
wire net_9746;
wire net_16411;
wire net_21654;
wire net_13027;
wire net_12797;
wire net_7274;
wire net_17866;
wire net_17274;
wire net_14641;
wire net_11459;
wire net_8571;
wire net_5915;
wire net_21658;
wire net_19056;
wire net_18738;
wire net_5184;
wire net_21478;
wire net_17401;
wire net_16189;
wire net_5788;
wire net_11920;
wire net_8472;
wire net_773;
wire net_4759;
wire net_11770;
wire net_9590;
wire net_20942;
wire net_19900;
wire net_16653;
wire net_11796;
wire net_11622;
wire net_8537;
wire net_12098;
wire net_15976;
wire net_3727;
wire net_15887;
wire net_13986;
wire net_6766;
wire net_13269;
wire net_6355;
wire net_5052;
wire net_14400;
wire net_9997;
wire x5505;
wire net_8305;
wire net_54;
wire net_14091;
wire net_4205;
wire net_834;
wire net_10298;
wire net_694;
wire net_13615;
wire net_13556;
wire net_18528;
wire net_13794;
wire net_5925;
wire net_9950;
wire net_7609;
wire net_8778;
wire net_8946;
wire net_8409;
wire net_1570;
wire net_13385;
wire net_4645;
wire net_11100;
wire net_17415;
wire net_12204;
wire net_9499;
wire net_11228;
wire net_111;
wire net_7320;
wire net_15811;
wire net_20382;
wire net_8779;
wire net_124;
wire net_252;
wire net_10497;
wire net_7693;
wire net_14897;
wire net_2399;
wire net_20541;
wire net_19951;
wire net_16325;
wire net_14508;
wire net_901;
wire net_6267;
wire net_7846;
wire net_3425;
wire net_16780;
wire net_410;
wire net_20082;
wire net_22493;
wire net_8134;
wire net_21343;
wire net_4243;
wire net_14940;
wire net_10539;
wire net_9136;
wire net_19846;
wire net_6798;
wire net_6607;
wire net_12470;
wire net_22417;
wire net_18956;
wire net_7886;
wire x5328;
wire net_17473;
wire net_20416;
wire net_7824;
wire net_2603;
wire net_5910;
wire net_1132;
wire net_14144;
wire net_5880;
wire net_10351;
wire net_2442;
wire net_20621;
wire net_22271;
wire net_3026;
wire net_7743;
wire net_13749;
wire net_12317;
wire net_9410;
wire net_5760;
wire net_18869;
wire net_5923;
wire net_22356;
wire net_21024;
wire net_2356;
wire net_3288;
wire net_971;
wire net_22533;
wire net_8194;
wire net_20994;
wire net_11734;
wire net_19702;
wire net_2184;
wire net_18278;
wire net_11824;
wire net_554;
wire net_16894;
wire net_14544;
wire net_13625;
wire net_18765;
wire net_4653;
wire net_21705;
wire net_14232;
wire net_11187;
wire net_8704;
wire net_3740;
wire net_15278;
wire net_14221;
wire net_8317;
wire net_19947;
wire net_6306;
wire net_584;
wire net_13753;
wire net_10446;
wire net_12656;
wire net_21070;
wire net_2411;
wire net_13104;
wire net_19726;
wire net_11511;
wire net_165;
wire net_9226;
wire net_16055;
wire net_14794;
wire net_18585;
wire net_3438;
wire net_3824;
wire net_21093;
wire net_8789;
wire net_4440;
wire net_8576;
wire net_20427;
wire net_18847;
wire net_13612;
wire net_10170;
wire net_21775;
wire net_16215;
wire net_12970;
wire net_3823;
wire net_21872;
wire net_20420;
wire net_9886;
wire net_17888;
wire net_8600;
wire net_18970;
wire net_22057;
wire net_16832;
wire net_17795;
wire net_9365;
wire net_13573;
wire net_3859;
wire net_8044;
wire net_21576;
wire net_15350;
wire net_7885;
wire net_21996;
wire net_3803;
wire net_17664;
wire net_8607;
wire net_11284;
wire net_16099;
wire net_15395;
wire net_14338;
wire net_20024;
wire net_14592;
wire net_8880;
wire net_8592;
wire net_7707;
wire net_3334;
wire net_6789;
wire net_3224;
wire net_21272;
wire net_1719;
wire net_17740;
wire net_15613;
wire net_15854;
wire x1471;
wire net_19695;
wire net_16068;
wire net_5715;
wire net_11562;
wire net_19884;
wire net_15739;
wire net_11464;
wire net_15426;
wire net_8786;
wire net_17917;
wire net_14448;
wire net_8034;
wire net_11598;
wire net_2440;
wire net_19683;
wire net_9386;
wire net_18995;
wire net_16077;
wire net_6809;
wire net_14043;
wire net_12800;
wire net_1379;
wire net_1322;
wire net_14437;
wire net_9538;
wire net_22373;
wire net_8526;
wire net_20132;
wire net_12143;
wire net_10373;
wire net_1301;
wire net_12066;
wire net_14258;
wire net_12487;
wire net_8749;
wire net_7596;
wire net_12756;
wire net_7247;
wire net_6932;
wire net_7116;
wire net_16575;
wire net_20553;
wire net_17456;
wire net_426;
wire net_5203;
wire net_16298;
wire net_6095;
wire net_19935;
wire net_14511;
wire net_414;
wire net_7793;
wire net_17611;
wire net_1048;
wire net_18249;
wire net_3048;
wire net_799;
wire net_5102;
wire net_21851;
wire net_5576;
wire net_18057;
wire net_20854;
wire net_15367;
wire net_22667;
wire net_20749;
wire net_5737;
wire net_12588;
wire net_2014;
wire net_21603;
wire net_16884;
wire net_22517;
wire net_19666;
wire net_16278;
wire x3354;
wire net_6747;
wire net_21781;
wire net_13487;
wire net_5999;
wire net_20548;
wire net_22088;
wire net_9845;
wire net_16952;
wire net_4742;
wire net_2454;
wire net_8917;
wire net_8716;
wire net_21448;
wire net_4761;
wire net_14709;
wire net_17547;
wire x2914;
wire net_22551;
wire net_18151;
wire net_7616;
wire net_15701;
wire net_16582;
wire net_6016;
wire net_18498;
wire net_17603;
wire net_10140;
wire net_15972;
wire net_12621;
wire net_247;
wire net_19553;
wire net_19321;
wire net_21886;
wire net_14630;
wire net_21632;
wire net_22362;
wire net_21984;
wire net_3413;
wire net_70;
wire net_14430;
wire net_9742;
wire net_20626;
wire net_8619;
wire net_19917;
wire net_12627;
wire net_1934;
wire net_14180;
wire net_13740;
wire net_12513;
wire net_6235;
wire net_11327;
wire net_1848;
wire net_639;
wire net_4724;
wire net_9583;
wire net_18363;
wire net_12309;
wire net_5697;
wire net_1238;
wire net_14923;
wire net_13697;
wire net_14074;
wire net_7599;
wire net_9483;
wire net_1033;
wire net_20928;
wire net_10604;
wire net_5560;
wire net_12458;
wire net_11333;
wire net_8333;
wire net_13149;
wire net_22267;
wire net_20680;
wire net_15163;
wire net_12005;
wire net_12302;
wire net_3107;
wire net_7069;
wire net_1686;
wire net_11860;
wire net_11481;
wire net_10686;
wire net_21433;
wire net_10263;
wire x16;
wire net_367;
wire net_3303;
wire net_17861;
wire net_17747;
wire net_6296;
wire net_19228;
wire net_20771;
wire net_10061;
wire net_1842;
wire net_19499;
wire net_9849;
wire net_13037;
wire net_8774;
wire net_3957;
wire net_1180;
wire net_20119;
wire net_8561;
wire net_1627;
wire net_10235;
wire net_5869;
wire net_20195;
wire net_2002;
wire net_1069;
wire net_20089;
wire net_2022;
wire net_9932;
wire net_12014;
wire net_5406;
wire net_18591;
wire net_2385;
wire net_3431;
wire x1373;
wire net_17118;
wire net_5829;
wire net_3565;
wire net_7009;
wire net_1416;
wire net_7656;
wire net_13484;
wire net_18167;
wire net_6065;
wire net_20228;
wire net_2433;
wire net_21400;
wire net_15111;
wire net_6726;
wire net_4029;
wire net_93;
wire net_1601;
wire net_6614;
wire net_4087;
wire net_4255;
wire net_9854;
wire net_17659;
wire net_13437;
wire net_8866;
wire net_348;
wire net_7398;
wire net_9667;
wire net_626;
wire net_10796;
wire net_15260;
wire net_20980;
wire net_5068;
wire net_22050;
wire net_16116;
wire net_11257;
wire net_1809;
wire net_686;
wire net_17904;
wire net_1615;
wire net_16521;
wire net_17266;
wire net_14037;
wire net_17192;
wire net_7859;
wire net_17495;
wire net_4578;
wire net_2112;
wire net_5072;
wire net_14505;
wire net_1828;
wire net_16063;
wire net_1466;
wire net_5320;
wire net_10438;
wire net_16182;
wire net_11268;
wire x4706;
wire net_157;
wire net_17074;
wire net_6695;
wire net_9006;
wire net_7759;
wire net_18139;
wire net_1205;
wire net_11627;
wire net_8154;
wire net_6978;
wire net_466;
wire net_9612;
wire net_1179;
wire net_18232;
wire net_21199;
wire net_15844;
wire net_15231;
wire net_18720;
wire net_7833;
wire net_13057;
wire net_16709;
wire net_11021;
wire net_16289;
wire net_1610;
wire net_3569;
wire net_6814;
wire net_13236;
wire net_4246;
wire net_8893;
wire net_4020;
wire net_16870;
wire net_21136;
wire net_8389;
wire net_4453;
wire net_17282;
wire net_16467;
wire net_15593;
wire net_11018;
wire net_20778;
wire net_7118;
wire net_644;
wire net_20455;
wire net_13495;
wire net_12111;
wire net_12063;
wire net_852;
wire net_11917;
wire net_11035;
wire net_15118;
wire net_14771;
wire net_7391;
wire net_8904;
wire net_8416;
wire net_8382;
wire net_11404;
wire net_18706;
wire net_14690;
wire net_14284;
wire net_10128;
wire net_8685;
wire net_20794;
wire net_11492;
wire net_9491;
wire net_8555;
wire x1845;
wire net_11410;
wire net_5871;
wire net_14061;
wire net_15243;
wire net_1693;
wire net_10707;
wire net_8853;
wire net_3779;
wire net_4252;
wire net_2068;
wire net_22698;
wire net_17880;
wire net_14659;
wire net_3705;
wire net_5907;
wire net_11821;
wire net_19864;
wire net_16673;
wire net_5930;
wire net_6371;
wire net_8939;
wire net_17584;
wire net_15692;
wire net_314;
wire net_5395;
wire net_17637;
wire net_19891;
wire net_19115;
wire net_15301;
wire net_18615;
wire net_11381;
wire net_9765;
wire net_18623;
wire net_21180;
wire net_12033;
wire net_19120;
wire net_14964;
wire net_8442;
wire net_4669;
wire net_13791;
wire net_5460;
wire net_12479;
wire net_4286;
wire net_9872;
wire net_3484;
wire net_16518;
wire net_945;
wire net_6532;
wire net_4380;
wire net_6971;
wire net_12266;
wire net_2101;
wire net_7738;
wire net_19086;
wire net_6863;
wire net_18572;
wire net_22466;
wire net_19172;
wire net_11451;
wire net_8875;
wire net_8376;
wire net_15246;
wire net_19686;
wire net_6582;
wire net_5800;
wire net_5601;
wire net_15312;
wire net_13426;
wire net_16851;
wire net_12251;
wire net_8808;
wire net_6340;
wire net_13256;
wire net_10516;
wire net_18823;
wire net_9099;
wire net_5174;
wire net_11343;
wire net_8943;
wire net_1784;
wire net_1296;
wire net_17253;
wire net_15738;
wire net_16823;
wire net_13081;
wire net_4326;
wire net_10245;
wire net_7159;
wire net_10762;
wire net_9735;
wire net_2424;
wire net_22455;
wire net_1968;
wire net_15364;
wire net_10746;
wire net_10407;
wire net_12291;
wire net_4488;
wire net_5092;
wire net_5295;
wire net_18534;
wire net_7713;
wire net_19283;
wire net_2507;
wire net_17024;
wire net_16791;
wire net_9633;
wire net_22481;
wire net_19364;
wire net_17335;
wire net_13908;
wire net_2685;
wire net_20617;
wire net_8340;
wire net_14264;
wire net_2898;
wire net_6197;
wire net_1391;
wire net_9334;
wire net_14933;
wire net_9926;
wire net_5132;
wire net_18203;
wire net_10304;
wire net_17235;
wire net_14847;
wire net_1772;
wire net_14552;
wire net_3529;
wire net_6128;
wire net_5437;
wire net_21995;
wire net_2498;
wire net_381;
wire net_9144;
wire net_6574;
wire net_6889;
wire net_10710;
wire net_15891;
wire net_3783;
wire net_22527;
wire net_1857;
wire net_7445;
wire net_11586;
wire net_11010;
wire net_19526;
wire net_12059;
wire net_6109;
wire net_15554;
wire net_14414;
wire net_9883;
wire net_17993;
wire net_16751;
wire net_1557;
wire net_6843;
wire x3701;
wire net_1514;
wire net_3852;
wire net_7668;
wire net_13072;
wire net_6825;
wire net_13874;
wire net_3092;
wire net_14407;
wire net_9209;
wire net_8802;
wire net_6995;
wire net_19103;
wire net_20031;
wire net_22746;
wire net_13240;
wire net_12241;
wire net_500;
wire net_5357;
wire net_1906;
wire net_17687;
wire net_9094;
wire net_20848;
wire net_8056;
wire net_5660;
wire net_15410;
wire net_22745;
wire net_11967;
wire net_19562;
wire net_22802;
wire net_14197;
wire net_10911;
wire net_14120;
wire net_17822;
wire net_14717;
wire net_10130;
wire net_11974;
wire net_16992;
wire net_19733;
wire net_4401;
wire net_18355;
wire net_15271;
wire net_3632;
wire net_2189;
wire net_2057;
wire net_1124;
wire net_13945;
wire net_7645;
wire net_16816;
wire net_21474;
wire net_13737;
wire x1176;
wire net_20473;
wire x2019;
wire net_5960;
wire net_5615;
wire net_143;
wire net_12434;
wire net_22767;
wire net_190;
wire net_4964;
wire net_1447;
wire net_1929;
wire net_9423;
wire net_19649;
wire net_3493;
wire net_2061;
wire net_13466;
wire net_5288;
wire net_15878;
wire net_13956;
wire net_14030;
wire net_13910;
wire net_13727;
wire net_14780;
wire net_22593;
wire net_13710;
wire net_1895;
wire net_5360;
wire net_509;
wire net_14983;
wire net_4975;
wire net_16157;
wire net_19559;
wire net_9983;
wire net_211;
wire net_21485;
wire net_16248;
wire net_22198;
wire net_13430;
wire net_10079;
wire net_6752;
wire net_14564;
wire net_19757;
wire net_18001;
wire net_5771;
wire net_13541;
wire net_3941;
wire net_6630;
wire net_12604;
wire net_22244;
wire net_20632;
wire net_17359;
wire net_8645;
wire net_2233;
wire net_22796;
wire net_22095;
wire net_2033;
wire net_18061;
wire net_12726;
wire net_12091;
wire net_8487;
wire net_15710;
wire net_2123;
wire net_21693;
wire net_10811;
wire net_12784;
wire net_19847;
wire net_12360;
wire net_9049;
wire net_5970;
wire net_16554;
wire net_2532;
wire net_18468;
wire net_12785;
wire net_13851;
wire net_11112;
wire net_1864;
wire net_20611;
wire net_15441;
wire net_14917;
wire net_11725;
wire net_6156;
wire net_12840;
wire net_2518;
wire net_14604;
wire net_6950;
wire net_10663;
wire net_4062;
wire net_22543;
wire net_21383;
wire net_17014;
wire net_12284;
wire net_14353;
wire net_7953;
wire x1330;
wire net_1646;
wire net_4115;
wire net_11437;
wire net_2776;
wire net_18433;
wire net_3389;
wire net_12938;
wire net_1562;
wire net_16743;
wire net_15225;
wire net_2522;
wire net_4178;
wire net_7267;
wire net_8671;
wire net_20316;
wire net_17928;
wire net_13878;
wire net_136;
wire net_12987;
wire net_1524;
wire net_16398;
wire net_18385;
wire net_10022;
wire net_9396;
wire net_17943;
wire net_15686;
wire net_12531;
wire net_9785;
wire net_11670;
wire net_15864;
wire net_16572;
wire net_6461;
wire net_21011;
wire net_2511;
wire net_2626;
wire net_2115;
wire net_4110;
wire net_4317;
wire net_2299;
wire net_21592;
wire net_21178;
wire net_9307;
wire net_10612;
wire net_16049;
wire x2659;
wire net_7123;
wire net_19806;
wire net_17837;
wire net_19604;
wire net_21051;
wire net_21018;
wire net_1405;
wire net_7726;
wire net_10072;
wire net_19630;
wire net_22778;
wire net_17902;
wire net_13518;
wire net_10881;
wire net_6555;
wire net_21461;
wire net_20335;
wire x622;
wire net_15102;
wire net_20805;
wire net_716;
wire net_5147;
wire net_13273;
wire net_13200;
wire net_10489;
wire net_11445;
wire net_1269;
wire net_19267;
wire net_16846;
wire net_13757;
wire net_8630;
wire net_20534;
wire net_3533;
wire net_3715;
wire net_5400;
wire net_36;
wire net_21558;
wire net_11805;
wire net_12406;
wire net_19894;
wire net_4293;
wire net_9176;
wire net_666;
wire net_20200;
wire net_19654;
wire net_13776;
wire net_4809;
wire net_11308;
wire net_18305;
wire net_12706;
wire net_12184;
wire net_6212;
wire net_9702;
wire net_15125;
wire net_3946;
wire net_10596;
wire net_19828;
wire net_19516;
wire net_19418;
wire x1238;
wire net_5522;
wire net_6319;
wire net_7636;
wire net_9024;
wire net_9824;
wire net_1657;
wire net_6063;
wire net_3084;
wire net_10689;
wire net_10863;
wire net_19010;
wire net_18894;
wire net_18477;
wire net_17380;
wire net_9859;
wire net_3994;
wire net_18790;
wire net_21868;
wire net_11764;
wire net_22257;
wire net_14213;
wire net_13645;
wire net_1976;
wire net_8510;
wire net_3169;
wire net_14734;
wire net_5647;
wire net_3792;
wire net_2758;
wire net_9972;
wire net_21145;
wire net_1826;
wire net_18327;
wire net_14634;
wire net_22635;
wire net_16531;
wire net_4609;
wire net_10337;
wire net_16860;
wire net_16160;
wire net_2142;
wire net_22345;
wire net_11841;
wire net_20618;
wire net_15335;
wire net_7332;
wire net_920;
wire net_22385;
wire net_22705;
wire net_3009;
wire net_12980;
wire net_5596;
wire net_21375;
wire net_15653;
wire net_4226;
wire net_820;
wire net_7137;
wire net_18656;
wire net_11249;
wire net_16530;
wire net_15765;
wire x697;
wire net_21966;
wire net_18901;
wire net_13447;
wire net_6137;
wire net_13465;
wire net_5959;
wire net_9681;
wire net_566;
wire net_5063;
wire net_7519;
wire x6110;
wire net_9768;
wire net_21356;
wire net_19296;
wire net_13173;
wire net_20051;
wire net_13811;
wire net_4735;
wire net_17771;
wire x2985;
wire net_18788;
wire net_17696;
wire net_2108;
wire net_2529;
wire net_19038;
wire net_6044;
wire net_4685;
wire net_19748;
wire net_4732;
wire net_9751;
wire net_8390;
wire net_5979;
wire net_7551;
wire net_19953;
wire net_11810;
wire net_20653;
wire net_18985;
wire net_18024;
wire net_14279;
wire net_21815;
wire net_4235;
wire net_21644;
wire net_20334;
wire net_19592;
wire net_15570;
wire net_14117;
wire net_11871;
wire net_14990;
wire net_13379;
wire net_21614;
wire net_9452;
wire net_4117;
wire net_1357;
wire net_15875;
wire net_13990;
wire net_3637;
wire net_5554;
wire net_19875;
wire net_18564;
wire net_17188;
wire net_21647;
wire net_14476;
wire net_8668;
wire net_18966;
wire net_4604;
wire net_7489;
wire net_6558;
wire net_12598;
wire net_419;
wire net_12463;
wire net_16974;
wire net_5658;
wire net_936;
wire net_15400;
wire net_9259;
wire net_8066;
wire net_7808;
wire net_17006;
wire net_819;
wire net_10969;
wire net_11954;
wire net_8241;
wire net_14121;
wire net_9106;
wire net_13653;
wire net_19583;
wire net_21963;
wire net_4070;
wire net_18256;
wire net_9327;
wire net_19251;
wire net_11173;
wire net_6272;
wire net_3141;
wire net_22611;
wire net_1670;
wire net_15939;
wire net_4274;
wire net_3265;
wire net_2801;
wire net_2932;
wire net_4951;
wire net_22201;
wire net_13342;
wire net_12420;
wire net_7928;
wire net_8277;
wire net_5812;
wire net_1264;
wire net_8077;
wire net_20841;
wire net_9852;
wire net_19855;
wire net_9300;
wire net_3148;
wire net_1229;
wire net_6316;
wire net_16148;
wire net_12746;
wire net_14385;
wire net_6277;
wire net_19332;
wire net_16125;
wire net_766;
wire net_1153;
wire net_21257;
wire net_3014;
wire net_8469;
wire net_10961;
wire net_9102;
wire net_20056;
wire net_9252;
wire net_6734;
wire net_5692;
wire net_14241;
wire x856;
wire net_18762;
wire net_18295;
wire net_3454;
wire net_5113;
wire net_9533;
wire net_13682;
wire net_12333;
wire net_3729;
wire net_20958;
wire net_10465;
wire net_18942;
wire net_14347;
wire net_9589;
wire net_2251;
wire net_12914;
wire net_8898;
wire net_9623;
wire net_19861;
wire net_7439;
wire net_10418;
wire net_9727;
wire net_955;
wire net_2585;
wire net_15670;
wire net_15952;
wire net_1996;
wire net_7046;
wire net_13635;
wire net_1029;
wire net_22704;
wire net_22344;
wire net_15702;
wire net_13664;
wire net_9812;
wire net_20881;
wire net_9066;
wire net_12566;
wire net_19101;
wire net_12762;
wire net_2986;
wire net_3162;
wire net_4034;
wire net_4791;
wire net_20155;
wire x1580;
wire net_13082;
wire net_11937;
wire net_3510;
wire net_16624;
wire net_11848;
wire net_10492;
wire net_3180;
wire net_3249;
wire net_20742;
wire net_15277;
wire net_14002;
wire net_6157;
wire net_16006;
wire net_734;
wire net_14152;
wire net_12564;
wire net_2544;
wire net_19767;
wire net_15801;
wire net_15957;
wire net_21742;
wire net_3186;
wire net_11314;
wire x2260;
wire net_8177;
wire net_21075;
wire net_13895;
wire net_20431;
wire net_16942;
wire net_21228;
wire net_5277;
wire net_17770;
wire net_14730;
wire net_7269;
wire net_4372;
wire net_15398;
wire net_1076;
wire net_14051;
wire net_10168;
wire net_8234;
wire net_10399;
wire net_9711;
wire net_4352;
wire net_15647;
wire net_19280;
wire net_681;
wire net_19303;
wire net_7346;
wire net_18864;
wire net_13136;
wire net_6533;
wire net_5252;
wire net_17260;
wire net_146;
wire net_9562;
wire net_20822;
wire net_20720;
wire net_16250;
wire net_5752;
wire net_21186;
wire net_4594;
wire net_15009;
wire net_4454;
wire net_6290;
wire net_20896;
wire x4980;
wire net_4624;
wire net_21289;
wire net_11522;
wire net_7621;
wire net_428;
wire net_16689;
wire net_9675;
wire net_10557;
wire net_14816;
wire net_7780;
wire net_20306;
wire net_4666;
wire net_16656;
wire net_2888;
wire net_17082;
wire net_12884;
wire net_22055;
wire net_14362;
wire net_888;
wire net_21574;
wire net_13066;
wire net_10772;
wire net_13212;
wire net_11298;
wire net_11095;
wire net_9526;
wire net_5191;
wire net_19506;
wire net_18833;
wire net_22821;
wire net_8480;
wire net_20303;
wire net_18378;
wire net_10513;
wire net_1023;
wire net_4814;
wire net_5233;
wire net_7499;
wire net_3623;
wire net_301;
wire net_2360;
wire net_3617;
wire net_7432;
wire net_1343;
wire net_18729;
wire net_7147;
wire net_2285;
wire net_19450;
wire net_16704;
wire net_12690;
wire net_7355;
wire net_16175;
wire net_20789;
wire net_16555;
wire net_590;
wire net_3879;
wire net_21622;
wire net_3240;
wire net_15150;
wire net_8229;
wire net_9342;
wire net_12135;
wire net_10094;
wire net_4194;
wire net_12361;
wire net_5464;
wire net_16136;
wire net_8335;
wire net_8530;
wire net_15059;
wire net_10145;
wire net_21267;
wire net_1736;
wire net_12807;
wire net_12258;
wire net_9814;
wire net_11660;
wire net_6947;
wire net_16363;
wire net_10314;
wire net_20687;
wire net_10574;
wire net_4148;
wire net_18854;
wire net_9155;
wire net_5048;
wire net_7869;
wire net_1669;
wire net_11505;
wire net_12408;
wire net_14096;
wire net_1041;
wire net_7628;
wire net_6385;
wire net_16804;
wire net_14027;
wire net_2950;
wire net_22679;
wire net_6056;
wire net_6108;
wire net_5851;
wire net_14350;
wire net_18340;
wire net_17051;
wire net_4778;
wire net_11211;
wire net_17207;
wire net_13159;
wire net_22327;
wire net_16638;
wire net_2364;
wire net_942;
wire net_12822;
wire net_8763;
wire net_22171;
wire net_22235;
wire net_17241;
wire net_17341;
wire net_17750;
wire net_13658;
wire net_10917;
wire net_6436;
wire net_15201;
wire net_1494;
wire net_18731;
wire net_4415;
wire net_18129;
wire net_2154;
wire net_1726;
wire net_5527;
wire net_4123;
wire net_7082;
wire net_5705;
wire net_16949;
wire net_12165;
wire net_3298;
wire net_3099;
wire net_17647;
wire net_10658;
wire net_16232;
wire net_15065;
wire net_19236;
wire net_6339;
wire net_7380;
wire net_1794;
wire net_18085;
wire net_9363;
wire net_12508;
wire net_6503;
wire net_5536;
wire net_1022;
wire net_4638;
wire net_22604;
wire net_11129;
wire net_6110;
wire net_16426;
wire net_21891;
wire net_8182;
wire net_15894;
wire net_16199;
wire net_17030;
wire x5957;
wire net_13960;
wire net_9270;
wire net_17446;
wire net_15401;
wire net_20664;
wire net_18122;
wire net_16089;
wire net_13152;
wire net_12439;
wire net_22576;
wire net_14673;
wire net_1122;
wire net_4911;
wire net_15679;
wire net_6228;
wire net_5505;
wire net_19465;
wire net_8540;
wire net_4534;
wire net_6252;
wire net_17206;
wire net_18692;
wire net_17303;
wire net_6491;
wire net_13898;
wire net_4713;
wire net_22646;
wire net_9709;
wire net_18091;
wire net_9002;
wire net_17284;
wire net_21711;
wire net_17434;
wire net_4307;
wire net_8292;
wire net_5513;
wire net_21533;
wire net_8248;
wire net_3962;
wire net_21412;
wire net_11834;
wire net_4553;
wire net_19545;
wire net_275;
wire net_12641;
wire net_9486;
wire net_4831;
wire net_2914;
wire net_22175;
wire net_15050;
wire net_11366;
wire net_2590;
wire net_22765;
wire net_10841;
wire net_7280;
wire net_13293;
wire net_13351;
wire net_1137;
wire net_7424;
wire net_4830;
wire net_5036;
wire net_12860;
wire net_13909;
wire net_4865;
wire net_16266;
wire net_11765;
wire net_9955;
wire net_14370;
wire net_11978;
wire net_11193;
wire net_12581;
wire net_11895;
wire net_5622;
wire net_18805;
wire net_20829;
wire net_3357;
wire net_9467;
wire net_14054;
wire net_21716;
wire net_9694;
wire net_8425;
wire net_17620;
wire net_8298;
wire net_16800;
wire net_19575;
wire net_21467;
wire net_14199;
wire net_14672;
wire net_943;
wire net_10413;
wire net_16736;
wire net_4392;
wire net_11330;
wire net_9435;
wire net_13088;
wire net_2542;
wire net_19224;
wire net_20154;
wire net_21196;
wire net_7594;
wire net_11996;
wire net_12537;
wire net_18035;
wire net_17009;
wire net_17642;
wire net_2256;
wire net_4934;
wire net_17779;
wire net_12809;
wire net_4122;
wire net_4315;
wire net_17418;
wire net_21222;
wire net_18365;
wire net_8503;
wire net_4996;
wire net_11190;
wire net_16442;
wire net_1064;
wire net_14016;
wire net_21674;
wire net_20738;
wire net_10165;
wire net_6227;
wire net_7173;
wire net_19157;
wire net_17819;
wire net_12907;
wire net_15734;
wire net_9784;
wire net_12704;
wire net_20172;
wire net_13544;
wire net_19338;
wire net_7191;
wire net_10988;
wire net_17175;
wire net_6037;
wire net_10554;
wire net_19069;
wire net_7283;
wire net_14609;
wire net_5627;
wire net_3817;
wire net_9441;
wire net_3281;
wire net_10659;
wire net_3949;
wire net_8185;
wire net_10215;
wire net_16171;
wire net_6231;
wire net_3434;
wire net_3818;
wire net_18067;
wire net_3756;
wire net_9464;
wire net_19685;
wire net_18341;
wire net_4169;
wire net_17059;
wire net_7845;
wire net_13451;
wire net_21620;
wire net_9957;
wire net_742;
wire net_11979;
wire net_19198;
wire net_5139;
wire net_20279;
wire net_18906;
wire net_6384;
wire net_18850;
wire net_12976;
wire net_16265;
wire net_7092;
wire net_2830;
wire net_18084;
wire net_4509;
wire net_22216;
wire net_21814;
wire net_883;
wire net_11605;
wire net_13476;
wire net_8124;
wire net_4108;
wire net_2957;
wire net_9970;
wire net_446;
wire net_1712;
wire net_20343;
wire net_3063;
wire net_1499;
wire net_21640;
wire x1765;
wire net_3295;
wire net_8242;
wire net_15060;
wire net_4379;
wire net_14985;
wire net_18943;
wire net_10000;
wire net_15141;
wire net_6114;
wire net_2303;
wire net_1735;
wire net_2210;
wire net_2176;
wire net_8249;
wire net_13191;
wire net_16592;
wire net_8563;
wire net_11933;
wire net_16130;
wire net_997;
wire net_17466;
wire net_10837;
wire net_12243;
wire net_11060;
wire net_256;
wire net_8762;
wire net_7490;
wire net_5797;
wire net_10931;
wire net_21719;
wire net_16104;
wire net_12891;
wire net_4835;
wire net_16662;
wire net_5342;
wire net_7463;
wire net_11124;
wire net_13216;
wire net_3987;
wire net_6557;
wire net_19737;
wire net_8468;
wire net_21324;
wire net_2219;
wire net_18418;
wire net_7343;
wire net_11166;
wire net_20139;
wire net_17264;
wire net_5680;
wire net_15657;
wire net_16176;
wire net_22107;
wire net_1876;
wire net_7483;
wire net_13130;
wire net_15567;
wire net_20945;
wire net_20414;
wire net_14611;
wire net_20179;
wire net_130;
wire net_9810;
wire net_5116;
wire net_15218;
wire net_19958;
wire net_369;
wire net_12051;
wire net_12709;
wire net_15756;
wire net_4358;
wire net_7543;
wire net_9835;
wire net_20990;
wire net_10495;
wire net_7959;
wire net_3935;
wire net_11290;
wire net_15551;
wire net_2809;
wire net_15273;
wire net_780;
wire net_3586;
wire net_3184;
wire net_19308;
wire net_6812;
wire net_12226;
wire x3635;
wire net_15979;
wire net_20311;
wire net_9272;
wire net_10095;
wire net_21182;
wire net_5263;
wire net_155;
wire net_11350;
wire net_9301;
wire net_11357;
wire net_12555;
wire net_16553;
wire net_10636;
wire net_20697;
wire net_3850;
wire net_9023;
wire net_9153;
wire net_349;
wire net_8222;
wire net_12923;
wire net_1409;
wire net_8547;
wire net_14367;
wire net_12576;
wire net_22826;
wire net_2977;
wire net_13140;
wire net_1428;
wire net_13679;
wire net_14629;
wire net_14518;
wire net_15297;
wire net_22303;
wire net_13137;
wire net_5222;
wire net_10510;
wire net_14340;
wire net_4238;
wire net_5844;
wire net_2350;
wire net_6293;
wire net_10506;
wire net_5740;
wire net_14763;
wire net_21621;
wire net_16697;
wire net_20747;
wire net_8950;
wire net_12366;
wire net_18226;
wire net_3143;
wire net_3226;
wire net_9819;
wire net_2757;
wire net_9531;
wire net_12776;
wire net_3629;
wire net_21058;
wire net_7315;
wire net_19502;
wire net_2038;
wire net_2369;
wire net_17731;
wire net_17491;
wire net_12878;
wire net_22099;
wire net_1676;
wire net_20194;
wire net_698;
wire net_14230;
wire net_12969;
wire net_14374;
wire net_5259;
wire net_17618;
wire net_8515;
wire net_4649;
wire net_2485;
wire net_6967;
wire net_13906;
wire net_19537;
wire net_3857;
wire net_21932;
wire net_18840;
wire net_749;
wire net_19456;
wire net_11729;
wire net_15053;
wire net_1948;
wire net_11500;
wire net_11898;
wire net_1006;
wire net_15922;
wire net_21683;
wire net_2781;
wire net_22774;
wire net_19801;
wire net_6767;
wire net_18264;
wire net_9724;
wire net_14695;
wire net_17694;
wire net_7839;
wire net_20408;
wire net_20204;
wire net_15950;
wire net_18536;
wire net_15253;
wire net_19548;
wire net_20463;
wire net_19052;
wire net_7544;
wire net_18392;
wire net_17395;
wire net_21517;
wire net_15955;
wire net_19176;
wire net_3056;
wire net_14050;
wire net_8710;
wire net_3614;
wire net_7624;
wire net_13007;
wire net_17399;
wire net_6792;
wire net_19494;
wire net_15600;
wire net_20964;
wire net_14991;
wire net_4496;
wire net_9525;
wire net_18748;
wire net_6067;
wire net_2127;
wire net_3407;
wire x3521;
wire net_8720;
wire net_13569;
wire net_17431;
wire net_737;
wire net_3656;
wire net_2284;
wire net_5865;
wire net_20005;
wire net_13372;
wire x5409;
wire net_17921;
wire net_15623;
wire net_5957;
wire net_20885;
wire net_20668;
wire net_11541;
wire net_11722;
wire net_5201;
wire net_12375;
wire net_1156;
wire net_15127;
wire net_14127;
wire net_16963;
wire net_1966;
wire net_13641;
wire net_13049;
wire net_14299;
wire net_12188;
wire net_4571;
wire net_11718;
wire net_16081;
wire net_12873;
wire net_5977;
wire net_16520;
wire net_19447;
wire net_326;
wire net_19743;
wire net_2381;
wire net_20453;
wire net_10286;
wire net_11012;
wire net_17142;
wire net_19668;
wire net_15393;
wire net_9504;
wire net_5403;
wire net_15932;
wire net_20984;
wire net_10242;
wire net_6668;
wire net_6735;
wire net_3175;
wire net_10076;
wire net_14918;
wire net_17865;
wire net_2829;
wire net_19244;
wire net_10288;
wire net_3142;
wire net_4099;
wire net_4815;
wire net_21092;
wire net_1219;
wire net_12826;
wire net_14410;
wire net_10886;
wire net_10871;
wire net_13815;
wire net_3884;
wire net_2877;
wire net_3736;
wire net_8745;
wire net_21021;
wire net_22793;
wire net_9352;
wire net_8334;
wire net_1632;
wire net_3796;
wire net_1661;
wire net_1236;
wire net_22150;
wire net_13627;
wire net_22637;
wire net_8987;
wire net_13771;
wire net_19022;
wire net_2700;
wire net_18444;
wire net_17778;
wire net_7996;
wire net_21189;
wire net_7868;
wire net_10307;
wire net_19413;
wire net_16514;
wire net_9548;
wire net_17701;
wire net_1488;
wire net_6273;
wire net_6841;
wire net_2812;
wire net_15406;
wire net_352;
wire net_5691;
wire net_12721;
wire net_18140;
wire net_9320;
wire net_21282;
wire net_3920;
wire net_19230;
wire net_6342;
wire net_7373;
wire net_15810;
wire net_7903;
wire net_1641;
wire net_7511;
wire net_16645;
wire net_19996;
wire net_19299;
wire net_22177;
wire net_4919;
wire net_22221;
wire net_20214;
wire net_1103;
wire net_18608;
wire net_17002;
wire net_767;
wire net_22800;
wire net_16742;
wire net_4557;
wire net_19470;
wire net_131;
wire net_9754;
wire net_21014;
wire net_5488;
wire net_8693;
wire net_2016;
wire net_4292;
wire net_7564;
wire net_14169;
wire net_17036;
wire net_7702;
wire net_10486;
wire net_16369;
wire net_3125;
wire net_13952;
wire net_21538;
wire net_10962;
wire net_12544;
wire net_6550;
wire net_18434;
wire net_22673;
wire net_9101;
wire net_13021;
wire net_9022;
wire net_19023;
wire net_10043;
wire net_15873;
wire net_16755;
wire net_21641;
wire net_13321;
wire net_21617;
wire net_7526;
wire net_14815;
wire net_468;
wire net_9308;
wire net_18916;
wire net_16433;
wire net_19081;
wire net_9257;
wire net_9372;
wire net_16596;
wire net_9738;
wire net_11654;
wire net_19975;
wire net_22194;
wire net_18077;
wire net_15573;
wire net_20054;
wire net_22653;
wire net_179;
wire net_16877;
wire net_9665;
wire net_22312;
wire net_10171;
wire net_62;
wire net_8677;
wire net_15898;
wire net_14871;
wire net_14722;
wire net_3261;
wire net_17100;
wire net_2289;
wire net_18145;
wire net_7300;
wire net_6759;
wire net_11244;
wire net_5919;
wire net_1868;
wire net_20059;
wire net_13942;
wire net_18345;
wire net_7205;
wire net_10110;
wire net_22357;
wire net_17900;
wire net_12684;
wire net_3863;
wire net_10538;
wire net_9856;
wire net_17280;
wire net_20389;
wire net_5778;
wire net_20107;
wire net_3382;
wire net_4257;
wire net_20809;
wire net_13756;
wire net_20355;
wire net_17944;
wire net_4872;
wire net_990;
wire net_7423;
wire net_11485;
wire net_11728;
wire net_10428;
wire net_21915;
wire net_10473;
wire net_11763;
wire net_19141;
wire net_3774;
wire net_1803;
wire net_13803;
wire net_8031;
wire net_20309;
wire net_1134;
wire net_363;
wire net_17025;
wire net_776;
wire net_4550;
wire net_44;
wire net_2508;
wire net_15358;
wire net_9624;
wire net_12118;
wire net_1650;
wire net_8451;
wire net_10353;
wire net_17018;
wire net_3149;
wire net_10717;
wire net_12696;
wire net_13574;
wire net_15174;
wire net_1675;
wire net_6454;
wire net_11253;
wire net_19019;
wire net_2247;
wire net_19657;
wire net_8115;
wire net_2291;
wire net_6525;
wire net_10531;
wire net_11108;
wire net_15220;
wire net_22395;
wire net_16045;
wire net_11096;
wire net_15558;
wire net_8414;
wire net_18802;
wire net_1201;
wire net_2525;
wire net_12404;
wire net_21104;
wire net_12073;
wire net_9701;
wire net_20013;
wire net_14331;
wire net_5106;
wire net_8074;
wire net_13852;
wire net_859;
wire net_1167;
wire net_7259;
wire net_8636;
wire net_19580;
wire net_1044;
wire net_20615;
wire net_18561;
wire net_4322;
wire net_10948;
wire net_10617;
wire net_22809;
wire net_2043;
wire net_19707;
wire net_18609;
wire net_6775;
wire net_10662;
wire net_15818;
wire net_3605;
wire net_14336;
wire net_6635;
wire net_10865;
wire net_12174;
wire net_22059;
wire net_4114;
wire net_7250;
wire net_11055;
wire net_17425;
wire net_14220;
wire net_22612;
wire net_865;
wire net_10330;
wire net_13500;
wire net_19753;
wire net_9896;
wire net_2621;
wire net_13326;
wire net_13832;
wire net_1223;
wire net_21530;
wire net_2750;
wire net_5816;
wire net_21599;
wire net_926;
wire net_11961;
wire net_19637;
wire net_4623;
wire net_7264;
wire net_7403;
wire net_17654;
wire net_6153;
wire net_14656;
wire net_8642;
wire net_7188;
wire net_10595;
wire net_12868;
wire net_9185;
wire net_6466;
wire net_2048;
wire net_18471;
wire net_4481;
wire net_3633;
wire net_7337;
wire net_21646;
wire net_7036;
wire net_14705;
wire net_3561;
wire net_1295;
wire net_1543;
wire net_10993;
wire net_13692;
wire net_9429;
wire net_5661;
wire net_2071;
wire net_1923;
wire net_1275;
wire net_13481;
wire net_11031;
wire net_13463;
wire net_940;
wire net_4411;
wire net_3719;
wire net_4857;
wire net_10572;
wire net_15681;
wire net_6061;
wire net_21062;
wire net_8311;
wire net_5350;
wire net_12330;
wire net_14329;
wire net_9627;
wire net_13631;
wire net_5335;
wire net_12849;
wire net_19569;
wire net_18578;
wire net_19035;
wire net_10133;
wire net_12438;
wire net_22492;
wire net_9485;
wire net_21858;
wire net_19906;
wire net_16786;
wire net_22747;
wire net_17503;
wire net_21811;
wire net_1454;
wire net_6949;
wire net_17793;
wire net_3342;
wire net_14711;
wire net_1550;
wire net_22485;
wire net_19084;
wire net_9642;
wire net_10069;
wire net_233;
wire net_18596;
wire net_5138;
wire net_18629;
wire net_3459;
wire net_16154;
wire net_13411;
wire net_1268;
wire net_11127;
wire net_3780;
wire net_13783;
wire net_1115;
wire net_4051;
wire net_11465;
wire net_22465;
wire net_17820;
wire net_6641;
wire net_961;
wire net_18886;
wire net_9643;
wire net_2106;
wire net_19602;
wire net_14691;
wire net_5175;
wire net_11909;
wire net_14196;
wire net_4894;
wire net_9424;
wire net_3327;
wire net_9480;
wire net_5091;
wire net_18189;
wire net_13719;
wire net_3456;
wire net_13700;
wire net_7627;
wire net_12250;
wire net_12453;
wire net_13220;
wire x7558;
wire net_9907;
wire net_4407;
wire net_13713;
wire net_16485;
wire net_1586;
wire net_14113;
wire net_5354;
wire x2160;
wire net_216;
wire net_13284;
wire net_22763;
wire net_10727;
wire net_18667;
wire net_2881;
wire net_22662;
wire net_12630;
wire net_4602;
wire net_15556;
wire net_12057;
wire net_5635;
wire net_9495;
wire net_16198;
wire net_8379;
wire net_8806;
wire net_11237;
wire net_21468;
wire net_9097;
wire net_12520;
wire net_1120;
wire net_5881;
wire net_2848;
wire net_20777;
wire net_7126;
wire net_973;
wire net_11832;
wire net_21135;
wire net_1139;
wire net_6998;
wire net_7394;
wire net_9337;
wire net_3902;
wire net_18291;
wire net_19174;
wire net_19105;
wire net_1574;
wire net_9008;
wire net_4842;
wire net_11576;
wire net_20044;
wire net_154;
wire net_8016;
wire net_3699;
wire net_19930;
wire net_16796;
wire net_13847;
wire net_22552;
wire net_12056;
wire net_14946;
wire net_1478;
wire net_14075;
wire net_587;
wire net_1696;
wire net_2179;
wire net_21050;
wire net_1262;
wire net_9163;
wire net_17892;
wire net_4027;
wire net_14106;
wire net_8750;
wire net_4213;
wire net_4505;
wire net_22090;
wire net_18170;
wire net_17517;
wire net_4131;
wire net_7396;
wire net_10779;
wire net_14937;
wire net_1907;
wire net_11323;
wire net_18898;
wire net_16201;
wire net_19786;
wire net_15420;
wire net_20717;
wire net_16982;
wire net_4164;
wire net_6312;
wire net_195;
wire net_21965;
wire net_20409;
wire net_10200;
wire net_18663;
wire net_10247;
wire net_21937;
wire net_16110;
wire net_19501;
wire net_10104;
wire net_17093;
wire net_22521;
wire net_8980;
wire net_19327;
wire net_13999;
wire net_18891;
wire net_22784;
wire net_8323;
wire net_9042;
wire net_7002;
wire net_3761;
wire net_9196;
wire net_13722;
wire net_21477;
wire net_242;
wire net_22052;
wire net_7076;
wire net_7719;
wire net_7722;
wire net_18724;
wire net_21415;
wire net_22073;
wire net_21675;
wire net_9543;
wire net_20220;
wire net_8938;
wire net_19195;
wire net_11384;
wire net_8336;
wire net_13514;
wire net_1311;
wire net_5939;
wire net_11230;
wire net_13307;
wire net_7068;
wire net_10207;
wire net_21968;
wire net_18732;
wire net_10549;
wire net_11911;
wire net_17278;
wire net_5937;
wire net_8208;
wire net_12314;
wire net_3558;
wire net_9678;
wire net_555;
wire net_16327;
wire net_1613;
wire net_7758;
wire net_13016;
wire net_15051;
wire net_790;
wire net_11938;
wire net_20655;
wire net_19132;
wire net_14665;
wire net_21997;
wire net_19059;
wire net_1417;
wire net_11466;
wire net_18501;
wire net_11520;
wire net_13423;
wire net_2386;
wire net_11063;
wire net_20339;
wire net_2166;
wire net_8359;
wire net_11588;
wire net_17918;
wire net_12830;
wire net_15846;
wire net_10650;
wire net_7150;
wire net_13699;
wire net_6537;
wire net_14873;
wire net_19882;
wire net_17497;
wire net_4416;
wire net_714;
wire net_5015;
wire net_1309;
wire net_2999;
wire net_9567;
wire net_683;
wire net_19146;
wire net_1771;
wire net_148;
wire net_4493;
wire net_12136;
wire net_13555;
wire x5723;
wire net_7220;
wire net_17544;
wire net_9171;
wire net_17950;
wire net_15852;
wire net_7449;
wire net_7751;
wire net_10362;
wire net_15799;
wire x5537;
wire net_21725;
wire net_14504;
wire net_5547;
wire net_9361;
wire net_15411;
wire net_9149;
wire net_5616;
wire net_7353;
wire x3153;
wire net_12117;
wire net_7113;
wire net_8588;
wire net_21897;
wire net_2403;
wire net_7740;
wire net_15173;
wire net_17957;
wire net_15582;
wire x3014;
wire net_20415;
wire net_21454;
wire net_14147;
wire net_7913;
wire net_15238;
wire net_18828;
wire net_16220;
wire net_8550;
wire net_14761;
wire net_16819;
wire net_394;
wire net_92;
wire net_810;
wire net_1548;
wire net_15861;
wire net_17159;
wire net_1189;
wire net_3778;
wire net_409;
wire net_20824;
wire net_7183;
wire net_15366;
wire net_21556;
wire net_3470;
wire net_21409;
wire net_11908;
wire net_16297;
wire net_88;
wire net_13354;
wire net_21743;
wire net_8036;
wire net_16790;
wire net_18393;
wire net_11509;
wire net_15113;
wire net_3419;
wire net_10754;
wire net_16021;
wire net_17807;
wire net_1254;
wire net_10733;
wire net_11417;
wire net_18708;
wire net_15616;
wire net_12793;
wire net_13171;
wire net_10533;
wire net_7240;
wire net_11862;
wire net_7365;
wire net_20071;
wire net_5361;
wire x912;
wire net_15496;
wire net_8703;
wire net_9383;
wire net_9841;
wire net_4675;
wire net_8378;
wire net_327;
wire net_3877;
wire net_21946;
wire net_21377;
wire net_16139;
wire net_16583;
wire net_353;
wire net_20878;
wire net_8052;
wire net_13799;
wire net_19322;
wire net_11730;
wire net_12322;
wire net_9584;
wire net_20138;
wire net_8552;
wire net_16620;
wire net_5730;
wire net_20551;
wire net_14209;
wire net_8770;
wire net_14140;
wire net_6927;
wire net_12628;
wire net_3046;
wire net_22599;
wire net_164;
wire net_6019;
wire net_4702;
wire net_22069;
wire net_7632;
wire net_19062;
wire net_15396;
wire net_17583;
wire net_3096;
wire net_1629;
wire net_8947;
wire net_14950;
wire net_19385;
wire net_11387;
wire net_14431;
wire net_805;
wire net_3277;
wire net_12032;
wire net_20117;
wire net_6740;
wire net_12093;
wire net_3590;
wire net_2151;
wire net_17198;
wire net_8521;
wire net_2688;
wire net_20329;
wire net_14304;
wire net_1622;
wire net_19461;
wire net_20582;
wire net_21202;
wire net_38;
wire net_20595;
wire net_22594;
wire net_13392;
wire net_5149;
wire net_6299;
wire net_11664;
wire net_16003;
wire net_17635;
wire net_7815;
wire net_7453;
wire net_14793;
wire net_20086;
wire net_12998;
wire net_22252;
wire net_11744;
wire net_13420;
wire net_20701;
wire net_18685;
wire net_2244;
wire net_12825;
wire net_15809;
wire net_11737;
wire x6797;
wire net_7826;
wire net_19944;
wire net_783;
wire net_11955;
wire x1526;
wire net_20410;
wire net_13686;
wire net_9211;
wire net_6305;
wire net_11703;
wire net_22000;
wire net_17549;
wire net_2605;
wire net_9469;
wire net_550;
wire net_9875;
wire net_10821;
wire net_5238;
wire net_12292;
wire net_17759;
wire net_9158;
wire net_3991;
wire net_5086;
wire x866;
wire net_10912;
wire net_461;
wire net_14516;
wire net_7778;
wire net_20733;
wire net_16517;
wire net_6879;
wire net_12962;
wire net_6657;
wire net_8524;
wire net_20230;
wire net_9284;
wire net_20075;
wire net_14185;
wire net_20247;
wire net_1512;
wire net_17744;
wire net_18636;
wire net_15370;
wire net_14593;
wire net_8047;
wire net_1330;
wire net_5025;
wire net_4275;
wire net_17586;
wire net_3015;
wire net_11011;
wire net_1785;
wire net_4771;
wire net_11077;
wire net_13507;
wire net_16062;
wire net_20921;
wire net_17132;
wire net_10680;
wire net_9516;
wire net_20450;
wire net_6870;
wire net_16752;
wire net_9655;
wire net_20322;
wire x1446;
wire net_5060;
wire net_12596;
wire net_15848;
wire net_5668;
wire net_10408;
wire net_985;
wire net_4679;
wire net_16492;
wire net_6719;
wire net_12190;
wire net_19310;
wire net_7061;
wire net_15494;
wire net_21529;
wire net_16609;
wire net_424;
wire net_6837;
wire net_19775;
wire net_22627;
wire net_1729;
wire net_3353;
wire net_12623;
wire net_16274;
wire net_4247;
wire net_21994;
wire net_17477;
wire net_5719;
wire net_17112;
wire net_21342;
wire net_3639;
wire net_14404;
wire net_15915;
wire net_8065;
wire net_12311;
wire net_12148;
wire net_11992;
wire net_3086;
wire net_21260;
wire x1159;
wire net_4585;
wire net_2058;
wire net_11110;
wire net_22277;
wire net_3045;
wire net_12206;
wire net_21835;
wire net_17669;
wire net_20815;
wire net_4875;
wire net_2018;
wire net_21636;
wire net_13100;
wire net_11731;
wire net_20255;
wire net_2510;
wire net_9952;
wire net_19837;
wire net_3808;
wire net_7881;
wire net_19261;
wire net_12941;
wire net_14631;
wire net_6243;
wire net_7882;
wire x2957;
wire net_6415;
wire x3117;
wire net_14393;
wire net_18316;
wire net_9201;
wire net_19699;
wire net_19554;
wire net_19434;
wire net_17666;
wire net_6302;
wire net_8916;
wire net_2279;
wire net_14048;
wire net_3447;
wire net_15633;
wire net_6174;
wire net_8401;
wire net_14588;
wire net_20289;
wire net_17812;
wire net_18487;
wire net_20122;
wire net_17408;
wire net_19211;
wire net_19073;
wire net_17224;
wire net_9267;
wire net_10826;
wire net_13893;
wire net_102;
wire net_8497;
wire net_22339;
wire net_18284;
wire net_17521;
wire net_10295;
wire net_7801;
wire net_3217;
wire net_21578;
wire net_1291;
wire net_4387;
wire net_6362;
wire net_1865;
wire net_21249;
wire net_19123;
wire net_13896;
wire net_18695;
wire net_5168;
wire net_6076;
wire net_5329;
wire net_21439;
wire net_18312;
wire net_14541;
wire net_22740;
wire net_19293;
wire net_10985;
wire net_17752;
wire net_8460;
wire net_10490;
wire net_2578;
wire net_8658;
wire net_16392;
wire net_1433;
wire net_10462;
wire net_18052;
wire net_17042;
wire net_11672;
wire net_13745;
wire net_15503;
wire net_19289;
wire net_14786;
wire net_8606;
wire net_5440;
wire net_9425;
wire net_2574;
wire net_5928;
wire net_14235;
wire net_3531;
wire net_3747;
wire net_18454;
wire net_5732;
wire net_12212;
wire net_8593;
wire net_18594;
wire net_20248;
wire net_1844;
wire net_389;
wire net_11512;
wire net_902;
wire net_19704;
wire net_13981;
wire net_11287;
wire net_15859;
wire net_15907;
wire net_13237;
wire net_736;
wire net_8771;
wire net_5462;
wire net_5282;
wire net_6498;
wire net_8372;
wire net_18767;
wire net_21861;
wire net_15737;
wire net_22609;
wire net_21447;
wire net_6262;
wire net_17713;
wire net_19511;
wire net_10905;
wire net_15379;
wire net_19005;
wire net_12517;
wire net_18400;
wire x3079;
wire net_14092;
wire net_10034;
wire net_7249;
wire net_18137;
wire net_15152;
wire net_21782;
wire net_20083;
wire net_21275;
wire net_19804;
wire net_5717;
wire net_869;
wire net_3714;
wire net_12144;
wire net_20558;
wire net_8308;
wire net_11280;
wire net_4077;
wire net_2441;
wire net_21163;
wire net_18825;
wire net_20492;
wire net_4749;
wire net_5828;
wire net_6799;
wire net_20421;
wire net_20624;
wire net_21072;
wire net_8775;
wire net_12092;
wire net_13774;
wire net_19641;
wire net_2459;
wire net_15512;
wire net_10394;
wire net_19981;
wire net_14434;
wire net_5422;
wire net_6629;
wire net_6704;
wire net_12395;
wire net_15329;
wire net_19002;
wire net_16415;
wire net_19646;
wire net_6508;
wire net_15832;
wire net_18968;
wire net_2075;
wire net_2548;
wire net_20338;
wire net_3359;
wire net_5848;
wire net_15883;
wire net_10085;
wire net_12296;
wire net_20187;
wire net_9069;
wire net_15900;
wire net_7548;
wire net_12889;
wire net_14866;
wire net_6165;
wire net_4795;
wire net_511;
wire net_9263;
wire net_19452;
wire net_12759;
wire net_3967;
wire net_20899;
wire net_19489;
wire net_2654;
wire net_1819;
wire net_2911;
wire net_11791;
wire net_8258;
wire net_15509;
wire net_21794;
wire net_12821;
wire net_19764;
wire net_12763;
wire net_19742;
wire net_17404;
wire net_19096;
wire net_7236;
wire net_17271;
wire net_11379;
wire net_13181;
wire net_9031;
wire net_18508;
wire net_13661;
wire net_11083;
wire net_989;
wire net_8446;
wire net_17629;
wire net_458;
wire net_18512;
wire net_20294;
wire net_11748;
wire net_7442;
wire net_8322;
wire net_14471;
wire net_9030;
wire net_10998;
wire net_16686;
wire net_10957;
wire net_21049;
wire net_14183;
wire net_13333;
wire net_4616;
wire net_11408;
wire net_13096;
wire net_16186;
wire net_4786;
wire net_19162;
wire net_16212;
wire net_8616;
wire net_21305;
wire net_18779;
wire net_5893;
wire net_7872;
wire net_10542;
wire net_17287;
wire net_10891;
wire net_2111;
wire net_3410;
wire net_14954;
wire net_5525;
wire net_8162;
wire net_12496;
wire net_16867;
wire net_21128;
wire net_21044;
wire net_21367;
wire net_5610;
wire net_14894;
wire net_16627;
wire net_14278;
wire net_20874;
wire net_13045;
wire net_2535;
wire net_3191;
wire net_13165;
wire net_19239;
wire net_13822;
wire net_14396;
wire net_15106;
wire net_10355;
wire net_12865;
wire net_19727;
wire net_18093;
wire net_12125;
wire net_20949;
wire net_20647;
wire net_2983;
wire net_21160;
wire net_12916;
wire net_14617;
wire net_22335;
wire net_10024;
wire net_1647;
wire net_198;
wire net_12460;
wire net_10058;
wire net_7509;
wire net_4756;
wire net_20252;
wire net_5196;
wire net_13280;
wire net_15293;
wire net_19346;
wire net_16255;
wire net_18476;
wire net_2892;
wire net_13263;
wire net_15646;
wire net_18711;
wire net_13077;
wire net_4444;
wire net_848;
wire net_22587;
wire net_9550;
wire net_20069;
wire net_1080;
wire net_12022;
wire net_10641;
wire net_16705;
wire net_1890;
wire net_21522;
wire net_13648;
wire net_21122;
wire net_18755;
wire net_11293;
wire net_22205;
wire net_2357;
wire net_4501;
wire net_12449;
wire net_13319;
wire net_11114;
wire net_19720;
wire net_18736;
wire net_19356;
wire net_20180;
wire net_5492;
wire net_11772;
wire net_17875;
wire net_12383;
wire net_11372;
wire net_10199;
wire net_20737;
wire net_6536;
wire net_15728;
wire net_4363;
wire net_7417;
wire net_16016;
wire net_606;
wire net_623;
wire net_3906;
wire net_663;
wire net_12503;
wire net_1891;
wire net_5180;
wire net_579;
wire net_3998;
wire net_16443;
wire net_9490;
wire net_8597;
wire net_21881;
wire net_2062;
wire net_18074;
wire net_13666;
wire net_9828;
wire net_22600;
wire net_18380;
wire x1134;
wire net_22690;
wire net_6418;
wire net_10844;
wire net_19678;
wire net_17678;
wire net_20524;
wire net_4834;
wire net_7296;
wire net_17673;
wire net_8061;
wire net_9317;
wire net_4067;
wire net_20511;
wire net_4717;
wire net_20661;
wire net_1518;
wire net_17682;
wire net_4618;
wire net_1437;
wire net_1194;
wire net_18273;
wire net_15837;
wire net_22758;
wire net_5517;
wire net_17576;
wire net_21580;
wire net_17150;
wire net_6770;
wire net_7587;
wire net_11923;
wire net_20530;
wire net_1664;
wire net_17345;
wire net_13651;
wire net_15718;
wire net_16227;
wire net_705;
wire net_10326;
wire x585;
wire x2666;
wire net_2948;
wire net_10523;
wire net_19184;
wire net_17055;
wire net_1036;
wire net_18186;
wire net_5608;
wire net_6052;
wire net_7497;
wire net_11966;
wire net_4537;
wire net_1196;
wire net_3973;
wire net_6331;
wire net_21712;
wire net_22210;
wire net_6762;
wire net_9077;
wire net_5531;
wire net_20919;
wire net_6085;
wire net_6598;
wire net_20120;
wire net_5701;
wire net_11786;
wire net_3136;
wire net_21954;
wire net_4090;
wire net_12553;
wire net_21443;
wire net_6149;
wire net_20859;
wire net_19541;
wire net_9178;
wire net_10809;
wire net_3834;
wire net_10300;
wire net_13471;
wire net_3152;
wire net_20149;
wire net_14311;
wire net_3648;
wire net_1722;
wire net_16854;
wire net_2008;
wire net_6395;
wire net_18133;
wire net_11633;
wire net_2808;
wire net_18481;
wire x1987;
wire net_8265;
wire net_9055;
wire net_19349;
wire net_14008;
wire net_17761;
wire net_6575;
wire net_16907;
wire net_16654;
wire net_4707;
wire net_6432;
wire net_13918;
wire net_16119;
wire net_20676;
wire net_17932;
wire net_957;
wire net_12771;
wire net_15667;
wire net_18839;
wire net_1287;
wire net_10625;
wire net_14040;
wire net_2726;
wire net_19788;
wire net_77;
wire net_20285;
wire net_1340;
wire net_49;
wire net_20090;
wire net_7277;
wire net_21665;
wire net_7165;
wire net_9599;
wire net_12363;
wire net_22502;
wire net_2844;
wire net_12415;
wire net_9977;
wire net_5538;
wire net_19916;
wire net_4852;
wire net_6804;
wire net_9941;
wire net_10341;
wire net_14361;
wire net_4437;
wire net_10435;
wire net_51;
wire net_18281;
wire net_4028;
wire net_2860;
wire net_432;
wire net_4927;
wire net_6025;
wire net_6329;
wire net_10627;
wire net_1142;
wire net_14556;
wire net_3159;
wire net_5644;
wire net_67;
wire net_16380;
wire net_2240;
wire net_14600;
wire net_18859;
wire net_2416;
wire net_12882;
wire net_6404;
wire net_20518;
wire net_8727;
wire net_21758;
wire net_14354;
wire net_6185;
wire net_9713;
wire net_5383;
wire net_17833;
wire net_10540;
wire net_7487;
wire net_13520;
wire net_21218;
wire net_20354;
wire net_4013;
wire net_11517;
wire net_2144;
wire net_2236;
wire net_11057;
wire net_3443;
wire net_22240;
wire net_3945;
wire net_8824;
wire net_19399;
wire net_11529;
wire net_14622;
wire net_22188;
wire net_20581;
wire net_1505;
wire net_19530;
wire net_16476;
wire net_8279;
wire net_13836;
wire net_3669;
wire net_3952;
wire net_19836;
wire net_1861;
wire net_13448;
wire net_19440;
wire net_9999;
wire net_4388;
wire net_11852;
wire net_1594;
wire net_221;
wire net_5672;
wire net_20560;
wire net_18252;
wire x2382;
wire net_542;
wire net_14218;
wire net_17872;
wire net_13026;
wire net_12483;
wire net_20545;
wire x6631;
wire net_6487;
wire net_18818;
wire net_22254;
wire x3279;
wire net_4562;
wire net_9437;
wire net_2376;
wire net_1520;
wire net_6562;
wire net_6713;
wire net_18529;
wire net_15867;
wire net_16767;
wire net_8579;
wire net_9638;
wire net_22431;
wire net_16619;
wire net_15287;
wire net_19631;
wire net_8005;
wire net_3664;
wire net_3233;
wire net_5124;
wire net_14521;
wire net_9731;
wire net_19690;
wire net_16642;
wire net_7178;
wire net_10937;
wire net_17212;
wire net_11814;
wire net_9649;
wire net_1584;
wire net_16693;
wire net_13539;
wire net_22607;
wire net_20796;
wire net_20852;
wire net_12612;
wire net_2330;
wire net_7890;
wire net_3397;
wire net_16348;
wire net_9777;
wire net_5898;
wire net_18976;
wire net_6785;
wire net_15948;
wire net_4391;
wire net_7814;
wire net_11473;
wire net_22166;
wire net_9045;
wire net_12659;
wire net_6875;
wire net_20434;
wire net_2857;
wire net_8674;
wire net_2767;
wire net_9594;
wire net_6120;
wire net_16837;
wire net_11491;
wire net_6604;
wire net_12652;
wire net_22509;
wire net_825;
wire net_309;
wire x3989;
wire net_19902;
wire net_18522;
wire net_21175;
wire net_1366;
wire net_20960;
wire net_17185;
wire net_13054;
wire net_2615;
wire net_14978;
wire net_31;
wire net_14268;
wire net_9290;
wire net_16313;
wire net_7367;
wire net_8158;
wire net_1151;
wire net_16120;
wire net_21319;
wire net_5240;
wire net_5318;
wire net_9993;
wire net_11138;
wire net_17149;
wire net_8291;
wire net_15046;
wire net_21565;
wire net_2818;
wire net_3213;
wire net_7690;
wire net_580;
wire net_4173;
wire net_2136;
wire net_9805;
wire net_21957;
wire net_2339;
wire net_22548;
wire net_19409;
wire x4545;
wire net_7699;
wire net_8884;
wire net_4157;
wire net_19376;
wire net_1879;
wire net_14821;
wire net_20752;
wire net_6663;
wire net_12122;
wire net_19650;
wire net_13224;
wire net_8202;
wire net_22015;
wire net_19428;
wire net_19606;
wire net_21776;
wire net_4221;
wire net_4941;
wire net_17447;
wire net_6732;
wire net_12524;
wire net_12683;
wire net_19795;
wire net_22342;
wire net_17047;
wire net_5604;
wire net_11022;
wire net_11612;
wire net_8351;
wire net_21981;
wire net_21252;
wire net_19255;
wire net_18922;
wire net_4887;
wire net_15760;
wire net_18012;
wire net_13116;
wire net_21720;
wire net_763;
wire net_20375;
wire net_13704;
wire net_21709;
wire net_16285;
wire net_14088;
wire net_7762;
wire net_1740;
wire net_5639;
wire net_14495;
wire net_17217;
wire net_9455;
wire net_872;
wire net_22684;
wire net_20979;
wire net_9125;
wire net_22434;
wire net_10502;
wire net_21827;
wire net_8251;
wire net_3880;
wire net_5581;
wire net_21610;
wire net_20325;
wire net_18110;
wire net_16405;
wire net_4333;
wire net_21567;
wire net_11285;
wire net_14776;
wire net_18989;
wire net_5558;
wire net_7575;
wire net_22122;
wire net_21793;
wire net_22489;
wire net_4880;
wire net_1812;
wire net_8174;
wire net_12584;
wire net_4825;
wire net_10850;
wire net_18604;
wire net_8696;
wire net_4138;
wire net_3203;
wire net_21234;
wire net_12811;
wire net_11881;
wire net_21312;
wire net_2589;
wire net_2659;
wire net_7515;
wire net_12670;
wire net_591;
wire net_1700;
wire net_12739;
wire net_12985;
wire net_16766;
wire net_7557;
wire net_10188;
wire net_20302;
wire net_178;
wire net_18813;
wire net_18794;
wire net_11751;
wire net_20210;
wire net_15266;
wire net_9074;
wire net_2843;
wire net_22119;
wire net_6780;
wire net_14081;
wire net_22443;
wire net_7961;
wire net_10191;
wire net_15322;
wire net_3807;
wire net_10480;
wire net_21507;
wire net_809;
wire net_13995;
wire net_8393;
wire net_635;
wire net_1235;
wire net_266;
wire net_4279;
wire net_2691;
wire net_18041;
wire net_21328;
wire net_8610;
wire net_12600;
wire net_6622;
wire net_6007;
wire net_15520;
wire net_13205;
wire net_20953;
wire net_10176;
wire net_6549;
wire net_6542;
wire net_3460;
wire net_13091;
wire net_20038;
wire net_12859;
wire net_18811;
wire net_3198;
wire net_1626;
wire net_5720;
wire net_8366;
wire net_2822;
wire net_7317;
wire net_21206;
wire net_1258;
wire net_8413;
wire net_17857;
wire net_12041;
wire net_9866;
wire net_21903;
wire net_318;
wire net_10231;
wire net_19879;
wire net_3927;
wire net_10859;
wire net_1971;
wire net_8931;
wire net_2409;
wire net_1900;
wire net_3192;
wire net_1779;
wire net_21002;
wire net_2647;
wire net_21423;
wire net_5218;
wire net_21388;
wire net_8492;
wire net_22223;
wire net_7972;
wire net_228;
wire net_11886;
wire net_4737;
wire net_2640;
wire net_966;
wire net_13011;
wire net_21747;
wire net_7083;
wire net_3372;
wire net_4698;
wire net_2201;
wire net_6049;
wire net_2025;
wire net_2827;
wire net_16748;
wire net_20569;
wire net_2936;
wire net_7905;
wire net_5643;
wire net_9936;
wire net_20833;
wire net_19490;
wire net_5728;
wire net_13736;
wire net_16760;
wire net_17507;
wire net_8013;
wire net_17146;
wire net_20693;
wire net_10702;
wire net_12425;
wire net_10366;
wire net_20999;
wire net_16924;
wire net_14297;
wire net_21352;
wire net_11414;
wire net_10920;
wire net_11265;
wire net_12444;
wire net_15024;
wire net_22403;
wire net_22707;
wire net_12529;
wire net_10579;
wire net_16536;
wire net_7997;
wire net_4522;
wire net_11925;
wire net_8908;
wire net_14836;
wire net_3652;
wire net_8689;
wire net_2669;
wire net_6829;
wire net_22183;
wire net_22582;
wire net_18929;
wire net_4083;
wire net_1173;
wire net_1754;
wire net_2328;
wire net_7715;
wire net_11401;
wire net_16561;
wire x5244;
wire net_8080;
wire net_5571;
wire net_22129;
wire net_15302;
wire net_5805;
wire net_10205;
wire x5825;
wire net_12792;
wire net_7254;
wire net_22154;
wire net_13623;
wire net_7684;
wire net_17607;
wire net_16164;
wire net_12991;
wire net_10743;
wire net_9604;
wire net_13565;
wire net_13605;
wire net_14467;
wire net_6887;
wire net_18263;
wire net_9838;
wire net_15427;
wire net_4462;
wire net_15546;
wire net_11038;
wire net_1394;
wire net_2963;
wire net_5412;
wire net_5546;
wire net_6134;
wire net_1281;
wire net_9395;
wire net_2463;
wire net_9291;
wire net_8210;
wire net_15945;
wire net_16996;
wire net_21359;
wire net_8995;
wire net_11258;
wire net_8367;
wire net_4058;
wire net_8432;
wire net_16469;
wire net_21293;
wire net_3509;
wire net_1162;
wire net_13856;
wire net_17536;
wire net_2472;
wire net_2742;
wire net_2790;
wire net_13589;
wire net_13120;
wire net_22145;
wire net_5007;
wire net_10738;
wire net_10318;
wire net_15386;
wire net_22730;
wire net_10434;
wire net_13795;
wire net_20868;
wire net_22621;
wire net_8360;
wire net_11902;
wire net_6521;
wire net_10269;
wire net_17480;
wire net_22307;
wire net_3320;
wire net_10561;
wire net_17599;
wire net_16108;
wire net_5221;
wire net_3657;
wire net_5550;
wire net_1353;
wire net_14683;
wire net_21664;
wire net_11652;
wire net_15165;
wire net_5303;
wire net_3581;
wire net_20480;
wire net_18932;
wire net_14961;
wire net_4049;
wire net_19619;
wire net_1300;
wire net_18876;
wire net_18644;
wire net_14322;
wire net_12131;
wire net_22733;
wire net_16723;
wire net_14419;
wire net_21748;
wire net_16102;
wire net_17312;
wire net_13432;
wire net_547;
wire net_10941;
wire net_14026;
wire net_1098;
wire net_19523;
wire net_10049;
wire net_6683;
wire net_238;
wire net_20914;
wire net_3074;
wire x923;
wire net_5475;
wire net_8973;
wire net_7055;
wire net_11354;
wire net_2438;
wire net_7896;
wire net_1911;
wire net_19939;
wire net_6906;
wire net_17512;
wire net_22728;
wire net_649;
wire net_19138;
wire net_13597;
wire net_21582;
wire net_1374;
wire net_13887;
wire net_4843;
wire net_8959;
wire net_22087;
wire net_16887;
wire net_20447;
wire net_2494;
wire net_18671;
wire net_15747;
wire net_11217;
wire net_16989;
wire net_6819;
wire net_12274;
wire net_14811;
wire net_3700;
wire net_13349;
wire net_107;
wire net_530;
wire net_9140;
wire net_15155;
wire net_10529;
wire net_11839;
wire net_21338;
wire net_10004;
wire net_22739;
wire net_22423;
wire net_673;
wire net_4268;
wire net_7022;
wire net_7029;
wire net_12247;
wire net_2797;
wire net_6256;
wire net_9966;
wire net_3846;
wire net_12261;
wire net_3549;
wire net_9790;
wire net_1445;
wire net_8581;
wire net_10227;
wire net_6729;
wire net_13807;
wire net_19110;
wire net_16206;
wire net_9922;
wire net_22474;
wire net_7639;
wire net_10126;
wire net_11454;
wire net_11583;
wire net_5379;
wire net_13340;
wire net_3913;
wire net_9988;
wire net_11643;
wire net_3787;
wire net_17487;
wire net_1810;
wire net_1118;
wire net_10776;
wire net_21402;
wire net_21393;
wire net_372;
wire net_6858;
wire net_12235;
wire net_9882;
wire net_18678;
wire net_7086;
wire net_2990;
wire net_22386;
wire net_6324;
wire net_16145;
wire net_11749;
wire net_18741;
wire net_3595;
wire net_2788;
wire net_8923;
wire net_10383;
wire net_13787;
wire net_6899;
wire net_10142;
wire net_14490;
wire net_15774;
wire net_20275;
wire net_19925;
wire net_3489;
wire net_15346;
wire net_11184;
wire net_19047;
wire net_13581;
wire net_563;
wire net_7854;
wire net_1147;
wire net_13979;
wire net_18194;
wire net_13388;
wire net_15242;
wire net_15193;
wire x2027;
wire net_8815;
wire net_13452;
wire net_21456;
wire net_2158;
wire net_22830;
wire net_4366;
wire net_10234;
wire net_10175;
wire net_13936;
wire net_17997;
wire net_5009;
wire net_12254;
wire net_3684;
wire net_14677;
wire net_8418;
wire net_2428;
wire net_10695;
wire net_8652;
wire net_10814;
wire net_2895;
wire net_13299;
wire net_15488;
wire net_15985;
wire net_20600;
wire net_8238;
wire net_13418;
wire net_20110;
wire net_2477;
wire net_12957;
wire net_19421;
wire net_9927;
wire net_16238;
wire net_5653;
wire net_13819;
wire net_16770;
wire net_7664;
wire net_4188;
wire net_15451;
wire net_19889;
wire net_4040;
wire net_6146;
wire net_5433;
wire net_12766;
wire net_3759;
wire net_3511;
wire net_374;
wire net_12839;
wire net_14069;
wire net_8755;
wire net_17076;
wire x1103;
wire net_1987;
wire net_12816;
wire net_16242;
wire net_12910;
wire net_7011;
wire net_249;
wire net_3602;
wire net_16827;
wire net_13155;
wire net_22814;
wire net_19966;
wire net_17258;
wire net_9963;
wire net_17122;
wire net_5283;
wire net_21846;
wire net_18215;
wire net_9013;
wire net_8871;
wire net_15895;
wire net_6196;
wire net_4009;
wire net_10766;
wire net_13488;
wire net_17937;
wire net_7648;
wire net_8508;
wire net_13880;
wire x7584;
wire net_5993;
wire net_2632;
wire net_16028;
wire net_2547;
wire net_5076;
wire net_8634;
wire net_16487;
wire net_21731;
wire net_17167;
wire net_9084;
wire net_22719;
wire net_15440;
wire net_2295;
wire net_5831;
wire net_5628;
wire net_1817;
wire net_17962;
wire net_11009;
wire net_16078;
wire net_9348;
wire net_1381;
wire net_6445;
wire net_202;
wire net_3312;
wire net_13596;
wire net_17590;
wire net_1756;
wire net_7325;
wire net_18491;
wire net_2208;
wire net_6475;
wire net_918;
wire net_19367;
wire net_7727;
wire net_11204;
wire net_5397;
wire net_18573;
wire net_20972;
wire net_9204;
wire net_17374;
wire net_22619;
wire net_5901;
wire net_13610;
wire net_9356;
wire net_1129;
wire net_10780;
wire net_1056;
wire net_11345;
wire net_14689;
wire net_4908;
wire net_19823;
wire net_20506;
wire net_14561;
wire net_10896;
wire net_22553;
wire net_17969;
wire net_4781;
wire net_2044;
wire net_17458;
wire net_2181;
wire net_7402;
wire net_6913;
wire net_8626;
wire net_14782;
wire net_18414;
wire net_8406;
wire net_17508;
wire net_4530;
wire net_7379;
wire net_838;
wire net_21779;
wire net_6123;
wire net_10441;
wire net_18303;
wire net_16899;
wire net_11151;
wire net_14316;
wire net_14202;
wire net_22287;
wire net_11750;
wire net_5872;
wire net_20673;
wire net_20167;
wire net_4980;
wire net_7107;
wire net_20064;
wire net_17846;
wire net_11270;
wire net_15341;
wire net_3827;
wire net_16542;
wire net_8405;
wire x7607;
wire net_12072;
wire net_5308;
wire net_3515;
wire net_5033;
wire net_12747;
wire net_16059;
wire net_8085;
wire net_17171;
wire net_9720;
wire net_18153;
wire net_22323;
wire net_3398;
wire net_9223;
wire net_22334;
wire net_16721;
wire net_342;
wire net_13400;
wire net_612;
wire net_892;
wire net_16930;
wire net_8098;
wire net_4198;
wire net_12871;
wire net_22750;
wire net_21806;
wire net_10423;
wire net_20365;
wire net_5434;
wire net_11144;
wire net_10848;
wire net_14488;
wire net_20765;
wire net_8344;
wire net_12639;
wire net_19430;
wire net_6511;
wire net_10060;
wire net_19819;
wire net_1537;
wire net_11105;
wire net_13051;
wire x2855;
wire x511;
wire net_13399;
wire net_4074;
wire net_16730;
wire net_4000;
wire net_2214;
wire net_14913;
wire net_16073;
wire net_3338;
wire net_17973;
wire net_5987;
wire net_21490;
wire net_15468;
wire net_21975;
wire net_13238;
wire net_417;
wire net_9929;
wire net_21214;
wire net_17370;
wire x1192;
wire net_5387;
wire net_10634;
wire net_8217;
wire net_7467;
wire net_22199;
wire net_10758;
wire net_17191;
wire net_17011;
wire net_3337;
wire net_8287;
wire net_2662;
wire net_3752;
wire net_482;
wire net_5144;
wire net_10805;
wire net_3258;
wire net_20148;
wire net_10942;
wire net_149;
wire net_15437;
wire net_7790;
wire net_21600;
wire net_13107;
wire net_13127;
wire net_19596;
wire net_5160;
wire net_15995;
wire net_6494;
wire net_14137;
wire net_15035;
wire net_577;
wire net_3401;
wire net_13245;
wire net_10313;
wire net_2550;
wire net_797;
wire net_21738;
wire net_7747;
wire net_21818;
wire net_3545;
wire net_1799;
wire net_10150;
wire net_11224;
wire net_15132;
wire net_22410;
wire net_21916;
wire net_16092;
wire net_11859;
wire net_22564;
wire net_18544;
wire net_9218;
wire net_12909;
wire net_337;
wire net_10581;
wire net_13312;
wire net_4476;
wire net_20759;
wire net_690;
wire net_17729;
wire net_6820;
wire net_7933;
wire net_20396;
wire net_3743;
wire net_523;
wire net_21909;
wire net_11070;
wire net_6718;
wire net_7144;
wire net_21418;
wire net_20800;
wire net_3375;
wire net_6744;
wire net_9620;
wire net_18620;
wire net_22381;
wire net_4926;
wire net_19471;
wire net_3467;
wire net_16637;
wire net_9617;
wire net_15785;
wire net_21688;
wire net_8972;
wire net_9760;
wire net_20160;
wire net_17243;
wire net_16439;
wire net_4467;
wire net_20607;
wire net_21544;
wire net_12129;
wire net_5028;
wire net_4721;
wire net_18179;
wire net_5756;
wire net_18999;
wire net_1631;
wire net_4426;
wire net_16955;
wire net_1337;
wire net_21877;
wire net_5786;
wire net_1182;
wire net_14254;
wire net_17768;
wire net_7231;
wire net_16286;
wire net_13656;
wire net_14458;
wire net_18244;
wire net_1950;
wire net_9052;
wire net_15067;
wire net_18973;
wire net_9280;
wire x3163;
wire net_7039;
wire net_14803;
wire net_2421;
wire net_5684;
wire net_19152;
wire net_4901;
wire net_4804;
wire net_880;
wire net_1402;
wire net_18784;
wire net_18337;
wire net_4100;
wire net_18028;
wire net_8474;
wire net_17470;
wire net_16600;
wire net_8535;
wire net_20905;
wire net_19979;
wire net_5151;
wire net_21493;
wire net_21035;
wire net_16309;
wire net_13922;
wire net_2901;
wire net_11876;
wire net_15792;
wire net_21513;
wire net_4950;
wire net_13255;
wire net_4944;
wire net_18103;
wire net_20026;
wire net_18298;
wire net_20969;
wire net_4847;
wire net_12661;
wire net_3052;
wire net_6652;
wire net_10906;
wire net_7295;
wire net_11554;
wire net_6368;
wire net_16939;
wire net_14889;
wire net_487;
wire net_7992;
wire net_8861;
wire net_17785;
wire net_5056;
wire net_756;
wire net_7735;
wire net_13636;
wire net_22139;
wire net_4765;
wire net_17614;
wire net_14234;
wire net_7798;
wire net_10101;
wire net_12230;
wire net_17841;
wire net_5031;
wire net_11301;
wire net_15477;
wire net_17319;
wire net_72;
wire x603;
wire net_17724;
wire net_11845;
wire net_3537;
wire net_18447;
wire net_15541;
wire net_12897;
wire net_2225;
wire net_7659;
wire net_21978;
wire net_16356;
wire net_16342;
wire net_17104;
wire net_16917;
wire net_15257;
wire net_4741;
wire net_22630;
wire net_11687;
wire net_16334;
wire net_15720;
wire net_9402;
wire net_10469;
wire net_12852;
wire net_16501;
wire net_11420;
wire net_21009;
wire x668;
wire net_174;
wire net_7987;
wire net_7214;
wire net_15208;
wire net_1831;
wire net_6202;
wire net_11691;
wire net_1482;
wire net_19315;
wire net_17600;
wire net_3291;
wire net_2928;
wire net_3306;
wire net_14573;
wire net_21082;
wire net_17829;
wire net_7563;
wire net_14460;
wire net_1485;
wire net_4129;
wire net_9236;
wire net_10272;
wire net_10053;
wire net_3245;
wire net_13300;
wire net_16902;
wire net_9385;
wire net_7473;
wire net_6920;
wire net_21757;
wire net_7335;
wire net_14742;
wire net_22294;
wire net_7387;
wire net_19181;
wire net_11987;
wire net_10787;
wire net_12711;
wire net_12740;
wire net_13407;
wire net_13929;
wire net_745;
wire net_9651;
wire net_14737;
wire net_17774;
wire net_16352;
wire net_14271;
wire net_1244;
wire net_15919;
wire net_429;
wire net_10966;
wire net_12593;
wire net_20862;
wire net_356;
wire net_13701;
wire net_545;
wire net_11432;
wire net_2147;
wire net_11700;
wire net_10361;
wire net_560;
wire net_9253;
wire net_10098;
wire net_5148;
wire net_4603;
wire net_15120;
wire net_14017;
wire net_17705;
wire net_15586;
wire net_17984;
wire net_5510;
wire net_11951;
wire net_9359;
wire net_10500;
wire net_6709;
wire net_22446;
wire net_7310;
wire net_16874;
wire net_13151;
wire net_20846;
wire net_7522;
wire net_2872;
wire net_20542;
wire net_2432;
wire net_6833;
wire net_12780;
wire net_5401;
wire net_322;
wire net_420;
wire net_2322;
wire net_8944;
wire net_19874;
wire net_4344;
wire net_9109;
wire net_3341;
wire net_13376;
wire net_20682;
wire net_1072;
wire net_7136;
wire net_13738;
wire net_18737;
wire net_15527;
wire net_4510;
wire net_11113;
wire net_19014;
wire net_6278;
wire net_1730;
wire net_6311;
wire net_22797;
wire net_4575;
wire net_13501;
wire net_651;
wire net_15766;
wire net_18370;
wire net_14653;
wire net_2931;
wire net_12097;
wire net_6846;
wire net_21962;
wire net_18250;
wire net_17965;
wire net_598;
wire net_4967;
wire net_18709;
wire net_3455;
wire net_6317;
wire net_12011;
wire net_10068;
wire net_21734;
wire net_16421;
wire net_18438;
wire net_4818;
wire net_2820;
wire net_8690;
wire net_6091;
wire net_8348;
wire net_21698;
wire net_21613;
wire net_20586;
wire net_18914;
wire net_18689;
wire net_4404;
wire net_3068;
wire net_5973;
wire net_8585;
wire net_3892;
wire net_7921;
wire net_21702;
wire net_22437;
wire net_18183;
wire net_7080;
wire net_17911;
wire net_5978;
wire net_6739;
wire net_632;
wire net_21552;
wire net_20889;
wire net_843;
wire net_3860;
wire net_15652;
wire net_15603;
wire net_12720;
wire net_16759;
wire net_19245;
wire net_10063;
wire net_5484;
wire net_20574;
wire x7235;
wire net_2100;
wire net_11959;
wire net_2122;
wire net_19992;
wire net_6617;
wire net_12572;
wire net_18396;
wire net_19970;
wire net_1540;
wire net_20145;
wire net_22094;
wire net_9734;
wire net_11835;
wire net_18655;
wire net_1725;
wire net_10393;
wire net_22354;
wire net_3541;
wire net_16532;
wire net_18789;
wire net_21590;
wire net_5649;
wire net_3532;
wire net_13718;
wire net_12725;
wire net_17307;
wire net_5112;
wire net_18149;
wire net_17700;
wire net_21812;
wire net_5190;
wire net_9750;
wire net_10303;
wire x4139;
wire net_6554;
wire net_14712;
wire net_20372;
wire net_503;
wire net_7504;
wire net_19265;
wire net_16676;
wire net_13510;
wire net_18798;
wire net_5695;
wire net_2103;
wire net_1672;
wire net_11818;
wire net_996;
wire net_3091;
wire net_14165;
wire net_2994;
wire net_16510;
wire net_11617;
wire net_10838;
wire net_8327;
wire net_17504;
wire net_21059;
wire net_4004;
wire net_8767;
wire net_7706;
wire net_18705;
wire net_18605;
wire net_2973;
wire net_9304;
wire net_12342;
wire net_19065;
wire net_3106;
wire net_19895;
wire net_21191;
wire net_13792;
wire net_21010;
wire net_20659;
wire net_22397;
wire net_2503;
wire net_16683;
wire net_20804;
wire net_9705;
wire net_15170;
wire net_6646;
wire net_20055;
wire net_19584;
wire net_17834;
wire net_20514;
wire net_6469;
wire net_13578;
wire net_18565;
wire net_8330;
wire net_22657;
wire net_9821;
wire net_18889;
wire net_6211;
wire net_13670;
wire net_3721;
wire net_4606;
wire net_10556;
wire net_10982;
wire net_21245;
wire net_8894;
wire net_6572;
wire net_12397;
wire net_21595;
wire net_7416;
wire net_11677;
wire net_22190;
wire net_15064;
wire net_6901;
wire net_14726;
wire net_5051;
wire net_20634;
wire net_10688;
wire net_2469;
wire net_11214;
wire net_21172;
wire net_17229;
wire net_14819;
wire net_15938;
wire net_18545;
wire net_21961;
wire net_17421;
wire net_1404;
wire net_1012;
wire net_10458;
wire net_14824;
wire net_20093;
wire net_20201;
wire net_5807;
wire net_8809;
wire net_4694;
wire net_2036;
wire net_395;
wire net_15124;
wire net_12988;
wire net_15448;
wire net_22674;
wire net_8070;
wire net_9182;
wire net_10219;
wire net_17064;
wire net_8623;
wire net_2323;
wire net_3867;
wire net_16223;
wire net_3677;
wire net_4811;
wire net_15088;
wire net_22077;
wire net_16864;
wire net_5451;
wire net_20259;
wire net_15336;
wire net_4972;
wire net_10599;
wire net_10459;
wire net_19533;
wire net_17032;
wire net_1901;
wire net_4890;
wire net_8429;
wire net_3021;
wire net_22427;
wire net_3711;
wire net_21373;
wire net_19832;
wire net_7580;
wire net_19514;
wire net_602;
wire net_4580;
wire net_12605;
wire net_2379;
wire net_8273;
wire net_20988;
wire net_2918;
wire net_10932;
wire net_12288;
wire net_16084;
wire net_1497;
wire net_11658;
wire net_1800;
wire net_18590;
wire net_4634;
wire net_14480;
wire net_279;
wire net_21559;
wire net_19589;
wire net_3347;
wire net_12281;
wire net_18440;
wire net_4039;
wire net_4030;
wire net_11326;
wire net_10212;
wire net_6337;
wire net_10713;
wire net_15506;
wire net_19100;
wire net_14119;
wire net_4078;
wire net_14289;
wire net_2833;
wire net_2561;
wire net_12170;
wire net_21511;
wire net_15224;
wire net_17801;
wire net_18326;
wire net_18007;
wire net_13775;
wire net_20619;
wire net_17183;
wire net_22649;
wire net_3813;
wire net_16599;
wire net_18587;
wire net_20219;
wire net_1531;
wire net_1159;
wire net_21699;
wire net_10666;
wire net_19636;
wire net_861;
wire net_10334;
wire net_6755;
wire net_20385;
wire net_7217;
wire net_12645;
wire net_6696;
wire net_21230;
wire net_12400;
wire net_19611;
wire net_11102;
wire net_4914;
wire net_19288;
wire net_17658;
wire net_21316;
wire net_8544;
wire net_10882;
wire net_15814;
wire net_5213;
wire net_12951;
wire net_7696;
wire net_21986;
wire net_8567;
wire net_4552;
wire net_16946;
wire net_21534;
wire net_21771;
wire net_1527;
wire net_18963;
wire net_13270;
wire net_21100;
wire net_268;
wire net_11849;
wire net_21279;
wire net_3386;
wire net_48;
wire net_4134;
wire net_22805;
wire net_6631;
wire net_13324;
wire net_15627;
wire net_9406;
wire net_17135;
wire net_17117;
wire net_14536;
wire net_3638;
wire net_2570;
wire net_19040;
wire net_5793;
wire net_22207;
wire net_3354;
wire net_13195;
wire net_22113;
wire net_16558;
wire net_9468;
wire net_2712;
wire net_2005;
wire net_13976;
wire net_14827;
wire net_2771;
wire net_1123;
wire net_19192;
wire net_4897;
wire net_6040;
wire net_18947;
wire net_9343;
wire net_13911;
wire net_20565;
wire net_9980;
wire net_19359;
wire net_11241;
wire net_4838;
wire net_5958;
wire net_20965;
wire net_3363;
wire net_984;
wire net_11894;
wire net_5467;
wire net_6407;
wire net_7263;
wire net_10915;
wire net_22764;
wire net_13652;
wire net_1105;
wire net_22044;
wire net_12370;
wire x161;
wire net_20158;
wire net_2172;
wire net_11448;
wire net_19647;
wire net_14023;
wire net_15904;
wire x90;
wire net_16718;
wire net_7491;
wire net_18407;
wire net_4457;
wire net_9519;
wire net_22149;
wire net_1856;
wire net_830;
wire net_16205;
wire net_1279;
wire net_14642;
wire net_1047;
wire net_20244;
wire net_18019;
wire net_13003;
wire net_9475;
wire net_18523;
wire net_18080;
wire net_12642;
wire net_6394;
wire net_8439;
wire net_18698;
wire net_14553;
wire net_4688;
wire net_11425;
wire net_17339;
wire net_2631;
wire net_16129;
wire net_8101;
wire net_16906;
wire net_19579;
wire net_12386;
wire net_21668;
wire net_19778;
wire net_12926;
wire net_1467;
wire net_3181;
wire net_1061;
wire net_5623;
wire net_5951;
wire net_18121;
wire net_19841;
wire net_3837;
wire net_9096;
wire net_22556;
wire net_2288;
wire net_4839;
wire net_14843;
wire net_8718;
wire net_13752;
wire net_11189;
wire net_15213;
wire net_18763;
wire net_19311;
wire net_17414;
wire net_16320;
wire net_17681;
wire net_21017;
wire net_15200;
wire net_3983;
wire net_14378;
wire net_8121;
wire net_19331;
wire net_3814;
wire net_15730;
wire net_10534;
wire net_6266;
wire net_2072;
wire net_18691;
wire net_1872;
wire net_16233;
wire net_20743;
wire net_1716;
wire net_13926;
wire net_5003;
wire net_1607;
wire net_5247;
wire net_11768;
wire net_13472;
wire net_17222;
wire net_1263;
wire net_16377;
wire net_12331;
wire net_22360;
wire net_17924;
wire net_3452;
wire net_196;
wire net_4591;
wire net_8766;
wire net_11969;
wire net_14356;
wire net_2067;
wire net_8120;
wire net_14243;
wire net_8881;
wire net_5183;
wire net_7200;
wire net_21462;
wire net_18098;
wire net_1639;
wire net_16193;
wire net_5267;
wire net_4126;
wire net_4549;
wire net_7284;
wire net_3625;
wire net_11431;
wire net_22035;
wire net_14435;
wire net_4145;
wire net_7604;
wire net_20208;
wire net_22142;
wire net_15145;
wire net_2152;
wire net_732;
wire net_11981;
wire net_12880;
wire net_19661;
wire net_5286;
wire net_6105;
wire net_8285;
wire net_2088;
wire net_21892;
wire net_13083;
wire net_19189;
wire net_6423;
wire net_7572;
wire net_13963;
wire net_2689;
wire net_4217;
wire net_10655;
wire net_20528;
wire net_17646;
wire net_17121;
wire net_8422;
wire net_22219;
wire net_21831;
wire net_11678;
wire net_15399;
wire net_11092;
wire net_15935;
wire net_13970;
wire net_449;
wire net_5234;
wire net_8225;
wire net_11523;
wire net_1087;
wire net_15697;
wire net_18806;
wire net_4234;
wire net_11064;
wire net_3995;
wire net_21573;
wire net_733;
wire net_887;
wire net_8245;
wire net_5856;
wire net_18011;
wire net_18865;
wire net_6098;
wire net_20198;
wire net_7537;
wire net_11975;
wire net_21626;
wire net_6151;
wire net_10491;
wire net_2308;
wire net_6301;
wire net_19248;
wire net_9105;
wire net_19954;
wire x4319;
wire net_40;
wire net_4628;
wire net_2770;
wire net_19485;
wire net_2636;
wire net_1424;
wire net_4375;
wire net_19043;
wire net_21185;
wire net_4412;
wire net_22056;
wire net_16840;
wire net_9287;
wire net_17391;
wire net_18834;
wire net_21286;
wire net_21970;
wire net_8167;
wire net_4280;
wire net_10347;
wire net_9563;
wire net_19384;
wire net_950;
wire net_22174;
wire net_21397;
wire net_22822;
wire net_11441;
wire net_20623;
wire net_19680;
wire net_20725;
wire net_19414;
wire net_21550;
wire net_9839;
wire net_2816;
wire net_17435;
wire net_6610;
wire net_7651;
wire net_14507;
wire net_18959;
wire net_14344;
wire net_1214;
wire net_3641;
wire net_9529;
wire net_20175;
wire net_866;
wire net_12895;
wire net_20941;
wire x222;
wire net_4220;
wire net_12700;
wire net_15705;
wire net_10681;
wire net_18704;
wire net_18047;
wire net_1032;
wire net_567;
wire net_15563;
wire net_13985;
wire net_3726;
wire net_5255;
wire net_18506;
wire net_272;
wire net_5787;
wire net_13345;
wire net_8458;
wire net_13384;
wire net_3939;
wire net_14625;
wire net_1024;
wire net_12480;
wire net_21158;
wire net_21073;
wire net_1590;
wire net_22103;
wire net_14097;
wire net_18495;
wire net_1612;
wire net_17268;
wire net_814;
wire net_11121;
wire net_21729;
wire net_13685;
wire net_17320;
wire x2428;
wire net_5840;
wire net_8128;
wire net_22783;
wire net_6184;
wire net_12705;
wire net_12525;
wire net_17641;
wire net_14003;
wire net_3930;
wire net_4785;
wire net_10639;
wire net_9815;
wire net_3299;
wire net_2586;
wire net_15795;
wire net_1655;
wire net_10290;
wire net_6963;
wire net_2365;
wire net_15951;
wire net_17803;
wire net_18306;
wire net_17179;
wire net_22170;
wire net_19208;
wire net_21321;
wire net_4797;
wire net_9240;
wire net_10810;
wire net_2598;
wire net_2361;
wire net_18031;
wire net_11194;
wire net_14767;
wire net_17717;
wire net_2879;
wire net_1680;
wire net_14219;
wire net_16172;
wire net_16258;
wire net_3302;
wire net_20436;
wire net_17481;
wire net_7540;
wire net_15276;
wire net_15925;
wire net_11337;
wire net_3187;
wire net_15250;
wire net_2622;
wire net_84;
wire net_5966;
wire net_20599;
wire net_10514;
wire net_8294;
wire net_17690;
wire net_10997;
wire net_22506;
wire net_14500;
wire net_2262;
wire net_22716;
wire net_7505;
wire net_20757;
wire net_22367;
wire net_2087;
wire net_1002;
wire net_21943;
wire net_7620;
wire net_7224;
wire net_6118;
wire net_3188;
wire net_13308;
wire net_19276;
wire x1686;
wire net_17259;
wire net_1993;
wire net_8198;
wire net_11128;
wire net_8724;
wire net_2903;
wire net_8683;
wire net_11623;
wire net_8392;
wire net_9556;
wire net_4128;
wire net_16262;
wire net_4923;
wire net_21616;
wire net_3873;
wire net_11866;
wire net_6015;
wire net_2155;
wire net_6741;
wire net_168;
wire net_15056;
wire net_19070;
wire net_17194;
wire net_385;
wire net_2609;
wire net_13253;
wire net_14179;
wire net_5365;
wire net_5736;
wire net_5404;
wire net_5044;
wire net_14890;
wire net_8657;
wire net_10260;
wire net_8139;
wire net_10468;
wire net_6236;
wire net_11220;
wire net_7660;
wire net_13675;
wire net_2380;
wire net_3393;
wire net_4548;
wire net_19990;
wire net_8231;
wire net_20605;
wire net_16031;
wire net_9323;
wire x2344;
wire net_20234;
wire net_16135;
wire net_14797;
wire net_19779;
wire net_19055;
wire net_1412;
wire net_16524;
wire net_19808;
wire net_17816;
wire net_15402;
wire net_12327;
wire net_12965;
wire net_20629;
wire net_13357;
wire net_7358;
wire net_7211;
wire net_16666;
wire net_19088;
wire net_19948;
wire net_3040;
wire net_3557;
wire net_10825;
wire net_13762;
wire net_10609;
wire net_15975;
wire net_21820;
wire net_8801;
wire net_3004;
wire net_18453;
wire net_8014;
wire net_21990;
wire x3608;
wire net_12624;
wire net_7244;
wire net_17631;
wire net_7981;
wire net_10315;
wire net_16500;
wire net_3830;
wire net_9757;
wire net_8464;
wire net_22195;
wire net_19932;
wire net_17756;
wire net_22371;
wire net_12561;
wire net_12806;
wire net_10282;
wire net_18177;
wire net_833;
wire net_14044;
wire net_99;
wire net_12744;
wire net_6656;
wire net_17914;
wire x3178;
wire net_4758;
wire net_4249;
wire net_14512;
wire net_14757;
wire net_12931;
wire net_1399;
wire net_11349;
wire net_13681;
wire net_19591;
wire net_21750;
wire net_16270;
wire net_8529;
wire net_8667;
wire net_3350;
wire net_15877;
wire net_3553;
wire net_5161;
wire net_14489;
wire net_19158;
wire net_20521;
wire net_16578;
wire net_20705;
wire net_7623;
wire net_15416;
wire net_20363;
wire net_16277;
wire net_20087;
wire net_12751;
wire net_1781;
wire net_16067;
wire net_18998;
wire net_3049;
wire net_7457;
wire net_20351;
wire net_10299;
wire net_6918;
wire net_22270;
wire net_17572;
wire net_2514;
wire net_9250;
wire net_12183;
wire net_3474;
wire net_4775;
wire net_16754;
wire net_2013;
wire x4668;
wire net_5472;
wire net_15990;
wire net_7477;
wire net_13503;
wire net_20855;
wire net_97;
wire net_11262;
wire net_18556;
wire x539;
wire net_17869;
wire net_2028;
wire net_9758;
wire net_1889;
wire net_3766;
wire net_7361;
wire net_12065;
wire net_8717;
wire net_2981;
wire net_19972;
wire net_17895;
wire net_1164;
wire net_6810;
wire net_8912;
wire net_10817;
wire net_15528;
wire net_14449;
wire net_6923;
wire net_11148;
wire net_12500;
wire net_2583;
wire net_5708;
wire net_8854;
wire net_4665;
wire net_5824;
wire net_9366;
wire net_16525;
wire net_2706;
wire net_5163;
wire net_5580;
wire net_11842;
wire net_8304;
wire net_2602;
wire net_6366;
wire net_8449;
wire x532;
wire net_17970;
wire net_4484;
wire net_21309;
wire net_440;
wire net_21039;
wire net_22700;
wire net_8069;
wire net_8048;
wire net_10866;
wire net_17021;
wire net_5664;
wire net_14747;
wire net_21518;
wire net_16799;
wire net_4652;
wire net_14558;
wire net_718;
wire net_21470;
wire net_6178;
wire net_7773;
wire net_20018;
wire net_18023;
wire net_18243;
wire net_19538;
wire net_14193;
wire net_21302;
wire net_8707;
wire net_22458;
wire net_5714;
wire net_12995;
wire net_19216;
wire net_19723;
wire net_13367;
wire net_5838;
wire net_12215;
wire net_13946;
wire net_17579;
wire net_22451;
wire x132;
wire net_13545;
wire net_14078;
wire net_4448;
wire net_16985;
wire net_336;
wire net_9419;
wire net_15598;
wire net_10404;
wire net_14033;
wire net_1578;
wire net_14584;
wire x1204;
wire net_18464;
wire net_8417;
wire net_20113;
wire net_18206;
wire net_17097;
wire net_22167;
wire net_697;
wire net_2003;
wire net_5053;
wire net_22007;
wire net_19833;
wire net_18288;
wire net_17410;
wire net_3426;
wire x1718;
wire net_13008;
wire net_15632;
wire net_5095;
wire net_1333;
wire net_20549;
wire net_5325;
wire net_21034;
wire net_5924;
wire net_18483;
wire net_5107;
wire net_5593;
wire net_17662;
wire net_3082;
wire net_14422;
wire net_22279;
wire net_5859;
wire net_10802;
wire net_11503;
wire net_3676;
wire net_13521;
wire net_4185;
wire net_4204;
wire net_20828;
wire net_5630;
wire net_6072;
wire net_7591;
wire net_2054;
wire net_6682;
wire net_21065;
wire net_20925;
wire net_9880;
wire net_17665;
wire net_128;
wire net_6295;
wire net_20100;
wire net_9133;
wire net_19732;
wire net_14057;
wire net_10901;
wire net_14133;
wire net_15160;
wire net_2793;
wire net_18459;
wire net_1836;
wire net_14971;
wire net_4310;
wire net_8783;
wire net_10570;
wire net_20811;
wire net_5922;
wire net_13158;
wire net_14571;
wire net_3430;
wire net_11557;
wire net_8266;
wire net_6795;
wire net_15016;
wire net_21168;
wire net_4244;
wire net_14882;
wire net_18220;
wire net_7887;
wire net_15779;
wire net_6930;
wire net_4396;
wire net_6158;
wire net_21649;
wire net_21865;
wire net_9273;
wire net_21985;
wire net_22616;
wire net_16361;
wire net_2398;
wire x4888;
wire net_4581;
wire net_7811;
wire net_12140;
wire net_4431;
wire net_7821;
wire net_15374;
wire net_20620;
wire net_3315;
wire net_16580;
wire net_2455;
wire net_17624;
wire net_19077;
wire net_20554;
wire net_22499;
wire net_12732;
wire net_21789;
wire net_17400;
wire net_10753;
wire net_8493;
wire net_8744;
wire net_18124;
wire net_21473;
wire net_1386;
wire net_7841;
wire net_9431;
wire x346;
wire net_21346;
wire net_6546;
wire net_8949;
wire net_16150;
wire net_6115;
wire net_10550;
wire net_12805;
wire net_5991;
wire net_5101;
wire net_10252;
wire net_14968;
wire net_14989;
wire net_2186;
wire net_3696;
wire net_22418;
wire net_3473;
wire net_13551;
wire net_17231;
wire net_569;
wire net_12062;
wire net_13877;
wire net_16781;
wire net_12767;
wire net_21854;
wire net_20227;
wire net_19298;
wire net_8857;
wire x4496;
wire net_21139;
wire net_21290;
wire net_4018;
wire net_17439;
wire net_17281;
wire net_6826;
wire net_19128;
wire net_20863;
wire net_15249;
wire net_21450;
wire net_13696;
wire x2481;
wire net_18710;
wire net_3124;
wire net_1903;
wire net_2407;
wire x452;
wire net_13467;
wire net_10600;
wire net_13162;
wire net_7412;
wire net_13414;
wire net_17907;
wire net_2078;
wire net_779;
wire net_16511;
wire net_22469;
wire net_12473;
wire net_14438;
wire net_234;
wire net_20612;
wire x3463;
wire x1674;
wire net_4151;
wire net_12634;
wire net_5142;
wire net_13258;
wire net_17126;
wire net_16632;
wire net_15309;
wire net_5764;
wire net_7390;
wire net_11469;
wire net_17653;
wire net_7732;
wire net_20537;
wire net_6583;
wire net_19782;
wire net_19565;
wire net_9128;
wire net_491;
wire net_11460;
wire net_1299;
wire net_948;
wire net_6679;
wire net_19437;
wire net_18599;
wire net_11573;
wire net_20126;
wire net_17462;
wire net_17109;
wire net_2593;
wire net_876;
wire net_6479;
wire net_15841;
wire net_2162;
wire net_18820;
wire net_10833;
wire net_15424;
wire net_7154;
wire net_9646;
wire net_16041;
wire net_8601;
wire net_11960;
wire net_1458;
wire net_18160;
wire net_5587;
wire net_20712;
wire net_17160;
wire net_10184;
wire net_5933;
wire net_16977;
wire net_905;
wire net_10591;
wire net_14122;
wire net_20048;
wire net_142;
wire net_2229;
wire net_21107;
wire net_158;
wire net_5774;
wire net_10613;
wire net_13842;
wire net_7370;
wire net_3200;
wire net_14848;
wire net_19039;
wire net_19911;
wire net_16181;
wire net_15457;
wire net_5624;
wire net_16011;
wire net_2504;
wire net_11571;
wire net_2175;
wire net_3784;
wire net_5650;
wire net_18882;
wire net_10214;
wire net_15637;
wire net_21671;
wire net_2116;
wire net_4327;
wire net_14701;
wire net_11334;
wire net_22817;
wire net_8035;
wire net_16973;
wire net_8090;
wire net_9572;
wire net_1967;
wire net_22628;
wire net_21843;
wire x5053;
wire net_11565;
wire net_5171;
wire net_9333;
wire net_21060;
wire net_6860;
wire net_8754;
wire net_16481;
wire net_465;
wire x6764;
wire net_14676;
wire net_1883;
wire net_17948;
wire net_11233;
wire net_17381;
wire net_3058;
wire net_20159;
wire net_8484;
wire net_1315;
wire net_6994;
wire net_22134;
wire x1247;
wire net_5904;
wire net_20744;
wire net_5358;
wire net_10073;
wire net_15790;
wire net_19393;
wire net_19116;
wire net_5208;
wire net_9767;
wire net_22065;
wire net_5019;
wire net_13144;
wire net_6956;
wire net_9376;
wire net_9903;
wire net_19628;
wire net_4977;
wire net_10138;
wire net_5075;
wire net_11646;
wire net_7327;
wire net_293;
wire net_15117;
wire net_3666;
wire net_11890;
wire net_21141;
wire net_1938;
wire net_13303;
wire net_15677;
wire net_20915;
wire net_1823;
wire net_14660;
wire net_5081;
wire net_21431;
wire net_15516;
wire net_3576;
wire net_191;
wire net_21689;
wire net_558;
wire net_2069;
wire net_15021;
wire net_20458;
wire net_1618;
wire net_10910;
wire net_14399;
wire net_19622;
wire net_2497;
wire net_11594;
wire net_3562;
wire net_7006;
wire net_15319;
wire net_15110;
wire net_5885;
wire net_7112;
wire net_11905;
wire net_18893;
wire net_4023;
wire net_14720;
wire net_15853;
wire net_7755;
wire net_4450;
wire net_6881;
wire net_15610;
wire net_6942;
wire net_1984;
wire net_20763;
wire net_13959;
wire net_4670;
wire net_10734;
wire net_16436;
wire net_1944;
wire net_11545;
wire net_19142;
wire net_1775;
wire net_10112;
wire net_16993;
wire net_297;
wire net_346;
wire net_10158;
wire net_22378;
wire net_22408;
wire net_20272;
wire net_17956;
wire net_10693;
wire net_13725;
wire net_15982;
wire net_15870;
wire net_229;
wire net_14835;
wire net_4360;
wire net_4962;
wire net_19871;
wire net_687;
wire net_17334;
wire net_15073;
wire net_3266;
wire net_4160;
wire net_13339;
wire net_14702;
wire net_17265;
wire net_3888;
wire net_7072;
wire net_13949;
wire net_14303;
wire net_20472;
wire net_3566;
wire net_15263;
wire net_14945;
wire net_3596;
wire net_10143;
wire net_5021;
wire x7366;
wire net_13741;
wire net_9296;
wire net_9345;
wire net_5415;
wire net_1184;
wire net_13492;
wire x361;
wire net_4055;
wire net_5339;
wire net_18268;
wire net_6482;
wire net_18924;
wire net_6961;
wire net_14444;
wire net_19556;
wire net_21054;
wire net_7383;
wire net_15363;
wire net_10722;
wire net_5425;
wire net_1960;
wire net_9660;
wire net_19191;
wire net_15622;
wire net_7435;
wire net_12548;
wire net_15194;
wire net_828;
wire net_4256;
wire net_9145;
wire net_6222;
wire net_1603;
wire net_4490;
wire net_12222;
wire net_14349;
wire net_13031;
wire net_18728;
wire net_7446;
wire net_10009;
wire net_22085;
wire net_10108;
wire x577;
wire net_11017;
wire net_18981;
wire net_18321;
wire net_8385;
wire net_3521;
wire net_14877;
wire net_982;
wire net_14874;
wire net_9610;
wire net_19519;
wire net_21906;
wire net_1580;
wire net_19962;
wire net_3896;
wire net_5287;
wire net_4384;
wire net_6462;
wire net_9189;
wire net_19805;
wire net_17189;
wire net_9314;
wire net_19466;
wire net_9576;
wire net_4912;
wire net_6002;
wire net_14501;
wire net_15863;
wire net_5748;
wire net_12076;
wire net_15531;
wire net_8180;
wire net_5049;
wire net_10869;
wire net_11393;
wire net_17537;
wire net_11058;
wire net_19827;
wire net_8899;
wire net_225;
wire net_14927;
wire net_3128;
wire net_4733;
wire net_12937;
wire net_6524;
wire x779;
wire net_22011;
wire net_5313;
wire net_15334;
wire net_2611;
wire net_871;
wire net_11804;
wire net_14974;
wire net_390;
wire net_22678;
wire net_35;
wire net_20039;
wire net_1154;
wire net_22026;
wire net_11789;
wire net_6983;
wire net_6593;
wire net_20163;
wire net_11782;
wire net_20008;
wire net_16249;
wire net_4294;
wire net_22610;
wire net_5128;
wire net_6062;
wire net_15723;
wire net_12735;
wire net_7494;
wire net_12798;
wire net_19913;
wire net_19424;
wire net_280;
wire net_12132;
wire net_12027;
wire net_12715;
wire net_495;
wire net_13022;
wire net_16317;
wire net_10569;
wire net_2140;
wire net_13180;
wire net_6345;
wire net_13975;
wire net_15965;
wire net_16124;
wire net_13211;
wire net_2517;
wire net_20144;
wire net_8798;
wire net_2316;
wire net_12105;
wire net_8644;
wire net_6457;
wire net_14525;
wire net_6100;
wire net_6356;
wire net_2703;
wire net_19758;
wire net_11273;
wire net_13524;
wire net_14214;
wire net_1441;
wire net_18814;
wire net_969;
wire net_9154;
wire net_1525;
wire net_7097;
wire net_12710;
wire net_17443;
wire net_11458;
wire net_821;
wire net_4003;
wire net_13444;
wire net_4177;
wire net_9350;
wire net_18302;
wire net_8936;
wire net_8345;
wire net_2335;
wire net_11210;
wire net_19822;
wire net_3940;
wire net_14603;
wire net_21910;
wire net_18352;
wire net_11533;
wire net_11161;
wire net_14153;
wire net_19372;
wire net_2618;
wire net_4316;
wire net_19671;
wire net_6045;
wire net_20670;
wire net_6540;
wire net_21428;
wire net_14688;
wire net_16571;
wire net_7952;
wire net_20315;
wire net_16497;
wire net_12786;
wire net_8670;
wire net_20932;
wire net_5411;
wire net_19498;
wire net_12691;
wire net_21330;
wire net_1748;
wire net_3078;
wire net_2964;
wire net_11882;
wire net_9946;
wire net_16589;
wire net_2343;
wire net_2232;
wire net_726;
wire net_13241;
wire net_15349;
wire net_3237;
wire net_701;
wire net_808;
wire net_5553;
wire net_9121;
wire net_22680;
wire net_1704;
wire net_4821;
wire net_5026;
wire net_2738;
wire net_16432;
wire net_21256;
wire net_2944;
wire net_18624;
wire net_22526;
wire net_18259;
wire net_12079;
wire net_20842;
wire net_14384;
wire net_17709;
wire net_6662;
wire net_11176;
wire net_18417;
wire net_9451;
wire net_13058;
wire net_7927;
wire net_17247;
wire net_19268;
wire net_5654;
wire net_16845;
wire net_13034;
wire net_19250;
wire net_935;
wire net_8827;
wire net_19791;
wire net_3116;
wire net_1511;
wire net_645;
wire net_11436;
wire net_14649;
wire net_4071;
wire net_17005;
wire net_14242;
wire net_8825;
wire net_10862;
wire net_20102;
wire net_17428;
wire net_4533;
wire net_17963;
wire net_17145;
wire net_1816;
wire net_8076;
wire net_22544;
wire net_16149;
wire net_4195;
wire net_7909;
wire net_14085;
wire net_21154;
wire net_331;
wire net_12597;
wire net_17853;
wire net_20379;
wire net_4644;
wire net_19856;
wire net_8633;
wire net_2220;
wire net_4762;
wire net_2823;
wire net_19405;
wire x3001;
wire net_20034;
wire net_22640;
wire net_3728;
wire net_21562;
wire net_5724;
wire net_7138;
wire net_22634;
wire net_22703;
wire net_4884;
wire net_12981;
wire net_8000;
wire net_15537;
wire net_12541;
wire net_15764;
wire net_13808;
wire net_16399;
wire net_12841;
wire net_14333;
wire net_16615;
wire net_12199;
wire net_16928;
wire net_1259;
wire net_4753;
wire net_11207;
wire net_2839;
wire net_2143;
wire net_4225;
wire net_2196;
wire net_3791;
wire net_7676;
wire net_8059;
wire net_10478;
wire net_21503;
wire net_5275;
wire net_11611;
wire net_21089;
wire net_478;
wire net_16672;
wire net_22346;
wire net_6608;
wire net_11429;
wire net_4959;
wire net_5781;
wire net_8733;
wire net_1975;
wire net_19747;
wire net_8958;
wire net_8375;
wire net_13067;
wire net_11948;
wire net_13991;
wire net_5600;
wire net_17986;
wire net_7406;
wire net_17369;
wire net_7530;
wire net_20305;
wire net_7253;
wire net_3028;
wire net_18432;
wire net_17073;
wire net_22477;
wire net_19694;
wire net_21355;
wire net_11281;
wire net_1692;
wire net_7087;
wire net_21384;
wire net_5079;
wire net_12675;
wire net_2655;
wire net_2528;
wire net_22018;
wire net_16588;
wire net_18100;
wire net_10854;
wire net_9682;
wire net_1361;
wire net_21198;
wire net_16744;
wire net_2450;
wire net_9260;
wire net_14118;
wire net_19774;
wire x3209;
wire net_1208;
wire net_7948;
wire net_16161;
wire net_22573;
wire net_8920;
wire net_13201;
wire net_12162;
wire net_18600;
wire net_20333;
wire net_8560;
wire net_13769;
wire net_21146;
wire net_9279;
wire net_12954;
wire net_4710;
wire net_13378;
wire net_22819;
wire net_18780;
wire net_4808;
wire net_13810;
wire net_2889;
wire net_5506;
wire net_19161;
wire net_9537;
wire net_16731;
wire net_4544;
wire net_17887;
wire net_16504;
wire net_7340;
wire net_13901;
wire net_12187;
wire net_137;
wire net_6398;
wire net_3154;
wire net_4828;
wire net_19304;
wire net_15568;
wire net_16088;
wire net_15929;
wire net_9862;
wire net_3622;
wire net_13190;
wire net_9800;
wire net_10398;
wire net_21630;
wire net_2729;
wire net_10389;
wire net_19048;
wire net_4422;
wire net_16251;
wire net_10116;
wire net_19348;
wire net_302;
wire net_18954;
wire net_1131;
wire net_21651;
wire net_753;
wire net_20909;
wire net_17283;
wire net_15668;
wire net_9034;
wire net_5575;
wire net_20895;
wire net_18330;
wire net_9710;
wire net_12464;
wire net_13609;
wire net_8084;
wire net_4155;
wire net_13864;
wire net_6353;
wire net_11297;
wire net_19798;
wire net_6722;
wire net_22243;
wire net_8288;
wire net_6283;
wire net_12861;
wire net_19507;
wire net_5192;
wire net_12301;
wire net_13268;
wire net_1228;
wire net_10146;
wire net_7148;
wire net_17386;
wire net_7807;
wire net_2722;
wire net_13092;
wire net_16455;
wire net_9891;
wire net_19969;
wire net_12139;
wire net_6504;
wire net_9399;
wire net_8531;
wire net_12013;
wire net_13113;
wire net_16419;
wire net_15190;
wire net_8536;
wire net_11548;
wire net_11380;
wire net_17858;
wire net_13602;
wire net_11795;
wire net_1057;
wire net_2915;
wire net_17808;
wire net_7235;
wire net_15673;
wire net_20403;
wire net_20183;
wire net_5225;
wire net_10895;
wire net_22771;
wire net_6161;
wire net_19986;
wire x546;
wire net_6953;
wire net_2987;
wire net_10647;
wire net_15199;
wire net_18759;
wire net_2253;
wire net_22583;
wire net_1699;
wire net_21655;
wire net_9534;
wire net_4792;
wire net_12944;
wire net_13267;
wire net_15589;
wire x899;
wire net_19097;
wire net_11133;
wire net_11309;
wire net_16959;
wire net_18649;
wire net_2521;
wire net_6246;
wire net_12915;
wire net_21048;
wire net_11296;
wire net_19936;
wire net_1016;
wire net_16410;
wire net_6437;
wire x1457;
wire net_9035;
wire net_15256;
wire net_10017;
wire net_11315;
wire net_16970;
wire net_18248;
wire net_3977;
wire net_10323;
wire net_4567;
wire net_1744;
wire net_10201;
wire net_10417;
wire net_22130;
wire net_18664;
wire net_516;
wire net_17532;
wire net_3176;
wire net_3585;
wire net_11776;
wire net_12655;
wire net_12614;
wire net_956;
wire net_21229;
wire net_3963;
wire net_5799;
wire net_14383;
wire net_5496;
wire net_21076;
wire net_20293;
wire net_438;
wire net_15770;
wire net_8181;
wire net_18062;
wire net_8178;
wire net_18668;
wire net_19235;
wire net_2250;
wire net_12334;
wire net_3013;
wire net_5278;
wire net_5438;
wire net_19092;
wire net_13826;
wire net_3110;
wire net_2967;
wire net_19229;
wire net_21726;
wire net_21950;
wire net_19768;
wire net_10916;
wire net_8214;
wire net_13337;
wire net_17020;
wire net_7598;
wire net_6808;
wire net_18227;
wire net_10645;
wire net_13185;
wire net_20186;
wire net_17360;
wire net_21631;
wire net_22261;
wire net_15471;
wire net_22754;
wire net_3570;
wire net_15283;
wire net_17081;
wire x815;
wire net_19394;
wire net_15663;
wire net_15678;
wire net_5916;
wire net_9773;
wire net_21392;
wire net_18991;
wire net_19085;
wire net_19360;
wire net_2785;
wire net_21271;
wire net_9693;
wire net_10840;
wire net_8575;
wire net_473;
wire net_8274;
wire net_13169;
wire net_21297;
wire net_18467;
wire net_19166;
wire net_18745;
wire net_16012;
wire net_3599;
wire net_14426;
wire net_5099;
wire net_8350;
wire net_9512;
wire net_22268;
wire net_454;
wire x256;
wire net_5349;
wire net_6251;
wire net_15518;
wire net_16384;
wire net_18036;
wire net_709;
wire net_2484;
wire net_13535;
wire net_11342;
wire net_10791;
wire net_1066;
wire net_20488;
wire net_5514;
wire net_9956;
wire net_15095;
wire net_4304;
wire net_5847;
wire net_22647;
wire net_1344;
wire net_4560;
wire net_1084;
wire net_1500;
wire net_9778;
wire net_1136;
wire net_11376;
wire net_5418;
wire net_14010;
wire net_3008;
wire net_2763;
wire net_11707;
wire net_573;
wire net_22810;
wire net_18277;
wire net_9065;
wire net_20462;
wire net_12412;
wire net_6855;
wire net_13314;
wire net_15912;
wire net_17069;
wire net_3616;
wire net_11606;
wire net_9494;
wire net_19342;
wire net_17677;
wire net_21717;
wire net_5521;
wire net_8570;
wire net_13352;
wire net_5037;
wire net_19202;
wire net_3672;
wire net_6089;
wire net_11101;
wire net_9249;
wire net_21841;
wire net_14371;
wire net_11879;
wire net_5811;
wire net_21266;
wire net_20503;
wire net_941;
wire net_7560;
wire net_55;
wire net_6038;
wire net_22182;
wire net_13292;
wire net_14351;
wire net_14582;
wire net_8129;
wire net_22557;
wire net_2311;
wire net_17054;
wire net_9444;
wire net_4611;
wire net_7500;
wire net_17214;
wire net_1599;
wire net_6587;
wire net_10575;
wire net_15151;
wire net_11087;
wire net_17242;
wire net_3828;
wire net_3132;
wire net_11504;
wire net_9973;
wire net_12240;
wire net_3053;
wire net_19480;
wire net_9802;
wire net_15209;
wire net_20281;
wire net_9579;
wire net_7187;
wire net_20686;
wire net_19389;
wire net_7460;
wire net_6601;
wire net_2023;
wire net_8518;
wire net_123;
wire net_4523;
wire net_13923;
wire net_15041;
wire net_1668;
wire net_262;
wire net_527;
wire x975;
wire net_20298;
wire net_22300;
wire net_12151;
wire net_7552;
wire net_3139;
wire net_4063;
wire net_5388;
wire net_6399;
wire net_22234;
wire net_16362;
wire net_22661;
wire net_22202;
wire net_21494;
wire net_1793;
wire net_11714;
wire net_18092;
wire net_3786;
wire net_20898;
wire net_7161;
wire net_8261;
wire net_6215;
wire net_5706;
wire net_1859;
wire net_145;
wire net_12550;
wire net_22148;
wire net_15299;
wire net_8193;
wire net_10699;
wire net_10431;
wire net_2804;
wire net_4637;
wire net_11134;
wire net_21299;
wire net_188;
wire net_5535;
wire net_3753;
wire net_17699;
wire net_3319;
wire net_4353;
wire net_18855;
wire net_16425;
wire net_21497;
wire net_19960;
wire net_10160;
wire net_7141;
wire net_1077;
wire net_2924;
wire net_6520;
wire net_14163;
wire net_8969;
wire net_10050;
wire net_15700;
wire net_21929;
wire net_17638;
wire net_12318;
wire net_8022;
wire net_11825;
wire net_2410;
wire net_8281;
wire net_19696;
wire net_16913;
wire net_9208;
wire net_3108;
wire net_18423;
wire net_16895;
wire net_10975;
wire net_2185;
wire net_10445;
wire net_13103;
wire net_1321;
wire net_15780;
wire net_14263;
wire net_4441;
wire net_20243;
wire net_5392;
wire net_8741;
wire x4481;
wire net_4949;
wire net_14484;
wire net_1099;
wire net_18384;
wire net_21210;
wire net_20350;
wire net_7106;
wire net_14901;
wire net_19377;
wire net_17378;
wire net_7103;
wire net_14543;
wire net_9227;
wire net_9885;
wire net_22285;
wire net_18586;
wire net_404;
wire net_15185;
wire net_11683;
wire net_6033;
wire net_14941;
wire net_5455;
wire net_11624;
wire net_2666;
wire net_9276;
wire net_19810;
wire net_22560;
wire net_10929;
wire net_8402;
wire net_18715;
wire net_1239;
wire net_8663;
wire net_10246;
wire net_1463;
wire net_9743;
wire net_8793;
wire net_22058;
wire net_12257;
wire net_17825;
wire net_15833;
wire net_10081;
wire net_9266;
wire net_22338;
wire net_17325;
wire net_3822;
wire net_21766;
wire net_15139;
wire net_65;
wire net_17015;
wire net_16054;
wire net_6872;
wire net_484;
wire net_896;
wire net_18156;
wire net_7655;
wire net_3223;
wire net_21873;
wire x839;
wire net_5894;
wire net_11363;
wire net_20068;
wire net_11599;
wire net_16960;
wire net_20001;
wire net_15135;
wire net_10088;
wire net_9795;
wire net_18547;
wire net_12971;
wire net_13106;
wire net_22226;
wire net_11563;
wire net_20495;
wire net_11794;
wire net_13939;
wire net_15031;
wire net_7917;
wire net_11550;
wire net_13614;
wire net_1896;
wire net_1982;
wire net_14577;
wire net_13283;
wire net_12687;
wire net_16604;
wire net_16330;
wire net_8089;
wire net_12084;
wire net_10014;
wire net_15960;
wire net_20976;
wire net_11719;
wire net_6509;
wire net_12507;
wire net_3253;
wire net_10630;
wire net_20392;
wire net_6935;
wire net_20904;
wire net_5498;
wire net_13176;
wire net_1882;
wire net_12347;
wire net_12229;
wire net_12755;
wire net_7744;
wire net_21432;
wire net_16967;
wire net_413;
wire net_11072;
wire net_9613;
wire net_18540;
wire net_6141;
wire net_14982;
wire net_12666;
wire x1354;
wire net_2419;
wire net_7876;
wire net_10154;
wire net_22414;
wire net_5753;
wire net_14898;
wire net_7608;
wire net_12203;
wire net_14315;
wire net_18334;
wire net_19444;
wire net_253;
wire net_276;
wire net_11696;
wire net_9728;
wire net_14229;
wire net_17453;
wire net_8470;
wire net_12112;
wire net_13899;
wire net_15800;
wire net_6490;
wire net_10586;
wire net_16347;
wire net_9799;
wire net_13395;
wire net_20935;
wire net_22350;
wire net_616;
wire net_28;
wire net_17977;
wire net_18086;
wire net_1847;
wire net_18772;
wire net_17474;
wire net_17270;
wire net_15899;
wire net_2717;
wire net_20665;
wire net_793;
wire net_9137;
wire net_19220;
wire net_2353;
wire net_21364;
wire net_2272;
wire net_11919;
wire net_9231;
wire net_21604;
wire net_20381;
wire net_16934;
wire net_9708;
wire net_4104;
wire net_19815;
wire net_3287;
wire net_8133;
wire net_14922;
wire net_11305;
wire net_16465;
wire net_2866;
wire net_5866;
wire net_17787;
wire net_18651;
wire net_3025;
wire net_5407;
wire net_17568;
wire net_7673;
wire net_7309;
wire net_74;
wire net_6071;
wire net_10342;
wire net_17131;
wire net_6894;
wire net_205;
wire net_1286;
wire net_11702;
wire net_6427;
wire net_15204;
wire net_20721;
wire net_9764;
wire net_11872;
wire net_15290;
wire net_22298;
wire net_19475;
wire net_17780;
wire net_7617;
wire net_18955;
wire net_7533;
wire net_1952;
wire net_18497;
wire net_9214;
wire net_9846;
wire net_11495;
wire net_22317;
wire net_12512;
wire net_4620;
wire net_380;
wire net_5696;
wire net_14141;
wire net_2847;
wire net_6515;
wire net_7932;
wire net_1556;
wire net_12885;
wire net_5911;
wire net_6803;
wire x2219;
wire net_4337;
wire net_13548;
wire net_7976;
wire net_16292;
wire net_4745;
wire net_1270;
wire net_17610;
wire net_16657;
wire net_4905;
wire net_15345;
wire net_18613;
wire net_9717;
wire net_14178;
wire net_22290;
wire net_20021;
wire net_6094;
wire net_14454;
wire net_18375;
wire net_7712;
wire net_17043;
wire net_3878;
wire net_4940;
wire net_19109;
wire net_20981;
wire net_8132;
wire net_5585;
wire net_3241;
wire net_7273;
wire net_17748;
wire net_2555;
wire net_4864;
wire net_3504;
wire net_18490;
wire net_1687;
wire net_16857;
wire net_1762;
wire net_5243;
wire net_7407;
wire net_18910;
wire net_1181;
wire net_10685;
wire net_12299;
wire net_313;
wire net_932;
wire net_7472;
wire net_21241;
wire net_20734;
wire net_15577;
wire net_6082;
wire net_16446;
wire net_10783;
wire net_13403;
wire net_12488;
wire net_4767;
wire net_5271;
wire net_14257;
wire net_6771;
wire net_12814;
wire net_19746;
wire net_972;
wire net_7769;
wire net_20369;
wire net_21118;
wire net_17526;
wire net_9650;
wire net_15043;
wire net_20900;
wire net_4725;
wire net_15942;
wire net_6201;
wire net_11669;
wire net_14292;
wire net_22787;
wire net_7047;
wire net_1489;
wire net_13665;
wire net_15789;
wire net_4343;
wire net_10276;
wire net_19380;
wire net_20397;
wire net_16282;
wire net_22157;
wire net_7794;
wire net_2392;
wire net_7194;
wire net_17515;
wire net_10278;
wire net_8441;
wire x7088;
wire net_21852;
wire net_13064;
wire net_10266;
wire net_21449;
wire net_21547;
wire net_1040;
wire net_5947;
wire net_8978;
wire net_6781;
wire net_3089;
wire net_19684;
wire net_3037;
wire net_4472;
wire net_4463;
wire net_7331;
wire net_18115;
wire net_22666;
wire net_19759;
wire net_3686;
wire net_2907;
wire net_22567;
wire net_15607;
wire net_2243;
wire net_379;
wire x2186;
wire net_1569;
wire net_21086;
wire net_16951;
wire net_22372;
wire net_3133;
wire net_7795;
wire net_2559;
wire net_18614;
wire net_19527;
wire net_14451;
wire net_19114;
wire net_14475;
wire net_1358;
wire net_8477;
wire net_6815;
wire net_14708;
wire net_11405;
wire net_6888;
wire net_8927;
wire net_8421;
wire net_16409;
wire net_20440;
wire net_960;
wire net_3704;
wire x876;
wire net_20264;
wire net_17352;
wire net_8155;
wire net_10706;
wire net_22060;
wire net_14957;
wire net_11051;
wire net_14062;
wire net_16468;
wire net_12842;
wire net_13365;
wire net_9445;
wire net_13996;
wire net_6441;
wire net_22699;
wire net_4348;
wire net_4526;
wire net_7832;
wire net_22480;
wire net_581;
wire net_8991;
wire net_9909;
wire net_10564;
wire net_13967;
wire net_2899;
wire net_8799;
wire net_17881;
wire net_9609;
wire net_12421;
wire net_658;
wire net_18554;
wire x424;
wire net_7978;
wire net_14565;
wire net_13529;
wire net_2090;
wire net_18294;
wire net_16508;
wire net_7723;
wire net_9540;
wire net_12509;
wire net_18239;
wire net_19352;
wire net_12758;
wire net_10259;
wire net_5801;
wire net_21692;
wire net_7026;
wire net_8999;
wire net_15270;
wire net_5461;
wire net_1176;
wire net_2676;
wire net_14853;
wire net_6372;
wire net_19892;
wire net_4989;
wire net_7032;
wire net_11609;
wire net_15949;
wire net_1751;
wire net_13593;
wire net_6733;
wire net_16216;
wire net_3508;
wire net_21484;
wire net_16401;
wire net_2434;
wire net_2032;
wire net_118;
wire net_17843;
wire net_2467;
wire net_17741;
wire net_11524;
wire net_14499;
wire net_21407;
wire net_14415;
wire net_9916;
wire net_12008;
wire net_17496;
wire x288;
wire x4345;
wire net_7223;
wire net_8865;
wire net_17871;
wire net_18640;
wire net_246;
wire net_6613;
wire net_20348;
wire net_20570;
wire net_21113;
wire net_11269;
wire net_13041;
wire net_10121;
wire net_13436;
wire net_14914;
wire net_16140;
wire net_17347;
wire net_6725;
wire net_8968;
wire net_1378;
wire net_1600;
wire net_2531;
wire net_16339;
wire net_12440;
wire net_17720;
wire net_11971;
wire net_15743;
wire net_676;
wire net_11254;
wire net_12492;
wire net_6626;
wire net_4263;
wire net_15592;
wire net_2538;
wire net_17710;
wire net_20449;
wire net_5133;
wire net_21179;
wire net_5542;
wire net_20579;
wire net_5370;
wire net_4260;
wire net_3492;
wire net_2462;
wire net_6010;
wire net_12760;
wire net_9018;
wire net_9635;
wire net_8820;
wire net_3324;
wire net_13485;
wire net_18166;
wire net_16773;
wire x4172;
wire net_5426;
wire net_6450;
wire net_6138;
wire net_6979;
wire net_8398;
wire net_7893;
wire net_21763;
wire net_21586;
wire net_9600;
wire net_14463;
wire net_8112;
wire net_10429;
wire net_7939;
wire net_11274;
wire net_3207;
wire net_7810;
wire net_13920;
wire net_19609;
wire net_2204;
wire net_9668;
wire net_5088;
wire net_2492;
wire net_15485;
wire net_19121;
wire net_9088;
wire net_11188;
wire net_16871;
wire net_16727;
wire net_4045;
wire net_21263;
wire net_3843;
wire net_15228;
wire net_10223;
wire net_16048;
wire x1032;
wire net_19718;
wire net_6543;
wire net_7635;
wire net_19928;
wire net_11005;
wire net_3038;
wire net_2690;
wire net_13560;
wire net_3924;
wire net_7016;
wire net_9825;
wire net_5226;
wire net_10230;
wire net_22470;
wire net_8811;
wire net_1051;
wire net_10546;
wire net_18984;
wire net_10048;
wire net_10386;
wire x4734;
wire net_20643;
wire net_22162;
wire net_22779;
wire net_14770;
wire net_20783;
wire net_7644;
wire net_20793;
wire net_7858;
wire net_11034;
wire net_1515;
wire net_1573;
wire net_7669;
wire net_10356;
wire net_18844;
wire net_4983;
wire net_6869;
wire net_22382;
wire net_13932;
wire net_9984;
wire net_305;
wire net_7100;
wire net_4208;
wire net_4515;
wire net_12433;
wire net_12016;
wire net_15434;
wire net_12452;
wire net_9166;
wire net_16833;
wire net_1125;
wire net_14716;
wire net_18872;
wire net_10195;
wire net_15084;
wire net_10667;
wire net_17236;
wire net_17686;
wire net_12405;
wire net_6687;
wire net_8818;
wire net_15555;
wire net_19102;
wire net_13592;
wire net_20444;
wire net_19885;
wire net_17254;
wire net_18356;
wire x1623;
wire net_9175;
wire net_3485;
wire net_17483;
wire net_16168;
wire net_2886;
wire net_14408;
wire net_1921;
wire net_20468;
wire net_10945;
wire net_3853;
wire net_16472;
wire net_9962;
wire net_14781;
wire net_15462;
wire net_2135;
wire net_9091;
wire net_667;
wire net_18413;
wire net_853;
wire net_22074;
wire net_212;
wire net_12265;
wire net_914;
wire net_9508;
wire net_10254;
wire net_9923;
wire net_12835;
wire net_6320;
wire net_15245;
wire net_6448;
wire net_22766;
wire net_875;
wire net_17942;
wire net_5619;
wire net_14807;
wire net_22715;
wire net_21334;
wire net_1092;
wire net_627;
wire net_18937;
wire net_18570;
wire net_8759;
wire net_16115;
wire net_19618;
wire net_15313;
wire net_18388;
wire net_17358;
wire net_15989;
wire net_11042;
wire net_15444;
wire net_19173;
wire net_20133;
wire net_5636;
wire net_15469;
wire net_2473;
wire net_12231;
wire net_21925;
wire net_19284;
wire net_16034;
wire net_399;
wire net_8107;
wire net_15284;
wire net_5949;
wire net_5069;
wire net_19603;
wire net_1390;
wire net_10678;
wire net_5565;
wire net_7180;
wire net_16805;
wire net_10517;
wire net_19363;
wire net_1112;
wire net_10747;
wire net_21885;
wire net_15483;
wire net_5449;
wire net_8146;
wire net_19863;
wire net_11200;
wire net_12085;
wire net_18191;
wire net_3230;
wire net_13295;
wire net_14494;
wire net_10187;
wire net_8316;
wire net_13585;
wire net_14932;
wire net_5677;
wire net_11486;
wire net_17154;
wire net_5296;
wire net_1310;
wire net_14171;
wire net_9634;
wire net_6057;
wire net_15687;
wire net_18674;
wire net_1304;
wire net_7579;
wire net_4381;
wire net_9471;
wire net_6674;
wire net_11378;
wire net_11918;
wire net_7863;
wire net_13427;
wire net_11450;
wire net_11587;
wire net_10370;
wire net_6127;
wire net_21840;
wire net_6058;
wire net_13417;
wire net_10919;
wire net_6070;
wire net_2449;
wire net_17105;
wire net_6588;
wire net_416;
wire net_19890;
wire net_15986;
wire net_5629;
wire net_20867;
wire net_16326;
wire net_6896;
wire net_15851;
wire net_6642;
wire net_14814;
wire net_10760;
wire net_1786;
wire net_1377;
wire net_5620;
wire net_16239;
wire net_10253;
wire net_12031;
wire net_4513;
wire x3346;
wire net_10940;
wire net_14025;
wire net_5965;
wire net_14439;
wire net_5586;
wire net_11118;
wire net_13428;
wire net_5430;
wire net_17903;
wire net_1393;
wire net_20459;
wire net_13724;
wire net_17994;
wire net_2169;
wire net_22032;
wire net_1324;
wire net_8758;
wire net_7114;
wire net_12058;
wire net_8017;
wire net_6997;
wire net_4323;
wire net_9336;
wire net_3527;
wire net_1138;
wire net_8805;
wire net_17598;
wire net_10167;
wire net_20242;
wire net_18621;
wire net_3292;
wire net_1439;
wire net_8714;
wire net_13489;
wire net_1778;
wire net_508;
wire net_9700;
wire net_15428;
wire net_6907;
wire net_5098;
wire net_19931;
wire net_7438;
wire net_15617;
wire net_5355;
wire net_8149;
wire net_11453;
wire net_11962;
wire net_5413;
wire net_4434;
wire net_18128;
wire net_12068;
wire net_16197;
wire net_4744;
wire net_18178;
wire net_6636;
wire net_2896;
wire net_14707;
wire net_4258;
wire net_8371;
wire net_7443;
wire net_12838;
wire net_12454;
wire net_9985;
wire net_13833;
wire net_7301;
wire net_1555;
wire net_10594;
wire net_21732;
wire net_9349;
wire net_4480;
wire x323;
wire net_10131;
wire net_15454;
wire net_21783;
wire net_15153;
wire net_2171;
wire net_10233;
wire net_6338;
wire net_19328;
wire net_18025;
wire net_4521;
wire net_6112;
wire net_2425;
wire net_11245;
wire net_22045;
wire x2881;
wire net_13691;
wire net_18209;
wire net_8319;
wire net_19071;
wire net_10573;
wire net_2509;
wire net_22404;
wire net_17075;
wire net_2156;
wire net_9177;
wire net_14188;
wire net_8488;
wire net_6831;
wire net_13246;
wire net_4314;
wire net_20476;
wire net_11640;
wire net_19083;
wire net_10005;
wire net_20022;
wire net_3343;
wire net_18188;
wire net_3326;
wire net_11877;
wire net_2239;
wire net_16838;
wire net_3394;
wire net_12846;
wire net_17026;
wire net_4680;
wire net_18595;
wire net_3903;
wire net_15192;
wire net_22748;
wire net_8879;
wire net_4050;
wire net_16818;
wire net_1571;
wire net_16155;
wire net_11467;
wire net_9248;
wire net_18887;
wire net_5090;
wire net_10530;
wire net_850;
wire net_22454;
wire net_12511;
wire net_21476;
wire net_1168;
wire net_21459;
wire net_10118;
wire net_11008;
wire net_5545;
wire net_9631;
wire net_21792;
wire net_17685;
wire net_10744;
wire net_3090;
wire net_8747;
wire net_15052;
wire net_8387;
wire net_1009;
wire net_21077;
wire net_715;
wire net_11444;
wire net_18502;
wire net_13857;
wire net_14503;
wire net_16475;
wire net_8454;
wire net_16152;
wire net_2546;
wire net_11181;
wire net_7056;
wire net_12042;
wire net_19388;
wire net_15876;
wire net_16810;
wire net_6702;
wire net_20831;
wire net_312;
wire net_11130;
wire net_2627;
wire net_5386;
wire net_147;
wire net_21131;
wire net_17237;
wire net_7182;
wire net_12490;
wire net_16453;
wire net_8589;
wire net_12137;
wire net_7750;
wire net_12335;
wire net_2444;
wire net_17454;
wire net_13496;
wire net_21237;
wire net_5297;
wire net_8148;
wire net_12936;
wire net_9625;
wire net_17753;
wire net_10122;
wire net_20776;
wire net_14965;
wire net_8551;
wire net_19137;
wire net_10759;
wire net_14148;
wire net_7431;
wire net_5398;
wire net_21040;
wire net_18200;
wire net_2435;
wire net_245;
wire net_20321;
wire net_6990;
wire net_4858;
wire net_2383;
wire net_12177;
wire net_3491;
wire net_11013;
wire net_16296;
wire net_10829;
wire net_8380;
wire net_277;
wire net_16795;
wire net_4251;
wire net_1965;
wire net_21740;
wire net_89;
wire net_13886;
wire net_680;
wire net_16537;
wire net_17585;
wire net_338;
wire net_13230;
wire net_13435;
wire net_4494;
wire net_20006;
wire net_8397;
wire net_15672;
wire net_14597;
wire net_19410;
wire net_9971;
wire net_22061;
wire net_4089;
wire net_10705;
wire net_13721;
wire net_22008;
wire net_2009;
wire net_18134;
wire net_17604;
wire net_19945;
wire net_4026;
wire net_6697;
wire net_20879;
wire net_106;
wire net_1380;
wire net_14844;
wire net_22581;
wire net_14731;
wire net_20633;
wire net_22522;
wire net_9340;
wire net_21936;
wire net_5176;
wire net_20870;
wire net_5936;
wire net_18890;
wire net_11956;
wire net_19419;
wire net_8937;
wire net_6987;
wire net_18469;
wire net_14550;
wire net_1997;
wire x2127;
wire net_13206;
wire net_138;
wire net_14657;
wire net_20401;
wire net_19169;
wire net_15931;
wire net_21401;
wire net_7718;
wire net_8553;
wire net_6728;
wire net_13364;
wire net_13698;
wire net_11139;
wire net_18897;
wire net_14151;
wire net_6579;
wire net_15232;
wire net_19160;
wire net_14792;
wire net_1418;
wire net_8686;
wire net_13955;
wire net_5938;
wire net_21045;
wire net_19353;
wire net_6980;
wire net_5931;
wire net_8343;
wire net_22131;
wire net_15226;
wire net_20740;
wire net_1713;
wire net_12913;
wire net_4684;
wire net_11383;
wire net_8988;
wire net_2775;
wire net_7001;
wire net_14594;
wire net_12007;
wire net_17919;
wire net_14839;
wire net_7654;
wire net_163;
wire net_6022;
wire net_19799;
wire net_5802;
wire net_21029;
wire net_19542;
wire net_15736;
wire net_11037;
wire net_8037;
wire net_15843;
wire net_22622;
wire net_19046;
wire net_8444;
wire net_9830;
wire net_18169;
wire net_6135;
wire net_11580;
wire net_13863;
wire net_2193;
wire net_12595;
wire net_21341;
wire net_12002;
wire net_12293;
wire net_11159;
wire net_20709;
wire net_22696;
wire net_18102;
wire net_6304;
wire net_5574;
wire net_11704;
wire net_5258;
wire net_17133;
wire net_1886;
wire net_2604;
wire net_13689;
wire net_12191;
wire net_14115;
wire net_4678;
wire net_18593;
wire net_14307;
wire net_14256;
wire net_4866;
wire net_5652;
wire net_16256;
wire net_101;
wire net_2109;
wire net_1770;
wire net_21612;
wire net_9326;
wire net_4703;
wire net_20076;
wire net_22781;
wire net_21993;
wire net_17302;
wire net_22536;
wire net_14530;
wire net_19217;
wire net_4770;
wire net_7770;
wire net_378;
wire x6655;
wire net_14049;
wire net_14262;
wire net_3309;
wire net_20823;
wire net_5767;
wire net_20546;
wire net_16972;
wire net_10032;
wire net_18377;
wire net_4202;
wire net_11628;
wire net_18535;
wire net_1958;
wire net_21784;
wire net_1931;
wire net_15493;
wire net_14041;
wire net_1549;
wire net_6244;
wire net_10039;
wire net_16883;
wire net_7736;
wire net_2929;
wire net_20922;
wire net_7192;
wire net_20840;
wire net_16608;
wire net_7213;
wire net_5666;
wire x6043;
wire net_8527;
wire net_11227;
wire net_22411;
wire net_818;
wire net_15103;
wire x2139;
wire net_11275;
wire net_16855;
wire net_1211;
wire net_5448;
wire net_1183;
wire net_4248;
wire net_22191;
wire net_21817;
wire net_14537;
wire net_12337;
wire net_17979;
wire net_7241;
wire net_21417;
wire net_16035;
wire net_17190;
wire net_9753;
wire net_4674;
wire net_9203;
wire net_9551;
wire net_15495;
wire net_6791;
wire net_2017;
wire net_5154;
wire net_11508;
wire net_16138;
wire net_2735;
wire net_12145;
wire net_21947;
wire net_8780;
wire net_8377;
wire net_20072;
wire net_16466;
wire net_8800;
wire net_18747;
wire net_1621;
wire net_14432;
wire net_16661;
wire net_18247;
wire net_19524;
wire net_1035;
wire net_12253;
wire net_21924;
wire net_11331;
wire net_20368;
wire net_14076;
wire net_21884;
wire net_17509;
wire net_20550;
wire net_20413;
wire net_13035;
wire net_20882;
wire net_5597;
wire net_20027;
wire net_6914;
wire net_4656;
wire net_20817;
wire net_3593;
wire net_10264;
wire net_22039;
wire net_6748;
wire net_2641;
wire net_19462;
wire net_16584;
wire net_7711;
wire net_18972;
wire net_6688;
wire net_20342;
wire net_9389;
wire net_4035;
wire net_12321;
wire net_18058;
wire net_7816;
wire net_9362;
wire net_9881;
wire net_17697;
wire net_8948;
wire net_9092;
wire net_13464;
wire net_7919;
wire net_2882;
wire net_8131;
wire net_14440;
wire net_22253;
wire net_19736;
wire net_14191;
wire net_18785;
wire net_14253;
wire net_3064;
wire net_5731;
wire net_2276;
wire net_6369;
wire net_12748;
wire net_9302;
wire net_11639;
wire net_7748;
wire net_22591;
wire net_9426;
wire net_6745;
wire net_21203;
wire net_13716;
wire net_798;
wire net_14149;
wire net_14820;
wire net_18612;
wire net_16002;
wire net_2059;
wire net_18911;
wire net_15806;
wire net_15993;
wire net_19976;
wire net_9740;
wire net_8520;
wire net_6018;
wire net_8860;
wire net_21514;
wire x2767;
wire net_16074;
wire net_1336;
wire net_18905;
wire net_9915;
wire net_10033;
wire net_61;
wire net_6946;
wire net_11739;
wire net_19803;
wire net_14114;
wire net_20559;
wire net_11534;
wire net_11671;
wire net_3336;
wire net_903;
wire net_9561;
wire net_15502;
wire net_10025;
wire net_21919;
wire net_12069;
wire net_21274;
wire net_13796;
wire net_7354;
wire net_8407;
wire net_11395;
wire net_18387;
wire net_5986;
wire net_2378;
wire net_22276;
wire net_16896;
wire net_17290;
wire net_6261;
wire net_10461;
wire net_11758;
wire net_20533;
wire net_10319;
wire net_8046;
wire net_17974;
wire net_18238;
wire net_13746;
wire net_15378;
wire net_7125;
wire net_21874;
wire net_20388;
wire net_16393;
wire net_8605;
wire net_9865;
wire net_95;
wire net_10010;
wire net_14445;
wire net_5566;
wire net_5281;
wire net_8776;
wire net_19568;
wire net_2327;
wire net_1003;
wire net_8772;
wire net_10868;
wire net_17559;
wire net_15443;
wire net_17552;
wire net_7376;
wire net_11255;
wire net_10310;
wire net_14093;
wire net_19510;
wire net_5669;
wire net_6122;
wire net_6497;
wire net_6060;
wire net_11991;
wire net_13387;
wire net_22741;
wire net_16287;
wire net_22516;
wire net_11513;
wire net_13554;
wire net_3742;
wire net_21349;
wire net_445;
wire net_13398;
wire net_20084;
wire net_19555;
wire net_10773;
wire net_6673;
wire net_12319;
wire net_13637;
wire net_22608;
wire net_17828;
wire net_18583;
wire net_2213;
wire net_8307;
wire net_2575;
wire net_11986;
wire net_15880;
wire net_9219;
wire net_21836;
wire net_19006;
wire net_12142;
wire net_6921;
wire net_17099;
wire net_8445;
wire net_13517;
wire net_3713;
wire net_10876;
wire net_556;
wire net_21248;
wire net_19673;
wire net_18311;
wire net_4121;
wire net_3826;
wire net_620;
wire net_18157;
wire net_16096;
wire net_8702;
wire net_4659;
wire net_7321;
wire net_22086;
wire net_14529;
wire net_5997;
wire net_4779;
wire net_14392;
wire net_16954;
wire net_11150;
wire net_8156;
wire net_5129;
wire net_20638;
wire net_10444;
wire net_7883;
wire net_17471;
wire net_6414;
wire net_19262;
wire net_5393;
wire net_20233;
wire net_17327;
wire net_20816;
wire net_22328;
wire net_6937;
wire net_7825;
wire net_13613;
wire net_8855;
wire net_1493;
wire net_17407;
wire net_9167;
wire net_17459;
wire net_11143;
wire net_19728;
wire net_8498;
wire net_8897;
wire net_4179;
wire net_2579;
wire net_19074;
wire net_21038;
wire net_8235;
wire net_9581;
wire net_6013;
wire net_10296;
wire net_7307;
wire net_5873;
wire net_1866;
wire net_12990;
wire net_19294;
wire net_14852;
wire net_6934;
wire net_5761;
wire net_3211;
wire net_16552;
wire net_10820;
wire net_13060;
wire net_16798;
wire net_21869;
wire net_7634;
wire net_5927;
wire net_13894;
wire net_37;
wire net_11738;
wire x5015;
wire net_12754;
wire net_19259;
wire net_8625;
wire net_16680;
wire net_8342;
wire net_11732;
wire net_2516;
wire net_18480;
wire net_7553;
wire net_2807;
wire net_4687;
wire net_10676;
wire net_15908;
wire net_18694;
wire net_16655;
wire net_18342;
wire net_6321;
wire net_7584;
wire net_22233;
wire net_1288;
wire net_16382;
wire net_4708;
wire net_10511;
wire net_12554;
wire net_20616;
wire net_10559;
wire net_2300;
wire net_8119;
wire net_6710;
wire net_8426;
wire net_7091;
wire net_6383;
wire net_13915;
wire net_6434;
wire net_4816;
wire net_11428;
wire net_11604;
wire net_21684;
wire net_17760;
wire net_21628;
wire net_17058;
wire net_5524;
wire net_16381;
wire net_4937;
wire net_4199;
wire net_1043;
wire net_11897;
wire net_16543;
wire net_15086;
wire net_18764;
wire net_18846;
wire net_9737;
wire net_6389;
wire net_16806;
wire net_7493;
wire net_1630;
wire net_22213;
wire net_2956;
wire net_18094;
wire net_1082;
wire net_11170;
wire net_15645;
wire net_10405;
wire net_16516;
wire net_16365;
wire net_15407;
wire net_18282;
wire net_11861;
wire net_3296;
wire net_257;
wire net_8543;
wire net_10096;
wire net_11407;
wire net_5500;
wire net_9978;
wire net_19177;
wire net_5770;
wire net_18682;
wire net_6576;
wire net_958;
wire net_12646;
wire net_4556;
wire net_6400;
wire net_11447;
wire net_12407;
wire net_6199;
wire net_22624;
wire net_1734;
wire net_10189;
wire net_17205;
wire net_11175;
wire net_5534;
wire net_4308;
wire net_22040;
wire net_10987;
wire net_17927;
wire net_17041;
wire net_16424;
wire net_7166;
wire net_13450;
wire net_14510;
wire net_19773;
wire net_3050;
wire net_1728;
wire net_20301;
wire net_5963;
wire net_12883;
wire net_15394;
wire net_20091;
wire net_3956;
wire net_16441;
wire net_12426;
wire net_10218;
wire net_8467;
wire net_8761;
wire net_22641;
wire net_425;
wire net_17818;
wire net_5204;
wire net_17417;
wire net_22603;
wire net_22108;
wire net_2205;
wire net_20739;
wire net_13154;
wire net_19061;
wire net_16123;
wire net_8108;
wire net_20131;
wire net_11344;
wire net_17621;
wire net_16087;
wire net_13667;
wire net_368;
wire net_8064;
wire net_19950;
wire net_4833;
wire net_52;
wire net_15914;
wire net_20153;
wire net_10670;
wire net_2000;
wire net_13089;
wire net_19765;
wire net_6226;
wire net_14799;
wire net_12502;
wire net_18313;
wire net_2984;
wire net_1020;
wire net_10603;
wire net_21581;
wire net_15971;
wire net_18366;
wire net_3282;
wire net_3122;
wire net_13989;
wire net_17860;
wire net_8546;
wire net_20428;
wire net_10164;
wire net_10763;
wire net_16990;
wire net_8594;
wire net_12521;
wire net_18562;
wire net_19623;
wire net_2094;
wire net_11965;
wire net_7282;
wire net_2543;
wire net_8275;
wire net_760;
wire net_2083;
wire net_19330;
wire net_8318;
wire net_12050;
wire net_19581;
wire net_17223;
wire net_3851;
wire net_2488;
wire net_4536;
wire net_5034;
wire net_21850;
wire net_8192;
wire net_17767;
wire net_1870;
wire net_5200;
wire net_12772;
wire net_2063;
wire net_192;
wire net_17922;
wire net_1739;
wire net_2912;
wire net_4140;
wire net_22714;
wire net_18293;
wire net_13254;
wire net_735;
wire net_20171;
wire net_14269;
wire net_22258;
wire net_17060;
wire net_3809;
wire net_16824;
wire net_19665;
wire net_9442;
wire net_21713;
wire net_21577;
wire net_1081;
wire net_17636;
wire net_19238;
wire net_2037;
wire net_8163;
wire net_1237;
wire net_1420;
wire net_12478;
wire net_4789;
wire net_9112;
wire net_14921;
wire net_4064;
wire net_9587;
wire net_4237;
wire net_9712;
wire net_9542;
wire net_17486;
wire net_4559;
wire net_18265;
wire net_7782;
wire net_3144;
wire net_699;
wire net_359;
wire net_19271;
wire net_5239;
wire net_16940;
wire net_16065;
wire net_9068;
wire net_12862;
wire net_5827;
wire net_2819;
wire net_11316;
wire net_15901;
wire net_882;
wire net_15614;
wire net_6433;
wire net_1827;
wire net_14867;
wire net_4109;
wire net_12606;
wire net_15958;
wire net_8903;
wire net_3858;
wire net_19997;
wire net_7838;
wire net_10813;
wire net_14182;
wire net_21685;
wire net_16626;
wire net_15254;
wire net_2283;
wire net_1207;
wire net_20205;
wire net_10436;
wire net_2121;
wire net_8228;
wire net_14326;
wire net_20770;
wire net_14671;
wire net_2252;
wire net_4755;
wire net_18733;
wire net_20497;
wire net_7951;
wire net_17394;
wire net_2126;
wire x1747;
wire net_5022;
wire net_9931;
wire net_10449;
wire net_7342;
wire net_16947;
wire net_17657;
wire net_9524;
wire net_12461;
wire net_20193;
wire net_19549;
wire net_17398;
wire net_14616;
wire net_18944;
wire net_6952;
wire net_3655;
wire net_17432;
wire x4603;
wire net_2304;
wire net_14098;
wire net_12942;
wire net_7418;
wire net_19305;
wire net_1593;
wire net_8918;
wire net_3380;
wire net_10397;
wire net_19959;
wire net_16177;
wire net_15272;
wire net_20995;
wire net_18511;
wire net_12794;
wire net_14758;
wire net_11762;
wire net_5115;
wire net_14682;
wire net_4502;
wire x480;
wire net_15658;
wire x615;
wire net_16844;
wire net_12275;
wire net_2076;
wire net_12567;
wire net_13131;
wire net_6505;
wire net_4378;
wire net_2218;
wire net_19269;
wire net_6807;
wire net_10147;
wire net_21181;
wire net_15219;
wire net_20957;
wire net_1078;
wire net_9811;
wire net_12340;
wire net_9853;
wire net_6813;
wire net_14984;
wire net_6382;
wire net_14896;
wire net_5681;
wire net_13126;
wire net_10635;
wire net_18930;
wire net_14341;
wire net_12269;
wire net_5197;
wire net_12703;
wire net_13059;
wire net_2355;
wire net_12856;
wire net_13825;
wire net_3262;
wire net_139;
wire net_19845;
wire net_22827;
wire net_22118;
wire net_20894;
wire net_4495;
wire net_12587;
wire net_16438;
wire net_12824;
wire net_7454;
wire net_16379;
wire net_4196;
wire net_3974;
wire net_13678;
wire net_4626;
wire net_20143;
wire net_8532;
wire net_19453;
wire net_8478;
wire net_19337;
wire net_2976;
wire net_15007;
wire net_13138;
wire net_988;
wire net_8221;
wire net_21188;
wire net_3621;
wire net_20202;
wire net_19183;
wire net_9820;
wire net_12441;
wire net_22687;
wire net_18917;
wire net_4091;
wire net_17448;
wire net_132;
wire net_12110;
wire net_18714;
wire net_2838;
wire net_21177;
wire net_5614;
wire net_5219;
wire net_1841;
wire net_20053;
wire net_1249;
wire net_22633;
wire net_17799;
wire net_4601;
wire net_22375;
wire net_21156;
wire net_18791;
wire net_7973;
wire x2835;
wire net_22363;
wire net_3163;
wire net_4928;
wire net_18479;
wire net_6221;
wire net_21642;
wire net_4417;
wire net_7145;
wire net_822;
wire net_7084;
wire net_20014;
wire net_15369;
wire net_21283;
wire net_15523;
wire net_17985;
wire net_21389;
wire net_6561;
wire net_21057;
wire net_16749;
wire net_13470;
wire net_6842;
wire net_15691;
wire net_7701;
wire net_1974;
wire net_8010;
wire net_4963;
wire net_9996;
wire net_11480;
wire net_9021;
wire net_22222;
wire net_1544;
wire net_22706;
wire net_15798;
wire net_7366;
wire net_20482;
wire net_4400;
wire net_10044;
wire net_18362;
wire net_15572;
wire net_22691;
wire net_10340;
wire net_17645;
wire net_7929;
wire net_1174;
wire net_15168;
wire net_6731;
wire net_6664;
wire net_1109;
wire net_12326;
wire net_4224;
wire net_13733;
wire net_22343;
wire net_20690;
wire net_3457;
wire net_9683;
wire net_10963;
wire net_21539;
wire net_5276;
wire net_11721;
wire net_4471;
wire net_1102;
wire net_16861;
wire net_5487;
wire net_13644;
wire net_4976;
wire net_5640;
wire net_5245;
wire net_18928;
wire net_18002;
wire net_11205;
wire net_18622;
wire net_14175;
wire net_2692;
wire x368;
wire net_3777;
wire net_11322;
wire net_19254;
wire net_18144;
wire net_14355;
wire net_13353;
wire net_10285;
wire net_6279;
wire net_14382;
wire net_15934;
wire net_7516;
wire x462;
wire net_7037;
wire net_1487;
wire net_4572;
wire net_2759;
wire net_10020;
wire net_19651;
wire net_5408;
wire net_8243;
wire net_3634;
wire net_12486;
wire net_14128;
wire net_13348;
wire net_16570;
wire x7467;
wire net_16117;
wire net_18533;
wire net_13705;
wire net_14215;
wire net_22121;
wire net_10338;
wire net_21557;
wire net_21200;
wire net_18650;
wire net_10349;
wire net_2564;
wire net_2821;
wire net_1658;
wire net_5688;
wire net_5481;
wire net_17891;
wire net_7318;
wire net_21313;
wire net_17823;
wire net_3007;
wire net_7554;
wire net_9505;
wire net_4487;
wire net_15412;
wire net_14998;
wire net_3174;
wire net_9122;
wire net_6966;
wire net_2876;
wire net_844;
wire net_1496;
wire net_325;
wire net_14470;
wire net_1820;
wire net_21896;
wire x1021;
wire net_8175;
wire net_14628;
wire net_5690;
wire net_13274;
wire net_10287;
wire net_16783;
wire net_5956;
wire net_5014;
wire net_7517;
wire net_4036;
wire net_11266;
wire x3863;
wire net_1521;
wire net_6274;
wire net_4182;
wire net_22794;
wire net_11813;
wire net_7908;
wire net_11727;
wire net_7179;
wire net_4734;
wire net_2991;
wire net_4276;
wire net_564;
wire net_10077;
wire net_14919;
wire net_19051;
wire net_6154;
wire net_10618;
wire net_22808;
wire net_2050;
wire net_4086;
wire net_9082;
wire net_13992;
wire net_21134;
wire net_813;
wire net_14105;
wire net_5609;
wire net_10661;
wire net_15279;
wire net_1027;
wire net_20433;
wire net_19629;
wire net_1408;
wire net_12403;
wire net_265;
wire net_15819;
wire net_8110;
wire net_11720;
wire net_8673;
wire net_11097;
wire net_13538;
wire net_6774;
wire net_10834;
wire net_9351;
wire net_1155;
wire net_9258;
wire net_14606;
wire net_9787;
wire net_22558;
wire net_7374;
wire net_12764;
wire net_16324;
wire net_864;
wire net_10331;
wire net_21645;
wire net_17186;
wire net_7691;
wire net_21777;
wire net_18569;
wire net_16340;
wire net_13004;
wire net_12787;
wire net_20037;
wire net_12285;
wire net_16706;
wire net_4113;
wire net_14992;
wire net_17148;
wire net_8850;
wire net_10365;
wire net_16591;
wire net_2298;
wire net_660;
wire net_14060;
wire net_19375;
wire net_9707;
wire net_21013;
wire net_21531;
wire net_6580;
wire net_1908;
wire net_7647;
wire net_9309;
wire net_22351;
wire net_3383;
wire net_18552;
wire net_13020;
wire net_7265;
wire net_12958;
wire net_21964;
wire net_6751;
wire net_20566;
wire net_19708;
wire net_3914;
wire x6912;
wire net_7607;
wire net_6531;
wire net_17084;
wire net_14104;
wire net_6463;
wire net_21967;
wire net_11973;
wire net_6455;
wire net_5777;
wire net_10610;
wire net_7576;
wire net_13449;
wire net_21598;
wire net_16595;
wire net_16916;
wire net_2145;
wire net_6488;
wire net_16529;
wire net_11109;
wire net_21270;
wire net_17101;
wire net_3311;
wire net_8874;
wire net_11020;
wire net_12729;
wire net_14036;
wire net_20808;
wire net_10887;
wire net_20722;
wire net_10454;
wire net_15310;
wire net_20561;
wire net_10716;
wire net_18346;
wire net_21940;
wire net_4853;
wire net_13943;
wire net_8699;
wire net_14775;
wire net_21061;
wire x5685;
wire net_20108;
wire x756;
wire net_10474;
wire net_13080;
wire net_3538;
wire net_11507;
wire net_22358;
wire net_17200;
wire net_22545;
wire net_20847;
wire net_17617;
wire net_21862;
wire net_22394;
wire net_1583;
wire net_15564;
wire net_9454;
wire net_4408;
wire net_19632;
wire net_1563;
wire net_3898;
wire net_4948;
wire net_13969;
wire net_7600;
wire net_16349;
wire net_5599;
wire net_13073;
wire net_3361;
wire net_10553;
wire net_13019;
wire net_8578;
wire net_14285;
wire net_15892;
wire net_21176;
wire net_18255;
wire net_21914;
wire net_1942;
wire net_11484;
wire net_10070;
wire net_12119;
wire net_13755;
wire net_20577;
wire net_7891;
wire net_18601;
wire net_1267;
wire net_14150;
wire net_6093;
wire net_3944;
wire net_3661;
wire net_11846;
wire net_12570;
wire net_9188;
wire net_4893;
wire net_18221;
wire net_12982;
wire net_6526;
wire net_5888;
wire net_5131;
wire net_19701;
wire net_2349;
wire net_18868;
wire net_22229;
wire net_11074;
wire net_1294;
wire net_10350;
wire net_14450;
wire net_14692;
wire net_3520;
wire net_5006;
wire net_18877;
wire net_1354;
wire net_15480;
wire net_2904;
wire net_1308;
wire net_7631;
wire net_18426;
wire net_4332;
wire net_12081;
wire net_15998;
wire net_1389;
wire net_9992;
wire net_12114;
wire net_19312;
wire net_13818;
wire net_4748;
wire net_19607;
wire net_3250;
wire net_5304;
wire net_10737;
wire net_17723;
wire net_548;
wire net_16931;
wire net_4985;
wire net_2402;
wire net_6529;
wire net_5902;
wire net_5082;
wire net_636;
wire net_10239;
wire net_4269;
wire net_18803;
wire net_8159;
wire net_18494;
wire net_8218;
wire net_8471;
wire net_17947;
wire net_21184;
wire net_12678;
wire net_4262;
wire net_4165;
wire net_19180;
wire net_16230;
wire net_4506;
wire net_1185;
wire net_10228;
wire net_13868;
wire net_5001;
wire net_22422;
wire net_16881;
wire net_21749;
wire net_7942;
wire net_11216;
wire net_9401;
wire net_22732;
wire net_4826;
wire net_21583;
wire net_1912;
wire net_9566;
wire net_11263;
wire net_11353;
wire net_17092;
wire net_11416;
wire net_9118;
wire net_19536;
wire net_11542;
wire net_9906;
wire net_15746;
wire net_15721;
wire net_18670;
wire net_1538;
wire net_14228;
wire net_9501;
wire net_21480;
wire net_20448;
wire net_11499;
wire net_13965;
wire net_1579;
wire net_13440;
wire net_6484;
wire net_10520;
wire net_1999;
wire net_6669;
wire net_1014;
wire net_1444;
wire net_2679;
wire net_21760;
wire net_17450;
wire net_6255;
wire net_4082;
wire net_11577;
wire net_14666;
wire net_21453;
wire net_538;
wire net_9083;
wire net_14746;
wire net_14864;
wire net_4130;
wire net_12994;
wire net_9965;
wire net_13306;
wire net_366;
wire net_20393;
wire net_1854;
wire net_1917;
wire net_21635;
wire net_1755;
wire net_1359;
wire net_21821;
wire net_16113;
wire net_2460;
wire net_8929;
wire net_13228;
wire net_19194;
wire net_21351;
wire net_19135;
wire net_14704;
wire net_11238;
wire net_22340;
wire net_15547;
wire net_11348;
wire net_13424;
wire net_12618;
wire net_14496;
wire net_209;
wire net_1282;
wire net_9242;
wire net_22711;
wire net_17804;
wire net_19857;
wire net_17883;
wire net_8211;
wire net_4041;
wire net_13291;
wire net_22264;
wire net_3204;
wire net_16406;
wire net_8996;
wire net_22109;
wire net_12315;
wire net_3471;
wire net_18723;
wire net_9677;
wire net_9692;
wire net_22066;
wire net_12354;
wire net_12966;
wire net_3512;
wire net_15387;
wire net_82;
wire net_8907;
wire net_9394;
wire net_11531;
wire net_10382;
wire net_20267;
wire net_19273;
wire net_2430;
wire net_10177;
wire net_22532;
wire net_4461;
wire net_8433;
wire net_19982;
wire net_17267;
wire net_7687;
wire net_13598;
wire net_3481;
wire net_11942;
wire net_1589;
wire net_14979;
wire net_17543;
wire net_19420;
wire net_8114;
wire net_2396;
wire net_9098;
wire net_19850;
wire net_19032;
wire net_13298;
wire net_15489;
wire net_16771;
wire net_8354;
wire net_5815;
wire x733;
wire net_2856;
wire x8;
wire net_787;
wire net_7777;
wire net_10789;
wire net_19924;
wire net_8125;
wire net_3603;
wire net_9656;
wire net_16029;
wire net_19438;
wire net_4187;
wire x4642;
wire net_8095;
wire net_20713;
wire net_16491;
wire net_12071;
wire net_14323;
wire net_22566;
wire net_8463;
wire net_11001;
wire net_6195;
wire net_20714;
wire net_10767;
wire net_22034;
wire net_16146;
wire net_3579;
wire net_18575;
wire x1662;
wire net_21251;
wire net_11069;
wire net_20256;
wire net_8870;
wire net_2139;
wire net_15638;
wire net_22554;
wire net_5332;
wire net_22720;
wire net_10250;
wire net_20041;
wire net_18633;
wire net_1910;
wire net_19213;
wire net_8103;
wire net_17158;
wire net_12689;
wire net_14891;
wire net_3544;
wire net_22718;
wire net_5229;
wire net_3034;
wire net_9517;
wire net_7895;
wire net_9488;
wire net_22315;
wire net_7938;
wire net_7610;
wire net_6285;
wire net_18866;
wire net_19826;
wire net_12817;
wire net_11030;
wire net_2493;
wire net_9664;
wire net_919;
wire net_11914;
wire net_9009;
wire net_11574;
wire net_7044;
wire net_6836;
wire net_6444;
wire net_4008;
wire net_12669;
wire net_15280;
wire net_2209;
wire net_1372;
wire net_1757;
wire net_11935;
wire net_22432;
wire net_15601;
wire net_21396;
wire net_5215;
wire net_8816;
wire net_13084;
wire net_13015;
wire x2011;
wire net_14547;
wire net_2682;
wire net_19474;
wire net_7151;
wire net_14936;
wire net_8053;
wire net_17500;
wire net_140;
wire net_14562;
wire net_11949;
wire net_6612;
wire net_7077;
wire net_8911;
wire net_3790;
wire net_17313;
wire net_9141;
wire net_15235;
wire net_4267;
wire net_15275;
wire net_12482;
wire net_18394;
wire net_7328;
wire net_19429;
wire net_20374;
wire net_2178;
wire net_20276;
wire net_5292;
wire net_22053;
wire net_3073;
wire net_10134;
wire net_22738;
wire net_21676;
wire net_8840;
wire net_7949;
wire net_13846;
wire net_18420;
wire net_804;
wire net_10541;
wire net_3548;
wire net_1314;
wire net_21337;
wire net_9400;
wire net_6325;
wire net_8845;
wire net_5376;
wire net_16484;
wire net_531;
wire net_8582;
wire net_499;
wire net_2752;
wire net_9126;
wire net_10701;
wire net_16165;
wire net_17792;
wire net_9476;
wire net_9699;
wire net_71;
wire net_19590;
wire net_22484;
wire net_4390;
wire net_3534;
wire net_8027;
wire net_13413;
wire net_17844;
wire net_1765;
wire net_12155;
wire net_8965;
wire net_18290;
wire net_10424;
wire net_14878;
wire net_11231;
wire net_6208;
wire net_6068;
wire net_2774;
wire net_2420;
wire net_12437;
wire net_13410;
wire net_1979;
wire net_5135;
wire net_19714;
wire net_13927;
wire net_19705;
wire net_1460;
wire net_1451;
wire net_13978;
wire net_12246;
wire net_18195;
wire net_17460;
wire net_5065;
wire net_5008;
wire net_6619;
wire net_8419;
wire net_15860;
wire net_4803;
wire net_22387;
wire net_14667;
wire net_20594;
wire net_17777;
wire net_15682;
wire net_203;
wire net_16890;
wire net_6597;
wire net_14589;
wire net_11071;
wire net_1602;
wire net_12213;
wire net_22001;
wire net_237;
wire net_613;
wire net_9919;
wire net_13239;
wire net_17561;
wire net_19811;
wire net_14236;
wire net_16070;
wire net_1095;
wire net_4729;
wire net_578;
wire net_20147;
wire net_12236;
wire net_15467;
wire net_15460;
wire net_14787;
wire net_22563;
wire net_16616;
wire net_11288;
wire net_8514;
wire net_18457;
wire net_18053;
wire net_14881;
wire net_2743;
wire net_2159;
wire net_388;
wire net_19143;
wire net_21491;
wire net_3647;
wire net_14360;
wire net_21114;
wire net_19572;
wire net_536;
wire net_1332;
wire net_17786;
wire net_18458;
wire net_3276;
wire net_10589;
wire net_393;
wire net_11980;
wire net_7468;
wire net_13525;
wire net_9130;
wire net_22155;
wire net_408;
wire net_22449;
wire net_16101;
wire net_10904;
wire net_15207;
wire net_16449;
wire net_3246;
wire net_10582;
wire net_1845;
wire net_18543;
wire net_10633;
wire net_12225;
wire net_17273;
wire net_17297;
wire net_9939;
wire net_15969;
wire net_15438;
wire net_21979;
wire x7443;
wire net_3390;
wire net_21081;
wire net_18740;
wire net_15446;
wire net_2372;
wire net_66;
wire net_12579;
wire net_12870;
wire net_868;
wire net_11223;
wire net_10979;
wire net_6079;
wire net_6821;
wire net_13750;
wire net_5029;
wire net_13871;
wire net_270;
wire net_522;
wire net_922;
wire net_20060;
wire net_2638;
wire net_17318;
wire net_9747;
wire net_13355;
wire net_19691;
wire net_5429;
wire net_15776;
wire net_4992;
wire net_6140;
wire net_5757;
wire net_2264;
wire net_977;
wire net_11632;
wire net_4780;
wire net_643;
wire net_11278;
wire net_6876;
wire net_6175;
wire net_11165;
wire net_13564;
wire net_15340;
wire net_3587;
wire net_3762;
wire net_10580;
wire net_17348;
wire net_3687;
wire net_19783;
wire net_10056;
wire net_5307;
wire net_10483;
wire net_12015;
wire net_4920;
wire net_3874;
wire net_2045;
wire net_9357;
wire net_21855;
wire net_11790;
wire net_11829;
wire net_2869;
wire net_22017;
wire net_21807;
wire net_3332;
wire net_3446;
wire net_1892;
wire net_18870;
wire net_1798;
wire net_4427;
wire net_7401;
wire net_29;
wire net_13109;
wire net_837;
wire net_13287;
wire net_3469;
wire net_10723;
wire net_9449;
wire net_20019;
wire net_927;
wire net_11686;
wire net_15838;
wire net_17375;
wire net_693;
wire net_1519;
wire net_12633;
wire net_17992;
wire net_16665;
wire net_6378;
wire net_20286;
wire net_11390;
wire net_17736;
wire net_3964;
wire net_13777;
wire net_12660;
wire net_4219;
wire net_19491;
wire net_9311;
wire net_15166;
wire net_9898;
wire net_11865;
wire x6280;
wire net_15816;
wire net_14632;
wire net_10847;
wire net_17847;
wire net_13391;
wire x1869;
wire net_10208;
wire net_11651;
wire net_488;
wire net_4909;
wire net_10460;
wire net_12009;
wire net_6034;
wire net_20908;
wire net_20123;
wire net_18287;
wire net_17170;
wire net_5452;
wire net_8088;
wire net_21410;
wire net_22324;
wire net_2319;
wire net_8324;
wire net_15717;
wire net_22751;
wire net_21608;
wire net_7102;
wire net_5458;
wire net_11785;
wire net_1532;
wire net_8440;
wire net_8971;
wire net_6653;
wire net_12308;
wire net_4475;
wire net_8207;
wire net_16981;
wire net_11595;
wire net_15478;
wire net_7765;
wire net_14639;
wire net_21800;
wire net_4958;
wire net_15215;
wire net_14719;
wire net_5057;
wire net_1093;
wire net_2592;
wire net_14947;
wire net_7680;
wire net_6230;
wire net_19755;
wire net_16343;
wire net_3580;
wire net_9876;
wire net_15505;
wire net_16641;
wire net_3259;
wire net_21008;
wire net_5260;
wire net_9877;
wire net_20246;
wire net_10057;
wire net_8833;
wire net_710;
wire net_8922;
wire net_14908;
wire net_17301;
wire net_18020;
wire net_17608;
wire net_21543;
wire net_14754;
wire net_15072;
wire net_3097;
wire net_14686;
wire net_5836;
wire net_6478;
wire net_16866;
wire net_14401;
wire net_17745;
wire net_19741;
wire net_18320;
wire net_3970;
wire net_3018;
wire net_173;
wire net_12516;
wire net_14317;
wire net_9237;
wire net_16264;
wire net_6203;
wire net_3006;
wire net_19513;
wire net_16778;
wire net_16273;
wire net_10970;
wire net_16131;
wire net_1681;
wire net_7936;
wire net_17632;
wire net_14468;
wire net_7998;
wire net_15511;
wire net_4272;
wire net_19212;
wire net_16726;
wire net_6512;
wire net_10532;
wire net_19316;
wire net_746;
wire net_13406;
wire net_6147;
wire net_5877;
wire net_17153;
wire net_1274;
wire net_1682;
wire net_11302;
wire net_5743;
wire net_10788;
wire net_7910;
wire net_14485;
wire net_19776;
wire net_18555;
wire net_10109;
wire net_3466;
wire net_16623;
wire net_15784;
wire net_21123;
wire net_4995;
wire net_7834;
wire net_20648;
wire net_22729;
wire net_1663;
wire net_629;
wire net_20845;
wire net_14579;
wire net_4209;
wire net_8666;
wire net_15326;
wire net_19263;
wire net_9382;
wire net_3019;
wire net_13784;
wire net_15017;
wire net_5579;
wire net_14710;
wire net_2351;
wire net_20730;
wire net_18950;
wire net_17244;
wire net_1350;
wire net_9628;
wire net_14457;
wire net_1648;
wire net_20505;
wire net_6219;
wire net_12594;
wire x5992;
wire net_631;
wire net_14201;
wire net_12128;
wire net_20948;
wire net_16603;
wire net_10086;
wire net_17811;
wire net_14988;
wire net_13143;
wire net_4007;
wire net_4499;
wire net_8566;
wire net_12100;
wire net_9910;
wire net_15733;
wire net_16306;
wire net_6928;
wire net_670;
wire net_19479;
wire net_15159;
wire net_6250;
wire net_2687;
wire net_9889;
wire net_7023;
wire net_22473;
wire net_21810;
wire net_10750;
wire net_9721;
wire net_9842;
wire net_22352;
wire net_12853;
wire net_20135;
wire net_22577;
wire net_16687;
wire net_3928;
wire net_13369;
wire net_19187;
wire net_14540;
wire net_7038;
wire net_3854;
wire x413;
wire net_21588;
wire net_22329;
wire net_6717;
wire net_9793;
wire net_9857;
wire net_5493;
wire net_13759;
wire net_755;
wire net_17522;
wire net_9557;
wire net_7754;
wire net_9285;
wire net_14981;
wire net_12545;
wire net_5892;
wire x3951;
wire net_16187;
wire net_13468;
wire net_20585;
wire net_3151;
wire net_14953;
wire net_6763;
wire net_12890;
wire net_6053;
wire net_3628;
wire net_18778;
wire net_12023;
wire net_18223;
wire net_14479;
wire net_12829;
wire net_16303;
wire net_20961;
wire net_1652;
wire net_11319;
wire net_16213;
wire net_1429;
wire net_11061;
wire net_14223;
wire net_14895;
wire net_7130;
wire net_18851;
wire net_15223;
wire net_2725;
wire net_3613;
wire net_13166;
wire net_8964;
wire net_4615;
wire net_727;
wire net_11242;
wire net_9804;
wire net_20218;
wire net_16259;
wire net_12559;
wire net_4955;
wire net_3190;
wire net_16022;
wire net_3757;
wire net_11457;
wire net_15750;
wire net_21111;
wire net_18836;
wire net_9224;
wire net_12658;
wire net_4445;
wire net_19090;
wire net_15142;
wire net_11115;
wire net_14247;
wire net_20422;
wire net_3951;
wire net_14614;
wire net_15054;
wire net_11635;
wire net_13010;
wire net_2259;
wire net_12124;
wire net_15079;
wire net_10651;
wire net_15107;
wire net_22488;
wire net_19905;
wire net_21958;
wire net_20834;
wire net_16319;
wire net_4095;
wire net_2739;
wire net_13330;
wire net_10113;
wire net_11715;
wire net_2110;
wire net_2919;
wire net_10642;
wire net_2893;
wire net_11435;
wire net_3227;
wire net_2358;
wire net_16335;
wire net_17465;
wire net_12651;
wire net_21306;
wire net_8682;
wire net_19206;
wire net_3057;
wire net_9039;
wire net_571;
wire net_22723;
wire net_21756;
wire net_10692;
wire net_10543;
wire net_7569;
wire net_16719;
wire net_21129;
wire net_14743;
wire net_19760;
wire net_10400;
wire net_4935;
wire net_3934;
wire net_12168;
wire net_17938;
wire net_10385;
wire net_19309;
wire net_1877;
wire net_16107;
wire net_720;
wire net_19225;
wire net_7653;
wire net_9038;
wire net_12152;
wire net_15978;
wire net_18752;
wire net_14005;
wire net_18509;
wire net_5209;
wire net_2199;
wire net_10628;
wire net_22295;
wire net_684;
wire net_2648;
wire net_16414;
wire net_7299;
wire net_7542;
wire net_22304;
wire net_3720;
wire net_510;
wire net_12922;
wire net_10909;
wire net_20314;
wire net_21041;
wire net_15808;
wire net_21120;
wire net_8885;
wire x4261;
wire net_2653;
wire net_19807;
wire net_2960;
wire net_9078;
wire net_8257;
wire net_6703;
wire net_12577;
wire net_7043;
wire net_2782;
wire net_494;
wire net_17364;
wire net_17693;
wire net_10999;
wire net_12877;
wire net_20429;
wire net_22540;
wire net_19488;
wire net_4283;
wire net_15726;
wire net_6592;
wire net_13830;
wire net_18095;
wire net_16044;
wire net_6084;
wire net_8953;
wire net_20094;
wire net_3461;
wire net_12365;
wire net_21955;
wire net_10327;
wire net_10956;
wire net_11747;
wire net_4610;
wire net_14366;
wire net_4459;
wire net_457;
wire net_2246;
wire net_8821;
wire net_12096;
wire net_772;
wire net_10180;
wire net_4371;
wire net_14375;
wire net_19249;
wire net_10190;
wire net_12773;
wire net_7966;
wire net_11807;
wire net_1277;
wire net_14567;
wire net_17712;
wire net_2661;
wire net_22112;
wire net_19675;
wire net_16496;
wire net_6113;
wire net_3893;
wire net_13459;
wire net_18988;
wire net_12467;
wire net_4075;
wire net_6421;
wire net_20597;
wire net_7385;
wire net_18589;
wire net_6051;
wire net_2852;
wire net_1721;
wire net_7851;
wire net_16370;
wire net_12975;
wire net_4633;
wire net_22495;
wire net_6605;
wire net_6249;
wire net_5843;
wire net_22501;
wire net_10626;
wire net_1073;
wire net_8073;
wire net_18064;
wire net_17626;
wire net_1947;
wire net_11932;
wire net_22215;
wire x3732;
wire net_19800;
wire net_141;
wire net_879;
wire net_7227;
wire net_2415;
wire x3007;
wire net_15034;
wire net_8738;
wire net_7312;
wire net_13225;
wire net_3197;
wire net_1348;
wire net_10740;
wire net_15707;
wire net_17371;
wire net_9774;
wire net_7276;
wire net_21215;
wire net_16997;
wire net_17388;
wire net_7201;
wire x3910;
wire net_18781;
wire net_16017;
wire net_19357;
wire net_3422;
wire net_199;
wire net_10151;
wire net_2789;
wire x5145;
wire net_7844;
wire net_16397;
wire net_3835;
wire net_431;
wire net_12903;
wire net_5783;
wire net_20260;
wire net_8250;
wire net_17874;
wire net_21703;
wire net_9373;
wire net_10898;
wire net_5186;
wire net_19688;
wire net_22618;
wire net_4362;
wire net_222;
wire net_13215;
wire net_17255;
wire net_4520;
wire net_15727;
wire net_7060;
wire net_3999;
wire net_7804;
wire net_1788;
wire net_16694;
wire net_4301;
wire net_12476;
wire net_21325;
wire net_2935;
wire net_20295;
wire net_6166;
wire x2272;
wire net_18841;
wire net_4345;
wire net_10507;
wire net_9318;
wire net_22759;
wire net_3516;
wire net_6547;
wire net_11799;
wire net_4588;
wire net_1438;
wire net_10374;
wire x5290;
wire net_4395;
wire net_8502;
wire net_20253;
wire net_21880;
wire net_1143;
wire net_14580;
wire net_15884;
wire net_1088;
wire net_6410;
wire net_9434;
wire net_20952;
wire net_19095;
wire net_19068;
wire net_13262;
wire net_3885;
wire net_706;
wire net_18015;
wire net_6373;
wire net_9298;
wire net_14376;
wire net_21845;
wire net_2768;
wire net_5125;
wire net_17575;
wire net_551;
wire net_12536;
wire net_13479;
wire net_5368;
wire net_7873;
wire net_4617;
wire net_20166;
wire net_13182;
wire net_15000;
wire x7642;
wire net_11033;
wire net_4168;
wire net_12419;
wire net_12376;
wire net_16979;
wire net_1199;
wire net_11371;
wire net_18081;
wire net_7986;
wire net_8930;
wire net_15675;
wire net_3627;
wire net_14764;
wire net_18032;
wire net_15087;
wire net_5530;
wire net_15296;
wire net_4869;
wire net_450;
wire net_289;
wire net_19021;
wire net_8041;
wire net_9046;
wire net_14204;
wire net_10972;
wire net_2614;
wire net_1642;
wire net_12158;
wire net_5322;
wire net_16958;
wire net_22165;
wire net_2524;
wire net_11490;
wire net_1224;
wire net_21902;
wire net_6786;
wire net_13804;
wire net_768;
wire net_22029;
wire net_11084;
wire net_14423;
wire net_14068;
wire net_908;
wire net_19028;
wire net_18969;
wire net_13189;
wire net_519;
wire net_9697;
wire net_11773;
wire net_19403;
wire net_22672;
wire net_11052;
wire net_2697;
wire net_22659;
wire net_15825;
wire net_9184;
wire net_10808;
wire x1497;
wire net_6282;
wire net_1204;
wire net_9190;
wire net_14082;
wire net_18216;
wire net_16312;
wire net_14089;
wire net_16923;
wire net_2342;
wire net_7336;
wire net_8331;
wire net_6628;
wire net_9969;
wire net_18719;
wire net_21564;
wire net_6778;
wire net_3214;
wire net_1986;
wire net_16679;
wire net_22098;
wire net_19754;
wire net_14972;
wire net_11472;
wire net_21103;
wire net_10864;
wire net_21878;
wire net_12881;
wire net_18405;
wire net_15321;
wire net_6467;
wire net_8203;
wire net_22014;
wire net_16528;
wire net_7527;
wire net_12613;
wire net_20795;
wire net_19897;
wire net_3406;
wire net_9012;
wire net_9164;
wire net_20991;
wire net_11657;
wire net_4229;
wire net_13110;
wire net_15624;
wire net_6474;
wire net_2130;
wire net_3362;
wire net_1148;
wire net_10198;
wire net_2382;
wire net_13620;
wire net_10698;
wire net_3442;
wire net_5942;
wire net_3864;
wire net_9271;
wire net_15357;
wire net_17063;
wire net_5796;
wire x339831;
wire net_9730;
wire net_20669;
wire net_14725;
wire net_9416;
wire net_6975;
wire net_19448;
wire net_16355;
wire net_4389;
wire net_11798;
wire net_13935;
wire net_19967;
wire net_10728;
wire net_10425;
wire net_4561;
wire net_11676;
wire net_22185;
wire net_14800;
wire net_1473;
wire net_15964;
wire net_41;
wire net_1674;
wire net_5582;
wire net_1651;
wire net_2375;
wire net_19658;
wire net_5109;
wire net_13582;
wire net_6422;
wire net_1806;
wire net_3234;
wire net_15666;
wire net_17578;
wire net_17211;
wire net_8746;
wire net_1363;
wire net_1869;
wire net_4053;
wire net_21424;
wire net_10526;
wire net_13029;
wire net_15713;
wire net_19980;
wire net_19018;
wire net_16863;
wire net_4012;
wire net_6169;
wire net_18975;
wire net_6647;
wire net_18503;
wire net_19291;
wire net_3681;
wire net_20685;
wire net_6621;
wire net_7902;
wire net_13097;
wire net_22078;
wire net_7503;
wire net_7857;
wire net_12717;
wire net_10015;
wire net_14522;
wire net_15180;
wire net_5246;
wire net_17982;
wire net_351;
wire x5637;
wire net_8558;
wire net_7761;
wire x5099;
wire net_19878;
wire net_12601;
wire net_6006;
wire net_10856;
wire net_4240;
wire net_7964;
wire net_15581;
wire net_2842;
wire net_21140;
wire net_21422;
wire net_3158;
wire net_1257;
wire net_939;
wire net_8365;
wire net_22248;
wire net_18810;
wire net_17424;
wire net_13781;
wire net_7984;
wire net_14411;
wire net_21003;
wire net_2791;
wire net_10479;
wire net_10111;
wire net_16513;
wire net_11023;
wire net_22442;
wire net_4271;
wire net_8795;
wire net_15047;
wire x2650;
wire net_9895;
wire net_11817;
wire net_317;
wire net_856;
wire net_17001;
wire net_11853;
wire net_9944;
wire net_7920;
wire net_3845;
wire net_16756;
wire net_2026;
wire net_19989;
wire net_16209;
wire net_5727;
wire net_11822;
wire net_21022;
wire net_18004;
wire net_16611;
wire net_5673;
wire net_12195;
wire net_3033;
wire net_16567;
wire net_14059;
wire net_19915;
wire net_18931;
wire net_17037;
wire net_3373;
wire net_20884;
wire net_5382;
wire net_17854;
wire net_2672;
wire net_11471;
wire net_5351;
wire net_22652;
wire net_588;
wire net_16648;
wire net_2200;
wire net_8641;
wire net_1157;
wire net_7486;
wire net_7785;
wire net_21157;
wire net_6001;
wire net_21639;
wire net_9378;
wire net_19080;
wire net_21523;
wire net_14198;
wire net_19796;
wire net_16922;
wire net_6350;
wire net_7993;
wire net_9840;
wire net_10560;
wire net_14270;
wire net_11800;
wire net_17704;
wire net_13604;
wire net_5603;
wire net_20983;
wire net_17830;
wire net_1065;
wire net_13117;
wire net_22464;
wire net_21721;
wire net_15831;
wire net_3795;
wire net_16245;
wire net_13046;
wire net_16450;
wire net_3100;
wire net_15696;
wire net_13375;
wire net_241;
wire net_9353;
wire net_13196;
wire net_12010;
wire net_13515;
wire net_13640;
wire net_21508;
wire x1121;
wire net_13350;
wire net_4597;
wire net_16291;
wire net_599;
wire net_13814;
wire net_20452;
wire net_4589;
wire net_22020;
wire net_21440;
wire net_4844;
wire net_21935;
wire net_21195;
wire net_5860;
wire net_3111;
wire net_19165;
wire net_18437;
wire net_20656;
wire net_21380;
wire net_10346;
wire net_11880;
wire net_13543;
wire net_16765;
wire net_9653;
wire net_21091;
wire net_8692;
wire net_13575;
wire net_8356;
wire net_18445;
wire net_3737;
wire net_18049;
wire net_6103;
wire net_15384;
wire net_18645;
wire net_12260;
wire net_15752;
wire net_19789;
wire net_15918;
wire net_20239;
wire net_9686;
wire net_17141;
wire net_2849;
wire net_12671;
wire net_18638;
wire net_10799;
wire net_15641;
wire net_15267;
wire net_12693;
wire net_5589;
wire net_17535;
wire net_4873;
wire net_10851;
wire net_16461;
wire net_4298;
wire net_20913;
wire net_16564;
wire net_21566;
wire net_11286;
wire net_15175;
wire net_20217;
wire net_18812;
wire net_16876;
wire net_7170;
wire net_8004;
wire net_11250;
wire net_4137;
wire net_8528;
wire net_5162;
wire net_9870;
wire net_20328;
wire net_17545;
wire net_7561;
wire net_5765;
wire net_3496;
wire net_15010;
wire net_20522;
wire net_4216;
wire net_13361;
wire net_20529;
wire net_98;
wire net_4889;
wire x1087;
wire net_19681;
wire net_10371;
wire net_151;
wire net_22330;
wire net_16950;
wire net_1625;
wire net_13638;
wire net_8784;
wire net_9930;
wire net_17915;
wire net_2513;
wire net_8662;
wire net_7360;
wire net_7142;
wire net_10291;
wire net_187;
wire net_21524;
wire net_3305;
wire net_14072;
wire net_21207;
wire net_20622;
wire net_14045;
wire net_18310;
wire net_160;
wire net_832;
wire net_12304;
wire net_19234;
wire net_7728;
wire net_6749;
wire net_5578;
wire net_18659;
wire net_13742;
wire net_6501;
wire net_17868;
wire net_16577;
wire net_9580;
wire net_5272;
wire net_20856;
wire net_6240;
wire net_3838;
wire net_7812;
wire net_7768;
wire net_21870;
wire net_22665;
wire net_11518;
wire net_19031;
wire net_6260;
wire net_120;
wire net_15116;
wire net_292;
wire net_12489;
wire net_5529;
wire net_96;
wire net_9384;
wire net_12141;
wire net_167;
wire net_12371;
wire net_21601;
wire net_7308;
wire net_6170;
wire x3820;
wire net_8864;
wire net_15325;
wire net_9847;
wire net_15849;
wire net_5735;
wire net_20352;
wire net_2806;
wire net_9679;
wire net_13163;
wire net_14624;
wire net_4924;
wire net_20483;
wire net_21634;
wire net_4483;
wire net_8391;
wire net_9367;
wire net_5045;
wire net_14441;
wire x2971;
wire net_17540;
wire net_6237;
wire net_11335;
wire net_2456;
wire net_2753;
wire net_1232;
wire net_10036;
wire net_14635;
wire net_4540;
wire net_9585;
wire net_19078;
wire net_5662;
wire net_3059;
wire net_11625;
wire net_13506;
wire net_10684;
wire net_12540;
wire net_5444;
wire net_17090;
wire net_13039;
wire net_22400;
wire net_17436;
wire net_464;
wire net_12003;
wire net_17286;
wire net_5699;
wire net_5089;
wire net_4200;
wire net_21828;
wire net_6300;
wire net_5867;
wire net_22316;
wire net_16629;
wire net_5362;
wire net_19599;
wire net_20002;
wire net_20628;
wire net_21435;
wire net_18539;
wire net_4658;
wire net_12625;
wire net_14195;
wire net_14602;
wire net_1256;
wire net_1413;
wire x339;
wire net_14252;
wire net_15262;
wire net_18997;
wire net_3556;
wire net_1840;
wire net_3041;
wire net_13872;
wire net_12602;
wire net_20926;
wire net_5637;
wire net_8015;
wire net_7167;
wire net_3427;
wire net_1031;
wire net_13170;
wire net_22695;
wire net_10265;
wire net_13394;
wire net_7245;
wire net_22173;
wire net_7458;
wire net_9744;
wire net_10467;
wire net_21888;
wire net_10991;
wire net_1688;
wire net_2020;
wire net_8523;
wire net_16787;
wire net_15968;
wire net_10794;
wire net_13522;
wire net_22415;
wire net_7665;
wire net_13383;
wire net_15858;
wire net_6126;
wire net_19731;
wire net_14056;
wire net_17527;
wire net_15076;
wire net_16684;
wire net_4324;
wire net_4159;
wire net_7322;
wire net_2374;
wire net_20347;
wire net_4203;
wire net_9911;
wire net_17663;
wire x6966;
wire net_20813;
wire net_20040;
wire net_16039;
wire net_10571;
wire net_250;
wire net_20827;
wire net_3600;
wire net_8655;
wire net_7260;
wire net_5882;
wire net_2055;
wire net_12929;
wire net_19625;
wire net_7420;
wire net_403;
wire net_10027;
wire net_3524;
wire net_6265;
wire net_13680;
wire net_12219;
wire net_15560;
wire net_18699;
wire net_14302;
wire net_22278;
wire net_9899;
wire net_19000;
wire net_12202;
wire net_12562;
wire net_8602;
wire net_14910;
wire net_794;
wire net_2397;
wire net_8136;
wire net_13277;
wire net_21839;
wire net_10537;
wire net_3433;
wire net_1468;
wire net_20812;
wire net_4774;
wire net_21138;
wire net_11767;
wire net_16360;
wire net_39;
wire net_7350;
wire net_8494;
wire net_6796;
wire net_1130;
wire net_5921;
wire net_14826;
wire net_8111;
wire net_8239;
wire net_9421;
wire net_19075;
wire x1259;
wire net_6451;
wire net_7918;
wire net_6493;
wire net_9281;
wire net_7745;
wire net_6309;
wire net_2318;
wire net_8787;
wire net_9207;
wire net_5562;
wire net_17166;
wire net_3449;
wire net_9004;
wire net_9134;
wire net_18463;
wire net_17475;
wire net_1039;
wire net_7822;
wire net_11972;
wire net_4651;
wire net_400;
wire net_8629;
wire net_15499;
wire net_20489;
wire net_14546;
wire net_1935;
wire net_11608;
wire net_19700;
wire net_13102;
wire net_2925;
wire net_9142;
wire net_11873;
wire net_18826;
wire x3242;
wire net_1855;
wire net_14956;
wire net_4882;
wire net_1163;
wire net_1177;
wire net_10206;
wire net_13890;
wire net_5466;
wire net_9521;
wire net_21099;
wire net_16053;
wire net_7840;
wire net_17029;
wire net_9215;
wire net_11494;
wire net_3273;
wire net_17978;
wire net_1559;
wire net_20425;
wire net_5665;
wire net_8706;
wire net_1620;
wire net_2608;
wire net_13966;
wire net_14266;
wire net_2813;
wire net_9763;
wire net_14856;
wire x2809;
wire net_14559;
wire net_719;
wire net_21345;
wire net_10878;
wire net_18234;
wire net_6873;
wire net_8068;
wire net_14032;
wire net_19648;
wire net_2571;
wire net_9888;
wire net_16892;
wire net_19258;
wire net_17886;
wire net_16066;
wire net_5703;
wire net_12264;
wire net_9418;
wire net_14325;
wire net_3479;
wire net_22512;
wire net_20384;
wire net_8609;
wire net_22412;
wire net_3222;
wire net_13617;
wire net_16134;
wire net_6393;
wire net_8410;
wire net_3552;
wire net_15314;
wire net_19834;
wire net_696;
wire net_7427;
wire net_5713;
wire net_10777;
wire net_10824;
wire net_14079;
wire net_17824;
wire net_13175;
wire net_22041;
wire net_10401;
wire net_13947;
wire net_16058;
wire net_12972;
wire net_12256;
wire net_10448;
wire net_15599;
wire net_16093;
wire net_9953;
wire net_15492;
wire net_22468;
wire net_21753;
wire net_17998;
wire net_3821;
wire net_16217;
wire net_9228;
wire net_14101;
wire net_8403;
wire net_4503;
wire net_10872;
wire net_20077;
wire net_6938;
wire net_19113;
wire net_3486;
wire net_7359;
wire net_15241;
wire net_19933;
wire net_17333;
wire net_5839;
wire net_7955;
wire net_8590;
wire net_11199;
wire net_19724;
wire net_8919;
wire net_9981;
wire net_8302;
wire net_1298;
wire net_296;
wire net_9733;
wire x315;
wire net_16040;
wire net_7004;
wire net_12053;
wire net_18574;
wire net_8941;
wire net_19886;
wire net_5435;
wire net_17461;
wire net_18071;
wire net_11461;
wire net_18568;
wire net_3020;
wire net_17233;
wire net_13720;
wire net_22461;
wire net_18205;
wire net_10518;
wire net_1339;
wire net_10608;
wire net_22450;
wire net_3781;
wire net_17169;
wire net_5685;
wire net_906;
wire net_15450;
wire net_2422;
wire net_5205;
wire net_21842;
wire net_13951;
wire net_652;
wire net_10185;
wire net_12955;
wire net_13958;
wire net_13707;
wire net_10590;
wire net_10211;
wire net_14840;
wire net_14513;
wire net_19366;
wire net_2505;
wire net_11185;
wire net_19290;
wire net_16988;
wire net_10748;
wire net_20049;
wire net_6139;
wire net_2683;
wire net_21069;
wire net_17516;
wire net_21106;
wire net_4812;
wire net_16180;
wire net_4253;
wire net_2165;
wire net_11943;
wire net_8315;
wire net_6861;
wire net_18821;
wire net_11049;
wire net_20735;
wire net_2562;
wire net_15417;
wire net_5134;
wire net_5293;
wire net_9129;
wire net_14931;
wire net_7195;
wire net_13841;
wire net_16079;
wire net_8151;
wire net_19985;
wire net_5172;
wire net_22743;
wire net_2182;
wire net_8145;
wire net_10092;
wire net_4718;
wire net_8032;
wire net_9928;
wire net_9295;
wire net_150;
wire net_19285;
wire net_6589;
wire net_21680;
wire net_16151;
wire net_11915;
wire net_4351;
wire net_6993;
wire net_10951;
wire net_12436;
wire net_15773;
wire net_22769;
wire net_7666;
wire net_1703;
wire net_12768;
wire net_11004;
wire net_7848;
wire net_9420;
wire net_22273;
wire net_9690;
wire net_3693;
wire net_19323;
wire net_9027;
wire net_5100;
wire net_4319;
wire net_14849;
wire net_18317;
wire net_16246;
wire net_3070;
wire net_13695;
wire net_3409;
wire net_9481;
wire net_17022;
wire net_4525;
wire net_16782;
wire net_1904;
wire net_3907;
wire net_9446;
wire x6071;
wire net_6332;
wire net_16493;
wire net_6584;
wire net_10001;
wire net_8617;
wire net_21464;
wire net_2187;
wire net_17639;
wire net_19919;
wire net_10764;
wire net_3387;
wire net_13242;
wire net_7157;
wire net_1479;
wire net_16127;
wire net_10268;
wire net_15611;
wire net_18532;
wire net_6895;
wire net_10066;
wire net_3094;
wire net_1927;
wire net_10243;
wire net_21920;
wire net_213;
wire net_6910;
wire net_19153;
wire net_9244;
wire net_947;
wire net_5359;
wire net_7970;
wire net_1126;
wire net_14715;
wire net_2004;
wire net_11538;
wire net_16636;
wire net_6943;
wire net_1325;
wire net_16474;
wire net_5094;
wire net_6298;
wire net_2567;
wire net_10258;
wire net_10944;
wire net_14029;
wire net_22525;
wire net_7643;
wire net_21372;
wire net_7411;
wire net_21679;
wire net_16445;
wire net_1303;
wire net_16158;
wire net_8050;
wire net_18029;
wire net_21472;
wire net_16834;
wire net_6334;
wire net_22491;
wire net_18260;
wire net_2102;
wire net_4451;
wire x1283;
wire net_1807;
wire net_11903;
wire net_20773;
wire net_20493;
wire net_1930;
wire net_1943;
wire net_21406;
wire net_20769;
wire net_17493;
wire net_16994;
wire net_20792;
wire net_22773;
wire net_19087;
wire net_17955;
wire net_20471;
wire net_16471;
wire net_12113;
wire net_4054;
wire net_11555;
wire net_5544;
wire net_18180;
wire net_113;
wire net_15842;
wire net_18744;
wire net_5054;
wire net_9674;
wire net_4848;
wire net_19993;
wire net_7791;
wire net_16114;
wire net_18165;
wire net_3889;
wire net_20405;
wire net_14899;
wire net_14039;
wire net_19528;
wire net_3567;
wire net_13717;
wire net_7831;
wire net_11525;
wire net_19557;
wire net_22539;
wire net_6483;
wire net_16323;
wire net_6616;
wire net_2448;
wire net_15285;
wire net_5424;
wire net_5541;
wire net_13234;
wire net_10719;
wire net_3400;
wire net_17601;
wire net_14925;
wire net_646;
wire net_5823;
wire net_2731;
wire net_20875;
wire net_19910;
wire net_2601;
wire net_11016;
wire net_8902;
wire net_8499;
wire net_520;
wire net_10159;
wire net_13482;
wire net_7237;
wire net_11201;
wire net_4722;
wire x6585;
wire net_14110;
wire net_20418;
wire net_16061;
wire net_21133;
wire net_3231;
wire net_21421;
wire net_981;
wire net_18961;
wire net_19721;
wire net_9636;
wire net_8895;
wire net_1566;
wire net_17941;
wire net_11584;
wire net_2354;
wire net_12156;
wire net_9393;
wire net_21430;
wire net_10378;
wire net_10709;
wire net_10440;
wire net_5018;
wire net_8858;
wire net_15676;
wire net_19561;
wire net_7369;
wire net_5013;
wire net_15856;
wire net_559;
wire net_11413;
wire net_16886;
wire net_3042;
wire net_12804;
wire net_7476;
wire net_1717;
wire net_6553;
wire net_398;
wire net_3399;
wire net_6976;
wire net_17072;
wire net_16943;
wire net_6693;
wire net_22135;
wire net_2117;
wire net_12834;
wire net_4085;
wire net_7393;
wire net_13493;
wire x2174;
wire net_10099;
wire net_17797;
wire net_12472;
wire net_18617;
wire net_20000;
wire net_5905;
wire net_9788;
wire net_15233;
wire net_17589;
wire net_6724;
wire net_6054;
wire net_18845;
wire net_18130;
wire net_1572;
wire net_11647;
wire net_9265;
wire net_5179;
wire net_2134;
wire net_15595;
wire net_20134;
wire net_5011;
wire net_316;
wire net_4250;
wire x719;
wire net_13439;
wire net_4961;
wire net_15303;
wire net_4184;
wire net_11462;
wire net_14736;
wire net_14398;
wire net_7033;
wire net_14962;
wire net_17906;
wire net_4647;
wire net_16523;
wire net_4022;
wire net_15649;
wire net_20718;
wire net_18553;
wire net_17490;
wire net_9618;
wire net_8347;
wire net_13282;
wire net_10040;
wire net_1695;
wire net_5932;
wire net_1617;
wire net_7005;
wire net_20457;
wire net_22457;
wire net_5969;
wire net_16815;
wire net_19866;
wire net_9332;
wire net_19887;
wire net_18892;
wire net_4579;
wire net_568;
wire net_13809;
wire net_4807;
wire net_1227;
wire net_6046;
wire net_1008;
wire net_5340;
wire net_21147;
wire net_18848;
wire net_21152;
wire net_12178;
wire net_19508;
wire net_4862;
wire net_3069;
wire net_3170;
wire net_12239;
wire net_22347;
wire net_20010;
wire net_22590;
wire net_4819;
wire net_21553;
wire net_17613;
wire net_17144;
wire net_14773;
wire net_14533;
wire net_19971;
wire net_15794;
wire net_469;
wire net_22355;
wire net_1978;
wire net_21280;
wire net_18307;
wire net_21053;
wire net_3167;
wire net_1170;
wire net_5656;
wire net_10144;
wire net_2280;
wire net_13202;
wire net_9174;
wire net_778;
wire net_2366;
wire net_21697;
wire net_21153;
wire net_1455;
wire net_2930;
wire net_20308;
wire net_9816;
wire net_15937;
wire net_14277;
wire net_20273;
wire net_15651;
wire net_16252;
wire net_16533;
wire net_5323;
wire net_22396;
wire net_12167;
wire net_6225;
wire net_18654;
wire net_6832;
wire net_5261;
wire net_4730;
wire net_6643;
wire net_11123;
wire net_17505;
wire net_15292;
wire net_20956;
wire net_19240;
wire net_4119;
wire net_18148;
wire net_16976;
wire net_9216;
wire net_9450;
wire net_13445;
wire net_18037;
wire net_10335;
wire x1362;
wire net_5645;
wire net_995;
wire net_15763;
wire net_8328;
wire net_17790;
wire net_7088;
wire net_7334;
wire net_12232;
wire x6145;
wire net_1246;
wire net_8957;
wire net_7705;
wire net_13325;
wire net_1774;
wire net_16162;
wire net_4228;
wire net_11402;
wire net_3060;
wire net_10712;
wire net_2568;
wire net_11103;
wire net_17008;
wire net_321;
wire net_5518;
wire net_9465;
wire net_17708;
wire net_19717;
wire net_2995;
wire net_16912;
wire net_3526;
wire net_15532;
wire net_22445;
wire net_934;
wire net_22804;
wire net_21535;
wire net_18795;
wire net_3103;
wire net_21096;
wire net_5941;
wire net_4896;
wire net_3630;
wire net_11952;
wire net_1824;
wire net_12037;
wire net_7603;
wire net_16008;
wire net_4763;
wire net_5074;
wire net_5694;
wire net_20058;
wire net_19395;
wire net_3166;
wire net_18983;
wire net_7065;
wire net_9104;
wire net_8079;
wire net_9831;
wire net_10861;
wire net_7513;
wire net_18272;
wire net_9652;
wire net_10665;
wire net_5552;
wire net_860;
wire net_20213;
wire net_16566;
wire net_19873;
wire net_9254;
wire net_2046;
wire net_14474;
wire net_7926;
wire net_11708;
wire net_2878;
wire net_2871;
wire net_9850;
wire net_18325;
wire net_21385;
wire net_3267;
wire net_20190;
wire net_2321;
wire net_9108;
wire net_21255;
wire net_817;
wire net_11667;
wire net_3414;
wire net_15006;
wire net_18349;
wire net_14804;
wire net_7058;
wire net_10967;
wire net_13502;
wire net_21025;
wire net_9766;
wire net_4576;
wire net_13655;
wire net_13344;
wire net_14123;
wire net_13278;
wire net_5483;
wire net_2012;
wire net_7139;
wire net_5557;
wire net_19201;
wire net_9890;
wire net_15178;
wire net_16690;
wire net_743;
wire net_3770;
wire net_14387;
wire net_1922;
wire net_9062;
wire net_15333;
wire net_14620;
wire net_17728;
wire net_6639;
wire net_12384;
wire net_8264;
wire net_2451;
wire net_13499;
wire net_14332;
wire net_17012;
wire net_17019;
wire net_4031;
wire net_1522;
wire net_22702;
wire net_20677;
wire net_2926;
wire net_12782;
wire net_15881;
wire net_16745;
wire net_8042;
wire net_12289;
wire net_17444;
wire net_13751;
wire net_18883;
wire net_6991;
wire net_4551;
wire net_5972;
wire net_13557;
wire net_18588;
wire net_12945;
wire net_3943;
wire net_9370;
wire net_14996;
wire net_21429;
wire net_19564;
wire net_22093;
wire net_15183;
wire net_17305;
wire net_7675;
wire net_4438;
wire net_56;
wire net_10839;
wire net_20371;
wire net_8557;
wire net_14154;
wire net_968;
wire net_17357;
wire net_13876;
wire net_13572;
wire net_9669;
wire net_10421;
wire net_12692;
wire net_19497;
wire net_16574;
wire net_17232;
wire net_18416;
wire net_2534;
wire net_6827;
wire net_4133;
wire net_15930;
wire net_22541;
wire net_3732;
wire net_17835;
wire net_16429;
wire net_2309;
wire net_502;
wire net_8647;
wire net_16047;
wire net_1564;
wire net_20861;
wire net_6632;
wire net_3804;
wire net_12282;
wire net_10883;
wire net_15353;
wire net_9398;
wire net_17106;
wire net_17046;
wire net_13271;
wire net_8290;
wire net_19570;
wire net_16707;
wire net_12209;
wire net_13858;
wire net_7990;
wire net_19896;
wire net_4112;
wire net_3868;
wire net_7121;
wire net_5887;
wire net_13233;
wire net_20996;
wire net_2628;
wire net_4512;
wire net_6535;
wire net_9305;
wire net_11692;
wire net_17449;
wire net_5145;
wire net_11439;
wire net_12757;
wire net_21987;
wire net_11160;
wire net_19550;
wire net_20803;
wire net_20726;
wire net_9047;
wire net_10494;
wire net_20613;
wire net_11078;
wire net_13837;
wire net_13800;
wire net_664;
wire net_20337;
wire net_19371;
wire net_6292;
wire net_4622;
wire net_22606;
wire net_4605;
wire net_4295;
wire net_10450;
wire net_10687;
wire net_12533;
wire net_15684;
wire x1291;
wire net_5773;
wire net_10614;
wire net_6405;
wire net_20033;
wire net_17085;
wire net_21960;
wire net_18448;
wire net_13550;
wire net_14779;
wire net_7469;
wire net_21691;
wire net_6210;
wire net_2952;
wire x592;
wire net_21866;
wire net_2035;
wire net_17429;
wire net_17403;
wire net_5070;
wire net_2826;
wire net_21998;
wire net_10451;
wire net_17173;
wire net_6847;
wire net_2141;
wire net_15123;
wire net_10830;
wire net_14211;
wire net_22677;
wire net_11803;
wire net_22651;
wire net_14818;
wire net_15866;
wire net_19012;
wire net_11213;
wire net_3453;
wire net_5702;
wire net_12648;
wire net_8632;
wire net_110;
wire net_9822;
wire net_10598;
wire net_15447;
wire net_6097;
wire net_1403;
wire net_4532;
wire net_2270;
wire net_1667;
wire net_7208;
wire net_22683;
wire net_8882;
wire net_1606;
wire net_3710;
wire net_15156;
wire net_3054;
wire net_7683;
wire net_21269;
wire net_17680;
wire net_8765;
wire net_3978;
wire net_16802;
wire net_4752;
wire net_12708;
wire net_15403;
wire net_15704;
wire net_2029;
wire net_5328;
wire net_3698;
wire net_11560;
wire net_4629;
wire net_2587;
wire net_20263;
wire net_2959;
wire net_1888;
wire net_11836;
wire net_9974;
wire net_4311;
wire net_18690;
wire net_22325;
wire net_12583;
wire net_16848;
wire net_1792;
wire net_2496;
wire net_4125;
wire net_17053;
wire net_10656;
wire net_22237;
wire net_3109;
wire net_1598;
wire net_17390;
wire net_14192;
wire net_21893;
wire net_731;
wire net_14369;
wire net_17221;
wire net_15063;
wire net_22203;
wire net_17698;
wire net_15896;
wire net_22496;
wire net_13042;
wire net_19467;
wire net_18185;
wire net_21463;
wire net_19955;
wire net_7287;
wire net_9704;
wire net_1733;
wire net_5853;
wire net_10576;
wire net_20689;
wire net_5511;
wire net_7590;
wire net_20580;
wire net_17737;
wire net_13962;
wire net_11093;
wire net_6708;
wire x6089;
wire x311;
wire net_10412;
wire net_20419;
wire net_18888;
wire net_4146;
wire net_20651;
wire net_22574;
wire net_1724;
wire net_6106;
wire net_3703;
wire net_12551;
wire net_19689;
wire net_17120;
wire net_12682;
wire net_20555;
wire net_17209;
wire net_12506;
wire net_22644;
wire x3021;
wire net_10843;
wire net_965;
wire net_20897;
wire net_12378;
wire net_15472;
wire net_17129;
wire net_22391;
wire net_16457;
wire net_2916;
wire net_5348;
wire net_421;
wire net_8184;
wire net_8314;
wire net_11976;
wire net_20197;
wire net_1104;
wire net_9783;
wire net_764;
wire net_18120;
wire net_4060;
wire net_5181;
wire net_13009;
wire net_20678;
wire net_18258;
wire net_5038;
wire net_12465;
wire net_7289;
wire net_1117;
wire net_13534;
wire net_16204;
wire net_15552;
wire net_7162;
wire net_6866;
wire net_19170;
wire net_3955;
wire net_13770;
wire net_14531;
wire net_16226;
wire net_5950;
wire net_11893;
wire net_8246;
wire net_20662;
wire net_18852;
wire net_9157;
wire net_18807;
wire net_7252;
wire net_5503;
wire net_2235;
wire net_8303;
wire net_20802;
wire net_11007;
wire net_11329;
wire net_5846;
wire net_21714;
wire net_2080;
wire net_3675;
wire net_6714;
wire net_2711;
wire net_18760;
wire net_2097;
wire net_6194;
wire net_11120;
wire net_3619;
wire net_20157;
wire x1068;
wire net_22242;
wire net_19207;
wire net_15362;
wire x1401;
wire net_1782;
wire net_16828;
wire net_8450;
wire net_11191;
wire net_4863;
wire net_273;
wire net_1278;
wire net_6430;
wire net_4714;
wire net_3182;
wire net_21787;
wire net_12643;
wire net_2098;
wire net_19662;
wire net_4232;
wire net_177;
wire net_3355;
wire net_4305;
wire net_18087;
wire net_7806;
wire net_19334;
wire net_17413;
wire net_19415;
wire net_8739;
wire net_2803;
wire net_3301;
wire net_6370;
wire x643;
wire net_12133;
wire net_6090;
wire net_17338;
wire net_953;
wire net_17640;
wire net_11600;
wire net_11171;
wire net_1074;
wire net_1058;
wire net_7186;
wire net_12728;
wire net_15911;
wire net_9535;
wire net_11295;
wire net_15954;
wire net_21329;
wire net_16658;
wire x6012;
wire net_22104;
wire net_6159;
wire x1215;
wire net_9064;
wire net_14004;
wire net_6962;
wire net_2489;
wire net_18063;
wire net_13829;
wire net_3160;
wire net_2125;
wire net_16173;
wire net_7622;
wire net_19586;
wire net_22301;
wire net_8179;
wire net_19769;
wire net_9546;
wire net_19849;
wire net_13078;
wire net_2623;
wire net_19669;
wire net_16210;
wire net_261;
wire net_8448;
wire net_17757;
wire net_10654;
wire net_15803;
wire net_20598;
wire net_2362;
wire net_12837;
wire net_8869;
wire net_18703;
wire net_4456;
wire net_4354;
wire net_5111;
wire net_1955;
wire net_8507;
wire net_8196;
wire net_12886;
wire net_9729;
wire net_21226;
wire net_18948;
wire net_20209;
wire net_3012;
wire net_21944;
wire net_13134;
wire net_22513;
wire net_6014;
wire net_5367;
wire net_3754;
wire net_10432;
wire net_17328;
wire net_6075;
wire net_9935;
wire net_18357;
wire net_3989;
wire net_11356;
wire net_21498;
wire net_13902;
wire net_7304;
wire net_10515;
wire net_22230;
wire net_5285;
wire net_10875;
wire net_11312;
wire net_1994;
wire net_10499;
wire x1948;
wire net_8574;
wire net_4668;
wire net_3897;
wire net_9288;
wire net_17262;
wire net_3960;
wire net_4374;
wire net_91;
wire net_15983;
wire net_20787;
wire net_16732;
wire net_6152;
wire net_3992;
wire net_15959;
wire net_17773;
wire net_22038;
wire net_21572;
wire net_19301;
wire net_2287;
wire net_4211;
wire net_14590;
wire net_18010;
wire net_21624;
wire net_448;
wire net_8224;
wire net_886;
wire net_3189;
wire net_18466;
wire net_2988;
wire net_18835;
wire net_6811;
wire net_4592;
wire net_20940;
wire net_16304;
wire net_5279;
wire net_19042;
wire net_3651;
wire net_12182;
wire net_21625;
wire net_16710;
wire net_9059;
wire net_14345;
wire net_21287;
wire net_1470;
wire net_11440;
wire net_13358;
wire net_14053;
wire net_4627;
wire net_4423;
wire net_20820;
wire net_15348;
wire net_14796;
wire net_15373;
wire net_13674;
wire net_16557;
wire net_4233;
wire net_18090;
wire net_22823;
wire net_7650;
wire net_4796;
wire net_15057;
wire net_8289;
wire net_2778;
wire net_13662;
wire net_15148;
wire net_2756;
wire net_12896;
wire net_21551;
wire net_22724;
wire net_20178;
wire net_9605;
wire net_21690;
wire net_1085;
wire net_19282;
wire net_592;
wire net_17228;
wire net_9528;
wire net_8983;
wire net_7531;
wire net_2266;
wire net_281;
wire net_8337;
wire net_12493;
wire net_14699;
wire net_17342;
wire net_5254;
wire net_5193;
wire net_5235;
wire net_22255;
wire net_16385;
wire net_18143;
wire net_5520;
wire net_15928;
wire net_21247;
wire net_15344;
wire net_10801;
wire net_10281;
wire net_13532;
wire net_526;
wire net_2718;
wire net_21363;
wire net_13123;
wire net_2747;
wire net_16331;
wire net_14365;
wire net_18016;
wire net_9232;
wire net_12271;
wire net_16192;
wire net_974;
wire net_12348;
wire net_22288;
wire net_11777;
wire net_16858;
wire net_923;
wire net_13853;
wire net_10947;
wire net_1707;
wire net_20362;
wire net_4566;
wire net_2190;
wire net_1881;
wire net_7014;
wire net_10487;
wire net_16607;
wire net_10900;
wire net_12925;
wire net_15788;
wire net_3323;
wire net_11697;
wire net_6347;
wire net_21495;
wire net_20467;
wire net_7867;
wire net_22320;
wire net_22196;
wire net_8961;
wire net_11073;
wire net_20509;
wire net_21971;
wire net_12221;
wire net_1492;
wire net_20799;
wire net_6179;
wire net_14312;
wire net_6363;
wire net_10585;
wire net_21414;
wire net_9275;
wire net_8267;
wire net_2537;
wire net_11088;
wire net_16966;
wire net_14904;
wire net_18211;
wire net_20903;
wire net_3767;
wire net_6919;
wire net_6408;
wire net_80;
wire net_18773;
wire net_4105;
wire net_11984;
wire net_11397;
wire net_5594;
wire net_6132;
wire net_9553;
wire net_9193;
wire net_4569;
wire net_5754;
wire net_34;
wire net_17379;
wire net_15829;
wire net_22505;
wire net_17553;
wire net_13000;
wire net_22438;
wire x1306;
wire net_6214;
wire net_9798;
wire net_15944;
wire net_2049;
wire net_2273;
wire net_11558;
wire net_617;
wire net_11026;
wire net_18158;
wire net_6030;
wire net_8656;
wire net_13456;
wire net_22004;
wire net_4176;
wire net_18486;
wire net_21085;
wire net_16935;
wire net_18402;
wire net_4032;
wire net_4154;
wire net_17565;
wire net_9294;
wire net_9413;
wire net_9794;
wire net_10420;
wire net_7877;
wire net_22282;
wire net_9000;
wire net_20756;
wire net_16505;
wire net_5917;
wire net_5709;
wire net_3870;
wire net_6254;
wire net_18269;
wire net_5456;
wire net_7105;
wire net_15662;
wire net_18383;
wire net_8310;
wire net_5946;
wire net_17296;
wire net_11662;
wire net_21928;
wire net_16281;
wire net_14481;
wire net_8742;
wire net_16984;
wire net_6854;
wire net_14132;
wire net_18271;
wire net_12216;
wire net_16560;
wire net_10082;
wire net_13766;
wire net_384;
wire net_4191;
wire net_3503;
wire net_17324;
wire net_17277;
wire net_16051;
wire net_18953;
wire net_5792;
wire net_13366;
wire net_2599;
wire net_15136;
wire net_2665;
wire net_17355;
wire net_3642;
wire net_9200;
wire net_2707;
wire net_19751;
wire net_7426;
wire net_15834;
wire net_21362;
wire x2468;
wire net_485;
wire x4099;
wire net_20762;
wire net_19108;
wire net_11179;
wire net_19203;
wire net_18106;
wire net_7772;
wire net_64;
wire net_21849;
wire net_15030;
wire net_21211;
wire x6494;
wire net_22158;
wire net_16394;
wire net_7348;
wire net_11364;
wire net_16669;
wire net_18718;
wire net_125;
wire net_11081;
wire net_11589;
wire net_9329;
wire net_22299;
wire net_13402;
wire net_15822;
wire net_1685;
wire x556;
wire net_4768;
wire net_17815;
wire net_12019;
wire net_13147;
wire net_14239;
wire net_2644;
wire net_6102;
wire net_12815;
wire net_18862;
wire net_16774;
wire net_13093;
wire net_21519;
wire net_12686;
wire net_21767;
wire net_286;
wire net_11668;
wire net_19745;
wire net_3584;
wire net_7051;
wire net_21541;
wire net_5588;
wire net_11591;
wire net_4999;
wire net_21656;
wire net_4340;
wire net_10275;
wire net_19463;
wire net_4954;
wire net_17971;
wire net_21119;
wire net_19159;
wire net_16268;
wire net_5878;
wire net_15588;
wire net_10277;
wire net_22141;
wire net_20644;
wire net_3475;
wire net_8423;
wire net_14142;
wire net_5832;
wire net_20223;
wire net_9070;
wire net_8232;
wire net_1951;
wire net_12608;
wire net_19973;
wire net_7292;
wire net_16200;
wire net_12724;
wire net_9759;
wire net_15608;
wire net_8976;
wire net_7661;
wire net_12000;
wire net_15576;
wire net_11869;
wire net_22291;
wire x3339;
wire net_5567;
wire net_2558;
wire net_2040;
wire x4916;
wire net_1508;
wire net_3379;
wire net_931;
wire net_4466;
wire net_20398;
wire net_18936;
wire net_5983;
wire net_18940;
wire net_2242;
wire net_8505;
wire net_22081;
wire net_19816;
wire net_7672;
wire net_6802;
wire net_759;
wire x675;
wire net_7852;
wire net_11711;
wire net_8832;
wire net_11155;
wire net_8083;
wire net_19991;
wire net_18376;
wire net_17781;
wire net_6742;
wire net_6428;
wire net_5242;
wire net_17788;
wire net_6924;
wire net_6516;
wire net_12573;
wire net_14585;
wire net_1341;
wire net_17689;
wire net_4541;
wire net_5210;
wire net_3242;
wire net_8138;
wire net_19998;
wire net_1835;
wire net_18324;
wire net_333;
wire net_15013;
wire net_14491;
wire net_22629;
wire net_9114;
wire net_9322;
wire net_15203;
wire net_22250;
wire net_4664;
wire net_15184;
wire net_18333;
wire net_5976;
wire net_13547;
wire net_20496;
wire net_3923;
wire net_10155;
wire net_21381;
wire net_8839;
wire net_7210;
wire net_20502;
wire net_2554;
wire net_16612;
wire net_12196;
wire net_17934;
wire net_4479;
wire net_15708;
wire net_16276;
wire net_7931;
wire net_14453;
wire x708;
wire net_9716;
wire net_14100;
wire net_22151;
wire net_6354;
wire net_9381;
wire net_13630;
wire net_10928;
wire net_22225;
wire net_10316;
wire net_7980;
wire net_204;
wire net_14885;
wire net_4596;
wire net_13065;
wire net_12932;
wire net_14750;
wire net_19927;
wire net_7626;
wire net_21802;
wire net_19642;
wire net_7382;
wire net_16431;
wire net_16402;
wire net_18641;
wire net_14942;
wire net_15461;
wire net_12045;
wire net_15239;
wire net_5416;
wire net_21972;
wire net_8142;
wire net_17096;
wire net_17161;
wire net_10784;
wire net_19503;
wire net_1916;
wire net_15941;
wire net_14808;
wire net_11419;
wire net_2468;
wire net_21661;
wire net_15306;
wire x659;
wire net_7073;
wire net_16141;
wire net_14416;
wire net_10953;
wire net_19441;
wire net_18412;
wire net_100;
wire net_20573;
wire net_2195;
wire net_11546;
wire net_3421;
wire net_11246;
wire net_1691;
wire net_10089;
wire net_19277;
wire net_9197;
wire net_22383;
wire net_18799;
wire net_595;
wire net_12312;
wire net_1320;
wire net_22331;
wire net_9461;
wire net_22476;
wire net_19853;
wire net_9573;
wire net_7434;
wire net_6960;
wire net_8960;
wire net_18050;
wire net_1710;
wire net_10994;
wire net_20065;
wire net_9017;
wire net_11456;
wire net_14274;
wire net_22426;
wire net_11922;
wire net_19612;
wire net_11443;
wire net_15742;
wire net_10524;
wire net_18192;
wire net_18619;
wire net_17625;
wire net_5988;
wire net_6969;
wire net_4336;
wire x610;
wire net_9601;
wire net_13030;
wire net_15699;
wire net_4161;
wire net_3039;
wire net_6207;
wire net_20318;
wire net_2217;
wire net_938;
wire net_20635;
wire net_1761;
wire net_12163;
wire net_5682;
wire net_4683;
wire x2745;
wire net_21504;
wire net_183;
wire net_21587;
wire net_1440;
wire net_21594;
wire net_7330;
wire net_18424;
wire net_20975;
wire net_6539;
wire net_19594;
wire net_1011;
wire net_8792;
wire net_7040;
wire net_1355;
wire net_9902;
wire net_800;
wire net_8420;
wire net_18231;
wire net_9221;
wire net_20015;
wire net_22062;
wire net_20237;
wire net_8847;
wire net_13586;
wire net_18964;
wire net_5992;
wire net_12750;
wire net_22586;
wire net_11648;
wire net_4046;
wire net_9405;
wire net_16733;
wire net_2580;
wire net_13834;
wire net_9696;
wire net_13997;
wire net_15994;
wire net_1643;
wire net_1385;
wire net_9961;
wire net_13302;
wire net_19119;
wire net_1534;
wire net_1919;
wire net_15029;
wire net_9836;
wire net_20837;
wire net_19007;
wire net_12843;
wire net_8992;
wire net_14162;
wire net_21144;
wire net_4876;
wire net_18566;
wire net_16234;
wire net_659;
wire net_9087;
wire net_14860;
wire net_8993;
wire net_14652;
wire net_19585;
wire net_899;
wire net_1010;
wire net_21358;
wire net_19150;
wire net_10224;
wire net_18873;
wire net_3654;
wire net_13883;
wire net_10139;
wire x1044;
wire net_15542;
wire net_15082;
wire net_18579;
wire net_19615;
wire net_2908;
wire net_14830;
wire net_4981;
wire net_14566;
wire x3491;
wire net_15020;
wire net_16083;
wire net_22105;
wire net_13594;
wire net_13780;
wire net_14576;
wire net_13813;
wire net_4449;
wire net_16720;
wire net_7339;
wire net_6458;
wire net_11929;
wire net_2675;
wire net_2794;
wire net_13528;
wire net_13567;
wire net_6986;
wire net_16633;
wire net_1752;
wire net_2527;
wire net_20477;
wire net_11906;
wire net_2091;
wire net_14478;
wire net_17594;
wire net_2406;
wire net_6289;
wire net_8722;
wire net_17157;
wire x6832;
wire net_19197;
wire net_18397;
wire net_807;
wire net_20830;
wire net_3405;
wire net_3270;
wire net_12422;
wire net_15456;
wire net_19270;
wire net_12665;
wire net_6880;
wire net_10238;
wire net_22407;
wire net_2474;
wire net_13931;
wire net_2530;
wire net_22798;
wire net_11578;
wire net_15824;
wire net_9472;
wire net_21825;
wire net_21000;
wire net_6192;
wire net_217;
wire net_7679;
wire net_18070;
wire net_14935;
wire net_22311;
wire net_5336;
wire net_12086;
wire net_915;
wire net_8844;
wire net_5634;
wire net_2226;
wire net_3849;
wire net_19190;
wire net_17016;
wire net_8099;
wire net_20866;
wire net_8909;
wire net_18637;
wire net_8028;
wire net_17306;
wire net_14700;
wire net_15479;
wire net_8369;
wire net_2863;
wire net_3507;
wire net_1165;
wire net_5167;
wire net_677;
wire net_1472;
wire net_20578;
wire net_18727;
wire net_2939;
wire net_20515;
wire net_1113;
wire net_13294;
wire net_20045;
wire net_9945;
wire net_17894;
wire net_11208;
wire net_11619;
wire net_15316;
wire net_21681;
wire net_18442;
wire net_7464;
wire net_8362;
wire net_11040;
wire net_22828;
wire net_22047;
wire net_5120;
wire net_15197;
wire net_14969;
wire net_5948;
wire net_5676;
wire net_15484;
wire net_8357;
wire net_2658;
wire net_2174;
wire net_14875;
wire net_784;
wire net_21672;
wire net_16460;
wire net_45;
wire net_8481;
wire net_21164;
wire net_8751;
wire net_6021;
wire net_18173;
wire net_20009;
wire net_2326;
wire net_11566;
wire net_3540;
wire net_8094;
wire net_11234;
wire x6740;
wire net_5375;
wire net_9489;
wire net_18431;
wire net_12078;
wire net_19036;
wire net_17125;
wire net_1318;
wire net_3238;
wire net_10677;
wire net_21262;
wire net_15227;
wire net_15486;
wire net_16480;
wire net_19710;
wire net_7155;
wire net_4349;
wire net_3575;
wire net_11195;
wire net_8023;
wire net_18240;
wire net_6440;
wire net_15039;
wire net_4984;
wire net_306;
wire net_18127;
wire net_4516;
wire net_5371;
wire net_9026;
wire net_5061;
wire net_6471;
wire net_2610;
wire net_4432;
wire net_4584;
wire net_1329;
wire net_14391;
wire net_362;
wire net_3127;
wire net_9959;
wire net_1052;
wire net_22776;
wire net_20127;
wire net_3831;
wire net_11180;
wire net_13974;
wire net_18163;
wire net_9477;
wire net_17966;
wire net_17004;
wire net_20784;
wire net_15083;
wire net_4859;
wire net_20536;
wire net_6413;
wire net_226;
wire net_18856;
wire net_18367;
wire net_7015;
wire net_9160;
wire net_16169;
wire net_2887;
wire net_4207;
wire net_15515;
wire net_21333;
wire net_19912;
wire net_7741;
wire net_19124;
wire net_1983;
wire net_8735;
wire net_10129;
wire net_10248;
wire net_3030;
wire net_10251;
wire net_20118;
wire net_3842;
wire net_15433;
wire net_4266;
wire net_20700;
wire net_1553;
wire net_13421;
wire net_2491;
wire net_8819;
wire net_10563;
wire net_3208;
wire net_2704;
wire net_10933;
wire net_15591;
wire net_5819;
wire net_14663;
wire net_3910;
wire net_1851;
wire net_21444;
wire net_13684;
wire net_3445;
wire net_10976;
wire net_18470;
wire net_8709;
wire net_2941;
wire net_477;
wire net_3348;
wire net_17368;
wire net_2943;
wire net_9377;
wire net_3861;
wire net_10892;
wire net_6758;
wire net_6905;
wire net_2315;
wire net_8325;
wire net_85;
wire net_2231;
wire net_15501;
wire net_22615;
wire net_17582;
wire net_14646;
wire net_3812;
wire net_1200;
wire net_9595;
wire net_17136;
wire net_9509;
wire net_18429;
wire net_22570;
wire net_12329;
wire net_7558;
wire x1731;
wire net_11135;
wire net_11487;
wire net_13980;
wire net_16675;
wire net_3437;
wire net_19672;
wire x1808;
wire net_18391;
wire net_19266;
wire net_19024;
wire net_472;
wire net_1510;
wire net_14286;
wire net_14022;
wire net_3077;
wire net_19838;
wire net_19963;
wire net_18401;
wire net_8639;
wire net_4829;
wire net_13608;
wire net_9430;
wire net_4171;
wire net_1528;
wire net_12676;
wire net_13579;
wire net_15628;
wire net_1749;
wire net_3367;
wire net_4915;
wire net_21068;
wire net_4784;
wire net_8386;
wire net_12355;
wire net_601;
wire net_20931;
wire net_1362;
wire net_4385;
wire net_2346;
wire net_829;
wire net_9315;
wire net_13025;
wire net_12396;
wire net_2294;
wire net_11856;
wire net_13867;
wire net_4978;
wire net_14174;
wire net_2393;
wire net_18646;
wire net_3917;
wire net_15171;
wire net_8539;
wire net_8812;
wire net_3376;
wire net_13671;
wire net_7979;
wire net_16351;
wire net_13845;
wire net_14926;
wire net_21190;
wire net_22161;
wire net_15090;
wire net_17983;
wire net_17174;
wire net_7218;
wire net_5319;
wire net_22595;
wire net_11045;
wire net_6357;
wire x7042;
wire net_3750;
wire x3106;
wire net_12637;
wire net_5314;
wire x3220;
wire net_5749;
wire net_20103;
wire net_2696;
wire net_9687;
wire net_10464;
wire net_12736;
wire net_6026;
wire net_14168;
wire net_8457;
wire net_10457;
wire net_22189;
wire net_21561;
wire net_19425;
wire net_1449;
wire net_16222;
wire net_20356;
wire net_6984;
wire net_5618;
wire net_15740;
wire net_5310;
wire net_9725;
wire net_8620;
wire net_13114;
wire net_22025;
wire net_1220;
wire net_12989;
wire net_14729;
wire net_21487;
wire net_17420;
wire net_12343;
wire net_21899;
wire net_4693;
wire net_4017;
wire net_11394;
wire net_22075;
wire net_10194;
wire net_6346;
wire net_12716;
wire x833;
wire net_19679;
wire net_11781;
wire net_4945;
wire net_19406;
wire net_18046;
wire net_15097;
wire net_14208;
wire net_2334;
wire net_17213;
wire net_1367;
wire net_7943;
wire net_16644;
wire net_17531;
wire net_20987;
wire net_7960;
wire net_18817;
wire net_4079;
wire net_12104;
wire net_1371;
wire net_12542;
wire net_13511;
wire net_21619;
wire net_117;
wire net_16769;
wire net_5002;
wire net_8054;
wire net_18441;
wire net_6609;
wire net_7837;
wire net_16420;
wire net_16261;
wire net_6517;
wire net_4704;
wire net_15526;
wire net_5782;
wire net_9843;
wire net_7864;
wire net_11885;
wire net_22126;
wire net_19659;
wire net_10359;
wire net_11826;
wire net_1461;
wire net_18008;
wire net_17859;
wire net_12799;
wire net_7512;
wire net_16762;
wire net_3177;
wire net_15769;
wire net_19390;
wire net_8270;
wire net_11325;
wire x184;
wire net_10011;
wire net_12556;
wire net_14526;
wire net_20888;
wire net_7222;
wire net_9459;
wire net_15921;
wire net_19246;
wire net_8891;
wire net_10360;
wire net_10475;
wire net_437;
wire net_10568;
wire net_3573;
wire net_13208;
wire net_16926;
wire net_9861;
wire net_10390;
wire net_11477;
wire net_21278;
wire net_7371;
wire net_9071;
wire net_10855;
wire net_12498;
wire net_22483;
wire net_7140;
wire net_17113;
wire net_624;
wire net_2148;
wire net_15669;
wire net_22220;
wire net_11616;
wire net_14427;
wire net_16295;
wire net_8517;
wire net_14063;
wire net_6005;
wire net_688;
wire net_21772;
wire net_21204;
wire net_8732;
wire net_5808;
wire net_8170;
wire net_3027;
wire net_12777;
wire net_16927;
wire net_17912;
wire net_5343;
wire net_14464;
wire net_22669;
wire net_6625;
wire net_15659;
wire net_15999;
wire net_9940;
wire net_15813;
wire net_5497;
wire net_4096;
wire net_7924;
wire net_21526;
wire net_22688;
wire net_16587;
wire net_5214;
wire net_4822;
wire net_3986;
wire x771;
wire net_11754;
wire net_7482;
wire net_1243;
wire net_19064;
wire net_6839;
wire net_1660;
wire net_12035;
wire net_1484;
wire net_5864;
wire net_19821;
wire net_3667;
wire net_6566;
wire net_9949;
wire net_6041;
wire net_21244;
wire net_1635;
wire net_6779;
wire net_5027;
wire net_4840;
wire net_12697;
wire net_7133;
wire net_7523;
wire net_8828;
wire net_7174;
wire net_6871;
wire net_10306;
wire net_22638;
wire net_7020;
wire net_3002;
wire net_16241;
wire net_854;
wire net_17850;
wire net_2619;
wire net_8713;
wire net_22656;
wire net_20936;
wire net_19792;
wire net_5559;
wire net_18351;
wire net_2221;
wire net_15585;
wire net_11424;
wire net_6959;
wire net_5264;
wire net_10369;
wire net_6447;
wire net_7789;
wire net_22010;
wire net_18606;
wire net_16873;
wire net_18625;
wire net_9181;
wire net_5746;
wire net_16366;
wire net_4643;
wire net_332;
wire net_1745;
wire net_13601;
wire net_1679;
wire net_7364;
wire net_4883;
wire net_9058;
wire net_13739;
wire net_656;
wire net_5723;
wire net_4800;
wire net_8489;
wire net_18371;
wire net_17180;
wire x5605;
wire net_8935;
wire net_4284;
wire net_7027;
wire net_16316;
wire net_3113;
wire net_17033;
wire net_10924;
wire net_14157;
wire net_8826;
wire net_6816;
wire net_22770;
wire net_8614;
wire net_15974;
wire net_3969;
wire net_21322;
wire net_20169;
wire net_7232;
wire net_13266;
wire net_14768;
wire net_6602;
wire net_9873;
wire net_11164;
wire net_12615;
wire net_7688;
wire net_17732;
wire net_15198;
wire net_6162;
wire net_17765;
wire net_21737;
wire net_1698;
wire net_5897;
wire net_18756;
wire net_1017;
wire net_12391;
wire net_20525;
wire net_14309;
wire net_14379;
wire net_18722;
wire net_21931;
wire net_22368;
wire net_13334;
wire net_14293;
wire net_412;
wire net_4798;
wire net_8887;
wire net_16090;
wire net_9869;
wire net_20404;
wire net_1873;
wire net_22786;
wire net_3801;
wire net_453;
wire net_7547;
wire net_22519;
wire net_20290;
wire net_10209;
wire net_17139;
wire net_5835;
wire net_18450;
wire net_2263;
wire net_10439;
wire net_20487;
wire net_6181;
wire net_3624;
wire net_7967;
wire net_9391;
wire net_951;
wire net_2086;
wire net_11596;
wire net_21853;
wire net_21296;
wire net_17382;
wire net_4930;
wire net_18665;
wire net_21727;
wire net_17252;
wire net_16715;
wire net_12278;
wire net_12869;
wire net_7272;
wire net_20184;
wire net_7096;
wire net_8977;
wire net_12654;
wire net_19091;
wire net_18517;
wire net_10222;
wire net_14389;
wire net_10648;
wire net_12350;
wire net_12121;
wire net_21951;
wire net_2966;
wire net_15146;
wire net_19439;
wire net_1253;
wire net_13186;
wire net_21952;
wire net_2500;
wire net_9808;
wire net_10508;
wire net_17716;
wire net_13971;
wire net_22116;
wire net_3900;
wire net_21982;
wire net_13315;
wire net_19221;
wire net_15889;
wire net_3153;
wire net_22833;
wire net_16456;
wire net_6721;
wire net_5471;
wire net_5155;
wire net_19484;
wire net_3598;
wire net_16418;
wire net_3938;
wire net_8676;
wire net_7534;
wire net_11289;
wire net_15757;
wire net_9592;
wire net_18669;
wire net_20694;
wire net_1502;
wire x6404;
wire net_11282;
wire net_20966;
wire net_6596;
wire net_11065;
wire net_10329;
wire net_11306;
wire net_640;
wire net_10117;
wire net_12138;
wire net_7508;
wire net_775;
wire net_21638;
wire net_752;
wire net_10903;
wire net_18114;
wire x1005;
wire net_3716;
wire net_498;
wire net_535;
wire net_17387;
wire net_21652;
wire net_2721;
wire net_8900;
wire net_2637;
wire net_15380;
wire net_20892;
wire net_20589;
wire net_6768;
wire net_4902;
wire net_5419;
wire net_299;
wire net_12228;
wire net_18266;
wire x4815;
wire net_12894;
wire net_7413;
wire net_12387;
wire net_20918;
wire net_2024;
wire net_11755;
wire net_3254;
wire net_11549;
wire net_9569;
wire net_19058;
wire net_9779;
wire net_22308;
wire net_9040;
wire net_3725;
wire net_17809;
wire net_15569;
wire net_9111;
wire net_19400;
wire net_6088;
wire net_5857;
wire net_5041;
wire net_15161;
wire net_20944;
wire net_407;
wire net_19532;
wire net_21832;
wire net_4405;
wire net_16903;
wire net_11793;
wire net_20282;
wire net_18884;
wire net_19840;
wire net_19457;
wire net_20299;
wire net_8723;
wire net_9801;
wire net_2312;
wire net_21797;
wire net_16547;
wire net_21124;
wire net_8586;
wire net_19961;
wire net_2073;
wire net_8189;
wire net_9146;
wire net_4057;
wire net_5105;
wire net_14244;
wire net_6081;
wire net_14975;
wire net_14863;
wire x6600;
wire net_21298;
wire net_16374;
wire net_5507;
wire net_12173;
wire net_12526;
wire net_7565;
wire net_15339;
wire net_1981;
wire net_4302;
wire net_6245;
wire net_1218;
wire net_22239;
wire net_10606;
wire net_15042;
wire net_22361;
wire net_16128;
wire net_3286;
wire net_19909;
wire net_27;
wire net_11430;
wire net_15604;
wire net_1398;
wire net_12432;
wire net_13219;
wire net_10503;
wire net_4399;
wire net_19478;
wire net_8197;
wire net_6117;
wire net_1144;
wire net_8297;
wire net_19188;
wire net_16373;
wire net_17571;
wire net_10646;
wire net_2260;
wire net_2865;
wire net_3606;
wire net_9770;
wire net_17116;
wire net_702;
wire net_4328;
wire net_1477;
wire net_3195;
wire net_3210;
wire net_16013;
wire net_3318;
wire net_13221;
wire net_7800;
wire net_8188;
wire net_17674;
wire net_8122;
wire net_7571;
wire x353;
wire net_11682;
wire net_12948;
wire net_12904;
wire net_22755;
wire net_15214;
wire net_1193;
wire x4444;
wire net_12979;
wire net_9412;
wire net_1425;
wire net_17331;
wire net_17068;
wire net_8436;
wire net_10790;
wire net_22660;
wire net_20378;
wire net_1813;
wire net_10622;
wire net_18406;
wire net_10673;
wire net_7945;
wire net_17363;
wire net_12411;
wire net_22269;
wire net_983;
wire net_18992;
wire net_16651;
wire net_355;
wire net_21165;
wire net_7258;
wire net_13702;
wire net_9513;
wire net_8102;
wire net_19576;
wire net_12427;
wire net_15534;
wire net_7311;
wire net_723;
wire net_11341;
wire net_7614;
wire net_2483;
wire net_18068;
wire net_16080;
wire net_12026;
wire net_14608;
wire net_10202;
wire net_10501;
wire net_20604;
wire net_15096;
wire net_20162;
wire net_10547;
wire net_19013;
wire net_16388;
wire net_3948;
wire net_6142;
wire net_22218;
wire net_13475;
wire net_13455;
wire net_12414;
wire net_12872;
wire net_9493;
wire net_8254;
wire net_20097;
wire net_11945;
wire net_21707;
wire net_3819;
wire net_15640;
wire net_254;
wire net_1501;
wire net_22811;
wire net_3003;
wire net_12103;
wire net_574;
wire net_11375;

// Start cells
OAI21_X2 inst_1783 ( .ZN(net_14659), .A(net_13437), .B2(net_11934), .B1(net_11588) );
INV_X4 inst_17321 ( .A(net_655), .ZN(net_583) );
INV_X2 inst_18950 ( .ZN(net_5642), .A(net_5641) );
INV_X4 inst_17160 ( .A(net_8556), .ZN(net_7284) );
NOR3_X2 inst_2685 ( .ZN(net_14373), .A3(net_12578), .A1(net_12051), .A2(net_8143) );
NAND4_X2 inst_5359 ( .ZN(net_15320), .A2(net_13725), .A3(net_13438), .A1(net_12219), .A4(net_11386) );
INV_X4 inst_16895 ( .ZN(net_11311), .A(net_4430) );
INV_X4 inst_13828 ( .ZN(net_12036), .A(net_6051) );
NAND3_X2 inst_6439 ( .ZN(net_11817), .A3(net_11816), .A2(net_10178), .A1(net_8110) );
NAND4_X2 inst_5306 ( .ZN(net_19706), .A1(net_18973), .A3(net_13901), .A2(net_11008), .A4(net_5460) );
OAI21_X2 inst_2205 ( .A(net_10383), .ZN(net_8538), .B1(net_8537), .B2(net_7009) );
INV_X4 inst_17222 ( .ZN(net_7597), .A(net_733) );
NOR2_X4 inst_2858 ( .ZN(net_11769), .A2(net_8766), .A1(net_7240) );
NAND2_X2 inst_8981 ( .ZN(net_14499), .A2(net_12740), .A1(net_10920) );
NAND4_X2 inst_5488 ( .ZN(net_12288), .A1(net_12287), .A4(net_12286), .A2(net_10111), .A3(net_7647) );
INV_X2 inst_19257 ( .ZN(net_3198), .A(net_3197) );
INV_X2 inst_19173 ( .ZN(net_11260), .A(net_3822) );
AOI21_X2 inst_20505 ( .ZN(net_14637), .B1(net_14636), .B2(net_12082), .A(net_7692) );
INV_X4 inst_13926 ( .ZN(net_9578), .A(net_6871) );
INV_X4 inst_15089 ( .ZN(net_3644), .A(net_3255) );
XNOR2_X2 inst_214 ( .ZN(net_17540), .A(net_17537), .B(net_6372) );
CLKBUF_X2 inst_21381 ( .A(net_21246), .Z(net_21253) );
INV_X2 inst_19279 ( .A(net_3717), .ZN(net_2939) );
INV_X4 inst_13990 ( .A(net_9006), .ZN(net_6536) );
INV_X4 inst_18233 ( .A(net_21208), .ZN(net_15588) );
INV_X4 inst_15915 ( .ZN(net_1746), .A(net_1745) );
NAND2_X2 inst_9115 ( .ZN(net_13573), .A2(net_12377), .A1(net_9733) );
XNOR2_X2 inst_548 ( .B(net_16921), .A(net_9255), .ZN(net_723) );
CLKBUF_X2 inst_22931 ( .A(net_22644), .Z(net_22803) );
INV_X4 inst_16093 ( .ZN(net_1524), .A(net_1523) );
NOR2_X2 inst_4372 ( .A2(net_11292), .ZN(net_7221), .A1(net_5448) );
INV_X4 inst_18084 ( .A(net_21081), .ZN(net_739) );
NAND2_X4 inst_7191 ( .ZN(net_13170), .A2(net_8644), .A1(net_7860) );
INV_X4 inst_12796 ( .ZN(net_17269), .A(net_17268) );
INV_X4 inst_14747 ( .ZN(net_6962), .A(net_4080) );
NAND2_X2 inst_8488 ( .ZN(net_16960), .A2(net_16959), .A1(net_516) );
INV_X4 inst_14178 ( .ZN(net_7462), .A(net_5988) );
INV_X4 inst_17516 ( .ZN(net_4865), .A(net_1848) );
INV_X4 inst_14148 ( .ZN(net_9696), .A(net_7815) );
INV_X4 inst_13127 ( .ZN(net_15296), .A(net_14960) );
NAND3_X2 inst_6406 ( .ZN(net_11972), .A1(net_11971), .A2(net_11970), .A3(net_7932) );
CLKBUF_X2 inst_21454 ( .A(net_21325), .Z(net_21326) );
INV_X2 inst_18400 ( .A(net_16571), .ZN(net_16522) );
INV_X8 inst_12400 ( .ZN(net_174), .A(net_87) );
OR2_X2 inst_1228 ( .ZN(net_2136), .A2(net_2135), .A1(net_1431) );
NAND2_X2 inst_8913 ( .ZN(net_14969), .A2(net_13662), .A1(net_5755) );
INV_X4 inst_13185 ( .ZN(net_14232), .A(net_13634) );
NOR2_X2 inst_4221 ( .A1(net_12551), .ZN(net_6628), .A2(net_6627) );
XNOR2_X2 inst_521 ( .A(net_21210), .ZN(net_4440), .B(net_4439) );
NAND3_X2 inst_6534 ( .A1(net_20439), .ZN(net_10584), .A2(net_7571), .A3(net_4424) );
NAND3_X2 inst_5947 ( .ZN(net_14889), .A1(net_13719), .A2(net_12958), .A3(net_8550) );
NOR2_X2 inst_4473 ( .A1(net_13206), .ZN(net_7283), .A2(net_4406) );
OAI21_X2 inst_1685 ( .ZN(net_15451), .A(net_15450), .B2(net_14381), .B1(net_12407) );
OAI211_X2 inst_2511 ( .B(net_14442), .ZN(net_12460), .C2(net_10847), .A(net_7833), .C1(net_6682) );
INV_X8 inst_12320 ( .ZN(net_1344), .A(net_973) );
NAND2_X2 inst_9038 ( .A1(net_15224), .ZN(net_14060), .A2(net_11838) );
NAND2_X4 inst_6910 ( .A2(net_19295), .A1(net_19294), .ZN(net_17881) );
NOR2_X2 inst_3578 ( .ZN(net_12699), .A2(net_11014), .A1(net_8337) );
NAND2_X2 inst_9257 ( .A1(net_13605), .ZN(net_12643), .A2(net_8016) );
INV_X4 inst_15477 ( .ZN(net_6404), .A(net_1591) );
INV_X4 inst_14731 ( .ZN(net_11925), .A(net_4117) );
NAND2_X2 inst_9938 ( .ZN(net_9135), .A2(net_7095), .A1(net_6669) );
INV_X8 inst_12238 ( .ZN(net_5109), .A(net_2879) );
NAND3_X2 inst_5940 ( .ZN(net_14905), .A2(net_14904), .A1(net_14181), .A3(net_13046) );
INV_X4 inst_17892 ( .A(net_2585), .ZN(net_66) );
INV_X4 inst_18107 ( .A(net_21141), .ZN(net_726) );
INV_X4 inst_14010 ( .ZN(net_10251), .A(net_6309) );
INV_X4 inst_13236 ( .ZN(net_14825), .A(net_13469) );
AOI22_X2 inst_19978 ( .ZN(net_15482), .B1(net_15481), .A2(net_14606), .B2(net_8558), .A1(net_2434) );
NAND2_X2 inst_10825 ( .ZN(net_14933), .A2(net_5526), .A1(net_5486) );
CLKBUF_X2 inst_22829 ( .A(net_22700), .Z(net_22701) );
NOR2_X2 inst_3392 ( .ZN(net_18998), .A2(net_15834), .A1(net_15601) );
INV_X2 inst_18376 ( .ZN(net_17203), .A(net_17202) );
NAND3_X2 inst_6232 ( .ZN(net_13223), .A2(net_11161), .A3(net_11132), .A1(net_10721) );
OAI21_X2 inst_2342 ( .ZN(net_4663), .A(net_2866), .B1(net_2021), .B2(net_712) );
AOI21_X2 inst_20314 ( .ZN(net_15975), .B1(net_15864), .B2(net_15593), .A(net_9546) );
INV_X4 inst_15849 ( .ZN(net_7116), .A(net_1830) );
NAND2_X2 inst_9143 ( .ZN(net_13410), .A2(net_10509), .A1(net_1927) );
OAI21_X2 inst_1617 ( .A(net_20856), .ZN(net_16075), .B2(net_15534), .B1(net_11539) );
INV_X4 inst_12553 ( .ZN(net_18319), .A(net_18271) );
XNOR2_X2 inst_151 ( .ZN(net_17985), .A(net_17909), .B(net_17600) );
OAI21_X2 inst_2256 ( .A(net_8179), .ZN(net_7259), .B2(net_7258), .B1(net_2188) );
CLKBUF_X2 inst_22023 ( .A(net_21894), .Z(net_21895) );
AOI21_X2 inst_20440 ( .ZN(net_15125), .B2(net_13223), .A(net_13057), .B1(net_652) );
INV_X2 inst_18916 ( .ZN(net_5963), .A(net_5962) );
NAND2_X4 inst_7519 ( .A1(net_19826), .ZN(net_3024), .A2(net_129) );
NOR2_X2 inst_4880 ( .ZN(net_4975), .A1(net_2183), .A2(net_2164) );
NAND2_X2 inst_11637 ( .A2(net_7676), .ZN(net_2513), .A1(net_836) );
NAND2_X2 inst_10370 ( .ZN(net_7400), .A1(net_7399), .A2(net_4540) );
NOR2_X2 inst_3867 ( .A2(net_9397), .ZN(net_9377), .A1(net_5033) );
OAI21_X2 inst_2072 ( .B1(net_13355), .A(net_12226), .ZN(net_10601), .B2(net_5279) );
OAI21_X2 inst_1603 ( .ZN(net_16154), .B2(net_15730), .B1(net_12941), .A(net_1850) );
NAND2_X2 inst_9634 ( .ZN(net_11690), .A1(net_10405), .A2(net_8358) );
XNOR2_X2 inst_340 ( .ZN(net_16964), .B(net_16648), .A(net_16451) );
INV_X4 inst_18322 ( .ZN(net_20536), .A(net_20529) );
INV_X4 inst_14978 ( .ZN(net_5945), .A(net_3416) );
NAND2_X2 inst_8109 ( .A2(net_20443), .ZN(net_19206), .A1(net_17029) );
NAND2_X2 inst_11075 ( .ZN(net_11164), .A1(net_4478), .A2(net_3506) );
NOR2_X2 inst_4280 ( .ZN(net_9597), .A2(net_6100), .A1(net_5866) );
NAND2_X2 inst_8171 ( .ZN(net_17954), .A1(net_17901), .A2(net_17803) );
NAND2_X4 inst_7493 ( .ZN(net_3879), .A1(net_3350), .A2(net_2315) );
NAND4_X2 inst_5411 ( .ZN(net_14588), .A1(net_12429), .A3(net_11435), .A2(net_11171), .A4(net_9996) );
INV_X2 inst_18543 ( .A(net_11705), .ZN(net_10984) );
INV_X4 inst_14279 ( .A(net_5719), .ZN(net_5653) );
NOR2_X2 inst_4244 ( .ZN(net_11295), .A2(net_4654), .A1(net_2985) );
CLKBUF_X2 inst_22354 ( .A(net_22225), .Z(net_22226) );
OAI21_X4 inst_1490 ( .ZN(net_20459), .A(net_13080), .B1(net_9627), .B2(net_9539) );
CLKBUF_X2 inst_22460 ( .A(net_21899), .Z(net_22332) );
AND2_X4 inst_21223 ( .A2(net_12915), .A1(net_8991), .ZN(net_8641) );
INV_X4 inst_15421 ( .A(net_16051), .ZN(net_15971) );
NOR2_X2 inst_4559 ( .A1(net_11296), .A2(net_8714), .ZN(net_5532) );
NOR2_X2 inst_3709 ( .ZN(net_11035), .A2(net_11034), .A1(net_9161) );
NAND2_X2 inst_10934 ( .A1(net_11893), .ZN(net_8415), .A2(net_5209) );
NAND3_X2 inst_6319 ( .ZN(net_12562), .A3(net_12561), .A1(net_6404), .A2(net_2098) );
SDFF_X2 inst_827 ( .Q(net_21189), .SI(net_17546), .SE(net_945), .CK(net_22324), .D(x6381) );
INV_X2 inst_18560 ( .ZN(net_10799), .A(net_10798) );
INV_X4 inst_15309 ( .ZN(net_14078), .A(net_7295) );
NAND2_X2 inst_11477 ( .ZN(net_4071), .A2(net_2453), .A1(net_36) );
INV_X4 inst_17498 ( .ZN(net_6788), .A(net_693) );
NAND2_X2 inst_9573 ( .ZN(net_10955), .A2(net_6213), .A1(net_3805) );
INV_X4 inst_15231 ( .ZN(net_4319), .A(net_2839) );
NAND2_X2 inst_10730 ( .ZN(net_5827), .A1(net_4470), .A2(net_3428) );
NAND2_X2 inst_10574 ( .ZN(net_6693), .A1(net_6692), .A2(net_4948) );
NAND2_X4 inst_7140 ( .ZN(net_12737), .A2(net_9812), .A1(net_9785) );
NOR2_X4 inst_3040 ( .ZN(net_5098), .A1(net_4409), .A2(net_733) );
AOI211_X2 inst_21011 ( .ZN(net_19494), .C1(net_15688), .C2(net_15030), .B(net_14957), .A(net_6529) );
INV_X4 inst_12937 ( .ZN(net_17485), .A(net_16985) );
NOR2_X2 inst_3870 ( .A1(net_11365), .ZN(net_9370), .A2(net_7866) );
INV_X4 inst_16707 ( .ZN(net_15501), .A(net_12275) );
NAND3_X2 inst_5675 ( .ZN(net_20227), .A3(net_16154), .A2(net_15288), .A1(net_11732) );
AND2_X4 inst_21155 ( .A1(net_15457), .ZN(net_14304), .A2(net_14298) );
INV_X4 inst_17052 ( .ZN(net_10447), .A(net_6668) );
NOR2_X2 inst_4640 ( .ZN(net_3411), .A1(net_3410), .A2(net_1572) );
XOR2_X2 inst_18 ( .A(net_21144), .Z(net_16980), .B(net_16979) );
NAND3_X2 inst_6047 ( .ZN(net_19814), .A3(net_14215), .A2(net_12364), .A1(net_8605) );
AOI21_X2 inst_20952 ( .A(net_21238), .ZN(net_5368), .B2(net_5367), .B1(net_1974) );
NOR2_X2 inst_4128 ( .A2(net_10630), .ZN(net_6964), .A1(net_6963) );
NAND2_X2 inst_9040 ( .ZN(net_14058), .A1(net_12877), .A2(net_12037) );
NAND2_X2 inst_10154 ( .ZN(net_8270), .A2(net_6310), .A1(net_1670) );
NOR2_X2 inst_4861 ( .A1(net_8241), .ZN(net_3734), .A2(net_2258) );
NAND4_X4 inst_5183 ( .A4(net_18957), .A1(net_18956), .ZN(net_17330), .A3(net_14955), .A2(net_12167) );
AOI211_X2 inst_21023 ( .ZN(net_14884), .B(net_13598), .C2(net_11492), .A(net_6726), .C1(net_5759) );
NOR2_X2 inst_3936 ( .ZN(net_8699), .A2(net_8625), .A1(net_6892) );
INV_X4 inst_13738 ( .ZN(net_9234), .A(net_7646) );
INV_X4 inst_17866 ( .A(net_108), .ZN(net_88) );
NAND3_X2 inst_6069 ( .ZN(net_14127), .A3(net_10707), .A1(net_9826), .A2(net_9475) );
INV_X4 inst_17612 ( .A(net_1790), .ZN(net_388) );
NAND3_X2 inst_6675 ( .ZN(net_7758), .A1(net_6265), .A2(net_5914), .A3(net_5445) );
NAND3_X2 inst_6020 ( .ZN(net_14382), .A3(net_13159), .A2(net_12369), .A1(net_5697) );
CLKBUF_X2 inst_22803 ( .A(net_21359), .Z(net_22675) );
INV_X4 inst_12739 ( .ZN(net_17444), .A(net_17443) );
INV_X4 inst_14663 ( .ZN(net_5599), .A(net_4336) );
CLKBUF_X2 inst_22346 ( .A(net_22217), .Z(net_22218) );
NAND2_X2 inst_9217 ( .A1(net_13367), .ZN(net_12986), .A2(net_8855) );
NAND3_X2 inst_6475 ( .ZN(net_11286), .A3(net_11285), .A2(net_7590), .A1(net_3313) );
NAND2_X4 inst_7364 ( .ZN(net_10442), .A1(net_6394), .A2(net_5743) );
NAND3_X2 inst_5816 ( .ZN(net_15620), .A2(net_15211), .A3(net_14504), .A1(net_6923) );
INV_X4 inst_18259 ( .A(net_20903), .ZN(net_163) );
NOR3_X2 inst_2695 ( .ZN(net_14098), .A3(net_10463), .A2(net_8482), .A1(net_7307) );
INV_X4 inst_13801 ( .ZN(net_9190), .A(net_7552) );
INV_X4 inst_18158 ( .A(net_21080), .ZN(net_440) );
AOI21_X4 inst_20230 ( .B1(net_20036), .ZN(net_13477), .B2(net_10759), .A(net_6036) );
INV_X4 inst_14833 ( .A(net_13651), .ZN(net_3870) );
INV_X4 inst_12515 ( .ZN(net_19057), .A(net_18598) );
INV_X4 inst_13635 ( .ZN(net_8214), .A(net_8213) );
INV_X4 inst_14980 ( .ZN(net_8448), .A(net_5351) );
AOI21_X2 inst_20365 ( .ZN(net_15638), .B2(net_14432), .A(net_11851), .B1(net_2488) );
NAND2_X2 inst_10692 ( .ZN(net_6082), .A1(net_6081), .A2(net_4594) );
INV_X4 inst_14150 ( .ZN(net_7495), .A(net_6045) );
CLKBUF_X2 inst_22944 ( .A(net_22815), .Z(net_22816) );
INV_X4 inst_13228 ( .ZN(net_13522), .A(net_12514) );
NOR2_X2 inst_3521 ( .ZN(net_13751), .A1(net_13578), .A2(net_5771) );
NAND2_X2 inst_8969 ( .ZN(net_19169), .A2(net_12892), .A1(net_2355) );
NOR2_X2 inst_3440 ( .ZN(net_19014), .A2(net_14543), .A1(net_11569) );
AOI22_X2 inst_19992 ( .ZN(net_14735), .B1(net_14734), .A1(net_13517), .A2(net_12234), .B2(net_9962) );
NAND3_X2 inst_5802 ( .ZN(net_15705), .A3(net_14982), .A2(net_13279), .A1(net_13094) );
CLKBUF_X2 inst_22064 ( .A(net_21935), .Z(net_21936) );
NOR2_X2 inst_4001 ( .ZN(net_8177), .A1(net_6298), .A2(net_3874) );
INV_X2 inst_19492 ( .A(net_8851), .ZN(net_1297) );
INV_X8 inst_12249 ( .A(net_3797), .ZN(net_2621) );
NAND2_X2 inst_7897 ( .ZN(net_18485), .A2(net_18386), .A1(net_17813) );
NAND2_X2 inst_9188 ( .ZN(net_20387), .A1(net_13128), .A2(net_13127) );
NAND3_X2 inst_6184 ( .A2(net_20314), .A1(net_20313), .ZN(net_20240), .A3(net_3728) );
NAND2_X2 inst_10958 ( .A2(net_19461), .ZN(net_5078), .A1(net_3350) );
CLKBUF_X2 inst_22738 ( .A(net_22609), .Z(net_22610) );
INV_X2 inst_18869 ( .A(net_8351), .ZN(net_6279) );
INV_X4 inst_14388 ( .ZN(net_8318), .A(net_5140) );
INV_X4 inst_14922 ( .A(net_14515), .ZN(net_14075) );
NAND2_X2 inst_10106 ( .ZN(net_8443), .A1(net_5548), .A2(net_5396) );
SDFF_X2 inst_1027 ( .QN(net_21071), .D(net_489), .SE(net_263), .CK(net_21707), .SI(x1891) );
NAND2_X2 inst_8432 ( .A1(net_17441), .ZN(net_17176), .A2(net_17175) );
OR2_X2 inst_1143 ( .ZN(net_11112), .A2(net_10407), .A1(net_8330) );
NAND2_X2 inst_11336 ( .A1(net_9843), .ZN(net_3694), .A2(net_2960) );
AND2_X2 inst_21351 ( .ZN(net_2194), .A1(net_2193), .A2(net_2192) );
CLKBUF_X2 inst_21913 ( .A(net_21784), .Z(net_21785) );
NAND2_X2 inst_12024 ( .ZN(net_1664), .A2(net_1025), .A1(net_61) );
NAND2_X2 inst_10457 ( .ZN(net_7027), .A1(net_7026), .A2(net_7025) );
INV_X4 inst_12679 ( .ZN(net_17731), .A(net_17730) );
NAND2_X2 inst_11824 ( .ZN(net_2377), .A1(net_1790), .A2(net_1789) );
NAND2_X2 inst_8503 ( .ZN(net_17058), .A2(net_16598), .A1(net_16463) );
AND2_X4 inst_21242 ( .ZN(net_2843), .A2(net_2842), .A1(net_1870) );
INV_X2 inst_18874 ( .ZN(net_12574), .A(net_7900) );
NOR2_X2 inst_4147 ( .A2(net_8442), .A1(net_6990), .ZN(net_6909) );
OAI21_X2 inst_1538 ( .ZN(net_17910), .A(net_17716), .B2(net_17715), .B1(net_17046) );
INV_X4 inst_15273 ( .ZN(net_2758), .A(net_2631) );
NAND2_X2 inst_10349 ( .ZN(net_7504), .A2(net_7503), .A1(net_5551) );
INV_X4 inst_12525 ( .ZN(net_18462), .A(net_18461) );
NAND3_X2 inst_6465 ( .ZN(net_11361), .A3(net_10629), .A2(net_10619), .A1(net_3798) );
NAND3_X2 inst_6312 ( .ZN(net_12747), .A3(net_12746), .A2(net_4895), .A1(net_3925) );
OAI21_X2 inst_2179 ( .B2(net_20225), .ZN(net_19350), .B1(net_9801), .A(net_6635) );
AOI21_X2 inst_20561 ( .ZN(net_14253), .A(net_14009), .B1(net_12242), .B2(net_7999) );
OAI211_X2 inst_2578 ( .ZN(net_7685), .B(net_7669), .C1(net_5201), .C2(net_4959), .A(net_3198) );
NAND2_X4 inst_7514 ( .ZN(net_2138), .A2(net_2137), .A1(net_2058) );
OAI21_X2 inst_1996 ( .ZN(net_11905), .B2(net_11832), .B1(net_10279), .A(net_7053) );
AOI21_X4 inst_20185 ( .ZN(net_15252), .A(net_14159), .B1(net_13555), .B2(net_13463) );
INV_X4 inst_12838 ( .ZN(net_17250), .A(net_17146) );
NOR2_X2 inst_3340 ( .ZN(net_20692), .A2(net_18823), .A1(net_17163) );
NOR2_X2 inst_4683 ( .ZN(net_3831), .A1(net_3201), .A2(net_1857) );
INV_X4 inst_17414 ( .ZN(net_773), .A(net_507) );
CLKBUF_X2 inst_22421 ( .A(x7698), .Z(net_22293) );
AOI21_X2 inst_20634 ( .ZN(net_19808), .B2(net_19589), .B1(net_19588), .A(net_696) );
OAI21_X4 inst_1380 ( .B2(net_20123), .B1(net_20122), .ZN(net_18969), .A(net_16368) );
INV_X4 inst_15890 ( .ZN(net_9418), .A(net_4457) );
CLKBUF_X2 inst_22672 ( .A(net_21271), .Z(net_22544) );
NOR2_X2 inst_3891 ( .ZN(net_9232), .A2(net_5322), .A1(net_1342) );
NAND2_X2 inst_11298 ( .A1(net_3886), .ZN(net_3793), .A2(net_2945) );
INV_X4 inst_12484 ( .ZN(net_18679), .A(net_18678) );
NAND2_X2 inst_8318 ( .ZN(net_17636), .A2(net_17343), .A1(net_17226) );
INV_X2 inst_19643 ( .ZN(net_19439), .A(net_2479) );
INV_X4 inst_17924 ( .A(net_20922), .ZN(net_146) );
NOR2_X2 inst_4834 ( .ZN(net_7140), .A2(net_3393), .A1(net_1775) );
NOR2_X2 inst_3472 ( .ZN(net_14455), .A1(net_14454), .A2(net_12776) );
NAND2_X2 inst_8736 ( .A1(net_16385), .ZN(net_16026), .A2(net_15719) );
NAND2_X2 inst_9933 ( .ZN(net_19850), .A1(net_8029), .A2(net_7152) );
INV_X2 inst_19402 ( .ZN(net_3530), .A(net_2011) );
CLKBUF_X2 inst_22532 ( .A(net_22403), .Z(net_22404) );
CLKBUF_X2 inst_21906 ( .A(net_21488), .Z(net_21778) );
OAI21_X2 inst_2322 ( .ZN(net_5663), .A(net_5299), .B1(net_4259), .B2(net_1968) );
XNOR2_X2 inst_513 ( .A(net_21185), .ZN(net_5793), .B(net_5792) );
INV_X4 inst_17725 ( .ZN(net_3201), .A(net_196) );
INV_X4 inst_14340 ( .ZN(net_7851), .A(net_5375) );
OAI21_X2 inst_1630 ( .A(net_16395), .ZN(net_16022), .B2(net_15415), .B1(net_14774) );
OAI21_X2 inst_1586 ( .A(net_20960), .ZN(net_16262), .B2(net_15930), .B1(net_12584) );
INV_X4 inst_16624 ( .ZN(net_2252), .A(net_974) );
NAND2_X2 inst_9318 ( .A1(net_13512), .ZN(net_12343), .A2(net_12342) );
INV_X2 inst_18584 ( .ZN(net_10289), .A(net_10288) );
CLKBUF_X2 inst_21517 ( .A(net_21388), .Z(net_21389) );
CLKBUF_X2 inst_22689 ( .A(net_22560), .Z(net_22561) );
INV_X4 inst_13954 ( .A(net_12805), .ZN(net_6757) );
NAND3_X2 inst_6083 ( .ZN(net_20699), .A3(net_11154), .A1(net_7039), .A2(net_3545) );
NOR2_X2 inst_4256 ( .A1(net_6433), .ZN(net_6324), .A2(net_6323) );
INV_X2 inst_18416 ( .ZN(net_15838), .A(net_15672) );
NAND2_X2 inst_10773 ( .ZN(net_5622), .A1(net_5621), .A2(net_4257) );
AOI21_X2 inst_20386 ( .ZN(net_15490), .B2(net_14580), .A(net_13975), .B1(net_828) );
INV_X2 inst_18556 ( .ZN(net_20349), .A(net_10882) );
OAI21_X2 inst_1508 ( .B2(net_20692), .B1(net_20691), .ZN(net_18866), .A(net_18582) );
OR2_X2 inst_1222 ( .ZN(net_5376), .A2(net_2986), .A1(net_1790) );
NAND2_X2 inst_9151 ( .ZN(net_13397), .A1(net_12401), .A2(net_10585) );
NAND2_X2 inst_11366 ( .ZN(net_6098), .A2(net_3590), .A1(net_1501) );
NOR2_X2 inst_3407 ( .ZN(net_15767), .A2(net_15243), .A1(net_13575) );
OR2_X4 inst_1073 ( .ZN(net_13747), .A1(net_10445), .A2(net_8333) );
OAI21_X2 inst_2323 ( .ZN(net_5654), .A(net_2545), .B1(net_2288), .B2(net_1167) );
NOR2_X2 inst_3741 ( .ZN(net_19728), .A1(net_8737), .A2(net_7332) );
INV_X4 inst_14643 ( .ZN(net_6088), .A(net_2956) );
OAI21_X4 inst_1449 ( .ZN(net_20224), .B2(net_19360), .B1(net_19359), .A(net_15690) );
DFF_X1 inst_19884 ( .D(net_17114), .CK(net_21750), .Q(x90) );
NAND3_X2 inst_5657 ( .ZN(net_17000), .A2(net_16349), .A3(net_16283), .A1(net_12856) );
NAND2_X2 inst_11614 ( .ZN(net_5315), .A1(net_3368), .A2(net_2595) );
NAND2_X2 inst_7872 ( .ZN(net_18544), .A1(net_18468), .A2(net_17758) );
XNOR2_X2 inst_187 ( .B(net_18211), .ZN(net_17757), .A(net_17334) );
XNOR2_X2 inst_206 ( .B(net_21184), .ZN(net_17579), .A(net_17578) );
INV_X4 inst_16449 ( .ZN(net_9768), .A(net_1229) );
NOR2_X2 inst_3739 ( .ZN(net_10698), .A2(net_8447), .A1(net_2407) );
XNOR2_X2 inst_405 ( .ZN(net_16651), .A(net_16650), .B(net_1677) );
NAND3_X2 inst_6436 ( .ZN(net_11829), .A2(net_11828), .A3(net_10503), .A1(net_6938) );
NOR2_X2 inst_4788 ( .ZN(net_5091), .A2(net_2011), .A1(net_85) );
NAND2_X2 inst_10505 ( .ZN(net_8258), .A2(net_6908), .A1(net_1197) );
NAND3_X2 inst_6166 ( .ZN(net_13633), .A3(net_13632), .A2(net_13605), .A1(net_10931) );
INV_X4 inst_17734 ( .ZN(net_10319), .A(net_6078) );
INV_X4 inst_12833 ( .A(net_17416), .ZN(net_17415) );
INV_X4 inst_15868 ( .ZN(net_1801), .A(net_1393) );
NAND3_X2 inst_6776 ( .ZN(net_4513), .A2(net_4512), .A3(net_4511), .A1(net_2544) );
INV_X4 inst_13087 ( .ZN(net_19275), .A(net_15912) );
NAND3_X2 inst_5645 ( .A3(net_19124), .A1(net_19123), .ZN(net_17339), .A2(net_16269) );
INV_X4 inst_18140 ( .A(net_21139), .ZN(net_557) );
INV_X4 inst_13046 ( .ZN(net_16423), .A(net_16393) );
OAI21_X2 inst_2176 ( .A(net_10066), .ZN(net_8873), .B2(net_5007), .B1(net_4098) );
NOR2_X4 inst_2892 ( .A1(net_19319), .ZN(net_10941), .A2(net_9458) );
NAND3_X2 inst_6339 ( .ZN(net_12274), .A2(net_12273), .A3(net_9386), .A1(net_9015) );
INV_X4 inst_13024 ( .A(net_16476), .ZN(net_16416) );
INV_X2 inst_19027 ( .A(net_4923), .ZN(net_4922) );
CLKBUF_X2 inst_22368 ( .A(net_22239), .Z(net_22240) );
INV_X4 inst_18001 ( .A(net_21054), .ZN(net_509) );
CLKBUF_X2 inst_22124 ( .A(net_21809), .Z(net_21996) );
INV_X4 inst_14929 ( .ZN(net_4436), .A(net_3552) );
INV_X4 inst_15082 ( .ZN(net_3624), .A(net_3264) );
NAND2_X2 inst_11663 ( .ZN(net_8384), .A1(net_3988), .A2(net_2337) );
NAND2_X2 inst_7804 ( .ZN(net_18695), .A2(net_18662), .A1(net_18646) );
INV_X4 inst_14968 ( .ZN(net_19784), .A(net_5042) );
NAND2_X2 inst_9795 ( .ZN(net_14237), .A1(net_13375), .A2(net_9710) );
NAND4_X2 inst_5365 ( .A4(net_19789), .A1(net_19788), .ZN(net_19320), .A3(net_13265), .A2(net_13087) );
INV_X4 inst_15889 ( .ZN(net_11345), .A(net_9733) );
OAI211_X2 inst_2482 ( .ZN(net_13484), .B(net_13483), .C2(net_12454), .A(net_10743), .C1(net_4386) );
NOR2_X4 inst_2957 ( .ZN(net_12147), .A2(net_9571), .A1(net_6807) );
INV_X4 inst_15606 ( .ZN(net_3268), .A(net_3109) );
NAND2_X2 inst_10880 ( .ZN(net_7305), .A1(net_5414), .A2(net_5270) );
INV_X4 inst_15551 ( .A(net_2520), .ZN(net_2341) );
NOR3_X2 inst_2711 ( .ZN(net_13642), .A3(net_13641), .A1(net_11570), .A2(net_9905) );
INV_X4 inst_12808 ( .ZN(net_17472), .A(net_17348) );
NOR2_X2 inst_3531 ( .ZN(net_13559), .A2(net_12271), .A1(net_2423) );
NOR3_X2 inst_2753 ( .ZN(net_11814), .A2(net_11813), .A1(net_8819), .A3(net_7982) );
INV_X4 inst_16525 ( .ZN(net_2961), .A(net_1181) );
NOR2_X2 inst_3672 ( .ZN(net_19011), .A2(net_11150), .A1(net_9177) );
INV_X4 inst_14329 ( .ZN(net_8945), .A(net_5421) );
INV_X4 inst_16329 ( .ZN(net_1770), .A(net_1309) );
XNOR2_X2 inst_132 ( .ZN(net_18234), .A(net_18157), .B(net_16798) );
CLKBUF_X2 inst_22277 ( .A(net_21916), .Z(net_22149) );
INV_X2 inst_18927 ( .ZN(net_5905), .A(net_5904) );
INV_X4 inst_15484 ( .ZN(net_4361), .A(net_2031) );
NAND2_X2 inst_10353 ( .ZN(net_7471), .A1(net_7449), .A2(net_3279) );
INV_X4 inst_13900 ( .ZN(net_7965), .A(net_5429) );
NAND2_X2 inst_11502 ( .ZN(net_3066), .A2(net_2860), .A1(net_2663) );
INV_X4 inst_17092 ( .ZN(net_1074), .A(net_802) );
INV_X4 inst_12619 ( .ZN(net_18012), .A(net_18011) );
INV_X4 inst_17000 ( .ZN(net_1608), .A(net_870) );
NAND2_X2 inst_10369 ( .ZN(net_7402), .A2(net_7401), .A1(net_5576) );
NAND2_X2 inst_7935 ( .ZN(net_18433), .A2(net_18321), .A1(net_18274) );
NAND3_X2 inst_6149 ( .ZN(net_13682), .A1(net_12531), .A2(net_10781), .A3(net_8665) );
NOR2_X2 inst_3545 ( .ZN(net_13123), .A2(net_10199), .A1(net_8783) );
CLKBUF_X2 inst_21889 ( .A(net_21760), .Z(net_21761) );
INV_X4 inst_16982 ( .ZN(net_885), .A(net_420) );
INV_X4 inst_15681 ( .ZN(net_4188), .A(net_1498) );
NOR2_X2 inst_3611 ( .ZN(net_12397), .A2(net_12396), .A1(net_10726) );
INV_X4 inst_12612 ( .ZN(net_18084), .A(net_18079) );
AOI21_X2 inst_20917 ( .B2(net_9913), .ZN(net_7312), .B1(net_1920), .A(net_948) );
INV_X4 inst_16964 ( .ZN(net_1228), .A(net_222) );
INV_X2 inst_18476 ( .ZN(net_12632), .A(net_12631) );
CLKBUF_X2 inst_22554 ( .A(net_22425), .Z(net_22426) );
AND2_X2 inst_21322 ( .A2(net_10429), .ZN(net_6785), .A1(net_6784) );
CLKBUF_X2 inst_22926 ( .A(net_22797), .Z(net_22798) );
INV_X4 inst_17968 ( .A(net_20947), .ZN(net_154) );
INV_X4 inst_15083 ( .ZN(net_5792), .A(net_3262) );
NOR2_X2 inst_3975 ( .A2(net_9971), .ZN(net_8401), .A1(net_5618) );
CLKBUF_X2 inst_21628 ( .A(net_21428), .Z(net_21500) );
NAND2_X2 inst_11025 ( .A1(net_9984), .ZN(net_4786), .A2(net_4785) );
NAND2_X2 inst_10976 ( .ZN(net_6566), .A2(net_3537), .A1(net_1376) );
XNOR2_X2 inst_327 ( .B(net_21210), .ZN(net_17023), .A(net_17022) );
CLKBUF_X2 inst_21589 ( .A(net_21248), .Z(net_21461) );
NAND2_X2 inst_8874 ( .ZN(net_15254), .A2(net_14742), .A1(net_2547) );
NAND2_X2 inst_7801 ( .ZN(net_18699), .A2(net_18672), .A1(net_16876) );
AOI21_X2 inst_20900 ( .B2(net_20576), .A(net_9516), .ZN(net_7719), .B1(net_2162) );
AOI21_X2 inst_20931 ( .B1(net_9461), .ZN(net_7069), .B2(net_4297), .A(net_2122) );
NAND2_X2 inst_9431 ( .ZN(net_11604), .A1(net_11603), .A2(net_11602) );
NOR2_X2 inst_3853 ( .ZN(net_10960), .A2(net_7553), .A1(net_7115) );
NAND2_X2 inst_8044 ( .ZN(net_18235), .A2(net_18223), .A1(net_17490) );
INV_X4 inst_15132 ( .ZN(net_5605), .A(net_3127) );
NAND3_X2 inst_6702 ( .A2(net_12409), .A3(net_11995), .ZN(net_7359), .A1(net_2040) );
INV_X4 inst_14304 ( .ZN(net_6015), .A(net_5520) );
INV_X8 inst_12421 ( .A(net_20931), .ZN(net_703) );
NAND2_X2 inst_7905 ( .ZN(net_18476), .A2(net_18398), .A1(net_18334) );
CLKBUF_X2 inst_21566 ( .A(net_21437), .Z(net_21438) );
INV_X4 inst_17415 ( .ZN(net_1242), .A(net_1025) );
NAND2_X2 inst_10739 ( .A1(net_8205), .ZN(net_5747), .A2(net_4227) );
NOR2_X2 inst_3661 ( .ZN(net_20030), .A2(net_11593), .A1(net_9999) );
INV_X4 inst_16758 ( .ZN(net_18003), .A(net_2524) );
INV_X4 inst_13678 ( .A(net_8710), .ZN(net_8000) );
INV_X4 inst_14244 ( .A(net_9236), .ZN(net_7341) );
INV_X4 inst_15963 ( .ZN(net_12884), .A(net_9968) );
NAND2_X2 inst_9001 ( .ZN(net_14287), .A2(net_13484), .A1(net_11651) );
NAND2_X2 inst_11836 ( .ZN(net_7663), .A1(net_1747), .A2(net_225) );
AOI21_X4 inst_20180 ( .B1(net_19621), .ZN(net_15394), .B2(net_15121), .A(net_12850) );
NOR2_X4 inst_3221 ( .ZN(net_5515), .A1(net_2636), .A2(net_2265) );
INV_X4 inst_16251 ( .ZN(net_2535), .A(net_1346) );
INV_X4 inst_14585 ( .A(net_8500), .ZN(net_4487) );
INV_X4 inst_16209 ( .ZN(net_14367), .A(net_10398) );
INV_X8 inst_12335 ( .A(net_1192), .ZN(net_1159) );
XNOR2_X2 inst_357 ( .ZN(net_16890), .A(net_16504), .B(net_551) );
NAND2_X2 inst_11083 ( .ZN(net_8571), .A1(net_4430), .A2(net_4429) );
NAND2_X4 inst_6969 ( .A2(net_20232), .A1(net_20231), .ZN(net_17411) );
NAND2_X2 inst_10028 ( .ZN(net_19981), .A2(net_10523), .A1(net_8744) );
DFF_X1 inst_19915 ( .D(net_16625), .CK(net_21806), .Q(x1159) );
NAND3_X2 inst_6173 ( .ZN(net_13550), .A3(net_9214), .A2(net_6011), .A1(net_5164) );
NOR2_X2 inst_4092 ( .A1(net_10765), .A2(net_9045), .ZN(net_8729) );
INV_X4 inst_13865 ( .A(net_12968), .ZN(net_7453) );
NAND2_X2 inst_10098 ( .ZN(net_14596), .A2(net_8649), .A1(net_8618) );
NOR2_X2 inst_3980 ( .ZN(net_8387), .A2(net_7151), .A1(net_5515) );
CLKBUF_X2 inst_22879 ( .A(net_22750), .Z(net_22751) );
DFF_X1 inst_19889 ( .D(net_16981), .CK(net_22790), .Q(x1275) );
NAND2_X2 inst_11438 ( .ZN(net_4391), .A2(net_3118), .A1(net_454) );
NOR2_X2 inst_3758 ( .ZN(net_10358), .A2(net_9422), .A1(net_7320) );
SDFF_X2 inst_912 ( .Q(net_21205), .SI(net_16623), .SE(net_125), .CK(net_22413), .D(x5957) );
INV_X4 inst_18087 ( .A(net_21155), .ZN(net_16775) );
INV_X4 inst_15653 ( .A(net_2399), .ZN(net_2106) );
NAND2_X2 inst_10065 ( .A1(net_10031), .ZN(net_8671), .A2(net_8631) );
INV_X4 inst_15923 ( .ZN(net_3118), .A(net_1738) );
AOI21_X2 inst_20407 ( .ZN(net_15331), .B2(net_13683), .A(net_9088), .B1(net_1613) );
INV_X2 inst_18516 ( .ZN(net_11565), .A(net_11564) );
INV_X2 inst_18451 ( .ZN(net_14829), .A(net_13440) );
INV_X4 inst_12724 ( .A(net_17690), .ZN(net_17524) );
NAND3_X2 inst_5872 ( .A3(net_20817), .A1(net_20816), .ZN(net_15307), .A2(net_13508) );
AOI22_X2 inst_20015 ( .B1(net_20531), .A1(net_12669), .ZN(net_11734), .A2(net_11733), .B2(net_11230) );
INV_X4 inst_16735 ( .A(net_10183), .ZN(net_8020) );
NAND2_X4 inst_6988 ( .A2(net_21126), .ZN(net_20050), .A1(net_17287) );
NOR2_X2 inst_4188 ( .A2(net_8039), .ZN(net_6741), .A1(net_81) );
INV_X4 inst_14888 ( .ZN(net_6369), .A(net_2914) );
INV_X4 inst_14405 ( .A(net_6421), .ZN(net_6245) );
NOR2_X2 inst_4169 ( .ZN(net_20292), .A1(net_6550), .A2(net_4981) );
INV_X4 inst_16755 ( .A(net_2137), .ZN(net_1651) );
NAND2_X2 inst_9894 ( .ZN(net_12944), .A1(net_9363), .A2(net_154) );
AOI211_X2 inst_20997 ( .ZN(net_19970), .C1(net_15666), .B(net_15549), .C2(net_15434), .A(net_14913) );
INV_X2 inst_19563 ( .A(net_1328), .ZN(net_804) );
NAND2_X4 inst_6863 ( .ZN(net_18378), .A1(net_18268), .A2(net_18229) );
AOI21_X2 inst_20296 ( .A(net_20952), .B2(net_20093), .B1(net_20092), .ZN(net_16147) );
INV_X4 inst_18149 ( .A(net_20963), .ZN(net_809) );
NAND4_X2 inst_5346 ( .ZN(net_20290), .A1(net_14555), .A3(net_13546), .A4(net_13071), .A2(net_12287) );
CLKBUF_X2 inst_22507 ( .A(net_21906), .Z(net_22379) );
NOR2_X2 inst_4181 ( .A2(net_13840), .ZN(net_8102), .A1(net_6889) );
NAND2_X2 inst_10865 ( .ZN(net_11731), .A1(net_10286), .A2(net_5709) );
OAI21_X2 inst_2008 ( .ZN(net_11396), .A(net_11395), .B1(net_7411), .B2(net_4808) );
INV_X4 inst_16786 ( .ZN(net_1209), .A(net_1019) );
XNOR2_X2 inst_641 ( .A(net_16743), .B(net_16607), .ZN(net_408) );
XNOR2_X2 inst_498 ( .ZN(net_9003), .A(net_9002), .B(net_2511) );
INV_X4 inst_17902 ( .ZN(net_294), .A(net_115) );
INV_X4 inst_17623 ( .A(net_20851), .ZN(net_8369) );
OAI21_X2 inst_1988 ( .B1(net_20121), .ZN(net_12045), .A(net_11195), .B2(net_1963) );
NAND2_X2 inst_8374 ( .ZN(net_19854), .A1(net_19451), .A2(net_17357) );
INV_X8 inst_12346 ( .ZN(net_1692), .A(net_63) );
NAND2_X2 inst_8287 ( .A2(net_20464), .ZN(net_17621), .A1(net_17446) );
NAND2_X2 inst_11971 ( .ZN(net_6899), .A1(net_1345), .A2(net_112) );
NAND4_X2 inst_5517 ( .A1(net_11746), .ZN(net_9888), .A2(net_9887), .A4(net_6591), .A3(net_6105) );
CLKBUF_X2 inst_22229 ( .A(net_22100), .Z(net_22101) );
OAI21_X2 inst_1912 ( .B1(net_20497), .ZN(net_13068), .A(net_12203), .B2(net_9729) );
INV_X4 inst_14478 ( .ZN(net_8187), .A(net_4879) );
OAI21_X2 inst_1831 ( .ZN(net_19093), .B1(net_11237), .B2(net_10450), .A(net_784) );
INV_X4 inst_13438 ( .ZN(net_11677), .A(net_9817) );
NAND3_X2 inst_6714 ( .ZN(net_7095), .A2(net_7094), .A3(net_7093), .A1(net_3950) );
NAND3_X2 inst_6683 ( .A2(net_13542), .A3(net_8567), .ZN(net_7716), .A1(net_4423) );
INV_X4 inst_14339 ( .ZN(net_5829), .A(net_5380) );
INV_X4 inst_13671 ( .A(net_11594), .ZN(net_8052) );
NOR2_X2 inst_3468 ( .ZN(net_14590), .A2(net_13277), .A1(net_12205) );
OAI211_X2 inst_2395 ( .ZN(net_16129), .A(net_15859), .B(net_15670), .C2(net_11843), .C1(net_5186) );
XNOR2_X2 inst_231 ( .ZN(net_17453), .A(net_17034), .B(net_306) );
NAND2_X2 inst_9024 ( .ZN(net_14089), .A2(net_12158), .A1(net_11893) );
NOR2_X4 inst_3309 ( .A2(net_20876), .ZN(net_1090), .A1(net_796) );
NAND2_X2 inst_9952 ( .A1(net_11713), .A2(net_11589), .ZN(net_8936) );
NAND3_X2 inst_5676 ( .ZN(net_16366), .A3(net_16148), .A2(net_14003), .A1(net_12750) );
AOI222_X2 inst_20063 ( .C1(net_20447), .ZN(net_14187), .A1(net_14186), .B1(net_14185), .C2(net_12320), .A2(net_9077), .B2(net_5290) );
INV_X4 inst_15459 ( .ZN(net_11783), .A(net_7822) );
OAI21_X2 inst_2317 ( .ZN(net_19705), .A(net_12382), .B2(net_5683), .B1(net_2169) );
NAND2_X2 inst_11365 ( .ZN(net_6130), .A2(net_3595), .A1(net_1100) );
INV_X4 inst_15816 ( .ZN(net_3864), .A(net_1872) );
NAND3_X2 inst_6756 ( .A2(net_11751), .ZN(net_5704), .A3(net_4284), .A1(net_2596) );
INV_X4 inst_15208 ( .ZN(net_3670), .A(net_2900) );
NOR2_X2 inst_5000 ( .A1(net_3713), .ZN(net_2844), .A2(net_780) );
NOR2_X2 inst_4077 ( .ZN(net_10290), .A2(net_7448), .A1(net_90) );
NOR2_X4 inst_3139 ( .ZN(net_6700), .A2(net_3820), .A1(net_911) );
INV_X4 inst_12801 ( .ZN(net_17747), .A(net_17590) );
OAI211_X2 inst_2558 ( .ZN(net_9934), .C1(net_8836), .A(net_8515), .C2(net_8505), .B(net_5195) );
INV_X2 inst_18591 ( .ZN(net_10153), .A(net_10152) );
XNOR2_X2 inst_352 ( .ZN(net_16936), .A(net_16935), .B(net_16335) );
XNOR2_X2 inst_286 ( .B(net_21202), .ZN(net_17153), .A(net_16806) );
INV_X4 inst_17452 ( .ZN(net_4183), .A(net_86) );
INV_X4 inst_13354 ( .A(net_12989), .ZN(net_10985) );
NAND2_X2 inst_10112 ( .A1(net_9018), .ZN(net_8426), .A2(net_5207) );
NAND2_X4 inst_6880 ( .ZN(net_18202), .A1(net_18125), .A2(net_18110) );
INV_X4 inst_15328 ( .A(net_11858), .ZN(net_3397) );
INV_X4 inst_15663 ( .ZN(net_2069), .A(net_2068) );
NAND2_X2 inst_10447 ( .ZN(net_11728), .A1(net_7155), .A2(net_3551) );
INV_X4 inst_14959 ( .ZN(net_6000), .A(net_3490) );
INV_X4 inst_12984 ( .A(net_17517), .ZN(net_16994) );
INV_X4 inst_15524 ( .ZN(net_14319), .A(net_10292) );
INV_X4 inst_13006 ( .ZN(net_16748), .A(net_16584) );
NAND2_X2 inst_7961 ( .ZN(net_20154), .A2(net_18390), .A1(net_16999) );
CLKBUF_X2 inst_21865 ( .A(net_21736), .Z(net_21737) );
INV_X4 inst_16900 ( .ZN(net_1279), .A(net_532) );
NAND3_X2 inst_6792 ( .A3(net_5836), .ZN(net_4019), .A2(net_4018), .A1(net_1496) );
INV_X4 inst_16361 ( .ZN(net_13542), .A(net_1291) );
INV_X4 inst_15058 ( .A(net_15542), .ZN(net_3306) );
NOR2_X2 inst_3841 ( .ZN(net_9598), .A2(net_9597), .A1(net_6037) );
NAND2_X2 inst_9555 ( .ZN(net_13746), .A2(net_10952), .A1(net_9014) );
CLKBUF_X2 inst_22777 ( .A(net_22566), .Z(net_22649) );
NAND2_X2 inst_7737 ( .ZN(net_18810), .A2(net_18778), .A1(net_17723) );
NAND2_X4 inst_6972 ( .ZN(net_17406), .A1(net_16975), .A2(net_16817) );
INV_X8 inst_12203 ( .ZN(net_11135), .A(net_7631) );
NAND2_X2 inst_9427 ( .ZN(net_11616), .A2(net_9670), .A1(net_2484) );
AOI21_X2 inst_20613 ( .ZN(net_19614), .B2(net_10901), .A(net_8414), .B1(net_7316) );
DFF_X1 inst_19817 ( .QN(net_21175), .D(net_17836), .CK(net_22473) );
NAND3_X2 inst_5887 ( .ZN(net_15228), .A3(net_14126), .A2(net_10462), .A1(net_3157) );
INV_X2 inst_19438 ( .ZN(net_1720), .A(net_956) );
NAND2_X2 inst_11598 ( .ZN(net_2667), .A2(net_2039), .A1(net_1848) );
AND2_X2 inst_21362 ( .ZN(net_1486), .A2(net_108), .A1(net_61) );
AOI211_X2 inst_21045 ( .ZN(net_12893), .C2(net_9490), .C1(net_7573), .B(net_3899), .A(net_2755) );
INV_X4 inst_13452 ( .ZN(net_9731), .A(net_9730) );
CLKBUF_X2 inst_22339 ( .A(net_22210), .Z(net_22211) );
NAND2_X2 inst_12001 ( .ZN(net_1179), .A1(net_1013), .A2(net_879) );
INV_X4 inst_17809 ( .A(net_525), .ZN(net_118) );
XNOR2_X2 inst_425 ( .A(net_16506), .ZN(net_16503), .B(net_1517) );
CLKBUF_X2 inst_22174 ( .A(net_22045), .Z(net_22046) );
CLKBUF_X2 inst_21688 ( .A(net_21442), .Z(net_21560) );
NAND2_X2 inst_8416 ( .A2(net_17245), .ZN(net_17226), .A1(net_16990) );
AOI21_X4 inst_20118 ( .B2(net_19055), .B1(net_19054), .A(net_16395), .ZN(net_16253) );
INV_X4 inst_15298 ( .ZN(net_5208), .A(net_2078) );
OAI211_X2 inst_2572 ( .C1(net_20549), .ZN(net_8996), .B(net_8995), .A(net_8486), .C2(net_3177) );
INV_X4 inst_13764 ( .ZN(net_11435), .A(net_7608) );
NAND2_X2 inst_9380 ( .ZN(net_11938), .A1(net_9470), .A2(net_8930) );
NAND3_X2 inst_6755 ( .A1(net_10091), .A2(net_8376), .ZN(net_5710), .A3(net_5709) );
INV_X4 inst_13111 ( .ZN(net_19987), .A(net_15409) );
NOR2_X2 inst_3365 ( .A2(net_17416), .ZN(net_17145), .A1(net_17144) );
NOR2_X4 inst_3254 ( .ZN(net_7144), .A1(net_1666), .A2(net_412) );
INV_X4 inst_17885 ( .ZN(net_1435), .A(net_75) );
SDFF_X2 inst_983 ( .QN(net_20987), .D(net_2313), .SE(net_263), .CK(net_21842), .SI(x3209) );
NOR2_X2 inst_4980 ( .ZN(net_2127), .A1(net_1491), .A2(net_1236) );
NAND2_X2 inst_8026 ( .ZN(net_20719), .A2(net_18202), .A1(net_17362) );
AOI22_X2 inst_20004 ( .A1(net_15372), .ZN(net_13311), .B1(net_13310), .A2(net_9919), .B2(net_5597) );
NAND2_X2 inst_7773 ( .ZN(net_18739), .A1(net_18738), .A2(net_18737) );
CLKBUF_X2 inst_22572 ( .A(net_21660), .Z(net_22444) );
INV_X4 inst_17426 ( .ZN(net_1991), .A(net_504) );
NAND2_X2 inst_11291 ( .ZN(net_11264), .A2(net_2367), .A1(net_1650) );
NAND2_X2 inst_11196 ( .A1(net_8457), .ZN(net_5158), .A2(net_2150) );
NOR2_X2 inst_4776 ( .ZN(net_2910), .A1(net_2909), .A2(net_2908) );
NAND3_X2 inst_6237 ( .ZN(net_13210), .A3(net_13209), .A2(net_11925), .A1(net_9769) );
NOR3_X4 inst_2633 ( .ZN(net_19250), .A1(net_10479), .A2(net_8391), .A3(net_4215) );
NAND2_X4 inst_6947 ( .A2(net_19656), .A1(net_19655), .ZN(net_17615) );
NAND3_X2 inst_6274 ( .ZN(net_12920), .A2(net_12245), .A3(net_10949), .A1(net_4766) );
CLKBUF_X2 inst_22459 ( .A(net_22330), .Z(net_22331) );
NAND2_X4 inst_7029 ( .A2(net_20744), .A1(net_20743), .ZN(net_17060) );
OAI21_X2 inst_2130 ( .ZN(net_9996), .B1(net_8120), .B2(net_5039), .A(net_948) );
NOR2_X2 inst_4388 ( .ZN(net_6328), .A2(net_3667), .A1(net_809) );
SDFF_X2 inst_1055 ( .QN(net_21051), .D(net_350), .SE(net_263), .CK(net_22482), .SI(x2174) );
INV_X4 inst_13114 ( .ZN(net_15614), .A(net_15347) );
OAI21_X2 inst_2100 ( .A(net_10158), .ZN(net_10069), .B2(net_10068), .B1(net_3668) );
INV_X4 inst_16813 ( .ZN(net_4464), .A(net_3151) );
OAI21_X2 inst_2284 ( .ZN(net_6546), .A(net_6545), .B2(net_1875), .B1(net_1852) );
INV_X4 inst_16028 ( .ZN(net_3235), .A(net_1136) );
NOR2_X2 inst_4829 ( .ZN(net_2480), .A2(net_1609), .A1(net_790) );
INV_X4 inst_16032 ( .ZN(net_11007), .A(net_5712) );
INV_X4 inst_16505 ( .ZN(net_9667), .A(net_5217) );
INV_X2 inst_19041 ( .ZN(net_4769), .A(net_4768) );
SDFF_X2 inst_923 ( .Q(net_21170), .D(net_16532), .SE(net_263), .CK(net_22412), .SI(x4888) );
NAND2_X1 inst_12153 ( .ZN(net_9851), .A1(net_9847), .A2(net_6434) );
NAND2_X2 inst_8671 ( .A2(net_19423), .ZN(net_16466), .A1(net_16465) );
NAND2_X2 inst_8599 ( .A1(net_21198), .A2(net_19431), .ZN(net_19129) );
INV_X4 inst_17569 ( .ZN(net_1562), .A(net_227) );
NAND2_X2 inst_11604 ( .A2(net_8184), .ZN(net_2635), .A1(net_2634) );
INV_X4 inst_13470 ( .A(net_10269), .ZN(net_9649) );
NAND2_X4 inst_6975 ( .A1(net_17353), .ZN(net_17241), .A2(net_17239) );
NAND2_X2 inst_11819 ( .ZN(net_3543), .A1(net_2563), .A2(net_1818) );
NAND2_X4 inst_7564 ( .A2(net_20580), .ZN(net_1877), .A1(net_169) );
NAND2_X4 inst_7109 ( .ZN(net_11517), .A2(net_11174), .A1(net_10987) );
INV_X1 inst_19746 ( .ZN(net_17306), .A(net_17305) );
INV_X4 inst_16073 ( .A(net_8455), .ZN(net_1560) );
NAND3_X2 inst_5890 ( .ZN(net_15221), .A3(net_14118), .A2(net_11152), .A1(net_9684) );
INV_X2 inst_18764 ( .A(net_9793), .ZN(net_7615) );
NAND2_X2 inst_8793 ( .ZN(net_18945), .A1(net_15742), .A2(net_15382) );
INV_X2 inst_19634 ( .A(net_19422), .ZN(net_19420) );
INV_X4 inst_12946 ( .ZN(net_16783), .A(net_16630) );
NOR2_X2 inst_3766 ( .ZN(net_14293), .A2(net_11807), .A1(net_2520) );
INV_X4 inst_12480 ( .ZN(net_18691), .A(net_18690) );
NAND3_X2 inst_5935 ( .ZN(net_14924), .A3(net_13474), .A1(net_9370), .A2(net_2612) );
NAND2_X4 inst_7704 ( .ZN(net_511), .A2(net_265), .A1(net_153) );
OAI211_X2 inst_2536 ( .A(net_20592), .ZN(net_11237), .C1(net_6886), .B(net_6243), .C2(net_5719) );
NAND2_X2 inst_11730 ( .A2(net_3688), .A1(net_3350), .ZN(net_2223) );
INV_X4 inst_13103 ( .ZN(net_19336), .A(net_15646) );
NAND2_X2 inst_9389 ( .ZN(net_11788), .A2(net_10029), .A1(net_8779) );
CLKBUF_X2 inst_21743 ( .A(net_21614), .Z(net_21615) );
NAND2_X4 inst_7100 ( .ZN(net_13555), .A2(net_13554), .A1(net_13553) );
NAND2_X2 inst_9618 ( .A1(net_10930), .ZN(net_10692), .A2(net_8471) );
INV_X4 inst_14036 ( .ZN(net_9807), .A(net_5137) );
NAND2_X4 inst_6870 ( .ZN(net_19391), .A1(net_18231), .A2(net_18142) );
CLKBUF_X2 inst_22848 ( .A(net_22399), .Z(net_22720) );
INV_X4 inst_13300 ( .ZN(net_13589), .A(net_12322) );
NAND3_X2 inst_5915 ( .A2(net_20300), .A1(net_20299), .A3(net_19868), .ZN(net_19536) );
CLKBUF_X2 inst_22737 ( .A(net_22608), .Z(net_22609) );
NAND2_X2 inst_10998 ( .ZN(net_11029), .A2(net_3517), .A1(net_165) );
OAI21_X2 inst_1925 ( .ZN(net_13020), .B1(net_13019), .B2(net_13018), .A(net_11549) );
XOR2_X2 inst_40 ( .A(net_21121), .Z(net_590), .B(net_589) );
NOR2_X2 inst_4437 ( .ZN(net_4839), .A1(net_4838), .A2(net_4837) );
INV_X4 inst_16007 ( .ZN(net_13383), .A(net_1657) );
CLKBUF_X2 inst_22405 ( .A(net_21820), .Z(net_22277) );
AOI21_X2 inst_20899 ( .ZN(net_7721), .A(net_5028), .B2(net_3462), .B1(net_2411) );
NAND2_X2 inst_8765 ( .ZN(net_18951), .A2(net_15621), .A1(net_333) );
OAI21_X4 inst_1416 ( .A(net_20920), .ZN(net_20304), .B2(net_19936), .B1(net_19935) );
NAND2_X2 inst_12066 ( .A1(net_20545), .ZN(net_1886), .A2(net_61) );
CLKBUF_X2 inst_22281 ( .A(net_22152), .Z(net_22153) );
NAND2_X4 inst_7280 ( .ZN(net_9586), .A1(net_5806), .A2(net_3133) );
XNOR2_X2 inst_439 ( .B(net_17091), .A(net_16599), .ZN(net_16091) );
AOI21_X2 inst_20410 ( .ZN(net_20361), .B2(net_20149), .B1(net_20148), .A(net_12133) );
INV_X4 inst_17304 ( .ZN(net_9364), .A(net_3816) );
INV_X4 inst_16582 ( .A(net_1219), .ZN(net_1151) );
NAND2_X2 inst_11567 ( .ZN(net_2796), .A1(net_2795), .A2(net_1201) );
NOR2_X2 inst_4529 ( .ZN(net_7035), .A1(net_4056), .A2(net_1891) );
INV_X4 inst_17445 ( .A(net_20889), .ZN(net_750) );
INV_X4 inst_15216 ( .ZN(net_6541), .A(net_2482) );
CLKBUF_X2 inst_22121 ( .A(net_21992), .Z(net_21993) );
NAND2_X2 inst_8280 ( .A1(net_21120), .ZN(net_20243), .A2(net_17613) );
INV_X4 inst_16816 ( .ZN(net_1505), .A(net_1007) );
INV_X4 inst_13309 ( .A(net_13140), .ZN(net_11692) );
INV_X4 inst_13475 ( .ZN(net_12923), .A(net_9616) );
INV_X4 inst_17009 ( .A(net_1821), .ZN(net_1341) );
NAND2_X2 inst_9478 ( .ZN(net_14312), .A1(net_11460), .A2(net_10893) );
INV_X2 inst_19614 ( .A(net_20871), .ZN(net_45) );
INV_X2 inst_18643 ( .A(net_10160), .ZN(net_9372) );
XNOR2_X2 inst_654 ( .B(net_17097), .A(net_543), .ZN(net_360) );
INV_X4 inst_17077 ( .ZN(net_14174), .A(net_1000) );
AND2_X2 inst_21299 ( .ZN(net_19842), .A2(net_10116), .A1(net_9623) );
INV_X4 inst_16152 ( .ZN(net_4669), .A(net_1063) );
INV_X4 inst_13616 ( .ZN(net_9815), .A(net_8371) );
AOI21_X2 inst_20834 ( .ZN(net_9326), .A(net_9325), .B2(net_7672), .B1(net_4527) );
INV_X4 inst_16284 ( .A(net_11460), .ZN(net_10151) );
INV_X4 inst_16486 ( .ZN(net_3205), .A(net_1200) );
INV_X4 inst_13656 ( .ZN(net_8146), .A(net_8145) );
INV_X4 inst_17130 ( .ZN(net_770), .A(net_769) );
INV_X4 inst_16574 ( .ZN(net_1933), .A(net_1797) );
OAI21_X2 inst_1708 ( .ZN(net_15203), .B1(net_15202), .B2(net_14087), .A(net_13687) );
INV_X4 inst_15264 ( .A(net_5671), .ZN(net_5088) );
CLKBUF_X2 inst_22657 ( .A(net_22528), .Z(net_22529) );
INV_X4 inst_15096 ( .ZN(net_5215), .A(net_2223) );
NAND2_X2 inst_11997 ( .ZN(net_1191), .A2(net_915), .A1(net_400) );
NAND2_X2 inst_10440 ( .A1(net_9516), .A2(net_8704), .ZN(net_7191) );
NAND2_X2 inst_11004 ( .A1(net_10015), .ZN(net_4886), .A2(net_3176) );
INV_X4 inst_17469 ( .ZN(net_7071), .A(net_6377) );
NOR3_X2 inst_2738 ( .ZN(net_12772), .A2(net_12771), .A3(net_12770), .A1(net_10308) );
INV_X4 inst_16164 ( .ZN(net_9943), .A(net_6150) );
XNOR2_X2 inst_634 ( .B(net_16775), .ZN(net_436), .A(net_435) );
CLKBUF_X2 inst_22714 ( .A(net_22585), .Z(net_22586) );
NOR2_X4 inst_3122 ( .ZN(net_6672), .A2(net_3333), .A1(net_85) );
INV_X4 inst_15229 ( .ZN(net_2853), .A(net_2852) );
NAND2_X2 inst_9090 ( .A1(net_14363), .ZN(net_13794), .A2(net_12472) );
INV_X4 inst_16989 ( .ZN(net_1233), .A(net_90) );
INV_X4 inst_17184 ( .ZN(net_903), .A(net_252) );
NAND2_X2 inst_9232 ( .ZN(net_12759), .A2(net_10099), .A1(net_7529) );
NAND2_X2 inst_10420 ( .ZN(net_20265), .A2(net_8995), .A1(net_7232) );
INV_X4 inst_18202 ( .A(net_21041), .ZN(net_496) );
AND2_X2 inst_21316 ( .A2(net_9037), .ZN(net_7177), .A1(net_7074) );
INV_X2 inst_19540 ( .ZN(net_2576), .A(net_1784) );
OAI21_X4 inst_1477 ( .ZN(net_14699), .A(net_14663), .B2(net_12191), .B1(net_11517) );
INV_X4 inst_13774 ( .ZN(net_11054), .A(net_9553) );
NAND2_X2 inst_9263 ( .ZN(net_14272), .A2(net_12305), .A1(net_11270) );
NAND2_X4 inst_7043 ( .ZN(net_16701), .A2(net_16376), .A1(net_16363) );
NAND2_X2 inst_9813 ( .ZN(net_18992), .A1(net_9666), .A2(net_9665) );
XNOR2_X2 inst_529 ( .B(net_21106), .ZN(net_4406), .A(net_1352) );
OAI21_X2 inst_1528 ( .ZN(net_18016), .A(net_17971), .B1(net_17970), .B2(net_17969) );
NAND2_X2 inst_11192 ( .ZN(net_7041), .A1(net_4088), .A2(net_4087) );
INV_X4 inst_17122 ( .A(net_6951), .ZN(net_6274) );
INV_X4 inst_15921 ( .ZN(net_13703), .A(net_12522) );
INV_X4 inst_15705 ( .ZN(net_3646), .A(net_3053) );
INV_X4 inst_16333 ( .ZN(net_11614), .A(net_8286) );
NAND3_X2 inst_5788 ( .ZN(net_15773), .A3(net_15132), .A2(net_13377), .A1(net_12704) );
NAND2_X2 inst_11788 ( .A2(net_2232), .ZN(net_1974), .A1(net_90) );
INV_X4 inst_17562 ( .A(net_937), .ZN(net_363) );
INV_X4 inst_15460 ( .ZN(net_2688), .A(net_2476) );
INV_X4 inst_14267 ( .A(net_8019), .ZN(net_5720) );
NAND2_X2 inst_11030 ( .ZN(net_4763), .A1(net_3106), .A2(net_2190) );
XNOR2_X2 inst_675 ( .ZN(net_18870), .B(net_18138), .A(net_11863) );
NOR2_X2 inst_4068 ( .ZN(net_9096), .A2(net_7695), .A1(net_732) );
NAND2_X2 inst_11953 ( .ZN(net_10587), .A2(net_8097), .A1(net_293) );
INV_X4 inst_13706 ( .ZN(net_9404), .A(net_7868) );
NAND3_X2 inst_5729 ( .ZN(net_16104), .A3(net_16009), .A1(net_15856), .A2(net_13379) );
NOR3_X2 inst_2705 ( .ZN(net_13909), .A2(net_12915), .A1(net_12046), .A3(net_3141) );
INV_X2 inst_19210 ( .A(net_4828), .ZN(net_3510) );
INV_X2 inst_19192 ( .A(net_5106), .ZN(net_3647) );
INV_X4 inst_16662 ( .ZN(net_12330), .A(net_948) );
INV_X4 inst_13291 ( .ZN(net_13571), .A(net_12390) );
INV_X4 inst_12902 ( .ZN(net_16707), .A(net_16552) );
INV_X4 inst_12924 ( .A(net_16689), .ZN(net_16658) );
NAND3_X2 inst_5737 ( .ZN(net_19950), .A3(net_15467), .A1(net_14478), .A2(net_14390) );
NAND4_X2 inst_5332 ( .ZN(net_15557), .A4(net_14618), .A2(net_13990), .A1(net_11581), .A3(net_11117) );
CLKBUF_X2 inst_22267 ( .A(net_22138), .Z(net_22139) );
INV_X2 inst_19382 ( .ZN(net_19522), .A(net_3065) );
NAND2_X2 inst_11144 ( .A1(net_6702), .ZN(net_4730), .A2(net_2024) );
NAND2_X2 inst_9078 ( .A1(net_15248), .ZN(net_13831), .A2(net_13820) );
AOI21_X2 inst_20344 ( .A(net_20904), .B2(net_19199), .B1(net_19198), .ZN(net_15763) );
NOR2_X2 inst_3751 ( .ZN(net_10413), .A2(net_10190), .A1(net_8581) );
INV_X2 inst_19503 ( .ZN(net_1252), .A(net_1251) );
INV_X4 inst_17272 ( .A(net_1384), .ZN(net_1354) );
AOI21_X2 inst_20285 ( .B2(net_19717), .B1(net_19716), .A(net_16390), .ZN(net_16251) );
INV_X4 inst_12463 ( .ZN(net_18824), .A(net_18823) );
NAND3_X2 inst_6735 ( .ZN(net_6475), .A2(net_6474), .A1(net_3455), .A3(net_2832) );
NAND3_X2 inst_6643 ( .A3(net_9046), .ZN(net_8944), .A1(net_6699), .A2(net_2767) );
AOI21_X2 inst_20862 ( .ZN(net_8757), .B2(net_7906), .B1(net_3569), .A(net_761) );
INV_X4 inst_16538 ( .ZN(net_6639), .A(net_3293) );
NAND2_X2 inst_9123 ( .ZN(net_13539), .A1(net_13538), .A2(net_11078) );
OAI21_X2 inst_2222 ( .B2(net_9887), .ZN(net_8510), .A(net_7791), .B1(net_6743) );
NOR2_X2 inst_4578 ( .ZN(net_4835), .A2(net_3850), .A1(net_209) );
AOI21_X4 inst_20254 ( .ZN(net_6500), .B1(net_5211), .B2(net_3416), .A(net_890) );
AOI21_X2 inst_20819 ( .ZN(net_10016), .B1(net_10015), .B2(net_6851), .A(net_5938) );
NAND2_X2 inst_12102 ( .ZN(net_476), .A2(net_265), .A1(net_80) );
NOR2_X2 inst_4059 ( .ZN(net_9344), .A2(net_7833), .A1(net_6750) );
CLKBUF_X2 inst_22049 ( .A(net_21920), .Z(net_21921) );
OAI21_X2 inst_1755 ( .ZN(net_20844), .A(net_14791), .B2(net_13259), .B1(net_9694) );
CLKBUF_X2 inst_21495 ( .A(net_21366), .Z(net_21367) );
INV_X2 inst_19508 ( .ZN(net_1218), .A(net_1217) );
AOI21_X2 inst_20655 ( .ZN(net_13037), .B2(net_9749), .B1(net_5322), .A(net_1611) );
AOI21_X4 inst_20203 ( .B2(net_19251), .B1(net_19250), .ZN(net_14797), .A(net_14714) );
INV_X4 inst_15390 ( .ZN(net_5582), .A(net_2549) );
AOI211_X2 inst_21029 ( .ZN(net_14540), .B(net_11752), .A(net_11324), .C1(net_10947), .C2(net_9040) );
INV_X4 inst_15027 ( .ZN(net_15519), .A(net_10947) );
CLKBUF_X2 inst_22707 ( .A(net_21683), .Z(net_22579) );
INV_X4 inst_12715 ( .A(net_17550), .ZN(net_17549) );
SDFF_X2 inst_806 ( .Q(net_20855), .SE(net_18864), .SI(net_17936), .D(net_347), .CK(net_22612) );
INV_X1 inst_19751 ( .A(net_11425), .ZN(net_10901) );
INV_X2 inst_18851 ( .ZN(net_6596), .A(net_6595) );
NAND2_X4 inst_7119 ( .ZN(net_11019), .A1(net_10240), .A2(net_7922) );
NAND2_X4 inst_7232 ( .ZN(net_12266), .A1(net_6656), .A2(net_86) );
XNOR2_X2 inst_491 ( .A(net_16093), .ZN(net_9239), .B(net_4440) );
NAND2_X2 inst_10485 ( .ZN(net_12233), .A1(net_6945), .A2(net_6944) );
NAND3_X2 inst_6027 ( .A3(net_19750), .ZN(net_19593), .A1(net_12633), .A2(net_6642) );
NOR2_X2 inst_4943 ( .ZN(net_2237), .A2(net_1320), .A1(net_85) );
INV_X4 inst_13219 ( .ZN(net_13631), .A(net_12785) );
INV_X4 inst_13515 ( .ZN(net_11582), .A(net_9398) );
NAND2_X2 inst_10987 ( .ZN(net_4941), .A2(net_4181), .A1(net_2431) );
NAND2_X2 inst_12097 ( .A2(net_1271), .ZN(net_882), .A1(net_550) );
NAND2_X2 inst_9441 ( .ZN(net_20162), .A2(net_11554), .A1(net_9983) );
NOR2_X4 inst_3086 ( .ZN(net_6781), .A1(net_4081), .A2(net_2585) );
NOR3_X2 inst_2791 ( .A2(net_9768), .ZN(net_4509), .A3(net_4508), .A1(net_3715) );
NAND2_X2 inst_12090 ( .A1(net_1097), .ZN(net_978), .A2(net_664) );
NAND3_X4 inst_5583 ( .A2(net_19329), .A1(net_19328), .ZN(net_15529), .A3(net_14718) );
INV_X4 inst_16514 ( .ZN(net_3947), .A(net_1689) );
NAND2_X2 inst_10243 ( .ZN(net_10202), .A1(net_9301), .A2(net_5119) );
INV_X4 inst_15633 ( .ZN(net_3380), .A(net_1388) );
INV_X4 inst_14814 ( .A(net_14751), .ZN(net_3943) );
CLKBUF_X2 inst_21853 ( .A(net_21724), .Z(net_21725) );
NOR2_X2 inst_4419 ( .ZN(net_6319), .A2(net_5211), .A1(net_4990) );
INV_X4 inst_16342 ( .ZN(net_1937), .A(net_1003) );
NAND2_X4 inst_6850 ( .ZN(net_18536), .A2(net_18482), .A1(net_18454) );
NAND3_X2 inst_6698 ( .ZN(net_7611), .A2(net_7610), .A1(net_4485), .A3(net_2795) );
OAI221_X2 inst_1349 ( .C1(net_13785), .C2(net_11338), .ZN(net_10782), .B2(net_10781), .B1(net_8991), .A(net_8661) );
AOI21_X2 inst_20676 ( .B1(net_13080), .ZN(net_12482), .B2(net_11053), .A(net_6230) );
INV_X2 inst_18390 ( .A(net_16792), .ZN(net_16633) );
NAND2_X4 inst_7012 ( .A2(net_18972), .A1(net_18971), .ZN(net_17138) );
INV_X4 inst_12744 ( .ZN(net_17431), .A(net_17430) );
NOR2_X2 inst_3745 ( .A2(net_12105), .ZN(net_11999), .A1(net_8967) );
AOI21_X2 inst_20970 ( .A(net_5950), .ZN(net_4909), .B2(net_4908), .B1(net_1540) );
INV_X4 inst_15345 ( .ZN(net_12542), .A(net_7396) );
NOR2_X2 inst_4347 ( .ZN(net_5626), .A1(net_5625), .A2(net_2984) );
INV_X4 inst_16404 ( .ZN(net_10864), .A(net_8674) );
NAND3_X2 inst_5962 ( .ZN(net_20011), .A3(net_13445), .A2(net_11653), .A1(net_8170) );
OAI21_X2 inst_2224 ( .ZN(net_12229), .B2(net_8483), .B1(net_5596), .A(net_60) );
NAND2_X2 inst_10002 ( .A2(net_8942), .ZN(net_8818), .A1(net_8481) );
NAND2_X2 inst_10185 ( .ZN(net_20322), .A1(net_8179), .A2(net_4899) );
CLKBUF_X2 inst_21427 ( .A(net_21249), .Z(net_21299) );
NAND4_X4 inst_5226 ( .A4(net_19316), .A1(net_19315), .ZN(net_16336), .A2(net_16108), .A3(net_15734) );
INV_X4 inst_13012 ( .ZN(net_16742), .A(net_16574) );
NAND4_X2 inst_5310 ( .ZN(net_15794), .A2(net_14801), .A1(net_14004), .A4(net_11528), .A3(net_8167) );
INV_X2 inst_19687 ( .A(net_20532), .ZN(net_20531) );
NAND2_X2 inst_8412 ( .ZN(net_19855), .A1(net_19452), .A2(net_17231) );
CLKBUF_X2 inst_22662 ( .A(net_22533), .Z(net_22534) );
NOR2_X2 inst_4996 ( .ZN(net_1371), .A1(net_1370), .A2(net_1369) );
OAI21_X2 inst_1890 ( .A(net_14195), .ZN(net_13420), .B1(net_10669), .B2(net_5971) );
OAI21_X2 inst_2308 ( .A(net_11572), .ZN(net_5753), .B2(net_5752), .B1(net_2191) );
NOR2_X2 inst_4093 ( .A1(net_8748), .ZN(net_7241), .A2(net_6770) );
NOR2_X4 inst_2879 ( .ZN(net_10147), .A1(net_10146), .A2(net_8226) );
INV_X2 inst_19397 ( .ZN(net_2048), .A(net_2047) );
DFF_X1 inst_19786 ( .D(net_18681), .CK(net_22131), .Q(x539) );
INV_X4 inst_14676 ( .ZN(net_4311), .A(net_4310) );
NAND2_X4 inst_7482 ( .ZN(net_3333), .A1(net_1708), .A2(net_1041) );
OAI21_X2 inst_2338 ( .ZN(net_4680), .B2(net_3695), .B1(net_3595), .A(net_3482) );
NOR2_X2 inst_3475 ( .ZN(net_14451), .A2(net_12780), .A1(net_12144) );
INV_X4 inst_13170 ( .ZN(net_20143), .A(net_14124) );
INV_X4 inst_15547 ( .A(net_3224), .ZN(net_2353) );
NAND2_X2 inst_7818 ( .ZN(net_18658), .A2(net_18639), .A1(net_16762) );
NAND2_X2 inst_11431 ( .ZN(net_5607), .A1(net_4286), .A2(net_3374) );
INV_X4 inst_18319 ( .A(net_20529), .ZN(net_20528) );
INV_X2 inst_18977 ( .ZN(net_5172), .A(net_5171) );
CLKBUF_X2 inst_21755 ( .A(net_21626), .Z(net_21627) );
NAND3_X2 inst_6516 ( .ZN(net_19410), .A3(net_13323), .A2(net_9661), .A1(net_6344) );
NAND2_X2 inst_8649 ( .A1(net_16734), .ZN(net_16563), .A2(net_16562) );
NAND4_X4 inst_5198 ( .A2(net_19068), .A1(net_19067), .A3(net_19049), .ZN(net_17483), .A4(net_16280) );
NAND3_X2 inst_5909 ( .ZN(net_15056), .A3(net_12964), .A1(net_11649), .A2(net_7191) );
CLKBUF_X2 inst_22607 ( .A(net_21697), .Z(net_22479) );
INV_X2 inst_19003 ( .ZN(net_5040), .A(net_5039) );
AOI21_X2 inst_20328 ( .ZN(net_15834), .A(net_15833), .B2(net_15279), .B1(net_13033) );
INV_X4 inst_16341 ( .ZN(net_14738), .A(net_14689) );
INV_X4 inst_15934 ( .A(net_2260), .ZN(net_1726) );
OAI21_X2 inst_2016 ( .A(net_13984), .ZN(net_11369), .B1(net_11368), .B2(net_4400) );
INV_X4 inst_15679 ( .A(net_13418), .ZN(net_13353) );
INV_X4 inst_12723 ( .ZN(net_17530), .A(net_17529) );
INV_X2 inst_19393 ( .ZN(net_2057), .A(net_2056) );
INV_X4 inst_16431 ( .ZN(net_1422), .A(net_1248) );
NOR2_X2 inst_4012 ( .ZN(net_8073), .A2(net_5948), .A1(net_4913) );
NAND2_X2 inst_8385 ( .ZN(net_17432), .A2(net_17047), .A1(net_16900) );
INV_X4 inst_15152 ( .ZN(net_13651), .A(net_3067) );
NAND2_X2 inst_9289 ( .ZN(net_12462), .A2(net_9420), .A1(net_8200) );
NAND2_X4 inst_7630 ( .ZN(net_1479), .A1(net_1192), .A2(net_282) );
NAND2_X2 inst_9920 ( .ZN(net_9280), .A1(net_5069), .A2(net_2684) );
XNOR2_X2 inst_393 ( .ZN(net_16767), .A(net_16766), .B(net_13292) );
AND2_X2 inst_21344 ( .A1(net_2747), .ZN(net_2719), .A2(net_2718) );
NAND3_X2 inst_5969 ( .A3(net_19904), .A1(net_19903), .ZN(net_19685), .A2(net_11396) );
OAI21_X2 inst_1813 ( .ZN(net_14178), .B1(net_10795), .B2(net_6939), .A(net_4300) );
XNOR2_X2 inst_92 ( .ZN(net_18562), .A(net_18463), .B(net_17159) );
INV_X4 inst_15405 ( .ZN(net_2531), .A(net_1950) );
NAND2_X2 inst_11168 ( .A1(net_5482), .ZN(net_4165), .A2(net_4164) );
XNOR2_X2 inst_345 ( .ZN(net_16953), .A(net_16952), .B(net_10803) );
INV_X4 inst_16386 ( .A(net_14600), .ZN(net_1277) );
NAND2_X2 inst_9086 ( .ZN(net_13799), .A1(net_13544), .A2(net_12489) );
NAND2_X2 inst_11856 ( .A1(net_20495), .ZN(net_1671), .A2(net_883) );
CLKBUF_X2 inst_22160 ( .A(net_22031), .Z(net_22032) );
NAND2_X2 inst_10233 ( .ZN(net_13458), .A1(net_10445), .A2(net_8047) );
NAND2_X2 inst_10087 ( .A1(net_8854), .ZN(net_8627), .A2(net_6386) );
NAND3_X2 inst_6362 ( .A3(net_13914), .ZN(net_12082), .A2(net_5928), .A1(net_5218) );
INV_X2 inst_18377 ( .ZN(net_17062), .A(net_17060) );
NAND2_X2 inst_8076 ( .ZN(net_18159), .A2(net_18158), .A1(net_16655) );
INV_X4 inst_13806 ( .ZN(net_12563), .A(net_7544) );
NAND2_X2 inst_11009 ( .ZN(net_9867), .A2(net_4928), .A1(net_4876) );
NAND2_X2 inst_10585 ( .A1(net_6877), .ZN(net_6663), .A2(net_6662) );
XNOR2_X2 inst_57 ( .ZN(net_18867), .A(net_18850), .B(net_17130) );
INV_X4 inst_15928 ( .ZN(net_9490), .A(net_6999) );
INV_X4 inst_16717 ( .ZN(net_6150), .A(net_1358) );
AOI21_X2 inst_20337 ( .ZN(net_19985), .B1(net_19785), .A(net_10197), .B2(net_750) );
NAND2_X2 inst_9312 ( .ZN(net_12356), .A2(net_10761), .A1(net_10515) );
OAI22_X2 inst_1307 ( .A2(net_9967), .ZN(net_9904), .A1(net_9903), .B1(net_7901), .B2(net_7712) );
NAND2_X2 inst_7759 ( .ZN(net_18762), .A2(net_18710), .A1(net_18686) );
NAND2_X2 inst_10878 ( .ZN(net_5420), .A2(net_5419), .A1(net_955) );
NAND2_X2 inst_8565 ( .ZN(net_16744), .A2(net_16742), .A1(net_5789) );
NAND3_X2 inst_6789 ( .ZN(net_5187), .A1(net_4110), .A3(net_2827), .A2(net_2597) );
INV_X4 inst_16842 ( .ZN(net_8067), .A(net_975) );
INV_X4 inst_12960 ( .A(net_17526), .ZN(net_16683) );
INV_X4 inst_16925 ( .ZN(net_3086), .A(net_1056) );
NAND2_X4 inst_7124 ( .ZN(net_13644), .A1(net_10894), .A2(net_9667) );
NAND2_X2 inst_8616 ( .A2(net_16912), .ZN(net_16611), .A1(net_5788) );
SDFF_X2 inst_851 ( .Q(net_21182), .SI(net_17252), .SE(net_125), .CK(net_22303), .D(x6571) );
SDFF_X2 inst_831 ( .Q(net_21191), .SI(net_17454), .SE(net_125), .CK(net_22238), .D(x6320) );
AOI21_X2 inst_20496 ( .ZN(net_14732), .B1(net_14319), .B2(net_13654), .A(net_13457) );
INV_X4 inst_18024 ( .A(net_21198), .ZN(net_9193) );
NAND3_X2 inst_5824 ( .ZN(net_15568), .A2(net_15567), .A1(net_14811), .A3(net_13511) );
NOR2_X2 inst_4264 ( .A1(net_9514), .ZN(net_6226), .A2(net_6225) );
CLKBUF_X2 inst_21827 ( .A(net_21297), .Z(net_21699) );
INV_X4 inst_17259 ( .ZN(net_1272), .A(net_795) );
INV_X2 inst_19620 ( .A(net_20958), .ZN(net_38) );
INV_X4 inst_17668 ( .A(net_303), .ZN(net_245) );
AOI21_X2 inst_20585 ( .A(net_15452), .ZN(net_14024), .B2(net_10394), .B1(net_10077) );
NAND2_X2 inst_11448 ( .A1(net_9575), .ZN(net_3271), .A2(net_1994) );
NOR2_X2 inst_4430 ( .ZN(net_4897), .A2(net_4758), .A1(net_955) );
AND2_X2 inst_21337 ( .ZN(net_8524), .A2(net_3462), .A1(net_2624) );
INV_X4 inst_15007 ( .ZN(net_7787), .A(net_2626) );
NAND2_X2 inst_11174 ( .ZN(net_7054), .A1(net_4158), .A2(net_4157) );
OAI21_X4 inst_1497 ( .B1(net_19601), .A(net_14642), .ZN(net_12030), .B2(net_8222) );
INV_X2 inst_19663 ( .A(net_20470), .ZN(net_20469) );
NAND3_X2 inst_5706 ( .ZN(net_16202), .A3(net_15857), .A2(net_14649), .A1(net_14294) );
SDFF_X2 inst_1002 ( .QN(net_21069), .D(net_793), .SE(net_263), .CK(net_21720), .SI(x1932) );
CLKBUF_X2 inst_22314 ( .A(net_22185), .Z(net_22186) );
NAND2_X2 inst_12076 ( .ZN(net_1615), .A1(net_801), .A2(net_438) );
NAND2_X2 inst_8057 ( .ZN(net_18206), .A1(net_18205), .A2(net_18204) );
INV_X4 inst_13179 ( .ZN(net_14340), .A(net_13861) );
XNOR2_X2 inst_478 ( .A(net_11876), .ZN(net_11873), .B(net_11872) );
INV_X2 inst_18985 ( .A(net_10361), .ZN(net_5122) );
INV_X4 inst_18113 ( .A(net_20939), .ZN(net_955) );
NAND2_X2 inst_8630 ( .A1(net_19438), .ZN(net_16593), .A2(net_16465) );
INV_X4 inst_15832 ( .ZN(net_3410), .A(net_2047) );
NAND3_X2 inst_5666 ( .A3(net_19823), .A1(net_19822), .ZN(net_16397), .A2(net_14220) );
INV_X2 inst_19229 ( .A(net_14751), .ZN(net_3378) );
INV_X2 inst_18788 ( .ZN(net_10924), .A(net_8744) );
INV_X4 inst_18219 ( .A(net_20877), .ZN(net_132) );
DFF_X1 inst_19904 ( .D(net_16805), .CK(net_22345), .Q(x899) );
INV_X2 inst_19544 ( .A(net_3148), .ZN(net_944) );
INV_X4 inst_13953 ( .ZN(net_6761), .A(net_6760) );
INV_X8 inst_12173 ( .ZN(net_17754), .A(net_17660) );
INV_X4 inst_14126 ( .ZN(net_9688), .A(net_4968) );
NAND4_X2 inst_5378 ( .ZN(net_15163), .A4(net_13783), .A2(net_11811), .A1(net_7400), .A3(net_7282) );
NAND3_X2 inst_5665 ( .A3(net_19169), .A1(net_19168), .ZN(net_16398), .A2(net_14223) );
NOR2_X2 inst_4931 ( .ZN(net_10054), .A1(net_3805), .A2(net_1021) );
NAND2_X2 inst_11540 ( .ZN(net_20815), .A1(net_9345), .A2(net_969) );
INV_X4 inst_15111 ( .ZN(net_14346), .A(net_9762) );
NAND2_X4 inst_7334 ( .ZN(net_6067), .A1(net_3565), .A2(net_3226) );
SDFF_X2 inst_799 ( .Q(net_20919), .SE(net_18577), .SI(net_17985), .D(net_371), .CK(net_21271) );
INV_X4 inst_12906 ( .ZN(net_19768), .A(net_16703) );
NOR2_X2 inst_3481 ( .ZN(net_14362), .A2(net_13134), .A1(net_7245) );
SDFF_X2 inst_738 ( .Q(net_20907), .SE(net_18585), .SI(net_18552), .D(net_13661), .CK(net_22702) );
AOI21_X2 inst_20604 ( .ZN(net_13759), .B2(net_11105), .B1(net_5784), .A(net_702) );
INV_X4 inst_13666 ( .A(net_8098), .ZN(net_8089) );
AOI21_X2 inst_20265 ( .B2(net_20912), .ZN(net_19473), .B1(net_15953), .A(net_15242) );
NAND3_X2 inst_6481 ( .ZN(net_11241), .A2(net_11240), .A3(net_7404), .A1(net_2801) );
AOI22_X2 inst_20038 ( .ZN(net_7654), .B2(net_7653), .A2(net_6088), .B1(net_690), .A1(net_154) );
INV_X4 inst_14284 ( .ZN(net_7084), .A(net_6851) );
XNOR2_X2 inst_255 ( .B(net_21108), .ZN(net_17289), .A(net_16963) );
NOR3_X2 inst_2726 ( .ZN(net_13248), .A1(net_10531), .A3(net_9605), .A2(net_4985) );
NAND2_X2 inst_10555 ( .ZN(net_6722), .A2(net_6721), .A1(net_3031) );
NOR3_X2 inst_2674 ( .ZN(net_20310), .A1(net_13581), .A3(net_12396), .A2(net_9338) );
INV_X4 inst_14471 ( .ZN(net_11192), .A(net_4903) );
NAND2_X2 inst_10390 ( .A1(net_13444), .ZN(net_10747), .A2(net_5604) );
NAND2_X2 inst_10279 ( .ZN(net_7953), .A2(net_7952), .A1(net_3049) );
NAND3_X2 inst_6686 ( .ZN(net_7710), .A3(net_5621), .A1(net_3708), .A2(net_2620) );
NAND2_X2 inst_8784 ( .A1(net_16385), .ZN(net_15761), .A2(net_15400) );
OR2_X4 inst_1113 ( .ZN(net_2204), .A2(net_1697), .A1(net_193) );
CLKBUF_X2 inst_22190 ( .A(net_22061), .Z(net_22062) );
INV_X1 inst_19757 ( .A(net_7449), .ZN(net_5816) );
INV_X8 inst_12438 ( .A(net_20464), .ZN(net_20463) );
NOR2_X2 inst_4206 ( .A1(net_6672), .ZN(net_6671), .A2(net_6670) );
NAND4_X2 inst_5415 ( .ZN(net_14582), .A4(net_12156), .A3(net_11157), .A1(net_9959), .A2(net_8500) );
INV_X2 inst_18398 ( .ZN(net_16442), .A(net_16441) );
NAND2_X2 inst_8101 ( .ZN(net_20280), .A2(net_18118), .A1(net_17262) );
OAI21_X2 inst_2191 ( .A(net_14308), .ZN(net_8663), .B1(net_5011), .B2(net_4839) );
NAND4_X2 inst_5296 ( .ZN(net_15922), .A4(net_15165), .A2(net_14138), .A1(net_12188), .A3(net_10713) );
OR2_X4 inst_1127 ( .ZN(net_2964), .A2(net_170), .A1(net_90) );
INV_X8 inst_12184 ( .ZN(net_16864), .A(net_16496) );
XNOR2_X2 inst_362 ( .A(net_16885), .ZN(net_16880), .B(net_16879) );
INV_X4 inst_17013 ( .ZN(net_5097), .A(net_1138) );
AOI21_X2 inst_20327 ( .ZN(net_20172), .B2(net_15308), .A(net_14260), .B1(net_1402) );
INV_X2 inst_19036 ( .ZN(net_7811), .A(net_4926) );
INV_X2 inst_19336 ( .ZN(net_2475), .A(net_2474) );
XNOR2_X2 inst_306 ( .ZN(net_17094), .A(net_17086), .B(net_14420) );
NAND2_X2 inst_8662 ( .A2(net_20766), .ZN(net_18972), .A1(net_3433) );
CLKBUF_X2 inst_21412 ( .A(net_21248), .Z(net_21284) );
INV_X4 inst_13499 ( .A(net_10116), .ZN(net_9436) );
NAND2_X2 inst_9460 ( .ZN(net_11495), .A1(net_11494), .A2(net_9521) );
NOR2_X4 inst_3095 ( .ZN(net_4973), .A2(net_2828), .A1(net_2609) );
CLKBUF_X2 inst_21676 ( .A(net_21547), .Z(net_21548) );
NAND2_X2 inst_9884 ( .ZN(net_9426), .A2(net_9425), .A1(net_6592) );
OAI21_X2 inst_1715 ( .ZN(net_15190), .B2(net_13917), .B1(net_7243), .A(net_652) );
NAND3_X2 inst_6396 ( .ZN(net_11994), .A3(net_11837), .A1(net_9610), .A2(net_7935) );
AND2_X4 inst_21265 ( .ZN(net_4690), .A2(net_874), .A1(net_120) );
INV_X4 inst_16245 ( .ZN(net_2701), .A(net_1362) );
NAND2_X4 inst_7355 ( .ZN(net_13620), .A1(net_6445), .A2(net_3988) );
XNOR2_X2 inst_267 ( .ZN(net_17251), .A(net_16768), .B(net_360) );
INV_X4 inst_16630 ( .ZN(net_15744), .A(net_14476) );
INV_X4 inst_16100 ( .ZN(net_15659), .A(net_333) );
SDFF_X2 inst_716 ( .Q(net_20888), .SE(net_18863), .SI(net_18770), .D(net_395), .CK(net_22011) );
OAI21_X2 inst_1906 ( .ZN(net_13124), .B1(net_12370), .A(net_9914), .B2(net_6988) );
SDFF_X2 inst_792 ( .Q(net_20854), .SE(net_18577), .SI(net_18016), .D(net_600), .CK(net_22618) );
OAI21_X2 inst_2024 ( .ZN(net_11327), .A(net_10709), .B2(net_5802), .B1(net_5550) );
AOI21_X2 inst_20332 ( .ZN(net_15820), .B1(net_15706), .B2(net_14920), .A(net_8984) );
NAND2_X2 inst_9984 ( .ZN(net_8852), .A1(net_8851), .A2(net_6503) );
NAND2_X2 inst_9061 ( .ZN(net_13992), .A2(net_11990), .A1(net_1641) );
INV_X4 inst_16359 ( .ZN(net_12326), .A(net_6589) );
NAND2_X2 inst_10476 ( .ZN(net_10565), .A1(net_6981), .A2(net_6980) );
NAND2_X2 inst_8933 ( .ZN(net_14856), .A2(net_14146), .A1(net_10056) );
INV_X4 inst_16692 ( .A(net_3436), .ZN(net_1659) );
OAI21_X2 inst_2216 ( .ZN(net_8522), .A(net_8521), .B1(net_5752), .B2(net_4846) );
NOR2_X4 inst_2988 ( .ZN(net_8592), .A1(net_5934), .A2(net_5173) );
INV_X4 inst_15043 ( .A(net_4313), .ZN(net_4048) );
NOR2_X2 inst_4494 ( .ZN(net_4953), .A2(net_4041), .A1(net_222) );
OR2_X2 inst_1199 ( .ZN(net_3843), .A1(net_3842), .A2(net_3841) );
NAND2_X2 inst_11520 ( .A1(net_20542), .ZN(net_8164), .A2(net_2988) );
OAI21_X2 inst_1662 ( .A(net_20889), .ZN(net_15758), .B2(net_15057), .B1(net_11428) );
NAND2_X4 inst_7508 ( .ZN(net_4677), .A1(net_2535), .A2(net_1327) );
CLKBUF_X2 inst_22321 ( .A(net_22160), .Z(net_22193) );
CLKBUF_X2 inst_22146 ( .A(net_22017), .Z(net_22018) );
DFF_X1 inst_19893 ( .D(net_16941), .CK(net_21319), .Q(x205) );
INV_X4 inst_13240 ( .A(net_13562), .ZN(net_13398) );
NAND2_X2 inst_11251 ( .ZN(net_3917), .A1(net_2585), .A2(net_2323) );
OAI22_X2 inst_1285 ( .ZN(net_20685), .A1(net_14706), .A2(net_12477), .B2(net_5862), .B1(net_5557) );
XNOR2_X2 inst_380 ( .A(net_16846), .B(net_16833), .ZN(net_16830) );
AND2_X4 inst_21161 ( .ZN(net_13779), .A2(net_13778), .A1(net_10242) );
INV_X4 inst_14711 ( .ZN(net_14974), .A(net_14511) );
CLKBUF_X2 inst_22433 ( .A(net_22304), .Z(net_22305) );
INV_X4 inst_13508 ( .ZN(net_12991), .A(net_9411) );
INV_X2 inst_18688 ( .ZN(net_8609), .A(net_7185) );
NAND2_X4 inst_7423 ( .ZN(net_5914), .A2(net_4221), .A1(net_3009) );
NOR2_X2 inst_4970 ( .ZN(net_3757), .A2(net_1572), .A1(net_1330) );
INV_X4 inst_12583 ( .ZN(net_18299), .A(net_18183) );
SDFF_X2 inst_706 ( .Q(net_20894), .SE(net_18858), .SI(net_18831), .D(net_542), .CK(net_21313) );
INV_X4 inst_16137 ( .ZN(net_1917), .A(net_1474) );
INV_X4 inst_14692 ( .ZN(net_19267), .A(net_15027) );
NAND2_X2 inst_10874 ( .A1(net_12053), .ZN(net_5427), .A2(net_2958) );
NAND2_X2 inst_9834 ( .ZN(net_10988), .A1(net_7950), .A2(net_6027) );
INV_X4 inst_13366 ( .A(net_12900), .ZN(net_10910) );
NAND2_X2 inst_7985 ( .ZN(net_19946), .A1(net_18332), .A2(net_17326) );
NOR2_X2 inst_4734 ( .ZN(net_4145), .A2(net_3069), .A1(net_3068) );
INV_X4 inst_15033 ( .ZN(net_11359), .A(net_3360) );
INV_X4 inst_13055 ( .ZN(net_18919), .A(net_16332) );
XNOR2_X2 inst_110 ( .ZN(net_18514), .A(net_18387), .B(net_17161) );
INV_X4 inst_17927 ( .A(net_21104), .ZN(net_8967) );
OAI21_X2 inst_2047 ( .ZN(net_11060), .B1(net_6273), .B2(net_5844), .A(net_4261) );
INV_X2 inst_19295 ( .ZN(net_2816), .A(net_2815) );
NOR2_X2 inst_4545 ( .ZN(net_6939), .A1(net_3890), .A2(net_2878) );
NOR2_X2 inst_3825 ( .ZN(net_20053), .A1(net_9764), .A2(net_8507) );
INV_X4 inst_17740 ( .ZN(net_970), .A(net_177) );
INV_X4 inst_16291 ( .ZN(net_1738), .A(net_1334) );
NAND2_X2 inst_7876 ( .ZN(net_18531), .A2(net_18480), .A1(net_18453) );
NAND2_X2 inst_10842 ( .ZN(net_6760), .A2(net_5476), .A1(net_5475) );
NAND2_X2 inst_11927 ( .ZN(net_2908), .A1(net_2012), .A2(net_1495) );
NAND2_X2 inst_7846 ( .ZN(net_18606), .A2(net_18604), .A1(net_16492) );
INV_X4 inst_16741 ( .ZN(net_15499), .A(net_15044) );
NOR2_X4 inst_2949 ( .ZN(net_8151), .A1(net_6837), .A2(net_5570) );
OAI211_X2 inst_2414 ( .ZN(net_15507), .C1(net_15214), .B(net_14631), .C2(net_13248), .A(net_11921) );
INV_X4 inst_18224 ( .A(net_20905), .ZN(net_100) );
CLKBUF_X2 inst_22202 ( .A(net_21912), .Z(net_22074) );
INV_X2 inst_19359 ( .ZN(net_2308), .A(net_1835) );
INV_X2 inst_19318 ( .A(net_4508), .ZN(net_2623) );
AOI211_X2 inst_21068 ( .C1(net_9579), .ZN(net_8436), .B(net_4860), .C2(net_3781), .A(net_3361) );
NAND2_X2 inst_10429 ( .ZN(net_12240), .A2(net_6560), .A1(net_1182) );
AOI21_X2 inst_20398 ( .ZN(net_15430), .B2(net_14370), .A(net_10200), .B1(net_278) );
NAND2_X2 inst_11132 ( .ZN(net_7182), .A1(net_4323), .A2(net_4089) );
NAND2_X2 inst_7901 ( .ZN(net_18481), .A2(net_18426), .A1(net_17903) );
CLKBUF_X2 inst_21883 ( .A(net_21754), .Z(net_21755) );
INV_X4 inst_15189 ( .A(net_4184), .ZN(net_2936) );
CLKBUF_X2 inst_22900 ( .A(net_22771), .Z(net_22772) );
NAND2_X4 inst_6981 ( .ZN(net_17493), .A1(net_16917), .A2(net_16733) );
NAND2_X2 inst_11695 ( .A1(net_2744), .ZN(net_2318), .A2(net_1480) );
INV_X4 inst_14648 ( .ZN(net_18856), .A(net_18025) );
NAND2_X4 inst_7316 ( .ZN(net_8398), .A1(net_4785), .A2(net_809) );
CLKBUF_X2 inst_22793 ( .A(net_21650), .Z(net_22665) );
INV_X4 inst_16619 ( .A(net_1608), .ZN(net_1117) );
AOI22_X2 inst_19986 ( .A1(net_20670), .ZN(net_15168), .B2(net_13300), .B1(net_11776), .A2(net_11407) );
INV_X1 inst_19754 ( .ZN(net_9097), .A(net_9096) );
INV_X4 inst_14440 ( .ZN(net_6281), .A(net_4994) );
SDFF_X2 inst_889 ( .Q(net_21196), .SI(net_16890), .SE(net_125), .CK(net_22145), .D(x6203) );
NAND2_X2 inst_8935 ( .ZN(net_14852), .A2(net_14150), .A1(net_10379) );
AOI21_X2 inst_20735 ( .ZN(net_11736), .B2(net_11735), .B1(net_11612), .A(net_7531) );
NAND2_X2 inst_8533 ( .A1(net_17025), .ZN(net_16862), .A2(net_16669) );
AND2_X4 inst_21179 ( .ZN(net_11600), .A2(net_11547), .A1(net_8826) );
INV_X4 inst_16302 ( .A(net_3086), .ZN(net_2321) );
INV_X8 inst_12457 ( .A(net_20778), .ZN(net_20776) );
NAND4_X4 inst_5188 ( .A4(net_19013), .A1(net_19012), .ZN(net_16579), .A3(net_16142), .A2(net_15440) );
OAI211_X4 inst_2379 ( .B(net_19901), .A(net_19900), .ZN(net_19762), .C1(net_15340), .C2(net_11363) );
AND2_X4 inst_21259 ( .ZN(net_4358), .A1(net_1660), .A2(net_573) );
NAND2_X2 inst_10358 ( .ZN(net_10623), .A1(net_6945), .A2(net_5850) );
NAND2_X2 inst_8774 ( .ZN(net_19256), .A2(net_15617), .A1(net_15569) );
AOI21_X2 inst_20905 ( .ZN(net_7694), .B2(net_4630), .A(net_2885), .B1(net_1846) );
NAND2_X2 inst_11754 ( .A1(net_4394), .ZN(net_3957), .A2(net_2109) );
NAND2_X2 inst_11244 ( .ZN(net_3927), .A2(net_2742), .A1(net_154) );
INV_X4 inst_15047 ( .ZN(net_4877), .A(net_3882) );
INV_X4 inst_16275 ( .ZN(net_15831), .A(net_15191) );
NAND2_X2 inst_10382 ( .ZN(net_9107), .A1(net_8868), .A2(net_4459) );
NOR2_X2 inst_4916 ( .A2(net_20489), .ZN(net_1888), .A1(net_1308) );
CLKBUF_X2 inst_22782 ( .A(net_22653), .Z(net_22654) );
AND2_X4 inst_21190 ( .ZN(net_19531), .A1(net_14092), .A2(net_10732) );
NAND2_X2 inst_8149 ( .ZN(net_18015), .A1(net_17968), .A2(net_17939) );
NOR2_X2 inst_3571 ( .ZN(net_19170), .A1(net_12345), .A2(net_11677) );
INV_X4 inst_15757 ( .ZN(net_14279), .A(net_10405) );
NAND3_X2 inst_6132 ( .ZN(net_13739), .A1(net_12883), .A2(net_11080), .A3(net_7926) );
OR2_X2 inst_1190 ( .A1(net_13080), .ZN(net_4352), .A2(net_4351) );
XNOR2_X2 inst_444 ( .B(net_21115), .ZN(net_15586), .A(net_15585) );
NAND2_X2 inst_8865 ( .ZN(net_15329), .A2(net_14497), .A1(net_12656) );
NAND2_X4 inst_7489 ( .A2(net_20559), .A1(net_19425), .ZN(net_6461) );
NAND2_X2 inst_8246 ( .ZN(net_17717), .A2(net_17708), .A1(net_16951) );
INV_X4 inst_12816 ( .ZN(net_17197), .A(net_17196) );
NAND2_X2 inst_9064 ( .ZN(net_13989), .A2(net_11982), .A1(net_10709) );
NAND2_X2 inst_10033 ( .A1(net_10728), .ZN(net_8728), .A2(net_8727) );
INV_X4 inst_14196 ( .ZN(net_11168), .A(net_4809) );
NAND2_X2 inst_8705 ( .A1(net_21228), .ZN(net_16304), .A2(net_16132) );
AOI211_X2 inst_21037 ( .C1(net_14166), .ZN(net_14120), .C2(net_11196), .A(net_9172), .B(net_5947) );
NAND2_X2 inst_11720 ( .A1(net_6617), .ZN(net_2256), .A2(net_2255) );
AND2_X4 inst_21182 ( .A2(net_12737), .ZN(net_11581), .A1(net_11580) );
INV_X2 inst_19410 ( .A(net_2899), .ZN(net_1975) );
INV_X2 inst_18612 ( .ZN(net_11048), .A(net_10254) );
AOI21_X2 inst_20667 ( .ZN(net_12912), .B1(net_12911), .B2(net_9429), .A(net_8276) );
NAND3_X2 inst_5833 ( .ZN(net_15514), .A2(net_14721), .A1(net_14646), .A3(net_14564) );
NAND2_X2 inst_12047 ( .ZN(net_1276), .A2(net_937), .A1(net_221) );
XNOR2_X2 inst_119 ( .B(net_20507), .ZN(net_18501), .A(net_18354) );
NOR2_X4 inst_3181 ( .ZN(net_5467), .A2(net_1872), .A1(net_170) );
SDFF_X2 inst_939 ( .QN(net_21045), .D(net_743), .SE(net_263), .CK(net_22531), .SI(x2249) );
NAND2_X2 inst_9722 ( .ZN(net_15211), .A1(net_10151), .A2(net_10150) );
INV_X4 inst_17912 ( .ZN(net_4268), .A(net_156) );
NAND2_X2 inst_10770 ( .A1(net_11050), .ZN(net_5630), .A2(net_4128) );
CLKBUF_X2 inst_22463 ( .A(net_22334), .Z(net_22335) );
INV_X2 inst_18609 ( .ZN(net_19783), .A(net_9711) );
NAND2_X2 inst_8205 ( .ZN(net_17915), .A2(net_17712), .A1(net_17619) );
INV_X2 inst_19425 ( .ZN(net_1817), .A(net_1142) );
INV_X4 inst_15389 ( .ZN(net_14962), .A(net_6934) );
SDFF_X2 inst_1019 ( .QN(net_21008), .D(net_565), .SE(net_263), .CK(net_21834), .SI(x2945) );
INV_X4 inst_17364 ( .A(net_949), .ZN(net_873) );
INV_X4 inst_13490 ( .A(net_12945), .ZN(net_9515) );
INV_X4 inst_16748 ( .ZN(net_2258), .A(net_1042) );
INV_X4 inst_15672 ( .ZN(net_2624), .A(net_2052) );
OAI21_X2 inst_1827 ( .B2(net_19797), .B1(net_19796), .ZN(net_19789), .A(net_816) );
NAND2_X2 inst_10830 ( .ZN(net_6772), .A1(net_5572), .A2(net_5451) );
SDFF_X2 inst_742 ( .Q(net_20970), .SE(net_18581), .SI(net_18543), .D(net_13663), .CK(net_22754) );
INV_X2 inst_19496 ( .A(net_1753), .ZN(net_1280) );
INV_X4 inst_13372 ( .ZN(net_14454), .A(net_10896) );
NOR2_X2 inst_4481 ( .ZN(net_4349), .A1(net_4348), .A2(net_4347) );
INV_X4 inst_17888 ( .ZN(net_10702), .A(net_10216) );
INV_X4 inst_13545 ( .ZN(net_10764), .A(net_9190) );
NAND2_X4 inst_7345 ( .ZN(net_7232), .A1(net_4840), .A2(net_3560) );
NAND4_X2 inst_5289 ( .A2(net_20645), .A1(net_20644), .ZN(net_15938), .A4(net_15416), .A3(net_14359) );
NAND2_X2 inst_9121 ( .A2(net_20078), .ZN(net_13557), .A1(net_13556) );
OAI21_X2 inst_1955 ( .A(net_20486), .ZN(net_12537), .B1(net_10080), .B2(net_9642) );
AOI211_X2 inst_21030 ( .ZN(net_14539), .B(net_11750), .A(net_11322), .C2(net_10564), .C1(net_5166) );
INV_X4 inst_18287 ( .A(net_20210), .ZN(net_20209) );
NOR2_X2 inst_3618 ( .ZN(net_12359), .A2(net_10744), .A1(net_7454) );
INV_X4 inst_17533 ( .ZN(net_1019), .A(net_884) );
INV_X4 inst_14807 ( .ZN(net_3975), .A(net_3974) );
INV_X4 inst_14430 ( .ZN(net_5030), .A(net_5029) );
INV_X4 inst_14945 ( .A(net_5013), .ZN(net_3518) );
NAND2_X2 inst_9181 ( .ZN(net_13318), .A1(net_10545), .A2(net_10363) );
NAND2_X2 inst_9781 ( .ZN(net_12957), .A2(net_9793), .A1(net_7075) );
NOR3_X2 inst_2704 ( .A3(net_15110), .ZN(net_13921), .A2(net_12546), .A1(net_12017) );
NAND2_X2 inst_8349 ( .A1(net_19453), .ZN(net_17473), .A2(net_17472) );
NAND2_X2 inst_11461 ( .ZN(net_5469), .A2(net_3194), .A1(net_2683) );
INV_X2 inst_18828 ( .ZN(net_6796), .A(net_6795) );
NAND3_X2 inst_5924 ( .ZN(net_14980), .A1(net_14050), .A3(net_13970), .A2(net_4684) );
INV_X4 inst_14551 ( .ZN(net_7167), .A(net_4591) );
INV_X4 inst_13327 ( .ZN(net_11239), .A(net_9924) );
NAND2_X2 inst_9508 ( .ZN(net_11329), .A2(net_8307), .A1(net_81) );
INV_X4 inst_16355 ( .ZN(net_1493), .A(net_1293) );
NAND2_X2 inst_9701 ( .A2(net_11943), .A1(net_11091), .ZN(net_10212) );
NAND4_X2 inst_5473 ( .ZN(net_13202), .A3(net_13201), .A2(net_12125), .A1(net_11029), .A4(net_6448) );
INV_X4 inst_15014 ( .ZN(net_16050), .A(net_15561) );
INV_X4 inst_18290 ( .ZN(net_20216), .A(net_20215) );
NOR2_X2 inst_4817 ( .ZN(net_3901), .A1(net_2563), .A2(net_2562) );
NOR2_X2 inst_4456 ( .ZN(net_5856), .A1(net_4672), .A2(net_1439) );
NOR2_X2 inst_4926 ( .ZN(net_2158), .A1(net_2001), .A2(net_1258) );
NAND2_X4 inst_6846 ( .A2(net_19766), .A1(net_19765), .ZN(net_18696) );
INV_X4 inst_13840 ( .A(net_7484), .ZN(net_7483) );
NOR2_X2 inst_4571 ( .ZN(net_4848), .A1(net_3865), .A2(net_3762) );
NOR2_X2 inst_5111 ( .A2(net_21219), .ZN(net_658), .A1(net_396) );
NOR2_X2 inst_3928 ( .A1(net_14881), .ZN(net_8745), .A2(net_8053) );
DFF_X1 inst_19875 ( .D(net_17020), .CK(net_22093), .Q(x452) );
INV_X8 inst_12212 ( .ZN(net_14642), .A(net_5098) );
NAND2_X2 inst_11849 ( .ZN(net_2836), .A1(net_1699), .A2(net_1636) );
NOR2_X2 inst_4017 ( .A1(net_13752), .ZN(net_8034), .A2(net_8033) );
NAND2_X4 inst_7121 ( .ZN(net_12614), .A1(net_11067), .A2(net_8369) );
INV_X2 inst_19054 ( .ZN(net_4731), .A(net_4730) );
INV_X4 inst_16917 ( .A(net_3886), .ZN(net_3805) );
AOI221_X2 inst_20088 ( .C1(net_16076), .ZN(net_15676), .B1(net_15481), .C2(net_14436), .B2(net_13187), .A(net_6667) );
INV_X2 inst_18723 ( .ZN(net_8106), .A(net_8105) );
NOR2_X2 inst_5135 ( .A2(net_525), .ZN(net_186), .A1(net_132) );
INV_X4 inst_17216 ( .ZN(net_2985), .A(net_2375) );
INV_X4 inst_12879 ( .ZN(net_16896), .A(net_16706) );
INV_X4 inst_13050 ( .A(net_16602), .ZN(net_16384) );
DFF_X1 inst_19787 ( .D(net_18660), .CK(net_21630), .Q(x522) );
NAND3_X2 inst_5760 ( .ZN(net_15980), .A3(net_15590), .A2(net_15111), .A1(net_14635) );
INV_X2 inst_19371 ( .ZN(net_2207), .A(net_2206) );
NAND2_X4 inst_7556 ( .ZN(net_2433), .A1(net_1730), .A2(net_299) );
NAND2_X2 inst_11513 ( .ZN(net_2999), .A2(net_1531), .A1(net_1235) );
CLKBUF_X2 inst_22631 ( .A(net_22033), .Z(net_22503) );
NAND2_X4 inst_7037 ( .A2(net_19963), .A1(net_19962), .ZN(net_17086) );
NAND2_X4 inst_7294 ( .ZN(net_11943), .A1(net_5574), .A2(net_4288) );
NOR2_X2 inst_5095 ( .ZN(net_1291), .A2(net_734), .A1(net_222) );
CLKBUF_X2 inst_21668 ( .A(net_21539), .Z(net_21540) );
INV_X4 inst_14591 ( .ZN(net_13157), .A(net_6295) );
INV_X4 inst_17760 ( .ZN(net_657), .A(net_159) );
INV_X4 inst_17905 ( .A(net_2274), .ZN(net_260) );
INV_X2 inst_18636 ( .A(net_12076), .ZN(net_9393) );
XNOR2_X2 inst_426 ( .ZN(net_16502), .A(net_16501), .B(net_1675) );
NAND3_X2 inst_6035 ( .ZN(net_14335), .A2(net_14334), .A3(net_14333), .A1(net_11507) );
INV_X4 inst_13856 ( .ZN(net_9137), .A(net_7463) );
NOR2_X2 inst_4302 ( .ZN(net_5939), .A2(net_3503), .A1(net_1182) );
NAND2_X2 inst_11654 ( .ZN(net_2440), .A2(net_253), .A1(x7413) );
NAND2_X2 inst_11068 ( .ZN(net_4515), .A2(net_3194), .A1(net_2641) );
NAND2_X2 inst_8092 ( .ZN(net_18130), .A2(net_18129), .A1(net_17526) );
CLKBUF_X2 inst_22385 ( .A(net_21947), .Z(net_22257) );
NAND3_X2 inst_6560 ( .ZN(net_10491), .A2(net_9911), .A1(net_7267), .A3(net_3809) );
NAND2_X2 inst_7725 ( .ZN(net_18831), .A2(net_18794), .A1(net_18779) );
AOI21_X2 inst_20528 ( .B1(net_15450), .ZN(net_14531), .B2(net_11825), .A(net_10110) );
NAND3_X2 inst_6341 ( .ZN(net_12253), .A1(net_9062), .A2(net_5760), .A3(net_1052) );
AOI21_X2 inst_20717 ( .ZN(net_19051), .A(net_8529), .B2(net_7708), .B1(net_1202) );
INV_X4 inst_16875 ( .ZN(net_14689), .A(net_320) );
AND2_X2 inst_21280 ( .ZN(net_13432), .A2(net_13431), .A1(net_7873) );
NAND2_X2 inst_11163 ( .ZN(net_9082), .A2(net_5327), .A1(net_952) );
NAND2_X2 inst_8544 ( .A1(net_20074), .ZN(net_19104), .A2(net_17370) );
NAND2_X2 inst_9247 ( .ZN(net_12671), .A2(net_10983), .A1(net_8732) );
AOI22_X2 inst_20047 ( .A1(net_8639), .ZN(net_4656), .B2(net_4655), .A2(net_4203), .B1(net_2219) );
NAND2_X2 inst_9904 ( .ZN(net_10880), .A2(net_7466), .A1(net_1187) );
INV_X4 inst_15182 ( .ZN(net_3873), .A(net_2298) );
INV_X4 inst_12558 ( .ZN(net_18365), .A(net_18310) );
NAND2_X2 inst_8136 ( .ZN(net_18034), .A1(net_18020), .A2(net_17999) );
INV_X4 inst_15645 ( .ZN(net_11902), .A(net_2116) );
INV_X2 inst_19055 ( .ZN(net_4728), .A(net_4727) );
NOR2_X2 inst_4211 ( .A1(net_9018), .ZN(net_7925), .A2(net_5113) );
AND4_X2 inst_21106 ( .ZN(net_11802), .A2(net_11801), .A3(net_11800), .A4(net_11799), .A1(net_7835) );
OAI21_X2 inst_1745 ( .ZN(net_14950), .A(net_14949), .B2(net_12727), .B1(net_11398) );
NOR2_X2 inst_3831 ( .ZN(net_9729), .A1(net_9728), .A2(net_9056) );
OAI21_X2 inst_2079 ( .B1(net_15950), .ZN(net_10537), .A(net_10536), .B2(net_6596) );
NAND2_X2 inst_10534 ( .A2(net_9558), .A1(net_8952), .ZN(net_6813) );
INV_X4 inst_15506 ( .A(net_3697), .ZN(net_3321) );
NAND3_X2 inst_6819 ( .A2(net_3493), .ZN(net_2857), .A3(net_1334), .A1(net_606) );
INV_X2 inst_19106 ( .ZN(net_4494), .A(net_4493) );
INV_X4 inst_18057 ( .A(net_20928), .ZN(net_16187) );
INV_X4 inst_14883 ( .ZN(net_3672), .A(net_3671) );
NAND2_X2 inst_9299 ( .ZN(net_12391), .A1(net_12330), .A2(net_9219) );
INV_X2 inst_19120 ( .A(net_14141), .ZN(net_4432) );
INV_X4 inst_14053 ( .ZN(net_9824), .A(net_8014) );
NAND3_X2 inst_6554 ( .ZN(net_10526), .A2(net_10525), .A3(net_10524), .A1(net_8578) );
NAND3_X4 inst_5615 ( .ZN(net_19235), .A2(net_9607), .A1(net_7959), .A3(net_7269) );
INV_X4 inst_14729 ( .ZN(net_13673), .A(net_4120) );
NAND2_X2 inst_12081 ( .A2(net_2919), .ZN(net_1633), .A1(net_195) );
OAI211_X2 inst_2596 ( .C2(net_5673), .C1(net_5616), .ZN(net_5253), .B(net_5252), .A(net_3907) );
INV_X2 inst_18575 ( .ZN(net_10657), .A(net_9095) );
NAND3_X2 inst_6599 ( .ZN(net_9893), .A2(net_7459), .A3(net_5587), .A1(net_4889) );
NAND3_X2 inst_6242 ( .A2(net_14145), .ZN(net_13180), .A3(net_13179), .A1(net_7225) );
NAND2_X2 inst_8579 ( .A2(net_16742), .ZN(net_16725), .A1(net_16724) );
NOR2_X4 inst_3022 ( .A2(net_6736), .ZN(net_6622), .A1(net_3873) );
NAND2_X1 inst_12133 ( .ZN(net_18209), .A1(net_18208), .A2(net_18168) );
XNOR2_X1 inst_680 ( .ZN(net_18193), .A(net_18192), .B(net_11880) );
NAND3_X2 inst_6575 ( .A3(net_10534), .ZN(net_10455), .A2(net_10454), .A1(net_4703) );
CLKBUF_X2 inst_22197 ( .A(net_22068), .Z(net_22069) );
CLKBUF_X2 inst_22741 ( .A(net_21882), .Z(net_22613) );
NAND2_X2 inst_10323 ( .ZN(net_11795), .A1(net_9591), .A2(net_6014) );
NOR2_X4 inst_3299 ( .A2(net_20559), .ZN(net_2144), .A1(net_1242) );
CLKBUF_X2 inst_21722 ( .A(net_21593), .Z(net_21594) );
INV_X4 inst_16565 ( .ZN(net_6682), .A(net_1790) );
NAND2_X2 inst_7820 ( .A1(net_21154), .ZN(net_19232), .A2(net_18648) );
NAND2_X4 inst_7065 ( .A2(net_20904), .A1(net_19470), .ZN(net_16246) );
INV_X4 inst_15717 ( .ZN(net_14554), .A(net_13070) );
NAND2_X4 inst_7643 ( .ZN(net_2045), .A2(net_1192), .A1(net_1158) );
AOI21_X4 inst_20174 ( .B2(net_20242), .B1(net_20241), .ZN(net_15545), .A(net_15362) );
CLKBUF_X2 inst_22288 ( .A(net_22159), .Z(net_22160) );
NAND2_X4 inst_7551 ( .A2(net_1934), .ZN(net_1863), .A1(net_1509) );
INV_X4 inst_12697 ( .ZN(net_19719), .A(net_17632) );
NOR2_X2 inst_3567 ( .ZN(net_12824), .A2(net_10224), .A1(net_8818) );
INV_X4 inst_16223 ( .ZN(net_10765), .A(net_6733) );
XNOR2_X2 inst_414 ( .ZN(net_16703), .A(net_16569), .B(net_16546) );
INV_X4 inst_18261 ( .A(net_19432), .ZN(net_19430) );
XNOR2_X2 inst_531 ( .ZN(net_2418), .A(net_979), .B(net_28) );
NAND2_X2 inst_9315 ( .A1(net_13752), .ZN(net_12351), .A2(net_9016) );
OAI21_X2 inst_1952 ( .ZN(net_12555), .A(net_11087), .B2(net_7535), .B1(net_3786) );
CLKBUF_X2 inst_22074 ( .A(net_21614), .Z(net_21946) );
NAND2_X2 inst_8827 ( .ZN(net_15540), .A1(net_15071), .A2(net_14862) );
NAND3_X2 inst_6060 ( .ZN(net_14194), .A2(net_14193), .A1(net_13425), .A3(net_8216) );
INV_X2 inst_19648 ( .A(net_19459), .ZN(net_19458) );
CLKBUF_X2 inst_21973 ( .A(net_21844), .Z(net_21845) );
NOR2_X2 inst_5023 ( .A1(net_3704), .ZN(net_1180), .A2(net_647) );
NAND3_X4 inst_5617 ( .ZN(net_19528), .A2(net_11984), .A1(net_11983), .A3(net_5930) );
NOR2_X2 inst_3698 ( .ZN(net_11137), .A2(net_7405), .A1(net_7035) );
NOR2_X2 inst_4155 ( .ZN(net_6894), .A2(net_6893), .A1(net_1458) );
NAND2_X4 inst_6962 ( .A2(net_19886), .A1(net_19885), .ZN(net_17430) );
NOR2_X2 inst_5118 ( .ZN(net_316), .A1(net_103), .A2(net_53) );
INV_X4 inst_14223 ( .ZN(net_9162), .A(net_7167) );
NAND2_X2 inst_9686 ( .ZN(net_11591), .A1(net_10248), .A2(net_10247) );
INV_X4 inst_15102 ( .A(net_9668), .ZN(net_3754) );
NAND2_X2 inst_10208 ( .ZN(net_13632), .A1(net_9324), .A2(net_7992) );
INV_X4 inst_16944 ( .ZN(net_1599), .A(net_919) );
INV_X4 inst_17771 ( .ZN(net_3842), .A(net_3789) );
NAND2_X2 inst_10699 ( .ZN(net_8919), .A2(net_6044), .A1(net_3818) );
NAND4_X2 inst_5338 ( .A4(net_20017), .A1(net_20016), .ZN(net_15504), .A2(net_11652), .A3(net_9492) );
XNOR2_X2 inst_570 ( .B(net_16839), .ZN(net_635), .A(net_634) );
AOI211_X2 inst_21075 ( .ZN(net_7680), .B(net_7679), .C2(net_4612), .C1(net_3027), .A(net_2777) );
OAI21_X2 inst_1570 ( .ZN(net_16403), .A(net_16402), .B2(net_16256), .B1(net_14064) );
INV_X4 inst_14697 ( .ZN(net_9623), .A(net_4266) );
INV_X4 inst_16424 ( .ZN(net_8785), .A(net_8361) );
NAND2_X2 inst_12055 ( .A2(net_4394), .ZN(net_1326), .A1(net_895) );
OAI21_X2 inst_1612 ( .B2(net_19595), .B1(net_19594), .A(net_16394), .ZN(net_16112) );
NOR2_X2 inst_4645 ( .ZN(net_6944), .A2(net_3986), .A1(net_3385) );
INV_X4 inst_16054 ( .ZN(net_2457), .A(net_1163) );
INV_X4 inst_12545 ( .ZN(net_18393), .A(net_18328) );
CLKBUF_X2 inst_22077 ( .A(net_21948), .Z(net_21949) );
INV_X4 inst_15649 ( .ZN(net_3819), .A(net_1419) );
INV_X4 inst_17295 ( .ZN(net_975), .A(net_673) );
CLKBUF_X2 inst_21561 ( .A(net_21432), .Z(net_21433) );
NAND2_X2 inst_11419 ( .ZN(net_3382), .A1(net_3381), .A2(net_3380) );
AOI21_X2 inst_20271 ( .ZN(net_19555), .B1(net_16404), .B2(net_16129), .A(net_16086) );
AOI21_X2 inst_20826 ( .ZN(net_9866), .B1(net_7915), .B2(net_5993), .A(net_3502) );
NOR2_X2 inst_3718 ( .ZN(net_19585), .A1(net_10976), .A2(net_10975) );
INV_X4 inst_12592 ( .ZN(net_18166), .A(net_18116) );
NOR2_X4 inst_3077 ( .A1(net_19671), .ZN(net_9974), .A2(net_4726) );
INV_X2 inst_18675 ( .ZN(net_9112), .A(net_9111) );
AND3_X2 inst_21146 ( .ZN(net_6442), .A1(net_6441), .A2(net_6440), .A3(net_6439) );
INV_X4 inst_15905 ( .ZN(net_2018), .A(net_1765) );
INV_X2 inst_19208 ( .A(net_5010), .ZN(net_3523) );
INV_X4 inst_12599 ( .ZN(net_18095), .A(net_18094) );
NAND4_X4 inst_5224 ( .A3(net_18945), .A1(net_18944), .ZN(net_16382), .A2(net_16109), .A4(net_16089) );
NAND2_X2 inst_8099 ( .A2(net_20217), .ZN(net_18121), .A1(net_16522) );
NAND2_X2 inst_9566 ( .A1(net_12100), .A2(net_11104), .ZN(net_10965) );
OAI21_X4 inst_1423 ( .A(net_20928), .B2(net_19354), .B1(net_19353), .ZN(net_16089) );
SDFF_X2 inst_1034 ( .QN(net_21076), .D(net_665), .SE(net_253), .CK(net_21703), .SI(x1781) );
INV_X4 inst_15448 ( .A(net_3030), .ZN(net_2770) );
NAND2_X2 inst_9855 ( .A1(net_20475), .ZN(net_9513), .A2(net_9512) );
OR2_X2 inst_1207 ( .ZN(net_20696), .A2(net_13002), .A1(net_7004) );
CLKBUF_X2 inst_22454 ( .A(net_22325), .Z(net_22326) );
INV_X4 inst_14492 ( .ZN(net_14145), .A(net_4846) );
XNOR2_X2 inst_613 ( .B(net_17294), .ZN(net_497), .A(net_496) );
NAND2_X2 inst_9945 ( .ZN(net_9036), .A1(net_9035), .A2(net_5695) );
NOR2_X2 inst_4275 ( .ZN(net_9654), .A2(net_6122), .A1(net_1958) );
NAND2_X2 inst_8694 ( .ZN(net_19111), .A1(net_16359), .A2(net_16197) );
NAND3_X2 inst_6444 ( .A2(net_13617), .ZN(net_11798), .A1(net_9440), .A3(net_8127) );
XNOR2_X2 inst_483 ( .A(net_16095), .ZN(net_10803), .B(net_5791) );
INV_X4 inst_16186 ( .ZN(net_1423), .A(net_1422) );
NOR2_X2 inst_5005 ( .A1(net_2071), .ZN(net_1667), .A2(net_1330) );
NAND2_X2 inst_9907 ( .A1(net_13938), .A2(net_12757), .ZN(net_9337) );
XNOR2_X2 inst_259 ( .B(net_21141), .ZN(net_17276), .A(net_17275) );
INV_X4 inst_17652 ( .ZN(net_6867), .A(net_270) );
NAND2_X4 inst_6845 ( .ZN(net_20210), .A1(net_18634), .A2(net_18619) );
INV_X4 inst_17659 ( .ZN(net_2955), .A(net_1655) );
NAND3_X2 inst_6812 ( .ZN(net_2390), .A1(net_2389), .A3(net_2388), .A2(net_1363) );
CLKBUF_X2 inst_22315 ( .A(net_21480), .Z(net_22187) );
NOR2_X2 inst_4707 ( .A1(net_3780), .ZN(net_3163), .A2(net_3162) );
NOR2_X2 inst_4846 ( .ZN(net_4339), .A1(net_1665), .A2(net_621) );
CLKBUF_X2 inst_22913 ( .A(net_21366), .Z(net_22785) );
NAND2_X2 inst_8621 ( .A1(net_21173), .ZN(net_16606), .A2(net_16605) );
NAND2_X4 inst_7592 ( .ZN(net_2038), .A2(net_212), .A1(net_123) );
INV_X4 inst_13197 ( .ZN(net_13950), .A(net_13949) );
NAND2_X2 inst_10517 ( .A1(net_10206), .ZN(net_8912), .A2(net_6875) );
CLKBUF_X2 inst_21471 ( .A(net_21342), .Z(net_21343) );
INV_X2 inst_19465 ( .A(net_6537), .ZN(net_1464) );
NAND2_X2 inst_10686 ( .A1(net_6930), .ZN(net_6120), .A2(net_6119) );
INV_X4 inst_16217 ( .ZN(net_1392), .A(net_1391) );
SDFF_X2 inst_894 ( .Q(net_21167), .SI(net_16891), .SE(net_125), .CK(net_21449), .D(x5015) );
INV_X2 inst_19083 ( .ZN(net_7503), .A(net_4583) );
OAI211_X2 inst_2425 ( .ZN(net_20661), .A(net_15211), .B(net_14091), .C2(net_2873), .C1(net_2368) );
CLKBUF_X2 inst_22619 ( .A(net_21344), .Z(net_22491) );
INV_X4 inst_16645 ( .A(net_4464), .ZN(net_4155) );
SDFF_X2 inst_994 ( .QN(net_21074), .D(net_671), .SE(net_263), .CK(net_21727), .SI(x1845) );
NAND2_X2 inst_9803 ( .ZN(net_20010), .A1(net_9695), .A2(net_6612) );
OAI21_X2 inst_1879 ( .ZN(net_13660), .B1(net_13659), .B2(net_13091), .A(net_7005) );
CLKBUF_X2 inst_22602 ( .A(net_22148), .Z(net_22474) );
OAI21_X2 inst_1863 ( .ZN(net_20834), .A(net_13343), .B1(net_11022), .B2(net_8001) );
OAI21_X2 inst_2135 ( .ZN(net_20247), .B1(net_9152), .B2(net_6940), .A(net_4032) );
INV_X4 inst_17439 ( .ZN(net_920), .A(net_267) );
INV_X4 inst_14082 ( .ZN(net_13966), .A(net_6217) );
INV_X2 inst_19235 ( .A(net_15926), .ZN(net_3338) );
SDFF_X2 inst_764 ( .Q(net_20867), .SE(net_18856), .SI(net_18514), .D(net_470), .CK(net_22333) );
INV_X4 inst_17764 ( .ZN(net_2746), .A(net_965) );
NAND2_X2 inst_10961 ( .A1(net_8674), .ZN(net_5072), .A2(net_5071) );
NAND2_X2 inst_12015 ( .ZN(net_1710), .A2(net_1142), .A1(net_1056) );
OAI21_X2 inst_1547 ( .ZN(net_17758), .A(net_17514), .B1(net_17513), .B2(net_17512) );
AOI21_X4 inst_20247 ( .B1(net_20409), .ZN(net_9873), .B2(net_6856), .A(net_3044) );
NAND2_X2 inst_11745 ( .ZN(net_4118), .A2(net_2141), .A1(net_1048) );
OAI211_X4 inst_2369 ( .C2(net_20960), .C1(net_19677), .ZN(net_17045), .B(net_16178), .A(net_9608) );
INV_X2 inst_18482 ( .ZN(net_12548), .A(net_11334) );
NAND3_X2 inst_6105 ( .ZN(net_13897), .A3(net_12129), .A1(net_11419), .A2(net_8235) );
OAI22_X2 inst_1274 ( .A2(net_16778), .ZN(net_16758), .B2(net_16757), .A1(net_11882), .B1(net_8774) );
NOR2_X2 inst_3838 ( .ZN(net_11574), .A2(net_7499), .A1(net_5415) );
INV_X4 inst_16444 ( .ZN(net_1802), .A(net_871) );
NAND4_X2 inst_5495 ( .ZN(net_12220), .A3(net_11659), .A2(net_11589), .A1(net_11167), .A4(net_8538) );
NAND4_X2 inst_5326 ( .ZN(net_20084), .A4(net_14970), .A2(net_14337), .A1(net_14072), .A3(net_13787) );
INV_X4 inst_14847 ( .A(net_5434), .ZN(net_5041) );
NAND2_X4 inst_7237 ( .A1(net_10034), .ZN(net_8832), .A2(net_6968) );
NOR2_X4 inst_2831 ( .ZN(net_19334), .A2(net_15597), .A1(net_15098) );
INV_X4 inst_12785 ( .A(net_17576), .ZN(net_17299) );
CLKBUF_X2 inst_22865 ( .A(net_22736), .Z(net_22737) );
OAI22_X2 inst_1300 ( .ZN(net_11267), .B1(net_10737), .A1(net_9276), .A2(net_5863), .B2(net_4077) );
NAND2_X2 inst_12022 ( .ZN(net_1029), .A2(net_809), .A1(net_114) );
NAND4_X2 inst_5317 ( .ZN(net_15775), .A1(net_15065), .A4(net_14977), .A3(net_14893), .A2(net_14474) );
INV_X4 inst_13698 ( .ZN(net_9455), .A(net_7919) );
AOI21_X2 inst_20639 ( .ZN(net_13273), .B1(net_10031), .B2(net_9982), .A(net_9560) );
INV_X4 inst_13693 ( .ZN(net_14214), .A(net_4822) );
AOI21_X4 inst_20101 ( .ZN(net_18974), .B1(net_16347), .A(net_16277), .B2(net_16231) );
NAND2_X4 inst_7309 ( .ZN(net_11984), .A2(net_7941), .A1(net_5521) );
INV_X4 inst_15284 ( .ZN(net_2724), .A(net_2723) );
OAI21_X2 inst_2279 ( .ZN(net_7126), .B2(net_7125), .A(net_5785), .B1(net_2282) );
INV_X4 inst_12572 ( .ZN(net_18295), .A(net_18258) );
CLKBUF_X2 inst_21704 ( .A(net_21575), .Z(net_21576) );
OAI21_X2 inst_2038 ( .ZN(net_11301), .A(net_11300), .B2(net_8476), .B1(net_4995) );
OAI21_X2 inst_2044 ( .B2(net_13442), .ZN(net_11187), .B1(net_11186), .A(net_6619) );
INV_X2 inst_19109 ( .ZN(net_4467), .A(net_4466) );
INV_X2 inst_19529 ( .ZN(net_1454), .A(net_1031) );
NAND2_X2 inst_7833 ( .ZN(net_18635), .A1(net_18633), .A2(net_18612) );
INV_X4 inst_15820 ( .A(net_4088), .ZN(net_2550) );
INV_X4 inst_15289 ( .ZN(net_14515), .A(net_14496) );
AND2_X2 inst_21287 ( .ZN(net_12685), .A2(net_12657), .A1(net_8973) );
INV_X4 inst_13630 ( .ZN(net_9756), .A(net_8303) );
CLKBUF_X2 inst_22606 ( .A(net_22477), .Z(net_22478) );
NAND3_X2 inst_6249 ( .ZN(net_13015), .A1(net_13014), .A3(net_11900), .A2(net_11126) );
INV_X2 inst_19712 ( .A(net_20713), .ZN(net_20712) );
INV_X4 inst_15245 ( .ZN(net_4641), .A(net_4256) );
INV_X4 inst_13711 ( .ZN(net_11813), .A(net_7857) );
AOI21_X4 inst_20177 ( .ZN(net_19745), .B1(net_18966), .A(net_14400), .B2(net_10082) );
NAND3_X2 inst_6610 ( .ZN(net_9284), .A2(net_7167), .A1(net_6107), .A3(net_3007) );
OAI211_X2 inst_2493 ( .ZN(net_13155), .B(net_13154), .A(net_12764), .C2(net_11278), .C1(net_9747) );
XNOR2_X2 inst_511 ( .ZN(net_6549), .B(net_6548), .A(net_1867) );
NAND2_X2 inst_9593 ( .ZN(net_10855), .A1(net_8836), .A2(net_7350) );
NAND2_X2 inst_8665 ( .A1(net_21163), .A2(net_16774), .ZN(net_16475) );
INV_X4 inst_14720 ( .ZN(net_10627), .A(net_2910) );
NOR3_X2 inst_2645 ( .ZN(net_15855), .A1(net_15614), .A3(net_15006), .A2(net_10543) );
OR2_X2 inst_1164 ( .A1(net_13343), .ZN(net_7158), .A2(net_7157) );
INV_X2 inst_18369 ( .ZN(net_17560), .A(net_17484) );
NOR2_X4 inst_3112 ( .ZN(net_4473), .A1(net_4027), .A2(net_1934) );
AND2_X2 inst_21365 ( .A1(net_2274), .ZN(net_2192), .A2(net_1645) );
INV_X4 inst_14025 ( .ZN(net_12483), .A(net_8122) );
NAND2_X2 inst_11410 ( .ZN(net_3427), .A1(net_3426), .A2(net_3211) );
INV_X4 inst_15994 ( .ZN(net_3224), .A(net_1210) );
NAND2_X4 inst_7276 ( .A1(net_19784), .ZN(net_8162), .A2(net_5658) );
INV_X4 inst_15340 ( .ZN(net_20291), .A(net_3164) );
INV_X4 inst_15501 ( .ZN(net_3298), .A(net_1654) );
INV_X4 inst_14613 ( .ZN(net_7979), .A(net_4422) );
INV_X2 inst_18742 ( .A(net_10524), .ZN(net_7907) );
NAND2_X2 inst_11416 ( .ZN(net_10042), .A1(net_7850), .A2(net_4331) );
INV_X4 inst_14596 ( .A(net_6862), .ZN(net_4451) );
OR2_X2 inst_1242 ( .A1(net_3867), .ZN(net_603), .A2(net_40) );
INV_X2 inst_19591 ( .ZN(net_19216), .A(net_295) );
INV_X4 inst_16558 ( .ZN(net_1167), .A(net_1166) );
INV_X4 inst_14915 ( .ZN(net_3571), .A(net_3570) );
INV_X4 inst_14578 ( .ZN(net_6217), .A(net_4528) );
INV_X2 inst_18849 ( .ZN(net_10634), .A(net_6615) );
INV_X4 inst_17838 ( .ZN(net_219), .A(net_101) );
INV_X4 inst_13363 ( .A(net_12816), .ZN(net_10935) );
NAND2_X2 inst_8362 ( .A1(net_21144), .A2(net_20714), .ZN(net_17397) );
AOI22_X2 inst_20013 ( .ZN(net_11777), .A1(net_11776), .A2(net_11775), .B2(net_9929), .B1(net_7903) );
XNOR2_X2 inst_388 ( .B(net_21123), .ZN(net_16773), .A(net_16769) );
AOI21_X2 inst_20796 ( .B2(net_12976), .A(net_12366), .ZN(net_10419), .B1(net_2911) );
INV_X8 inst_12374 ( .A(net_646), .ZN(net_264) );
INV_X4 inst_15119 ( .ZN(net_19213), .A(net_3181) );
XNOR2_X2 inst_489 ( .ZN(net_9257), .A(net_9256), .B(net_9255) );
NAND2_X2 inst_9278 ( .ZN(net_12590), .A2(net_10836), .A1(net_9981) );
NAND4_X2 inst_5502 ( .ZN(net_11821), .A2(net_11820), .A3(net_11819), .A1(net_11055), .A4(net_8299) );
NAND2_X4 inst_7153 ( .A1(net_13702), .ZN(net_10986), .A2(net_9575) );
NOR2_X2 inst_3622 ( .ZN(net_13584), .A1(net_12496), .A2(net_12310) );
AOI21_X2 inst_20888 ( .ZN(net_7799), .A(net_6788), .B2(net_4132), .B1(net_3464) );
INV_X4 inst_18041 ( .A(net_21088), .ZN(net_376) );
NAND2_X2 inst_11625 ( .ZN(net_4474), .A2(net_2726), .A1(net_90) );
XOR2_X2 inst_39 ( .A(net_21200), .Z(net_594), .B(net_593) );
NOR3_X4 inst_2627 ( .ZN(net_19580), .A3(net_19378), .A1(net_19377), .A2(net_13368) );
NAND2_X2 inst_8987 ( .ZN(net_14474), .A2(net_12914), .A1(net_1450) );
NOR2_X4 inst_3173 ( .ZN(net_3152), .A2(net_3109), .A1(net_252) );
XNOR2_X2 inst_125 ( .B(net_20794), .ZN(net_18382), .A(net_18315) );
CLKBUF_X2 inst_22923 ( .A(net_22794), .Z(net_22795) );
NOR2_X2 inst_4770 ( .ZN(net_5527), .A1(net_3101), .A2(net_2965) );
CLKBUF_X2 inst_22526 ( .A(net_22397), .Z(net_22398) );
AOI22_X2 inst_19982 ( .ZN(net_15373), .A1(net_15372), .A2(net_13886), .B2(net_9953), .B1(net_855) );
INV_X4 inst_15517 ( .ZN(net_11770), .A(net_5799) );
INV_X4 inst_17134 ( .ZN(net_15345), .A(net_652) );
NAND2_X4 inst_7696 ( .A1(net_880), .ZN(net_562), .A2(net_322) );
CLKBUF_X2 inst_22938 ( .A(net_22809), .Z(net_22810) );
INV_X4 inst_15233 ( .ZN(net_3586), .A(net_2268) );
NAND2_X2 inst_11919 ( .A1(net_20540), .A2(net_1751), .ZN(net_1541) );
INV_X4 inst_14753 ( .ZN(net_14226), .A(net_4070) );
INV_X4 inst_17557 ( .ZN(net_9367), .A(net_4805) );
XNOR2_X2 inst_430 ( .B(net_21171), .A(net_16482), .ZN(net_16481) );
CLKBUF_X2 inst_21554 ( .A(net_21425), .Z(net_21426) );
NAND2_X2 inst_11800 ( .A2(net_2606), .ZN(net_1920), .A1(net_1169) );
INV_X4 inst_16039 ( .ZN(net_10672), .A(net_5344) );
OAI211_X2 inst_2565 ( .ZN(net_9290), .C2(net_9289), .B(net_4644), .A(net_2680), .C1(net_1260) );
INV_X4 inst_17816 ( .A(net_824), .ZN(net_114) );
NAND2_X4 inst_7061 ( .A2(net_20872), .A1(net_19212), .ZN(net_16310) );
CLKBUF_X2 inst_22535 ( .A(net_21811), .Z(net_22407) );
INV_X2 inst_19679 ( .A(net_20514), .ZN(net_20513) );
NOR2_X4 inst_2945 ( .A2(net_8115), .ZN(net_6915), .A1(net_6914) );
INV_X2 inst_19283 ( .A(net_3656), .ZN(net_2922) );
XNOR2_X2 inst_642 ( .B(net_543), .ZN(net_407), .A(net_406) );
INV_X4 inst_13035 ( .A(net_16774), .ZN(net_16612) );
NOR2_X4 inst_2993 ( .A2(net_20491), .ZN(net_8061), .A1(net_5909) );
INV_X4 inst_14736 ( .ZN(net_4571), .A(net_4109) );
INV_X4 inst_13168 ( .ZN(net_14640), .A(net_14134) );
SDFF_X2 inst_1018 ( .QN(net_20998), .SE(net_2426), .D(net_1948), .CK(net_21836), .SI(x3058) );
INV_X4 inst_18104 ( .A(net_21217), .ZN(net_221) );
NAND2_X2 inst_10726 ( .ZN(net_5843), .A2(net_5835), .A1(net_887) );
NAND2_X2 inst_10655 ( .ZN(net_9849), .A1(net_6318), .A2(net_6317) );
INV_X4 inst_16416 ( .ZN(net_5289), .A(net_1515) );
INV_X4 inst_16227 ( .ZN(net_14636), .A(net_12326) );
INV_X4 inst_14160 ( .ZN(net_7323), .A(net_6018) );
SDFF_X2 inst_700 ( .Q(net_20958), .SE(net_18865), .SI(net_18842), .D(net_355), .CK(net_22271) );
INV_X4 inst_13507 ( .A(net_9414), .ZN(net_9413) );
INV_X8 inst_12295 ( .ZN(net_1092), .A(net_988) );
CLKBUF_X2 inst_22751 ( .A(net_22622), .Z(net_22623) );
INV_X4 inst_13323 ( .ZN(net_11413), .A(net_10083) );
NAND2_X2 inst_8107 ( .A2(net_20220), .ZN(net_18111), .A1(net_18081) );
NAND2_X2 inst_9152 ( .ZN(net_13395), .A1(net_12382), .A2(net_10584) );
NAND2_X2 inst_8555 ( .ZN(net_19865), .A2(net_16777), .A1(net_7341) );
INV_X4 inst_14457 ( .A(net_11090), .ZN(net_4947) );
SDFF_X2 inst_979 ( .QN(net_21024), .D(net_426), .SE(net_263), .CK(net_21896), .SI(x2618) );
CLKBUF_X2 inst_22113 ( .A(net_21984), .Z(net_21985) );
NOR2_X2 inst_4568 ( .A1(net_6177), .ZN(net_3880), .A2(net_3879) );
NAND3_X2 inst_5989 ( .ZN(net_19381), .A2(net_14535), .A1(net_13384), .A3(net_13335) );
NAND2_X2 inst_9785 ( .ZN(net_11106), .A2(net_7594), .A1(net_731) );
OAI21_X2 inst_2296 ( .B1(net_19439), .A(net_12406), .B2(net_6899), .ZN(net_6453) );
INV_X4 inst_13092 ( .ZN(net_20372), .A(net_15779) );
INV_X4 inst_12477 ( .ZN(net_18694), .A(net_18693) );
INV_X2 inst_18883 ( .ZN(net_6174), .A(net_6173) );
INV_X4 inst_17550 ( .A(net_10676), .ZN(net_5454) );
NAND2_X2 inst_12012 ( .ZN(net_1514), .A2(net_1289), .A1(net_236) );
NOR2_X2 inst_4964 ( .A2(net_2751), .ZN(net_2156), .A1(net_1755) );
NAND2_X2 inst_9587 ( .A1(net_12658), .ZN(net_10897), .A2(net_7347) );
INV_X4 inst_14133 ( .A(net_9885), .ZN(net_6106) );
AOI21_X2 inst_20513 ( .ZN(net_20680), .B1(net_14605), .B2(net_11719), .A(net_8214) );
INV_X4 inst_14912 ( .ZN(net_3575), .A(net_3574) );
INV_X4 inst_14919 ( .ZN(net_5806), .A(net_3563) );
INV_X4 inst_14802 ( .ZN(net_5029), .A(net_3982) );
NOR2_X2 inst_4258 ( .ZN(net_6268), .A2(net_6267), .A1(net_2144) );
NAND2_X2 inst_7889 ( .ZN(net_18509), .A2(net_18461), .A1(net_17702) );
NAND2_X2 inst_9607 ( .ZN(net_10729), .A1(net_10728), .A2(net_8804) );
NAND2_X2 inst_9764 ( .ZN(net_9830), .A2(net_9829), .A1(net_3450) );
NAND2_X2 inst_9018 ( .ZN(net_14189), .A1(net_14188), .A2(net_5427) );
CLKBUF_X2 inst_21653 ( .A(net_21524), .Z(net_21525) );
INV_X4 inst_17537 ( .ZN(net_19726), .A(net_955) );
NOR2_X2 inst_4040 ( .ZN(net_9441), .A1(net_7988), .A2(net_6055) );
AOI21_X2 inst_20517 ( .ZN(net_20370), .B1(net_19521), .A(net_7174), .B2(net_2408) );
OR3_X2 inst_1059 ( .A2(net_13018), .ZN(net_13006), .A3(net_13005), .A1(net_12890) );
CLKBUF_X2 inst_21729 ( .A(net_21298), .Z(net_21601) );
INV_X2 inst_18615 ( .A(net_11828), .ZN(net_9613) );
INV_X4 inst_13987 ( .ZN(net_7806), .A(net_5350) );
INV_X2 inst_19261 ( .A(net_15099), .ZN(net_3170) );
INV_X2 inst_19117 ( .ZN(net_4442), .A(net_4441) );
INV_X4 inst_16747 ( .ZN(net_7870), .A(net_154) );
INV_X4 inst_14227 ( .ZN(net_19157), .A(net_5834) );
NAND2_X2 inst_10215 ( .ZN(net_18892), .A1(net_8361), .A2(net_8086) );
INV_X4 inst_16237 ( .A(net_11407), .ZN(net_1850) );
NOR2_X2 inst_4328 ( .ZN(net_5803), .A1(net_3420), .A2(net_3393) );
CLKBUF_X2 inst_22694 ( .A(net_22565), .Z(net_22566) );
INV_X4 inst_15240 ( .A(net_3787), .ZN(net_2824) );
INV_X4 inst_15698 ( .ZN(net_2016), .A(net_1312) );
AOI21_X2 inst_20713 ( .B1(net_12551), .ZN(net_12044), .A(net_11388), .B2(net_7685) );
NOR2_X2 inst_4173 ( .A2(net_9956), .ZN(net_8158), .A1(net_6840) );
NAND3_X2 inst_6039 ( .ZN(net_14324), .A3(net_13211), .A2(net_11469), .A1(net_9531) );
INV_X4 inst_17934 ( .A(net_20934), .ZN(net_459) );
INV_X8 inst_12454 ( .A(net_20714), .ZN(net_20713) );
NAND3_X2 inst_6425 ( .A2(net_12406), .ZN(net_11931), .A3(net_8149), .A1(net_3684) );
OR2_X4 inst_1104 ( .ZN(net_10641), .A2(net_5248), .A1(net_952) );
INV_X4 inst_17486 ( .ZN(net_7428), .A(net_429) );
OAI21_X2 inst_2355 ( .ZN(net_2962), .A(net_2961), .B2(net_2960), .B1(net_2141) );
INV_X4 inst_17806 ( .ZN(net_20820), .A(net_123) );
INV_X4 inst_17756 ( .ZN(net_805), .A(net_161) );
NAND2_X2 inst_10886 ( .ZN(net_9037), .A2(net_5629), .A1(net_5448) );
NAND3_X2 inst_5753 ( .ZN(net_19682), .A1(net_15702), .A3(net_15390), .A2(net_11327) );
NAND2_X4 inst_7058 ( .A2(net_20928), .A1(net_19878), .ZN(net_16355) );
INV_X4 inst_15794 ( .A(net_4820), .ZN(net_1898) );
INV_X4 inst_12535 ( .ZN(net_18379), .A(net_18378) );
NAND2_X2 inst_9742 ( .ZN(net_10099), .A1(net_10098), .A2(net_9428) );
NAND2_X4 inst_7287 ( .ZN(net_8023), .A1(net_5537), .A2(net_4380) );
XNOR2_X2 inst_574 ( .B(net_9193), .A(net_675), .ZN(net_622) );
INV_X8 inst_12446 ( .ZN(net_20516), .A(net_20515) );
INV_X4 inst_17590 ( .ZN(net_15108), .A(net_934) );
NAND3_X4 inst_5552 ( .ZN(net_16530), .A1(net_16255), .A3(net_16158), .A2(net_15676) );
INV_X4 inst_14349 ( .A(net_15519), .ZN(net_13655) );
NAND2_X2 inst_8087 ( .ZN(net_20281), .A2(net_18140), .A1(net_16959) );
NOR2_X2 inst_4102 ( .A1(net_8502), .ZN(net_7215), .A2(net_7214) );
OR2_X2 inst_1229 ( .ZN(net_6830), .A1(net_2110), .A2(net_1825) );
NAND2_X2 inst_10512 ( .A1(net_11182), .A2(net_6917), .ZN(net_6882) );
INV_X4 inst_14725 ( .A(net_4189), .ZN(net_4135) );
INV_X2 inst_19031 ( .ZN(net_8047), .A(net_4883) );
AOI21_X2 inst_20359 ( .B1(net_19545), .ZN(net_19325), .B2(net_15664), .A(net_12258) );
NAND2_X4 inst_7545 ( .ZN(net_1829), .A2(net_1787), .A1(net_898) );
AND2_X2 inst_21313 ( .ZN(net_8379), .A1(net_8378), .A2(net_8377) );
INV_X4 inst_13780 ( .ZN(net_20184), .A(net_7576) );
INV_X4 inst_13604 ( .ZN(net_8574), .A(net_8573) );
NAND4_X4 inst_5219 ( .A4(net_19486), .A1(net_19485), .ZN(net_16369), .A3(net_14287), .A2(net_13830) );
CLKBUF_X2 inst_21994 ( .A(net_21334), .Z(net_21866) );
INV_X2 inst_19332 ( .ZN(net_3324), .A(net_2521) );
INV_X2 inst_18855 ( .ZN(net_6341), .A(net_6340) );
INV_X4 inst_15042 ( .ZN(net_6440), .A(net_3811) );
OAI21_X2 inst_2358 ( .A(net_2718), .ZN(net_2536), .B2(net_2535), .B1(net_2231) );
INV_X4 inst_13139 ( .ZN(net_20090), .A(net_14733) );
OAI21_X2 inst_2125 ( .ZN(net_10013), .A(net_10012), .B1(net_10011), .B2(net_10010) );
INV_X4 inst_15827 ( .ZN(net_8667), .A(net_5330) );
INV_X4 inst_17988 ( .A(net_20986), .ZN(net_2507) );
NAND2_X2 inst_11572 ( .ZN(net_8565), .A1(net_5984), .A2(net_2757) );
NAND2_X2 inst_10549 ( .ZN(net_15569), .A1(net_13026), .A2(net_5743) );
XNOR2_X2 inst_599 ( .B(net_16464), .ZN(net_545), .A(net_544) );
CLKBUF_X2 inst_22127 ( .A(net_21919), .Z(net_21999) );
INV_X4 inst_13382 ( .ZN(net_10784), .A(net_10783) );
XNOR2_X2 inst_541 ( .ZN(net_800), .A(net_799), .B(net_798) );
INV_X4 inst_16014 ( .ZN(net_2120), .A(net_1652) );
NOR2_X2 inst_4047 ( .ZN(net_9403), .A1(net_7816), .A2(net_6637) );
INV_X2 inst_18645 ( .ZN(net_9328), .A(net_9327) );
INV_X4 inst_13910 ( .ZN(net_8891), .A(net_5612) );
XNOR2_X2 inst_505 ( .ZN(net_8990), .B(net_5756), .A(net_2458) );
NAND3_X2 inst_6366 ( .A3(net_13054), .A2(net_12487), .ZN(net_12078), .A1(net_10414) );
OAI21_X4 inst_1365 ( .ZN(net_17841), .A(net_17597), .B2(net_17596), .B1(net_17062) );
NAND2_X4 inst_7247 ( .ZN(net_8931), .A2(net_5594), .A1(net_5021) );
INV_X4 inst_15722 ( .ZN(net_11858), .A(net_7975) );
NAND2_X2 inst_7936 ( .ZN(net_18432), .A2(net_18371), .A1(net_18317) );
XNOR2_X2 inst_198 ( .A(net_17675), .ZN(net_17671), .B(net_16266) );
INV_X4 inst_13624 ( .A(net_8829), .ZN(net_8332) );
NOR2_X2 inst_4125 ( .A1(net_14837), .ZN(net_7012), .A2(net_7011) );
OAI21_X4 inst_1371 ( .ZN(net_17231), .B1(net_16718), .A(net_16580), .B2(net_16579) );
NAND2_X2 inst_10809 ( .ZN(net_5529), .A2(net_5434), .A1(net_4726) );
NAND3_X4 inst_5622 ( .ZN(net_19610), .A1(net_10630), .A2(net_10629), .A3(net_7883) );
NOR2_X2 inst_4321 ( .A2(net_5908), .ZN(net_5867), .A1(net_5866) );
INV_X2 inst_19603 ( .A(net_337), .ZN(net_144) );
OAI21_X2 inst_1644 ( .ZN(net_19741), .A(net_16390), .B1(net_15177), .B2(net_15031) );
NAND3_X2 inst_6346 ( .ZN(net_18893), .A3(net_12240), .A1(net_8593), .A2(net_6123) );
INV_X2 inst_18531 ( .A(net_11499), .ZN(net_11081) );
INV_X4 inst_12645 ( .ZN(net_17882), .A(net_17881) );
CLKBUF_X2 inst_21718 ( .A(net_21589), .Z(net_21590) );
INV_X2 inst_18921 ( .ZN(net_5928), .A(net_5927) );
NAND2_X2 inst_8946 ( .A1(net_15345), .ZN(net_14728), .A2(net_13232) );
NAND2_X4 inst_7529 ( .A1(net_20201), .ZN(net_4232), .A2(net_1461) );
INV_X4 inst_13333 ( .A(net_11677), .ZN(net_11133) );
NAND2_X2 inst_9351 ( .ZN(net_18894), .A2(net_9901), .A1(net_7436) );
INV_X4 inst_16194 ( .A(net_7822), .ZN(net_2484) );
CLKBUF_X2 inst_22209 ( .A(net_21544), .Z(net_22081) );
CLKBUF_X2 inst_22338 ( .A(net_22209), .Z(net_22210) );
INV_X4 inst_15071 ( .ZN(net_14751), .A(net_11783) );
INV_X4 inst_17335 ( .A(net_3919), .ZN(net_1970) );
NOR2_X2 inst_3511 ( .ZN(net_13895), .A2(net_11987), .A1(net_4349) );
INV_X4 inst_18168 ( .A(net_20930), .ZN(net_152) );
NAND3_X2 inst_6726 ( .ZN(net_6503), .A1(net_5300), .A3(net_4951), .A2(net_4246) );
CLKBUF_X2 inst_22642 ( .A(net_22513), .Z(net_22514) );
NAND2_X2 inst_10363 ( .ZN(net_11300), .A1(net_7414), .A2(net_7401) );
NAND3_X2 inst_5693 ( .A3(net_19631), .A1(net_19630), .ZN(net_19466), .A2(net_14950) );
NAND2_X2 inst_9992 ( .A1(net_11771), .ZN(net_10328), .A2(net_8335) );
XNOR2_X2 inst_263 ( .ZN(net_17257), .A(net_16760), .B(net_622) );
CLKBUF_X2 inst_21826 ( .A(net_21697), .Z(net_21698) );
INV_X4 inst_18352 ( .A(net_20805), .ZN(net_20804) );
NAND2_X2 inst_10889 ( .ZN(net_7189), .A2(net_5409), .A1(net_3399) );
INV_X4 inst_15831 ( .ZN(net_3658), .A(net_1863) );
NAND2_X4 inst_7399 ( .ZN(net_4842), .A1(net_2800), .A2(net_2629) );
AND2_X4 inst_21215 ( .ZN(net_19664), .A1(net_7801), .A2(net_6347) );
NAND3_X2 inst_5953 ( .ZN(net_14875), .A2(net_14874), .A3(net_14873), .A1(net_8679) );
NAND3_X2 inst_6742 ( .A3(net_6971), .ZN(net_6403), .A2(net_6402), .A1(net_3709) );
AOI21_X2 inst_20455 ( .ZN(net_15052), .B1(net_13495), .B2(net_12959), .A(net_12631) );
NAND3_X2 inst_6307 ( .ZN(net_12781), .A2(net_11695), .A3(net_10210), .A1(net_8203) );
NAND2_X4 inst_7371 ( .ZN(net_5768), .A2(net_3187), .A1(net_3080) );
NAND2_X2 inst_10650 ( .A1(net_11549), .ZN(net_6352), .A2(net_6351) );
NAND2_X2 inst_10121 ( .ZN(net_9821), .A1(net_8376), .A2(net_8344) );
AOI21_X2 inst_20848 ( .A(net_9301), .ZN(net_9101), .B1(net_9100), .B2(net_9099) );
NAND2_X2 inst_11923 ( .ZN(net_1504), .A2(net_775), .A1(net_192) );
NOR2_X2 inst_4118 ( .A1(net_13091), .ZN(net_7047), .A2(net_7046) );
INV_X4 inst_13410 ( .ZN(net_10333), .A(net_10332) );
CLKBUF_X2 inst_21635 ( .A(net_21506), .Z(net_21507) );
NAND4_X2 inst_5440 ( .ZN(net_13913), .A3(net_12405), .A1(net_11033), .A4(net_10326), .A2(net_10065) );
NOR2_X2 inst_4849 ( .A1(net_8224), .ZN(net_2310), .A2(net_2309) );
INV_X4 inst_14689 ( .ZN(net_14222), .A(net_4291) );
CLKBUF_X2 inst_22953 ( .A(net_22824), .Z(net_22825) );
INV_X4 inst_17504 ( .A(net_9131), .ZN(net_5414) );
INV_X4 inst_16593 ( .ZN(net_2174), .A(net_1370) );
NAND2_X2 inst_8185 ( .ZN(net_17927), .A1(net_17926), .A2(net_17907) );
NAND2_X2 inst_11223 ( .ZN(net_7705), .A2(net_3410), .A1(net_809) );
INV_X4 inst_17647 ( .A(net_2274), .ZN(net_498) );
NAND2_X4 inst_7413 ( .A2(net_20559), .A1(net_19960), .ZN(net_4740) );
INV_X4 inst_15709 ( .A(net_2759), .ZN(net_1987) );
INV_X4 inst_14263 ( .ZN(net_7277), .A(net_5731) );
DFF_X1 inst_19833 ( .D(net_17434), .CK(net_22805), .Q(x1306) );
NAND2_X4 inst_7590 ( .ZN(net_2992), .A2(net_1752), .A1(net_1017) );
NAND2_X2 inst_8698 ( .A1(net_21236), .ZN(net_16324), .A2(net_16166) );
NOR2_X2 inst_5034 ( .ZN(net_10108), .A2(net_1133), .A1(net_888) );
NOR2_X2 inst_4853 ( .ZN(net_3055), .A2(net_2299), .A1(net_999) );
NAND3_X2 inst_6322 ( .ZN(net_12518), .A1(net_9275), .A3(net_7877), .A2(net_6158) );
INV_X2 inst_19587 ( .A(net_2121), .ZN(net_339) );
NOR2_X2 inst_3898 ( .ZN(net_9110), .A1(net_9109), .A2(net_5813) );
INV_X4 inst_17083 ( .A(net_1264), .ZN(net_1262) );
NAND4_X2 inst_5254 ( .A3(net_18910), .A1(net_18909), .ZN(net_16513), .A4(net_16234), .A2(net_14354) );
INV_X2 inst_18569 ( .ZN(net_10768), .A(net_10767) );
INV_X4 inst_18161 ( .A(net_21186), .ZN(net_16839) );
NAND2_X2 inst_9370 ( .A1(net_18025), .ZN(net_12085), .A2(net_9004) );
CLKBUF_X2 inst_22292 ( .A(net_21428), .Z(net_22164) );
NAND2_X2 inst_11949 ( .ZN(net_1421), .A2(net_1420), .A1(net_252) );
NOR2_X2 inst_3503 ( .A1(net_15995), .ZN(net_14032), .A2(net_11722) );
INV_X4 inst_13974 ( .ZN(net_8694), .A(net_6654) );
INV_X4 inst_15836 ( .ZN(net_3911), .A(net_1857) );
NAND2_X2 inst_7973 ( .ZN(net_18414), .A1(net_18255), .A2(net_18209) );
NOR2_X2 inst_4138 ( .ZN(net_6938), .A2(net_6878), .A1(net_4008) );
AOI21_X4 inst_20096 ( .B2(net_20936), .ZN(net_18600), .A(net_18590), .B1(net_15921) );
XOR2_X1 inst_52 ( .B(net_21158), .A(net_20523), .Z(net_18659) );
INV_X4 inst_12600 ( .A(net_18093), .ZN(net_18092) );
XNOR2_X2 inst_668 ( .A(net_21184), .B(net_21120), .ZN(net_188) );
INV_X4 inst_17799 ( .ZN(net_127), .A(net_126) );
NOR2_X4 inst_3049 ( .ZN(net_6171), .A1(net_5010), .A2(net_143) );
INV_X4 inst_15804 ( .ZN(net_12675), .A(net_7394) );
NAND2_X2 inst_11987 ( .A1(net_1730), .ZN(net_1263), .A2(net_863) );
INV_X4 inst_16015 ( .ZN(net_10395), .A(net_8326) );
INV_X4 inst_17571 ( .ZN(net_353), .A(net_352) );
NOR2_X2 inst_4159 ( .ZN(net_6887), .A1(net_6886), .A2(net_6885) );
AND2_X2 inst_21300 ( .ZN(net_15276), .A2(net_10218), .A1(net_10105) );
AOI21_X2 inst_20350 ( .ZN(net_15743), .B2(net_15097), .B1(net_14062), .A(net_2553) );
INV_X4 inst_12567 ( .ZN(net_18219), .A(net_18218) );
INV_X2 inst_19241 ( .ZN(net_3289), .A(net_1910) );
NOR2_X2 inst_3349 ( .ZN(net_17981), .A1(net_17947), .A2(net_17915) );
NAND2_X2 inst_11444 ( .ZN(net_3868), .A2(net_3246), .A1(net_225) );
CLKBUF_X2 inst_22555 ( .A(net_22135), .Z(net_22427) );
NAND2_X2 inst_10057 ( .A1(net_8798), .ZN(net_8687), .A2(net_8637) );
OAI211_X2 inst_2545 ( .ZN(net_10824), .B(net_9310), .A(net_7263), .C2(net_2880), .C1(net_1729) );
NAND2_X2 inst_8220 ( .ZN(net_17824), .A2(net_17652), .A1(net_17581) );
INV_X2 inst_18441 ( .ZN(net_19248), .A(net_12975) );
INV_X8 inst_12390 ( .A(net_234), .ZN(net_105) );
NAND2_X2 inst_10722 ( .ZN(net_19703), .A1(net_7676), .A2(net_3733) );
NAND2_X2 inst_7999 ( .ZN(net_18314), .A1(net_18313), .A2(net_18312) );
INV_X4 inst_13077 ( .ZN(net_16203), .A(net_16139) );
NOR3_X2 inst_2768 ( .ZN(net_9253), .A3(net_9252), .A2(net_4660), .A1(net_4399) );
CLKBUF_X2 inst_21373 ( .A(net_21244), .Z(net_21245) );
INV_X4 inst_14657 ( .ZN(net_4363), .A(net_4362) );
INV_X4 inst_17459 ( .A(net_6334), .ZN(net_2875) );
NAND2_X2 inst_9878 ( .ZN(net_9452), .A2(net_7418), .A1(net_1173) );
OAI21_X2 inst_1835 ( .ZN(net_14047), .A(net_14046), .B1(net_13081), .B2(net_8747) );
INV_X4 inst_16890 ( .ZN(net_7975), .A(net_4795) );
INV_X2 inst_19183 ( .ZN(net_3769), .A(net_3768) );
INV_X4 inst_15861 ( .ZN(net_9516), .A(net_8276) );
INV_X4 inst_13777 ( .ZN(net_7587), .A(net_7586) );
INV_X4 inst_15614 ( .ZN(net_7395), .A(net_2167) );
NOR2_X2 inst_4639 ( .ZN(net_4999), .A2(net_2006), .A1(net_143) );
INV_X8 inst_12399 ( .ZN(net_330), .A(net_203) );
NAND2_X2 inst_9670 ( .A1(net_11995), .ZN(net_10311), .A2(net_10310) );
NAND2_X2 inst_7797 ( .ZN(net_18705), .A1(net_18704), .A2(net_18679) );
INV_X4 inst_15410 ( .ZN(net_3371), .A(net_2529) );
INV_X4 inst_15176 ( .A(net_10993), .ZN(net_6360) );
XNOR2_X2 inst_621 ( .B(net_604), .ZN(net_474), .A(net_473) );
NAND2_X2 inst_7764 ( .ZN(net_18749), .A2(net_18720), .A1(net_18697) );
INV_X2 inst_18386 ( .A(net_16727), .ZN(net_16654) );
OAI211_X2 inst_2560 ( .ZN(net_9916), .B(net_9915), .C1(net_9914), .C2(net_9913), .A(net_6509) );
INV_X4 inst_17188 ( .ZN(net_4815), .A(net_718) );
INV_X1 inst_19765 ( .A(net_20874), .ZN(net_34) );
AOI21_X2 inst_20766 ( .ZN(net_10751), .B2(net_6713), .B1(net_1597), .A(net_178) );
INV_X4 inst_15224 ( .A(net_4041), .ZN(net_3600) );
INV_X8 inst_12236 ( .A(net_5136), .ZN(net_4578) );
INV_X2 inst_19670 ( .A(net_20485), .ZN(net_20484) );
NAND2_X2 inst_9651 ( .ZN(net_10356), .A1(net_10355), .A2(net_10354) );
INV_X4 inst_14435 ( .ZN(net_13481), .A(net_5039) );
OAI21_X4 inst_1387 ( .A(net_20944), .B2(net_19701), .B1(net_19700), .ZN(net_19238) );
INV_X4 inst_15138 ( .ZN(net_4053), .A(net_3304) );
INV_X4 inst_13687 ( .ZN(net_11397), .A(net_7965) );
OAI21_X1 inst_2365 ( .A(net_9324), .ZN(net_7148), .B1(net_7147), .B2(net_7146) );
INV_X2 inst_18367 ( .ZN(net_17864), .A(net_17863) );
INV_X4 inst_16851 ( .ZN(net_15649), .A(net_15300) );
NAND2_X2 inst_12094 ( .A2(net_896), .ZN(net_608), .A1(net_328) );
OAI21_X2 inst_2250 ( .A(net_8798), .ZN(net_7300), .B2(net_5526), .B1(net_3392) );
CLKBUF_X2 inst_22724 ( .A(net_22595), .Z(net_22596) );
INV_X4 inst_15190 ( .ZN(net_5211), .A(net_2259) );
NAND3_X2 inst_6629 ( .ZN(net_9022), .A1(net_9021), .A3(net_9020), .A2(net_5954) );
OAI21_X2 inst_2187 ( .ZN(net_8790), .A(net_5244), .B2(net_4965), .B1(net_4413) );
CLKBUF_X2 inst_21791 ( .A(net_21662), .Z(net_21663) );
INV_X4 inst_13221 ( .ZN(net_13626), .A(net_12775) );
NAND2_X2 inst_11215 ( .A1(net_5402), .ZN(net_5064), .A2(net_3121) );
NAND3_X2 inst_5747 ( .ZN(net_16013), .A1(net_15754), .A3(net_15151), .A2(net_11640) );
INV_X4 inst_14323 ( .ZN(net_5453), .A(net_5452) );
NAND2_X4 inst_7448 ( .ZN(net_4961), .A2(net_1794), .A1(net_1491) );
XOR2_X2 inst_25 ( .B(net_21170), .A(net_16530), .Z(net_16527) );
AOI21_X4 inst_20243 ( .B1(net_19276), .ZN(net_10600), .A(net_9525), .B2(net_5918) );
NAND2_X2 inst_9043 ( .ZN(net_14049), .A2(net_12021), .A1(net_10917) );
NAND4_X4 inst_5239 ( .ZN(net_15508), .A1(net_14686), .A4(net_14479), .A3(net_13020), .A2(net_12894) );
NOR2_X2 inst_5032 ( .ZN(net_5285), .A2(net_2872), .A1(net_1376) );
AOI21_X2 inst_20808 ( .ZN(net_10253), .A(net_10252), .B1(net_10251), .B2(net_4524) );
NAND4_X4 inst_5166 ( .A2(net_19884), .A1(net_19883), .A4(net_18955), .ZN(net_18083), .A3(net_15240) );
INV_X4 inst_16210 ( .ZN(net_7580), .A(net_1409) );
NAND2_X2 inst_9691 ( .ZN(net_10239), .A1(net_10238), .A2(net_10237) );
AOI21_X4 inst_20151 ( .ZN(net_15816), .B1(net_15697), .B2(net_14886), .A(net_14001) );
OAI211_X2 inst_2500 ( .C1(net_13569), .ZN(net_12855), .B(net_12854), .A(net_12414), .C2(net_6469) );
NAND2_X2 inst_12119 ( .A1(net_21230), .A2(net_1790), .ZN(net_429) );
NAND2_X2 inst_9734 ( .ZN(net_13846), .A2(net_11813), .A1(net_8983) );
NOR2_X2 inst_4395 ( .ZN(net_20760), .A1(net_12546), .A2(net_5194) );
NOR2_X2 inst_3434 ( .ZN(net_20248), .A2(net_14236), .A1(net_8034) );
NOR2_X2 inst_4296 ( .ZN(net_5971), .A2(net_5970), .A1(net_3098) );
CLKBUF_X2 inst_22518 ( .A(net_22389), .Z(net_22390) );
INV_X2 inst_19248 ( .ZN(net_4758), .A(net_3263) );
CLKBUF_X2 inst_21926 ( .A(net_21731), .Z(net_21798) );
AOI21_X2 inst_20800 ( .B2(net_10728), .ZN(net_10388), .B1(net_2863), .A(net_112) );
NOR2_X4 inst_3204 ( .ZN(net_3037), .A2(net_3036), .A1(net_1356) );
INV_X4 inst_14219 ( .ZN(net_11348), .A(net_7511) );
NOR2_X2 inst_3421 ( .ZN(net_20092), .A2(net_14762), .A1(net_13588) );
NOR2_X2 inst_4444 ( .ZN(net_4800), .A1(net_4799), .A2(net_4798) );
NAND2_X2 inst_12019 ( .ZN(net_1367), .A2(net_1056), .A1(net_140) );
NOR3_X2 inst_2679 ( .ZN(net_14585), .A3(net_12138), .A1(net_8461), .A2(net_5453) );
NAND2_X4 inst_6935 ( .ZN(net_19312), .A1(net_17557), .A2(net_17359) );
NOR2_X2 inst_3949 ( .ZN(net_8614), .A2(net_7966), .A1(net_3741) );
AND2_X2 inst_21349 ( .ZN(net_2496), .A2(net_2495), .A1(net_2060) );
INV_X4 inst_15731 ( .A(net_12366), .ZN(net_7396) );
INV_X4 inst_16727 ( .ZN(net_5884), .A(net_891) );
NOR2_X2 inst_4617 ( .ZN(net_4498), .A1(net_3646), .A2(net_1383) );
OAI21_X2 inst_1777 ( .ZN(net_14673), .A(net_12393), .B2(net_11935), .B1(net_10241) );
INV_X2 inst_18919 ( .ZN(net_5947), .A(net_5946) );
INV_X4 inst_14971 ( .ZN(net_13926), .A(net_4350) );
OR2_X4 inst_1068 ( .ZN(net_13120), .A2(net_13119), .A1(net_10129) );
SDFF_X2 inst_886 ( .Q(net_21208), .D(net_16934), .SE(net_263), .CK(net_21651), .SI(x5873) );
INV_X4 inst_12799 ( .ZN(net_17261), .A(net_17260) );
NAND2_X2 inst_11799 ( .ZN(net_6474), .A2(net_5884), .A1(net_1921) );
INV_X4 inst_16608 ( .ZN(net_2260), .A(net_1217) );
INV_X4 inst_12509 ( .ZN(net_18632), .A(net_18620) );
INV_X4 inst_15409 ( .ZN(net_15542), .A(net_15071) );
NAND4_X2 inst_5350 ( .ZN(net_20638), .A1(net_14666), .A3(net_14538), .A4(net_12171), .A2(net_10120) );
CLKBUF_X2 inst_21488 ( .A(net_21359), .Z(net_21360) );
INV_X2 inst_18620 ( .A(net_13458), .ZN(net_9585) );
INV_X4 inst_15251 ( .ZN(net_4914), .A(net_3937) );
INV_X4 inst_13319 ( .ZN(net_11567), .A(net_11566) );
NOR2_X2 inst_4468 ( .A1(net_21238), .ZN(net_12770), .A2(net_4474) );
NAND2_X2 inst_11740 ( .ZN(net_3992), .A2(net_2174), .A1(net_61) );
NAND2_X2 inst_11533 ( .A2(net_2952), .ZN(net_2930), .A1(net_1595) );
INV_X4 inst_14450 ( .ZN(net_6578), .A(net_4966) );
NAND2_X2 inst_11484 ( .ZN(net_19419), .A2(net_3089), .A1(net_107) );
INV_X4 inst_17520 ( .ZN(net_3047), .A(net_252) );
NAND2_X2 inst_11270 ( .ZN(net_3891), .A1(net_3890), .A2(net_2736) );
INV_X4 inst_15874 ( .ZN(net_1794), .A(net_1793) );
INV_X8 inst_12380 ( .ZN(net_328), .A(net_117) );
AOI21_X2 inst_20948 ( .ZN(net_5857), .B2(net_5649), .A(net_3665), .B1(net_1936) );
NAND2_X2 inst_8844 ( .ZN(net_15437), .A2(net_15025), .A1(net_13138) );
OAI21_X2 inst_1969 ( .B1(net_19731), .ZN(net_12255), .A(net_12254), .B2(net_4799) );
NAND2_X2 inst_7837 ( .A2(net_20521), .ZN(net_18630), .A1(net_16823) );
NAND2_X2 inst_11382 ( .ZN(net_5891), .A1(net_2224), .A2(net_2117) );
NAND2_X2 inst_9128 ( .ZN(net_20613), .A1(net_13530), .A2(net_10791) );
CLKBUF_X2 inst_21950 ( .A(net_21821), .Z(net_21822) );
INV_X4 inst_15631 ( .ZN(net_3312), .A(net_3025) );
CLKBUF_X2 inst_22299 ( .A(net_21694), .Z(net_22171) );
NAND2_X2 inst_9348 ( .ZN(net_12191), .A2(net_10038), .A1(net_9805) );
NAND2_X2 inst_8183 ( .ZN(net_17929), .A1(net_17900), .A2(net_17804) );
NAND2_X4 inst_6914 ( .A2(net_20596), .A1(net_20595), .ZN(net_17855) );
AOI21_X2 inst_20542 ( .ZN(net_14417), .A(net_14416), .B2(net_12565), .B1(net_3282) );
INV_X4 inst_15004 ( .ZN(net_14820), .A(net_12542) );
CLKBUF_X2 inst_22713 ( .A(net_22144), .Z(net_22585) );
INV_X2 inst_18993 ( .ZN(net_12508), .A(net_6841) );
NAND3_X2 inst_6540 ( .ZN(net_10574), .A2(net_10573), .A3(net_8736), .A1(net_4797) );
INV_X4 inst_14536 ( .ZN(net_4657), .A(net_3343) );
INV_X2 inst_18928 ( .ZN(net_5903), .A(net_5902) );
INV_X4 inst_13136 ( .ZN(net_15132), .A(net_14748) );
AOI21_X2 inst_20292 ( .B2(net_19394), .B1(net_19393), .A(net_16259), .ZN(net_16177) );
INV_X2 inst_19268 ( .A(net_3954), .ZN(net_3064) );
AND3_X4 inst_21126 ( .A2(net_13174), .ZN(net_12018), .A3(net_10465), .A1(net_4015) );
NOR2_X4 inst_3150 ( .ZN(net_20575), .A1(net_3355), .A2(net_3350) );
NAND2_X2 inst_10761 ( .ZN(net_6973), .A2(net_5649), .A1(net_1987) );
INV_X2 inst_18793 ( .ZN(net_7445), .A(net_7444) );
INV_X4 inst_15976 ( .ZN(net_14622), .A(net_8682) );
INV_X4 inst_12765 ( .ZN(net_17361), .A(net_17360) );
NAND2_X2 inst_8522 ( .ZN(net_16906), .A1(net_16664), .A2(net_16556) );
INV_X4 inst_14741 ( .ZN(net_6976), .A(net_2404) );
NAND3_X2 inst_6216 ( .ZN(net_20598), .A2(net_13002), .A1(net_9358), .A3(net_8740) );
NAND3_X2 inst_5791 ( .ZN(net_19935), .A1(net_15123), .A3(net_15001), .A2(net_5742) );
SDFF_X2 inst_866 ( .Q(net_21126), .D(net_17073), .SE(net_263), .CK(net_21465), .SI(x4172) );
NAND2_X2 inst_11061 ( .A2(net_4619), .ZN(net_4602), .A1(net_2887) );
OAI21_X4 inst_1439 ( .B2(net_20271), .B1(net_20270), .A(net_16357), .ZN(net_15885) );
AOI21_X2 inst_20466 ( .ZN(net_15000), .B1(net_13734), .B2(net_12993), .A(net_8904) );
NAND2_X4 inst_7214 ( .ZN(net_9409), .A2(net_7870), .A1(net_6015) );
NOR2_X2 inst_3640 ( .A1(net_20374), .ZN(net_12102), .A2(net_11538) );
INV_X8 inst_12367 ( .ZN(net_2001), .A(net_160) );
NAND2_X2 inst_8444 ( .ZN(net_19244), .A2(net_17126), .A1(net_16932) );
INV_X4 inst_17950 ( .A(net_21016), .ZN(net_392) );
INV_X4 inst_17200 ( .ZN(net_3402), .A(net_61) );
NAND3_X4 inst_5604 ( .A3(net_20056), .ZN(net_14406), .A2(net_14405), .A1(net_14333) );
XNOR2_X2 inst_248 ( .ZN(net_17315), .A(net_17308), .B(net_16093) );
NOR2_X4 inst_3107 ( .ZN(net_5160), .A2(net_4079), .A1(net_3179) );
AOI21_X2 inst_20743 ( .B2(net_11708), .ZN(net_11405), .A(net_11404), .B1(net_5798) );
OAI21_X2 inst_1919 ( .ZN(net_13028), .B2(net_11518), .A(net_7295), .B1(net_6345) );
INV_X4 inst_15747 ( .ZN(net_3255), .A(net_1559) );
INV_X2 inst_18442 ( .ZN(net_13689), .A(net_12924) );
INV_X8 inst_12222 ( .ZN(net_8867), .A(net_5175) );
AOI21_X2 inst_20871 ( .B2(net_12025), .ZN(net_8566), .B1(net_8565), .A(net_499) );
INV_X4 inst_18238 ( .A(net_20984), .ZN(net_382) );
NAND2_X2 inst_10528 ( .ZN(net_6833), .A1(net_6832), .A2(net_4944) );
CLKBUF_X2 inst_21761 ( .A(net_21632), .Z(net_21633) );
AOI21_X2 inst_20753 ( .ZN(net_11298), .B1(net_10183), .B2(net_9572), .A(net_6564) );
INV_X4 inst_15938 ( .ZN(net_3784), .A(net_1878) );
INV_X2 inst_18508 ( .ZN(net_11637), .A(net_10312) );
OAI21_X2 inst_1960 ( .ZN(net_12521), .B2(net_12520), .A(net_12495), .B1(net_7210) );
INV_X4 inst_15675 ( .A(net_11536), .ZN(net_10989) );
AND3_X2 inst_21135 ( .ZN(net_13224), .A1(net_13206), .A3(net_13205), .A2(net_13030) );
AOI22_X2 inst_20031 ( .ZN(net_9268), .B2(net_9267), .A1(net_6798), .B1(net_4312), .A2(net_3751) );
NAND2_X2 inst_8712 ( .A1(net_20944), .ZN(net_16236), .A2(net_16057) );
INV_X4 inst_13273 ( .ZN(net_12494), .A(net_11261) );
NAND2_X2 inst_11886 ( .ZN(net_6455), .A1(net_1604), .A2(net_187) );
NAND2_X2 inst_10283 ( .ZN(net_11834), .A2(net_7948), .A1(net_573) );
NAND2_X2 inst_10659 ( .A2(net_6336), .ZN(net_6306), .A1(net_4949) );
NAND2_X2 inst_10744 ( .A2(net_8696), .A1(net_5719), .ZN(net_5718) );
NOR2_X2 inst_4636 ( .ZN(net_6351), .A2(net_3492), .A1(net_154) );
XNOR2_X2 inst_302 ( .B(net_21125), .ZN(net_17108), .A(net_17107) );
XNOR2_X2 inst_673 ( .B(net_21167), .A(net_21135), .ZN(net_14915) );
CLKBUF_X2 inst_22241 ( .A(net_22112), .Z(net_22113) );
NOR2_X2 inst_3585 ( .ZN(net_12637), .A2(net_12636), .A1(net_6990) );
OR2_X2 inst_1151 ( .ZN(net_9767), .A2(net_9766), .A1(net_7230) );
INV_X4 inst_14952 ( .ZN(net_4538), .A(net_3506) );
NAND2_X2 inst_11399 ( .A2(net_10756), .ZN(net_3468), .A1(net_3467) );
AND2_X4 inst_21238 ( .ZN(net_8796), .A1(net_4212), .A2(net_4084) );
XNOR2_X2 inst_561 ( .A(net_21128), .B(net_11872), .ZN(net_680) );
INV_X4 inst_13417 ( .ZN(net_10273), .A(net_10272) );
INV_X4 inst_12999 ( .ZN(net_20186), .A(net_16420) );
NAND2_X2 inst_10903 ( .ZN(net_9075), .A1(net_7858), .A2(net_5071) );
OAI211_X2 inst_2505 ( .ZN(net_12766), .C2(net_12095), .B(net_10472), .C1(net_8952), .A(net_6813) );
NAND3_X2 inst_6504 ( .A3(net_20776), .ZN(net_10808), .A2(net_6122), .A1(net_3564) );
INV_X8 inst_12253 ( .ZN(net_9529), .A(net_2330) );
AOI21_X2 inst_20875 ( .ZN(net_20423), .B1(net_13080), .B2(net_6996), .A(net_4040) );
OAI21_X2 inst_1641 ( .A(net_16390), .ZN(net_15949), .B1(net_15250), .B2(net_14823) );
NAND3_X2 inst_6765 ( .A2(net_15833), .A3(net_13416), .A1(net_5618), .ZN(net_5324) );
INV_X2 inst_19167 ( .ZN(net_3860), .A(net_3859) );
INV_X4 inst_12524 ( .ZN(net_18468), .A(net_18467) );
INV_X4 inst_14620 ( .ZN(net_5826), .A(net_4408) );
NAND2_X2 inst_11749 ( .ZN(net_3245), .A1(net_2264), .A2(net_1350) );
XNOR2_X2 inst_196 ( .ZN(net_17674), .A(net_17673), .B(net_7650) );
OAI21_X2 inst_1567 ( .A(net_16743), .ZN(net_16433), .B2(net_16323), .B1(net_14065) );
INV_X2 inst_18661 ( .A(net_10903), .ZN(net_9197) );
INV_X4 inst_17542 ( .ZN(net_917), .A(net_380) );
INV_X4 inst_15161 ( .ZN(net_5481), .A(net_3028) );
NOR2_X2 inst_3451 ( .ZN(net_14887), .A1(net_13736), .A2(net_12980) );
OAI211_X2 inst_2417 ( .ZN(net_15420), .C1(net_15108), .A(net_14900), .C2(net_13642), .B(net_7199) );
INV_X4 inst_13481 ( .ZN(net_9584), .A(net_9583) );
INV_X4 inst_12828 ( .ZN(net_17537), .A(net_17143) );
AOI211_X2 inst_21008 ( .A(net_20364), .B(net_20363), .ZN(net_19481), .C1(net_15666), .C2(net_14776) );
INV_X2 inst_19556 ( .A(net_860), .ZN(net_859) );
NAND2_X2 inst_8405 ( .A1(net_17404), .ZN(net_17246), .A2(net_17245) );
INV_X4 inst_17960 ( .A(net_20954), .ZN(net_112) );
NAND3_X4 inst_5606 ( .ZN(net_19807), .A2(net_14361), .A3(net_13803), .A1(net_11453) );
INV_X4 inst_14371 ( .ZN(net_5183), .A(net_5182) );
XNOR2_X2 inst_298 ( .B(net_21115), .ZN(net_17118), .A(net_16624) );
OAI21_X2 inst_2180 ( .A(net_11776), .ZN(net_8853), .B2(net_8083), .B1(net_3394) );
OAI21_X2 inst_1856 ( .ZN(net_13987), .B1(net_13019), .A(net_10920), .B2(net_10112) );
NAND2_X2 inst_9379 ( .ZN(net_19329), .A1(net_14465), .A2(net_8617) );
NAND4_X2 inst_5507 ( .ZN(net_11246), .A2(net_11245), .A1(net_11244), .A4(net_11243), .A3(net_4789) );
INV_X4 inst_15993 ( .ZN(net_9330), .A(net_8020) );
NAND3_X2 inst_6594 ( .ZN(net_9924), .A2(net_9923), .A3(net_4723), .A1(net_2796) );
NAND2_X2 inst_11390 ( .ZN(net_3519), .A2(net_3328), .A1(net_924) );
NAND2_X2 inst_11124 ( .ZN(net_5471), .A2(net_4322), .A1(net_4286) );
NAND3_X2 inst_6180 ( .ZN(net_13500), .A1(net_11046), .A2(net_9181), .A3(net_7508) );
AOI21_X2 inst_20966 ( .ZN(net_5279), .A(net_5278), .B2(net_3632), .B1(net_3214) );
NOR2_X2 inst_3529 ( .ZN(net_13575), .A2(net_13574), .A1(net_2508) );
INV_X4 inst_14548 ( .ZN(net_4609), .A(net_4608) );
OAI21_X2 inst_2040 ( .ZN(net_13864), .A(net_11297), .B1(net_7424), .B2(net_7168) );
NAND2_X2 inst_10834 ( .ZN(net_10376), .A1(net_10037), .A2(net_3116) );
INV_X4 inst_17956 ( .A(net_21175), .ZN(net_17036) );
NAND2_X4 inst_7327 ( .A1(net_19375), .ZN(net_6224), .A2(net_1160) );
NOR2_X2 inst_4742 ( .A1(net_5454), .A2(net_4216), .ZN(net_3043) );
INV_X2 inst_18820 ( .A(net_9066), .ZN(net_6969) );
NAND3_X2 inst_6527 ( .A1(net_11640), .ZN(net_10611), .A2(net_10610), .A3(net_10609) );
NAND3_X2 inst_6099 ( .ZN(net_13912), .A3(net_13152), .A2(net_10948), .A1(net_7176) );
INV_X4 inst_12687 ( .ZN(net_17702), .A(net_17701) );
NOR2_X2 inst_4561 ( .ZN(net_12794), .A1(net_3908), .A2(net_3907) );
NAND2_X2 inst_11315 ( .ZN(net_4745), .A2(net_3730), .A1(net_1124) );
NAND2_X2 inst_9324 ( .ZN(net_12323), .A1(net_11691), .A2(net_9060) );
CLKBUF_X2 inst_22377 ( .A(net_22248), .Z(net_22249) );
NAND2_X2 inst_9611 ( .ZN(net_19830), .A2(net_8451), .A1(net_761) );
NAND3_X2 inst_6221 ( .ZN(net_13241), .A3(net_13126), .A2(net_6661), .A1(net_3271) );
NOR3_X2 inst_2743 ( .ZN(net_12751), .A1(net_10180), .A3(net_8109), .A2(net_6008) );
INV_X4 inst_17978 ( .A(net_20917), .ZN(net_972) );
AOI211_X4 inst_20988 ( .C1(net_20388), .ZN(net_16136), .B(net_15756), .A(net_14444), .C2(net_10182) );
OAI21_X2 inst_2083 ( .B1(net_11550), .ZN(net_10489), .B2(net_10488), .A(net_8365) );
AOI21_X4 inst_20237 ( .ZN(net_11205), .B1(net_11204), .A(net_7496), .B2(net_6437) );
AOI21_X4 inst_20124 ( .B2(net_19875), .B1(net_19874), .ZN(net_19837), .A(net_14522) );
INV_X4 inst_15144 ( .ZN(net_5547), .A(net_2356) );
OAI21_X4 inst_1470 ( .B2(net_19752), .B1(net_19751), .ZN(net_19273), .A(net_14755) );
INV_X4 inst_17493 ( .A(net_2214), .ZN(net_1215) );
NAND2_X2 inst_8019 ( .ZN(net_18279), .A2(net_18278), .A1(net_18208) );
INV_X4 inst_16198 ( .ZN(net_14986), .A(net_14709) );
INV_X4 inst_16294 ( .A(net_10096), .ZN(net_9914) );
OR2_X2 inst_1213 ( .A1(net_6334), .ZN(net_3008), .A2(net_3007) );
NOR2_X4 inst_3072 ( .ZN(net_5920), .A2(net_5595), .A1(net_4959) );
NAND2_X4 inst_7524 ( .ZN(net_3937), .A1(net_1861), .A2(net_1836) );
NAND2_X2 inst_12128 ( .ZN(net_1065), .A2(net_125), .A1(x7654) );
INV_X4 inst_14094 ( .ZN(net_9392), .A(net_5058) );
OAI211_X2 inst_2452 ( .ZN(net_14527), .C1(net_14186), .B(net_13962), .C2(net_10578), .A(net_4359) );
NAND2_X2 inst_11370 ( .ZN(net_3577), .A2(net_2846), .A1(net_2385) );
CLKBUF_X2 inst_22520 ( .A(net_22391), .Z(net_22392) );
INV_X4 inst_17243 ( .A(net_15301), .ZN(net_9656) );
XNOR2_X2 inst_428 ( .ZN(net_16483), .A(net_16482), .B(net_13296) );
NAND2_X2 inst_11821 ( .ZN(net_10046), .A2(net_7253), .A1(net_1815) );
INV_X4 inst_17842 ( .A(net_896), .ZN(net_284) );
NAND2_X2 inst_9093 ( .ZN(net_20312), .A1(net_13787), .A2(net_11521) );
INV_X4 inst_17043 ( .A(net_15959), .ZN(net_833) );
XNOR2_X2 inst_97 ( .ZN(net_18543), .A(net_18434), .B(net_16782) );
INV_X4 inst_15658 ( .ZN(net_4273), .A(net_1779) );
SDFF_X2 inst_775 ( .Q(net_20966), .SE(net_18859), .SI(net_18450), .D(net_642), .CK(net_22170) );
NAND2_X2 inst_8120 ( .ZN(net_18074), .A2(net_18064), .A1(net_7387) );
NOR2_X2 inst_4652 ( .ZN(net_3330), .A2(net_3287), .A1(net_1758) );
INV_X4 inst_16058 ( .ZN(net_2529), .A(net_1150) );
INV_X2 inst_18815 ( .ZN(net_7263), .A(net_7262) );
INV_X2 inst_18446 ( .A(net_14298), .ZN(net_13602) );
NAND2_X2 inst_11102 ( .ZN(net_7346), .A1(net_6201), .A2(net_4400) );
NAND2_X2 inst_11812 ( .ZN(net_5252), .A2(net_1837), .A1(net_1376) );
INV_X4 inst_14281 ( .ZN(net_6074), .A(net_3913) );
INV_X2 inst_19487 ( .A(net_3484), .ZN(net_1318) );
CLKBUF_X2 inst_22261 ( .A(net_22132), .Z(net_22133) );
AND4_X2 inst_21094 ( .ZN(net_15143), .A2(net_13276), .A3(net_10547), .A1(net_9426), .A4(net_8823) );
AOI211_X2 inst_21061 ( .C1(net_14186), .ZN(net_9950), .B(net_9949), .A(net_9485), .C2(net_2181) );
INV_X4 inst_17020 ( .ZN(net_1636), .A(net_472) );
INV_X4 inst_15124 ( .ZN(net_5573), .A(net_4206) );
OAI21_X2 inst_2242 ( .ZN(net_7381), .A(net_7380), .B1(net_3584), .B2(net_1437) );
INV_X4 inst_12954 ( .A(net_16748), .ZN(net_16540) );
OAI21_X2 inst_1671 ( .B2(net_19815), .B1(net_19814), .ZN(net_15617), .A(net_15616) );
NOR2_X2 inst_4581 ( .ZN(net_11212), .A2(net_7094), .A1(net_3836) );
NAND2_X2 inst_10044 ( .ZN(net_12194), .A2(net_12147), .A1(net_10098) );
INV_X4 inst_13203 ( .ZN(net_13858), .A(net_13175) );
NOR2_X4 inst_2884 ( .ZN(net_11664), .A1(net_8739), .A2(net_6145) );
XNOR2_X2 inst_600 ( .B(net_21155), .ZN(net_13284), .A(net_543) );
INV_X4 inst_13662 ( .ZN(net_11828), .A(net_8111) );
INV_X4 inst_15906 ( .ZN(net_2421), .A(net_1763) );
NAND4_X2 inst_5319 ( .A2(net_19643), .A1(net_19642), .ZN(net_15769), .A4(net_15002), .A3(net_8844) );
NOR2_X2 inst_4498 ( .A2(net_9289), .ZN(net_4643), .A1(net_3492) );
OR2_X2 inst_1194 ( .A1(net_11770), .ZN(net_7046), .A2(net_3169) );
AND2_X4 inst_21233 ( .A1(net_7912), .ZN(net_4168), .A2(net_4167) );
INV_X4 inst_14292 ( .ZN(net_13718), .A(net_10042) );
XOR2_X2 inst_49 ( .A(net_21184), .Z(net_423), .B(net_422) );
INV_X4 inst_14353 ( .ZN(net_9252), .A(net_5275) );
INV_X4 inst_17196 ( .ZN(net_962), .A(net_123) );
INV_X4 inst_14288 ( .ZN(net_7320), .A(net_5606) );
INV_X4 inst_15306 ( .A(net_11204), .ZN(net_9989) );
NOR2_X2 inst_4097 ( .ZN(net_7231), .A1(net_7230), .A2(net_7229) );
SDFF_X2 inst_693 ( .Q(net_20893), .SE(net_18865), .SI(net_18860), .D(net_484), .CK(net_21314) );
INV_X2 inst_18439 ( .ZN(net_14012), .A(net_13361) );
CLKBUF_X2 inst_21432 ( .A(net_21303), .Z(net_21304) );
INV_X4 inst_17246 ( .ZN(net_1445), .A(net_809) );
NAND2_X2 inst_10119 ( .A2(net_8933), .ZN(net_8382), .A1(net_4507) );
NAND2_X2 inst_8920 ( .ZN(net_14956), .A2(net_13740), .A1(net_10164) );
NAND3_X2 inst_6217 ( .A2(net_20772), .ZN(net_13257), .A1(net_9355), .A3(net_8742) );
NAND2_X4 inst_7383 ( .A2(net_20481), .ZN(net_5175), .A1(net_3256) );
NAND2_X4 inst_7390 ( .ZN(net_11702), .A1(net_9943), .A2(net_4188) );
INV_X4 inst_17402 ( .ZN(net_8341), .A(net_2274) );
NAND2_X2 inst_8303 ( .ZN(net_17597), .A2(net_17596), .A1(net_17061) );
INV_X2 inst_18605 ( .ZN(net_9783), .A(net_9782) );
INV_X4 inst_14987 ( .A(net_6363), .ZN(net_3404) );
SDFF_X2 inst_908 ( .Q(net_21204), .D(net_16803), .SE(net_263), .CK(net_22417), .SI(x5992) );
NAND2_X2 inst_11690 ( .A2(net_2331), .ZN(net_2330), .A1(net_2329) );
CLKBUF_X2 inst_22222 ( .A(net_21746), .Z(net_22094) );
INV_X4 inst_13731 ( .ZN(net_7768), .A(net_7767) );
NAND2_X2 inst_9227 ( .ZN(net_20605), .A2(net_10171), .A1(net_3474) );
XNOR2_X2 inst_218 ( .ZN(net_17594), .B(net_17526), .A(net_17339) );
NOR2_X2 inst_3647 ( .ZN(net_11680), .A2(net_11679), .A1(net_11134) );
INV_X4 inst_14773 ( .ZN(net_5679), .A(net_4048) );
AOI21_X2 inst_20523 ( .ZN(net_14560), .B2(net_11951), .A(net_8955), .B1(net_855) );
AOI22_X2 inst_19962 ( .ZN(net_16126), .A1(net_16125), .A2(net_15728), .B2(net_13166), .B1(net_3390) );
INV_X2 inst_19709 ( .A(net_20578), .ZN(net_20577) );
NAND2_X2 inst_11865 ( .A1(net_2327), .ZN(net_1653), .A2(net_997) );
INV_X4 inst_18094 ( .A(net_21042), .ZN(net_384) );
NAND2_X2 inst_11098 ( .A1(net_9943), .ZN(net_8881), .A2(net_4341) );
NAND2_X2 inst_8226 ( .ZN(net_17796), .A1(net_17692), .A2(net_17376) );
NAND2_X2 inst_10706 ( .A1(net_9591), .ZN(net_6023), .A2(net_2537) );
NAND3_X2 inst_6228 ( .ZN(net_13232), .A3(net_13231), .A2(net_9462), .A1(net_5628) );
INV_X4 inst_15877 ( .ZN(net_1931), .A(net_1182) );
AOI221_X2 inst_20079 ( .ZN(net_16099), .C2(net_15566), .B2(net_14357), .A(net_10135), .B1(net_9764), .C1(net_1052) );
NAND4_X4 inst_5236 ( .A1(net_20643), .ZN(net_15733), .A3(net_13630), .A2(net_13567), .A4(net_11584) );
INV_X4 inst_16602 ( .ZN(net_1132), .A(net_828) );
NAND4_X2 inst_5357 ( .ZN(net_20829), .A2(net_19053), .A1(net_19052), .A4(net_5276), .A3(net_4738) );
INV_X4 inst_12992 ( .A(net_16491), .ZN(net_16490) );
INV_X4 inst_14204 ( .ZN(net_12958), .A(net_5932) );
INV_X4 inst_16001 ( .ZN(net_2500), .A(net_1665) );
INV_X4 inst_14104 ( .A(net_6171), .ZN(net_6170) );
NAND2_X2 inst_9467 ( .ZN(net_11483), .A1(net_11482), .A2(net_11444) );
AND2_X4 inst_21206 ( .A2(net_9073), .A1(net_8995), .ZN(net_7294) );
INV_X4 inst_18277 ( .A(net_19462), .ZN(net_19461) );
INV_X4 inst_17403 ( .ZN(net_515), .A(net_103) );
INV_X8 inst_12231 ( .ZN(net_6077), .A(net_4826) );
NOR3_X2 inst_2682 ( .ZN(net_14559), .A1(net_12706), .A3(net_11812), .A2(net_11253) );
NAND2_X2 inst_8517 ( .ZN(net_16913), .A2(net_16912), .A1(net_16658) );
INV_X8 inst_12434 ( .ZN(net_20068), .A(net_16381) );
NOR2_X2 inst_4699 ( .A1(net_5479), .ZN(net_4143), .A2(net_3173) );
NAND2_X2 inst_10023 ( .A1(net_12708), .ZN(net_12007), .A2(net_8099) );
AOI21_X2 inst_20697 ( .ZN(net_12155), .A(net_11113), .B1(net_9966), .B2(net_8036) );
NOR2_X2 inst_4749 ( .A1(net_3148), .ZN(net_3021), .A2(net_3020) );
SDFF_X2 inst_964 ( .QN(net_21016), .D(net_392), .SE(net_263), .CK(net_21898), .SI(x2767) );
INV_X4 inst_16772 ( .ZN(net_1349), .A(net_1158) );
CLKBUF_X2 inst_21997 ( .A(net_21868), .Z(net_21869) );
NOR2_X2 inst_3372 ( .A2(net_17483), .ZN(net_16674), .A1(net_96) );
NAND2_X2 inst_7940 ( .ZN(net_18424), .A2(net_18366), .A1(net_18306) );
NAND2_X2 inst_10165 ( .A1(net_11345), .ZN(net_9724), .A2(net_8245) );
OAI21_X2 inst_2313 ( .ZN(net_5736), .A(net_5735), .B2(net_5629), .B1(net_2811) );
NAND3_X2 inst_6422 ( .ZN(net_20174), .A3(net_11941), .A1(net_9242), .A2(net_8316) );
CLKBUF_X2 inst_21648 ( .A(net_21519), .Z(net_21520) );
NAND2_X2 inst_10649 ( .ZN(net_6355), .A1(net_6354), .A2(net_6353) );
INV_X4 inst_14778 ( .ZN(net_7204), .A(net_5709) );
INV_X4 inst_12660 ( .ZN(net_17814), .A(net_17813) );
AOI21_X2 inst_20438 ( .ZN(net_15139), .B1(net_14972), .B2(net_13332), .A(net_8267) );
INV_X4 inst_12629 ( .ZN(net_17923), .A(net_17877) );
INV_X4 inst_14030 ( .ZN(net_11293), .A(net_6278) );
INV_X4 inst_12965 ( .A(net_16524), .ZN(net_16523) );
NAND3_X2 inst_6114 ( .ZN(net_19564), .A3(net_13103), .A1(net_11452), .A2(net_8772) );
INV_X4 inst_15359 ( .A(net_8618), .ZN(net_3383) );
NAND3_X2 inst_6193 ( .ZN(net_13315), .A3(net_9863), .A1(net_8405), .A2(net_4320) );
NOR2_X4 inst_3001 ( .ZN(net_9357), .A2(net_5875), .A1(net_5874) );
INV_X4 inst_18032 ( .A(net_20969), .ZN(net_888) );
INV_X4 inst_14111 ( .ZN(net_9710), .A(net_6156) );
INV_X4 inst_13741 ( .A(net_13442), .ZN(net_7642) );
NOR2_X4 inst_2818 ( .A2(net_19659), .A1(net_19658), .ZN(net_18941) );
NOR2_X4 inst_3198 ( .ZN(net_5560), .A2(net_3036), .A1(net_2955) );
INV_X4 inst_15893 ( .ZN(net_20298), .A(net_2293) );
NAND2_X2 inst_7979 ( .ZN(net_18345), .A2(net_18240), .A1(net_17192) );
NOR2_X4 inst_2904 ( .ZN(net_8922), .A2(net_6501), .A1(net_5233) );
NAND2_X2 inst_10075 ( .ZN(net_12120), .A2(net_7821), .A1(net_4340) );
INV_X2 inst_19092 ( .ZN(net_4554), .A(net_4553) );
OAI211_X2 inst_2383 ( .C2(net_20936), .ZN(net_18598), .C1(net_16015), .A(net_13828), .B(net_13798) );
OAI21_X2 inst_1701 ( .ZN(net_15313), .B1(net_15312), .A(net_14376), .B2(net_7726) );
INV_X4 inst_16933 ( .ZN(net_5153), .A(net_3108) );
INV_X4 inst_12853 ( .A(net_17571), .ZN(net_17376) );
AOI21_X2 inst_20765 ( .ZN(net_10766), .B1(net_10765), .B2(net_9151), .A(net_5349) );
INV_X4 inst_13853 ( .ZN(net_19281), .A(net_7466) );
NAND2_X2 inst_10401 ( .ZN(net_13122), .A1(net_10504), .A2(net_5540) );
INV_X4 inst_13577 ( .ZN(net_9116), .A(net_9115) );
AOI211_X4 inst_20992 ( .ZN(net_19136), .B(net_15548), .C2(net_15433), .A(net_15278), .C1(net_3306) );
NOR2_X2 inst_4987 ( .ZN(net_11651), .A2(net_1469), .A1(net_749) );
NAND2_X2 inst_9667 ( .ZN(net_10313), .A1(net_9174), .A2(net_8103) );
INV_X8 inst_12262 ( .ZN(net_3829), .A(net_2981) );
CLKBUF_X2 inst_21833 ( .A(net_21704), .Z(net_21705) );
NAND2_X2 inst_9838 ( .ZN(net_12254), .A2(net_7927), .A1(net_1187) );
NAND2_X2 inst_9627 ( .ZN(net_18885), .A2(net_7238), .A1(net_5469) );
NAND2_X2 inst_9163 ( .A1(net_14634), .ZN(net_13377), .A2(net_10576) );
CLKBUF_X2 inst_22636 ( .A(net_22507), .Z(net_22508) );
INV_X4 inst_13405 ( .ZN(net_13965), .A(net_8932) );
NAND2_X2 inst_8593 ( .A2(net_17815), .A1(net_16694), .ZN(net_16692) );
DFF_X2 inst_19775 ( .D(net_7354), .Q(net_27), .CK(net_22274) );
INV_X4 inst_14899 ( .ZN(net_3625), .A(net_3624) );
NAND2_X4 inst_7228 ( .ZN(net_10708), .A1(net_9061), .A2(net_5946) );
INV_X4 inst_12503 ( .ZN(net_18663), .A(net_18615) );
NAND2_X2 inst_9671 ( .A1(net_14321), .ZN(net_10307), .A2(net_10306) );
OR2_X2 inst_1135 ( .ZN(net_18983), .A2(net_12616), .A1(net_9176) );
AND2_X4 inst_21165 ( .ZN(net_19983), .A1(net_14537), .A2(net_10402) );
NAND2_X2 inst_8333 ( .ZN(net_19730), .A2(net_17334), .A1(net_16700) );
NAND2_X2 inst_11871 ( .ZN(net_2530), .A2(net_1636), .A1(net_683) );
INV_X4 inst_14419 ( .ZN(net_19945), .A(net_6716) );
NOR2_X4 inst_3127 ( .ZN(net_6740), .A1(net_3790), .A2(net_1991) );
NAND2_X2 inst_10945 ( .ZN(net_8348), .A2(net_5091), .A1(net_809) );
NAND2_X2 inst_8822 ( .ZN(net_19370), .A2(net_14831), .A1(net_13650) );
INV_X4 inst_17595 ( .A(net_6078), .ZN(net_884) );
NOR2_X4 inst_3243 ( .ZN(net_4341), .A1(net_3919), .A2(net_1905) );
INV_X4 inst_14039 ( .ZN(net_7621), .A(net_6269) );
NAND2_X2 inst_8605 ( .A2(net_20765), .ZN(net_19638), .A1(net_15519) );
NAND2_X2 inst_10564 ( .ZN(net_8769), .A1(net_7874), .A2(net_6841) );
INV_X2 inst_19223 ( .A(net_5037), .ZN(net_3443) );
OAI22_X2 inst_1266 ( .B1(net_21176), .ZN(net_17127), .B2(net_17126), .A1(net_16842), .A2(net_16640) );
NAND2_X2 inst_8904 ( .ZN(net_19518), .A2(net_14047), .A1(net_7775) );
NOR2_X2 inst_5102 ( .A2(net_1848), .ZN(net_768), .A1(net_152) );
NOR2_X2 inst_4872 ( .ZN(net_2222), .A2(net_2221), .A1(net_1406) );
INV_X4 inst_15781 ( .A(net_3023), .ZN(net_2834) );
NAND2_X4 inst_7216 ( .ZN(net_12076), .A2(net_6606), .A1(net_5823) );
NAND3_X2 inst_6287 ( .ZN(net_12843), .A3(net_12842), .A2(net_11598), .A1(net_9775) );
NOR2_X2 inst_4317 ( .A2(net_20783), .A1(net_10415), .ZN(net_5886) );
INV_X4 inst_13310 ( .A(net_13125), .ZN(net_11687) );
NAND2_X4 inst_7090 ( .A1(net_20135), .ZN(net_14960), .A2(net_13026) );
NAND2_X2 inst_11379 ( .ZN(net_4562), .A1(net_4110), .A2(net_2058) );
OAI21_X2 inst_1838 ( .A(net_14731), .ZN(net_14031), .B1(net_11144), .B2(net_8512) );
CLKBUF_X2 inst_22211 ( .A(net_22082), .Z(net_22083) );
NAND2_X2 inst_9414 ( .ZN(net_11652), .A1(net_11651), .A2(net_9297) );
OAI21_X4 inst_1454 ( .ZN(net_15348), .B2(net_13674), .B1(net_11694), .A(net_1402) );
NAND2_X2 inst_9438 ( .A2(net_13883), .A1(net_12987), .ZN(net_11570) );
CLKBUF_X2 inst_22541 ( .A(net_22357), .Z(net_22413) );
NOR2_X4 inst_3147 ( .ZN(net_4742), .A2(net_3187), .A1(net_1700) );
OAI21_X2 inst_1945 ( .ZN(net_12592), .B2(net_9120), .B1(net_6449), .A(net_855) );
INV_X4 inst_16643 ( .ZN(net_3592), .A(net_1100) );
NAND3_X4 inst_5564 ( .A3(net_20629), .A1(net_20628), .ZN(net_20358), .A2(net_13992) );
NOR3_X2 inst_2657 ( .ZN(net_15170), .A3(net_14996), .A1(net_14546), .A2(net_9555) );
CLKBUF_X2 inst_22527 ( .A(net_22398), .Z(net_22399) );
NAND3_X2 inst_5722 ( .ZN(net_19572), .A3(net_15654), .A2(net_15222), .A1(net_8317) );
CLKBUF_X2 inst_21963 ( .A(net_21244), .Z(net_21835) );
INV_X4 inst_14581 ( .ZN(net_7900), .A(net_4501) );
NAND2_X2 inst_7720 ( .ZN(net_18839), .A2(net_18818), .A1(net_18801) );
INV_X4 inst_13239 ( .ZN(net_13409), .A(net_12352) );
INV_X4 inst_13043 ( .ZN(net_19230), .A(net_16374) );
INV_X4 inst_12930 ( .ZN(net_17008), .A(net_17006) );
XNOR2_X2 inst_376 ( .A(net_17760), .ZN(net_16838), .B(net_1896) );
INV_X2 inst_19304 ( .A(net_6399), .ZN(net_2756) );
NAND2_X2 inst_10816 ( .ZN(net_20350), .A1(net_5509), .A2(net_2404) );
INV_X4 inst_15356 ( .ZN(net_14837), .A(net_10011) );
NOR2_X4 inst_3268 ( .ZN(net_3736), .A1(net_2597), .A2(net_1651) );
INV_X4 inst_14066 ( .ZN(net_9550), .A(net_6241) );
INV_X4 inst_17877 ( .A(net_1790), .ZN(net_226) );
NAND2_X2 inst_11676 ( .A1(net_20860), .A2(net_2402), .ZN(net_2354) );
INV_X4 inst_14840 ( .ZN(net_6893), .A(net_2560) );
MUX2_X2 inst_12167 ( .Z(net_20288), .S(net_15099), .A(net_12798), .B(net_11853) );
NAND2_X2 inst_7856 ( .ZN(net_18574), .A2(net_18562), .A1(net_18451) );
NAND2_X2 inst_10991 ( .A2(net_6445), .ZN(net_4929), .A1(net_90) );
NAND2_X2 inst_8897 ( .ZN(net_15105), .A1(net_15104), .A2(net_13887) );
NAND3_X2 inst_6299 ( .ZN(net_12811), .A3(net_12774), .A2(net_4771), .A1(net_3843) );
INV_X4 inst_18250 ( .A(net_21224), .ZN(net_222) );
INV_X4 inst_12627 ( .ZN(net_17951), .A(net_17950) );
CLKBUF_X2 inst_22306 ( .A(net_21855), .Z(net_22178) );
INV_X4 inst_13251 ( .ZN(net_12786), .A(net_11785) );
NAND2_X2 inst_10852 ( .ZN(net_7229), .A2(net_5433), .A1(net_809) );
NAND2_X2 inst_9951 ( .ZN(net_10421), .A1(net_8938), .A2(net_8937) );
NOR2_X2 inst_3880 ( .A1(net_14458), .ZN(net_9318), .A2(net_9317) );
NOR2_X4 inst_3100 ( .A1(net_6407), .ZN(net_5228), .A2(net_4183) );
NAND2_X2 inst_8359 ( .A2(net_19456), .ZN(net_17425), .A1(net_557) );
NOR2_X2 inst_4052 ( .ZN(net_7853), .A1(net_7852), .A2(net_4938) );
NAND2_X2 inst_8552 ( .ZN(net_16790), .A1(net_16789), .A2(net_16628) );
NOR2_X2 inst_4251 ( .A1(net_9733), .ZN(net_6371), .A2(net_4600) );
CLKBUF_X2 inst_22599 ( .A(net_22470), .Z(net_22471) );
NOR2_X2 inst_4487 ( .ZN(net_6581), .A2(net_3797), .A1(net_583) );
OAI21_X2 inst_1596 ( .A(net_20920), .ZN(net_16208), .B2(net_15854), .B1(net_9501) );
NOR2_X2 inst_4364 ( .ZN(net_5495), .A2(net_5494), .A1(net_3920) );
INV_X4 inst_15313 ( .ZN(net_3951), .A(net_2381) );
CLKBUF_X2 inst_21809 ( .A(net_21680), .Z(net_21681) );
INV_X4 inst_15788 ( .A(net_15666), .ZN(net_1906) );
NAND3_X2 inst_6400 ( .ZN(net_11989), .A3(net_11830), .A1(net_10783), .A2(net_5907) );
NAND2_X4 inst_7078 ( .A1(net_19637), .ZN(net_15832), .A2(net_15831) );
CLKBUF_X2 inst_22370 ( .A(net_21347), .Z(net_22242) );
INV_X4 inst_17145 ( .ZN(net_19670), .A(net_760) );
NAND2_X2 inst_10174 ( .ZN(net_8206), .A1(net_8205), .A2(net_8204) );
OAI21_X2 inst_2265 ( .ZN(net_7154), .A(net_7153), .B1(net_4003), .B2(net_3374) );
INV_X4 inst_13494 ( .ZN(net_11515), .A(net_9468) );
OAI21_X2 inst_1555 ( .ZN(net_17638), .B2(net_17571), .A(net_17347), .B1(net_17346) );
OAI22_X2 inst_1293 ( .ZN(net_12476), .A2(net_12475), .B2(net_12474), .B1(net_10993), .A1(net_10829) );
NAND2_X4 inst_7132 ( .ZN(net_14547), .A1(net_10206), .A2(net_9616) );
NOR2_X2 inst_3805 ( .ZN(net_9841), .A2(net_6301), .A1(net_5995) );
XNOR2_X2 inst_280 ( .ZN(net_17171), .A(net_17170), .B(net_13287) );
NAND2_X2 inst_11249 ( .ZN(net_20124), .A1(net_3919), .A2(net_3197) );
NOR2_X4 inst_3157 ( .ZN(net_6684), .A2(net_3861), .A1(net_3068) );
AOI21_X2 inst_20259 ( .A(net_18601), .ZN(net_18594), .B2(net_15492), .B1(net_13421) );
NAND2_X2 inst_9888 ( .ZN(net_10911), .A1(net_9418), .A2(net_8061) );
NAND2_X2 inst_11657 ( .ZN(net_4355), .A2(net_1718), .A1(net_222) );
INV_X4 inst_13648 ( .ZN(net_14391), .A(net_8157) );
NOR2_X2 inst_4676 ( .ZN(net_3473), .A1(net_3239), .A2(net_3238) );
INV_X4 inst_17340 ( .ZN(net_6884), .A(net_824) );
INV_X4 inst_16958 ( .ZN(net_11468), .A(net_904) );
INV_X4 inst_14071 ( .ZN(net_7577), .A(net_3421) );
INV_X2 inst_19129 ( .A(net_5611), .ZN(net_4281) );
INV_X4 inst_16729 ( .A(net_15468), .ZN(net_1051) );
NAND2_X2 inst_8110 ( .A2(net_20443), .ZN(net_18109), .A1(net_17139) );
NAND2_X2 inst_11556 ( .ZN(net_2838), .A2(net_2495), .A1(net_1601) );
INV_X4 inst_14789 ( .ZN(net_4559), .A(net_3097) );
NAND2_X2 inst_10344 ( .A1(net_7677), .ZN(net_7520), .A2(net_7519) );
INV_X2 inst_19361 ( .A(net_3138), .ZN(net_2287) );
NAND3_X2 inst_6586 ( .A3(net_11374), .ZN(net_10427), .A2(net_10426), .A1(net_5985) );
INV_X4 inst_15332 ( .ZN(net_3535), .A(net_2609) );
NAND2_X2 inst_11188 ( .ZN(net_10781), .A1(net_4707), .A2(net_4209) );
AOI21_X2 inst_20472 ( .ZN(net_14977), .B2(net_12826), .A(net_7200), .B1(net_449) );
INV_X4 inst_17284 ( .ZN(net_3185), .A(net_1614) );
NOR2_X2 inst_4393 ( .ZN(net_18987), .A1(net_13938), .A2(net_5197) );
AOI21_X2 inst_20784 ( .A(net_14022), .ZN(net_10554), .B1(net_10553), .B2(net_3468) );
NAND2_X2 inst_8299 ( .ZN(net_17601), .A2(net_17600), .A1(net_17411) );
INV_X4 inst_12743 ( .ZN(net_17433), .A(net_17432) );
INV_X4 inst_17677 ( .ZN(net_239), .A(net_238) );
INV_X4 inst_14780 ( .ZN(net_6862), .A(net_5114) );
INV_X4 inst_18348 ( .A(net_20789), .ZN(net_20788) );
OAI21_X4 inst_1359 ( .ZN(net_18098), .A(net_18075), .B2(net_18070), .B1(net_16133) );
AOI21_X2 inst_20443 ( .ZN(net_15122), .B1(net_15121), .B2(net_13181), .A(net_12135) );
NAND2_X2 inst_10345 ( .ZN(net_9174), .A2(net_7494), .A1(net_6876) );
NAND2_X4 inst_7499 ( .ZN(net_3566), .A1(net_2315), .A2(net_1765) );
INV_X4 inst_14522 ( .ZN(net_7163), .A(net_4778) );
INV_X2 inst_19460 ( .A(net_1876), .ZN(net_1497) );
INV_X4 inst_17209 ( .A(net_13030), .ZN(net_12928) );
NAND2_X2 inst_11328 ( .ZN(net_7025), .A1(net_3737), .A2(net_2155) );
NOR2_X2 inst_3797 ( .ZN(net_10024), .A1(net_6897), .A2(net_6787) );
XNOR2_X2 inst_100 ( .ZN(net_18535), .A(net_18428), .B(net_18335) );
NOR2_X2 inst_4352 ( .ZN(net_19149), .A1(net_6530), .A2(net_5689) );
XNOR2_X2 inst_279 ( .ZN(net_17172), .A(net_17166), .B(net_13294) );
INV_X2 inst_18468 ( .ZN(net_12719), .A(net_11662) );
NOR2_X2 inst_3387 ( .ZN(net_19498), .A2(net_16066), .A1(net_16029) );
NAND2_X2 inst_11683 ( .A1(net_3750), .ZN(net_3140), .A2(net_2075) );
NAND2_X2 inst_11014 ( .ZN(net_4856), .A1(net_4855), .A2(net_4854) );
NAND2_X2 inst_8271 ( .A2(net_20518), .ZN(net_17652), .A1(net_17651) );
XNOR2_X2 inst_81 ( .B(net_21156), .ZN(net_18657), .A(net_18642) );
NAND3_X2 inst_5806 ( .A3(net_19735), .A1(net_19734), .ZN(net_19595), .A2(net_13420) );
INV_X4 inst_13424 ( .ZN(net_19896), .A(net_8579) );
NAND2_X2 inst_9761 ( .ZN(net_19752), .A2(net_9314), .A1(net_4149) );
NAND2_X4 inst_7087 ( .A1(net_19593), .ZN(net_19023), .A2(net_15366) );
NAND2_X2 inst_9471 ( .ZN(net_11474), .A2(net_10906), .A1(net_9926) );
INV_X4 inst_14411 ( .ZN(net_11391), .A(net_6860) );
NAND2_X2 inst_12040 ( .A1(net_1848), .ZN(net_1129), .A2(net_954) );
AOI21_X2 inst_20594 ( .ZN(net_13930), .B2(net_11184), .A(net_8796), .B1(net_8674) );
CLKBUF_X2 inst_21768 ( .A(net_21607), .Z(net_21640) );
AOI21_X2 inst_20857 ( .ZN(net_8904), .B2(net_8057), .B1(net_3613), .A(net_761) );
AOI21_X2 inst_20644 ( .ZN(net_13189), .B1(net_12295), .B2(net_10249), .A(net_6569) );
NOR2_X4 inst_2954 ( .ZN(net_8721), .A2(net_5176), .A1(net_2585) );
CLKBUF_X2 inst_22118 ( .A(net_21989), .Z(net_21990) );
NAND2_X2 inst_9711 ( .ZN(net_10180), .A1(net_10179), .A2(net_10178) );
NAND2_X2 inst_12045 ( .ZN(net_1055), .A2(net_523), .A1(net_84) );
NAND2_X2 inst_11844 ( .A2(net_2744), .A1(net_1784), .ZN(net_1717) );
OAI21_X2 inst_2197 ( .A(net_10162), .ZN(net_8576), .B2(net_8575), .B1(net_3647) );
NAND2_X2 inst_7995 ( .ZN(net_18320), .A2(net_18319), .A1(net_17419) );
INV_X4 inst_13064 ( .ZN(net_19547), .A(net_16273) );
OAI211_X2 inst_2582 ( .ZN(net_7670), .B(net_7669), .C2(net_7133), .C1(net_5836), .A(net_4962) );
XNOR2_X2 inst_142 ( .B(net_21192), .ZN(net_18172), .A(net_18171) );
AOI21_X4 inst_20228 ( .ZN(net_19975), .B2(net_13619), .B1(net_12334), .A(net_6510) );
XNOR2_X2 inst_78 ( .B(net_20523), .ZN(net_18693), .A(net_18629) );
INV_X4 inst_13182 ( .ZN(net_14318), .A(net_13847) );
NAND2_X2 inst_7896 ( .ZN(net_18486), .A2(net_18435), .A1(net_17917) );
AOI22_X2 inst_19964 ( .ZN(net_16039), .B1(net_15537), .A2(net_15521), .B2(net_13158), .A1(net_5655) );
NOR2_X4 inst_2813 ( .ZN(net_17460), .A1(net_16827), .A2(net_16672) );
XNOR2_X2 inst_177 ( .B(net_21129), .ZN(net_17773), .A(net_17771) );
SDFF_X2 inst_783 ( .Q(net_20918), .SE(net_18804), .SI(net_18042), .D(net_682), .CK(net_21284) );
NAND2_X2 inst_7910 ( .ZN(net_18465), .A1(net_18412), .A2(net_17567) );
AND2_X4 inst_21184 ( .A1(net_15366), .ZN(net_11539), .A2(net_11538) );
NAND2_X2 inst_8450 ( .ZN(net_19220), .A2(net_17441), .A1(net_17099) );
NAND3_X2 inst_5696 ( .ZN(net_16254), .A3(net_15945), .A2(net_14856), .A1(net_12209) );
OAI21_X2 inst_2014 ( .ZN(net_11377), .A(net_11376), .B2(net_11295), .B1(net_5582) );
CLKBUF_X2 inst_22147 ( .A(net_22018), .Z(net_22019) );
INV_X4 inst_14610 ( .ZN(net_6046), .A(net_4431) );
NAND3_X2 inst_6122 ( .ZN(net_13844), .A2(net_13843), .A3(net_13842), .A1(net_5424) );
NAND2_X2 inst_10144 ( .ZN(net_8305), .A2(net_6180), .A1(net_4773) );
CLKBUF_X2 inst_22419 ( .A(net_22290), .Z(net_22291) );
INV_X4 inst_12821 ( .ZN(net_17186), .A(net_17185) );
NAND2_X2 inst_9999 ( .ZN(net_8827), .A2(net_8826), .A1(net_7227) );
INV_X2 inst_19531 ( .A(net_2976), .ZN(net_998) );
NOR2_X4 inst_2822 ( .ZN(net_16286), .A2(net_16153), .A1(net_16147) );
OAI211_X2 inst_2467 ( .B(net_20111), .A(net_20110), .ZN(net_19621), .C2(net_11915), .C1(net_10031) );
CLKBUF_X2 inst_22180 ( .A(net_21522), .Z(net_22052) );
NAND3_X2 inst_6176 ( .ZN(net_13543), .A1(net_13542), .A3(net_9186), .A2(net_2665) );
NAND2_X2 inst_10335 ( .ZN(net_20293), .A2(net_9252), .A1(net_7580) );
NAND2_X2 inst_8656 ( .ZN(net_19061), .A2(net_16397), .A1(net_16394) );
OAI21_X2 inst_2031 ( .ZN(net_20283), .A(net_11264), .B2(net_10467), .B1(net_9510) );
INV_X2 inst_18471 ( .ZN(net_12696), .A(net_12695) );
NOR2_X2 inst_4386 ( .ZN(net_8431), .A2(net_5208), .A1(net_761) );
INV_X4 inst_15367 ( .ZN(net_4044), .A(net_2575) );
INV_X4 inst_14797 ( .ZN(net_3996), .A(net_3995) );
NAND2_X2 inst_11282 ( .ZN(net_9875), .A2(net_2398), .A1(net_535) );
INV_X4 inst_16839 ( .ZN(net_7886), .A(net_4737) );
CLKBUF_X2 inst_22156 ( .A(net_22027), .Z(net_22028) );
NAND2_X2 inst_11527 ( .A1(net_7244), .ZN(net_2968), .A2(net_2967) );
NAND2_X2 inst_8525 ( .A2(net_20434), .ZN(net_19886), .A1(net_19430) );
INV_X4 inst_17937 ( .A(net_21014), .ZN(net_641) );
XNOR2_X2 inst_338 ( .ZN(net_16984), .A(net_16983), .B(net_16982) );
INV_X4 inst_16077 ( .ZN(net_6655), .A(net_1773) );
NAND3_X4 inst_5577 ( .A3(net_20631), .A1(net_20630), .ZN(net_15737), .A2(net_14726) );
NOR2_X2 inst_4005 ( .ZN(net_9605), .A1(net_9131), .A2(net_8100) );
NAND4_X2 inst_5424 ( .ZN(net_14192), .A4(net_12149), .A2(net_11165), .A3(net_8802), .A1(net_4710) );
NOR2_X2 inst_4323 ( .ZN(net_5863), .A2(net_3411), .A1(net_3344) );
INV_X4 inst_17235 ( .ZN(net_2490), .A(net_663) );
CLKBUF_X2 inst_21594 ( .A(net_21315), .Z(net_21466) );
INV_X4 inst_15212 ( .A(net_6400), .ZN(net_2890) );
NAND3_X2 inst_6468 ( .ZN(net_11356), .A3(net_7567), .A2(net_5002), .A1(net_3653) );
INV_X4 inst_17397 ( .ZN(net_5476), .A(net_655) );
OAI211_X2 inst_2474 ( .ZN(net_13653), .C1(net_13504), .B(net_11956), .C2(net_9286), .A(net_8258) );
XNOR2_X2 inst_579 ( .B(net_16646), .ZN(net_611), .A(net_610) );
NAND4_X4 inst_5247 ( .A2(net_20736), .A1(net_20735), .ZN(net_20670), .A3(net_11731), .A4(net_11106) );
CLKBUF_X2 inst_22364 ( .A(net_22235), .Z(net_22236) );
NAND2_X4 inst_7462 ( .ZN(net_5445), .A1(net_2746), .A2(net_2745) );
CLKBUF_X2 inst_22343 ( .A(net_22214), .Z(net_22215) );
SDFF_X2 inst_698 ( .Q(net_20863), .SI(net_18839), .SE(net_18576), .D(net_490), .CK(net_22041) );
INV_X4 inst_14378 ( .ZN(net_20618), .A(net_5174) );
NOR2_X2 inst_3964 ( .ZN(net_8422), .A1(net_8421), .A2(net_6556) );
NOR2_X2 inst_3944 ( .ZN(net_19479), .A2(net_8632), .A1(net_8631) );
NOR2_X2 inst_3394 ( .ZN(net_15985), .A2(net_15817), .A1(net_11961) );
INV_X4 inst_17280 ( .ZN(net_4110), .A(net_640) );
INV_X4 inst_17716 ( .ZN(net_405), .A(net_86) );
NAND3_X2 inst_5978 ( .ZN(net_14608), .A2(net_14226), .A3(net_13910), .A1(net_13243) );
NOR2_X4 inst_2863 ( .ZN(net_20308), .A2(net_11426), .A1(net_11425) );
NAND2_X2 inst_8401 ( .ZN(net_17386), .A1(net_16960), .A2(net_16797) );
INV_X4 inst_12882 ( .A(net_16919), .ZN(net_16822) );
INV_X4 inst_15565 ( .ZN(net_3883), .A(net_2295) );
NOR2_X2 inst_3897 ( .A2(net_10847), .ZN(net_9120), .A1(net_60) );
NAND3_X4 inst_5534 ( .A3(net_19152), .A1(net_19151), .ZN(net_18211), .A2(net_16118) );
INV_X4 inst_15897 ( .ZN(net_1772), .A(net_1771) );
NAND2_X2 inst_11458 ( .ZN(net_3218), .A2(net_3217), .A1(net_3095) );
NAND2_X2 inst_11693 ( .A2(net_9360), .ZN(net_2322), .A1(net_2321) );
NOR2_X2 inst_3754 ( .ZN(net_20057), .A2(net_10385), .A1(net_8370) );
NAND3_X2 inst_6160 ( .A3(net_20407), .ZN(net_13645), .A1(net_13644), .A2(net_10261) );
INV_X4 inst_15419 ( .ZN(net_4035), .A(net_3036) );
NAND2_X2 inst_10229 ( .ZN(net_9587), .A2(net_6220), .A1(net_6131) );
SDFF_X2 inst_837 ( .Q(net_21183), .SI(net_17453), .SE(net_125), .CK(net_21555), .D(x6544) );
NAND3_X2 inst_5716 ( .ZN(net_19992), .A3(net_15716), .A1(net_14614), .A2(net_14168) );
AOI21_X4 inst_20131 ( .B1(net_19708), .ZN(net_16092), .B2(net_15742), .A(net_14243) );
INV_X2 inst_19452 ( .ZN(net_1550), .A(net_238) );
INV_X4 inst_14425 ( .ZN(net_8288), .A(net_5046) );
CLKBUF_X2 inst_22488 ( .A(net_22359), .Z(net_22360) );
NAND2_X2 inst_8956 ( .ZN(net_14717), .A1(net_13452), .A2(net_13212) );
NAND3_X2 inst_6509 ( .ZN(net_10789), .A3(net_10733), .A2(net_6658), .A1(net_5636) );
NAND4_X2 inst_5457 ( .ZN(net_13435), .A3(net_11279), .A4(net_9987), .A2(net_9871), .A1(net_7020) );
NAND2_X4 inst_7025 ( .ZN(net_17235), .A1(net_16587), .A2(net_16459) );
INV_X4 inst_14997 ( .ZN(net_20024), .A(net_3537) );
NAND2_X2 inst_8785 ( .ZN(net_19176), .A1(net_15688), .A2(net_15379) );
NAND2_X2 inst_7798 ( .ZN(net_18776), .A2(net_18703), .A1(net_17632) );
NAND2_X2 inst_10497 ( .ZN(net_10428), .A1(net_7858), .A2(net_6946) );
NAND2_X4 inst_7664 ( .ZN(net_1230), .A2(net_1025), .A1(net_108) );
CLKBUF_X2 inst_21490 ( .A(net_21361), .Z(net_21362) );
XNOR2_X2 inst_65 ( .ZN(net_18806), .A(net_18750), .B(net_18650) );
INV_X8 inst_12443 ( .ZN(net_20502), .A(net_20501) );
NAND2_X2 inst_9563 ( .ZN(net_12373), .A2(net_11017), .A1(net_5799) );
NOR2_X2 inst_3592 ( .A1(net_14515), .ZN(net_12606), .A2(net_12605) );
NAND3_X1 inst_6822 ( .A3(net_12999), .ZN(net_12948), .A2(net_11984), .A1(net_4469) );
NOR2_X2 inst_5121 ( .A2(net_312), .ZN(net_292), .A1(net_291) );
NOR2_X2 inst_3732 ( .ZN(net_12635), .A2(net_10874), .A1(net_10395) );
INV_X4 inst_14931 ( .A(net_3931), .ZN(net_3545) );
AOI21_X2 inst_20377 ( .ZN(net_15564), .B2(net_14682), .A(net_9990), .B1(net_9080) );
NOR2_X2 inst_4503 ( .ZN(net_5381), .A1(net_4792), .A2(net_4248) );
AOI21_X2 inst_20651 ( .B2(net_20627), .B1(net_20626), .ZN(net_13052), .A(net_10699) );
NAND2_X2 inst_9658 ( .ZN(net_19906), .A1(net_10335), .A2(net_7758) );
NOR2_X2 inst_4907 ( .A1(net_4108), .ZN(net_1954), .A2(net_1953) );
NOR2_X4 inst_2926 ( .ZN(net_9414), .A2(net_7878), .A1(net_7877) );
CLKBUF_X2 inst_22841 ( .A(net_22712), .Z(net_22713) );
INV_X4 inst_16392 ( .A(net_15366), .ZN(net_15186) );
OR2_X2 inst_1158 ( .ZN(net_8108), .A1(net_8107), .A2(net_4671) );
INV_X2 inst_19314 ( .A(net_3410), .ZN(net_2654) );
INV_X4 inst_18312 ( .A(net_20508), .ZN(net_20507) );
NAND2_X2 inst_9059 ( .A1(net_14460), .ZN(net_13994), .A2(net_11993) );
OAI21_X2 inst_1870 ( .ZN(net_13711), .B2(net_13629), .A(net_11866), .B1(net_9726) );
INV_X4 inst_13445 ( .ZN(net_14410), .A(net_9771) );
INV_X2 inst_19408 ( .A(net_3546), .ZN(net_1979) );
NAND2_X4 inst_7038 ( .A2(net_20690), .A1(net_20689), .ZN(net_16979) );
NAND4_X2 inst_5270 ( .A2(net_19403), .A1(net_19402), .ZN(net_19217), .A4(net_15197), .A3(net_14235) );
AND2_X4 inst_21197 ( .ZN(net_10157), .A2(net_10156), .A1(net_9887) );
INV_X4 inst_15853 ( .ZN(net_2702), .A(net_1819) );
NAND2_X2 inst_8436 ( .ZN(net_17147), .A2(net_17146), .A1(net_17006) );
OAI211_X2 inst_2445 ( .ZN(net_14670), .B(net_14669), .C2(net_10776), .A(net_7501), .C1(net_6840) );
INV_X4 inst_16205 ( .ZN(net_2044), .A(net_1713) );
INV_X4 inst_14704 ( .ZN(net_6176), .A(net_4251) );
NOR2_X4 inst_3039 ( .ZN(net_8195), .A2(net_5107), .A1(net_5106) );
NAND4_X2 inst_5477 ( .A3(net_13010), .ZN(net_12839), .A2(net_12838), .A1(net_11707), .A4(net_11012) );
INV_X4 inst_17277 ( .A(net_14557), .ZN(net_14175) );
XNOR2_X2 inst_461 ( .B(net_16097), .ZN(net_13289), .A(net_9000) );
CLKBUF_X2 inst_22231 ( .A(net_21808), .Z(net_22103) );
NAND3_X2 inst_6092 ( .ZN(net_13935), .A2(net_13934), .A3(net_13862), .A1(net_12558) );
NAND2_X2 inst_8291 ( .ZN(net_17617), .A1(net_17616), .A2(net_17615) );
NAND3_X2 inst_6387 ( .A2(net_14321), .ZN(net_12015), .A3(net_10291), .A1(net_8141) );
OAI21_X2 inst_1973 ( .ZN(net_12199), .A(net_10087), .B2(net_7817), .B1(net_6900) );
NOR2_X4 inst_3051 ( .A1(net_8539), .ZN(net_6168), .A2(net_5008) );
NAND2_X2 inst_8326 ( .ZN(net_20666), .A2(net_17552), .A1(net_17520) );
NOR3_X2 inst_2668 ( .A3(net_19695), .A1(net_19694), .ZN(net_14831), .A2(net_10882) );
INV_X4 inst_14447 ( .ZN(net_6125), .A(net_3953) );
INV_X4 inst_14238 ( .ZN(net_5811), .A(net_5810) );
INV_X4 inst_17359 ( .ZN(net_5950), .A(net_4329) );
NAND3_X2 inst_5742 ( .ZN(net_19584), .A1(net_15669), .A3(net_15047), .A2(net_8108) );
INV_X2 inst_18862 ( .A(net_8197), .ZN(net_6308) );
NAND3_X2 inst_5775 ( .ZN(net_15891), .A3(net_15206), .A1(net_14760), .A2(net_12223) );
NOR2_X2 inst_4808 ( .A2(net_20493), .ZN(net_4017), .A1(net_4014) );
NOR2_X2 inst_4657 ( .A1(net_15108), .ZN(net_3802), .A2(net_81) );
OAI21_X2 inst_1669 ( .ZN(net_19828), .A(net_15366), .B2(net_14923), .B1(net_6961) );
NAND2_X4 inst_7456 ( .ZN(net_4749), .A2(net_1224), .A1(net_1034) );
INV_X2 inst_18973 ( .ZN(net_5222), .A(net_5221) );
INV_X4 inst_17695 ( .ZN(net_482), .A(net_219) );
INV_X4 inst_17690 ( .ZN(net_14563), .A(net_10087) );
INV_X8 inst_12195 ( .ZN(net_16721), .A(net_16380) );
INV_X2 inst_19411 ( .ZN(net_5272), .A(net_1973) );
INV_X2 inst_19082 ( .ZN(net_4585), .A(net_4584) );
NOR2_X4 inst_3162 ( .ZN(net_20211), .A2(net_3226), .A1(net_3225) );
CLKBUF_X2 inst_22165 ( .A(net_22036), .Z(net_22037) );
NOR2_X2 inst_3956 ( .ZN(net_8598), .A1(net_7989), .A2(net_6777) );
CLKBUF_X2 inst_22892 ( .A(net_22763), .Z(net_22764) );
AOI21_X2 inst_20733 ( .ZN(net_11740), .B2(net_11739), .B1(net_8338), .A(net_6118) );
OAI21_X2 inst_1801 ( .A(net_20897), .ZN(net_14480), .B2(net_11458), .B1(net_11190) );
INV_X4 inst_12777 ( .ZN(net_17446), .A(net_17320) );
CLKBUF_X2 inst_21391 ( .A(net_21262), .Z(net_21263) );
INV_X2 inst_19704 ( .A(net_20572), .ZN(net_20571) );
NAND2_X2 inst_9964 ( .ZN(net_8905), .A2(net_8211), .A1(net_5052) );
SDFF_X2 inst_720 ( .Q(net_20861), .SE(net_18837), .SI(net_18712), .D(net_794), .CK(net_22003) );
SDFF_X2 inst_958 ( .QN(net_20979), .D(net_2432), .SE(net_253), .CK(net_22674), .SI(x3332) );
INV_X8 inst_12412 ( .A(net_20893), .ZN(net_915) );
NAND2_X2 inst_10468 ( .ZN(net_11659), .A1(net_6999), .A2(net_6998) );
INV_X4 inst_13465 ( .A(net_11900), .ZN(net_9685) );
XNOR2_X2 inst_368 ( .ZN(net_16849), .A(net_16848), .B(net_13952) );
OAI21_X2 inst_1697 ( .ZN(net_19260), .A(net_14476), .B2(net_13675), .B1(net_11686) );
INV_X4 inst_14909 ( .A(net_4616), .ZN(net_3584) );
INV_X4 inst_14574 ( .ZN(net_6216), .A(net_5074) );
NAND2_X4 inst_6995 ( .ZN(net_17209), .A1(net_16739), .A2(net_16593) );
AND2_X2 inst_21292 ( .ZN(net_20629), .A1(net_11642), .A2(net_4445) );
INV_X4 inst_16269 ( .A(net_7975), .ZN(net_3700) );
AOI21_X2 inst_20723 ( .ZN(net_11977), .A(net_8101), .B2(net_7724), .B1(net_1721) );
CLKBUF_X2 inst_22702 ( .A(net_21272), .Z(net_22574) );
NOR2_X2 inst_3689 ( .ZN(net_11400), .A2(net_11399), .A1(net_4137) );
NOR2_X2 inst_3556 ( .ZN(net_13029), .A1(net_12635), .A2(net_10416) );
INV_X4 inst_17157 ( .A(net_1741), .ZN(net_1100) );
INV_X4 inst_17670 ( .ZN(net_916), .A(net_244) );
NAND2_X2 inst_8811 ( .ZN(net_15613), .A1(net_15612), .A2(net_14896) );
CLKBUF_X2 inst_22395 ( .A(net_21772), .Z(net_22267) );
OAI21_X2 inst_1966 ( .ZN(net_12258), .A(net_11597), .B2(net_8499), .B1(net_1245) );
NOR2_X2 inst_3914 ( .A2(net_13943), .ZN(net_10330), .A1(net_8722) );
CLKBUF_X2 inst_21921 ( .A(net_21792), .Z(net_21793) );
NOR2_X2 inst_4716 ( .A2(net_6237), .ZN(net_4411), .A1(net_3134) );
NAND2_X4 inst_6838 ( .ZN(net_18709), .A1(net_18671), .A2(net_18658) );
INV_X4 inst_18076 ( .A(net_21100), .ZN(net_632) );
OAI211_X2 inst_2435 ( .ZN(net_15006), .C2(net_12464), .B(net_9991), .A(net_8852), .C1(net_3067) );
INV_X4 inst_17946 ( .A(net_20995), .ZN(net_1866) );
INV_X4 inst_16673 ( .ZN(net_6636), .A(net_5008) );
INV_X4 inst_14078 ( .ZN(net_20753), .A(net_7899) );
CLKBUF_X2 inst_22013 ( .A(net_21884), .Z(net_21885) );
NAND2_X2 inst_10101 ( .ZN(net_8586), .A2(net_7029), .A1(net_816) );
INV_X4 inst_18210 ( .A(net_21047), .ZN(net_435) );
OAI21_X2 inst_1678 ( .B1(net_15636), .ZN(net_15491), .B2(net_14578), .A(net_10752) );
INV_X2 inst_19169 ( .ZN(net_5390), .A(net_5373) );
NAND2_X2 inst_11602 ( .A1(net_4794), .ZN(net_2658), .A2(net_2657) );
NAND2_X2 inst_10839 ( .ZN(net_8727), .A1(net_6091), .A2(net_5563) );
INV_X4 inst_15424 ( .ZN(net_2822), .A(net_2510) );
AOI21_X4 inst_20221 ( .B1(net_19610), .ZN(net_14099), .B2(net_14038), .A(net_7315) );
OAI21_X2 inst_2233 ( .ZN(net_7782), .A(net_7781), .B1(net_7780), .B2(net_1325) );
INV_X4 inst_17033 ( .ZN(net_1171), .A(net_843) );
NAND2_X4 inst_7266 ( .ZN(net_10610), .A1(net_6255), .A2(net_2744) );
CLKBUF_X2 inst_22003 ( .A(net_21582), .Z(net_21875) );
AOI22_X2 inst_20056 ( .B2(net_6696), .A1(net_5204), .ZN(net_2951), .A2(net_2950), .B1(net_1018) );
INV_X4 inst_14859 ( .ZN(net_3783), .A(net_3782) );
INV_X4 inst_13939 ( .ZN(net_6822), .A(net_6821) );
INV_X4 inst_13870 ( .A(net_9463), .ZN(net_9113) );
XNOR2_X2 inst_396 ( .A(net_16766), .ZN(net_16760), .B(net_16759) );
NOR2_X2 inst_3382 ( .A2(net_19835), .A1(net_19834), .ZN(net_19740) );
INV_X2 inst_19440 ( .ZN(net_1696), .A(net_1695) );
INV_X4 inst_15548 ( .ZN(net_2870), .A(net_2349) );
AOI21_X2 inst_20463 ( .ZN(net_15003), .B2(net_13009), .B1(net_10920), .A(net_7311) );
NOR2_X2 inst_3377 ( .ZN(net_19296), .A2(net_16388), .A1(net_13372) );
NOR2_X2 inst_5128 ( .ZN(net_2224), .A2(net_1848), .A1(net_703) );
CLKBUF_X2 inst_22451 ( .A(net_22322), .Z(net_22323) );
INV_X4 inst_14665 ( .ZN(net_4333), .A(net_4332) );
INV_X4 inst_14330 ( .A(net_8947), .ZN(net_5417) );
NAND2_X2 inst_10371 ( .ZN(net_7398), .A1(net_7397), .A2(net_4465) );
NAND2_X2 inst_11894 ( .ZN(net_3146), .A2(net_1420), .A1(net_903) );
INV_X2 inst_19324 ( .ZN(net_4942), .A(net_3977) );
INV_X4 inst_14992 ( .A(net_14395), .ZN(net_14264) );
AND2_X2 inst_21271 ( .ZN(net_18887), .A1(net_14535), .A2(net_12731) );
AOI21_X2 inst_20282 ( .B1(net_21228), .ZN(net_16264), .B2(net_15954), .A(net_15526) );
NOR2_X4 inst_2845 ( .ZN(net_20185), .A2(net_19567), .A1(net_19566) );
NAND2_X2 inst_7760 ( .ZN(net_18756), .A2(net_18702), .A1(net_16993) );
NOR2_X4 inst_2977 ( .ZN(net_9338), .A2(net_3500), .A1(net_3276) );
INV_X2 inst_19475 ( .A(net_2369), .ZN(net_1412) );
OR2_X4 inst_1092 ( .ZN(net_12072), .A2(net_5252), .A1(net_4715) );
NAND2_X2 inst_11181 ( .A2(net_4132), .ZN(net_4119), .A1(net_4118) );
NAND2_X2 inst_9843 ( .ZN(net_12774), .A2(net_7562), .A1(net_1253) );
NAND2_X4 inst_7492 ( .A1(net_19759), .ZN(net_2923), .A2(net_965) );
INV_X2 inst_18962 ( .A(net_9046), .ZN(net_5418) );
NAND2_X2 inst_11784 ( .A1(net_5169), .ZN(net_3114), .A2(net_1218) );
INV_X4 inst_15729 ( .ZN(net_4261), .A(net_1958) );
AND4_X2 inst_21111 ( .A4(net_9076), .A3(net_9033), .ZN(net_8447), .A1(net_8446), .A2(net_8035) );
INV_X2 inst_19170 ( .ZN(net_3832), .A(net_3831) );
NAND2_X2 inst_10011 ( .A1(net_12175), .ZN(net_8789), .A2(net_8788) );
INV_X4 inst_14231 ( .ZN(net_10847), .A(net_5826) );
AND3_X2 inst_21129 ( .ZN(net_16392), .A1(net_16297), .A2(net_14921), .A3(net_13879) );
INV_X4 inst_16637 ( .A(net_1349), .ZN(net_1105) );
INV_X4 inst_16920 ( .ZN(net_8533), .A(net_4430) );
NAND2_X2 inst_11356 ( .ZN(net_3618), .A1(net_2957), .A2(net_1841) );
AOI21_X2 inst_20289 ( .ZN(net_19822), .B1(net_18996), .A(net_15292), .B2(net_9656) );
NAND2_X2 inst_7780 ( .A1(net_21179), .ZN(net_18728), .A2(net_18721) );
CLKBUF_X2 inst_22401 ( .A(net_22037), .Z(net_22273) );
NOR2_X2 inst_4592 ( .A2(net_5517), .ZN(net_4767), .A1(net_2932) );
CLKBUF_X2 inst_21638 ( .A(net_21509), .Z(net_21510) );
INV_X4 inst_15696 ( .ZN(net_3355), .A(net_2018) );
XNOR2_X2 inst_451 ( .ZN(net_14421), .B(net_14420), .A(net_11889) );
NAND4_X2 inst_5478 ( .ZN(net_12837), .A2(net_12836), .A4(net_12835), .A1(net_11635), .A3(net_9923) );
OAI21_X2 inst_2166 ( .B1(net_11779), .ZN(net_9011), .B2(net_9010), .A(net_7051) );
INV_X2 inst_19536 ( .A(net_2388), .ZN(net_976) );
INV_X4 inst_16145 ( .ZN(net_1468), .A(net_1467) );
INV_X4 inst_14486 ( .ZN(net_6017), .A(net_4852) );
CLKBUF_X2 inst_21911 ( .A(net_21782), .Z(net_21783) );
INV_X4 inst_15377 ( .A(net_6528), .ZN(net_4034) );
NAND2_X2 inst_9910 ( .ZN(net_13561), .A1(net_11186), .A2(net_4822) );
NAND2_X4 inst_7471 ( .A1(net_20741), .ZN(net_20441), .A2(net_2629) );
NAND2_X4 inst_7221 ( .ZN(net_19196), .A2(net_7473), .A1(net_3586) );
INV_X4 inst_18193 ( .A(net_20952), .ZN(net_16359) );
NAND4_X2 inst_5295 ( .ZN(net_15923), .A4(net_15167), .A2(net_14137), .A1(net_13123), .A3(net_13088) );
NOR2_X2 inst_3657 ( .ZN(net_13789), .A2(net_11632), .A1(net_4452) );
NAND2_X4 inst_7319 ( .ZN(net_6154), .A1(net_5136), .A2(net_2744) );
NAND2_X4 inst_6896 ( .ZN(net_18010), .A2(net_17956), .A1(net_17932) );
CLKBUF_X2 inst_21734 ( .A(net_21605), .Z(net_21606) );
INV_X4 inst_14529 ( .ZN(net_8391), .A(net_4740) );
INV_X4 inst_17682 ( .A(net_310), .ZN(net_233) );
AND3_X4 inst_21118 ( .A3(net_13728), .ZN(net_13264), .A2(net_11743), .A1(net_10511) );
OAI21_X2 inst_1998 ( .ZN(net_11857), .B2(net_11856), .A(net_6991), .B1(net_1864) );
INV_X4 inst_17382 ( .ZN(net_1842), .A(net_539) );
NOR2_X4 inst_3302 ( .A2(net_19372), .ZN(net_1878), .A1(net_996) );
NAND2_X2 inst_11157 ( .ZN(net_8508), .A1(net_4194), .A2(net_2864) );
INV_X4 inst_16793 ( .ZN(net_10113), .A(net_9466) );
NOR2_X4 inst_2870 ( .A1(net_13324), .ZN(net_12616), .A2(net_9514) );
INV_X4 inst_14902 ( .ZN(net_11194), .A(net_6512) );
SDFF_X2 inst_874 ( .Q(net_21151), .SI(net_17043), .SE(net_125), .CK(net_21542), .D(x5669) );
CLKBUF_X2 inst_22512 ( .A(net_22383), .Z(net_22384) );
AND4_X4 inst_21087 ( .ZN(net_20187), .A3(net_15844), .A1(net_15603), .A4(net_12169), .A2(net_10107) );
INV_X4 inst_17991 ( .A(net_21166), .ZN(net_16759) );
OAI21_X2 inst_1681 ( .B2(net_19083), .B1(net_19082), .ZN(net_15466), .A(net_333) );
NAND2_X2 inst_10222 ( .ZN(net_14929), .A1(net_11088), .A2(net_8083) );
AOI21_X2 inst_20606 ( .ZN(net_13753), .B1(net_13752), .A(net_13586), .B2(net_6546) );
NAND2_X2 inst_9173 ( .A1(net_13651), .ZN(net_13347), .A2(net_10563) );
OAI21_X2 inst_1652 ( .A(net_16402), .ZN(net_15881), .B2(net_15313), .B1(net_13120) );
NAND2_X2 inst_9391 ( .ZN(net_11714), .A1(net_11713), .A2(net_11712) );
INV_X2 inst_19251 ( .ZN(net_4793), .A(net_3247) );
INV_X4 inst_15576 ( .A(net_7988), .ZN(net_2276) );
OAI21_X2 inst_1622 ( .A(net_16402), .ZN(net_16069), .B1(net_15541), .B2(net_15525) );
INV_X4 inst_13965 ( .ZN(net_7982), .A(net_6710) );
OAI21_X2 inst_1735 ( .ZN(net_20456), .B1(net_13505), .B2(net_10476), .A(net_828) );
OAI21_X2 inst_2050 ( .A(net_11118), .ZN(net_10852), .B2(net_6464), .B1(net_4039) );
NAND2_X2 inst_9516 ( .ZN(net_11145), .A2(net_7426), .A1(net_4142) );
NAND4_X2 inst_5458 ( .ZN(net_13434), .A3(net_10977), .A2(net_9874), .A1(net_8392), .A4(net_7126) );
NOR2_X2 inst_4555 ( .ZN(net_10950), .A2(net_3940), .A1(net_170) );
INV_X4 inst_16366 ( .A(net_1495), .ZN(net_1285) );
NAND2_X2 inst_8681 ( .A2(net_16562), .ZN(net_16452), .A1(net_16451) );
OR2_X2 inst_1189 ( .A2(net_7133), .ZN(net_4475), .A1(net_2244) );
INV_X4 inst_15762 ( .ZN(net_13565), .A(net_1986) );
OAI21_X2 inst_2360 ( .ZN(net_18874), .A(net_14600), .B1(net_11965), .B2(net_7756) );
INV_X4 inst_16847 ( .ZN(net_2855), .A(net_1491) );
CLKBUF_X2 inst_22762 ( .A(net_22633), .Z(net_22634) );
NAND2_X2 inst_11052 ( .ZN(net_11272), .A1(net_4704), .A2(net_2603) );
INV_X4 inst_16460 ( .ZN(net_6981), .A(net_809) );
CLKBUF_X2 inst_22410 ( .A(net_22132), .Z(net_22282) );
INV_X4 inst_16401 ( .ZN(net_14185), .A(net_10512) );
XOR2_X2 inst_33 ( .A(net_21210), .Z(net_717), .B(net_716) );
CLKBUF_X2 inst_21932 ( .A(net_21803), .Z(net_21804) );
OAI21_X2 inst_2107 ( .A(net_13348), .ZN(net_10051), .B2(net_10050), .B1(net_4067) );
INV_X4 inst_12756 ( .ZN(net_18715), .A(net_17406) );
XNOR2_X2 inst_232 ( .B(net_21147), .A(net_19457), .ZN(net_17447) );
INV_X2 inst_19377 ( .ZN(net_2162), .A(net_2161) );
INV_X4 inst_16764 ( .ZN(net_1052), .A(net_1030) );
NAND3_X2 inst_6253 ( .A3(net_19465), .ZN(net_18911), .A1(net_6330), .A2(net_4441) );
NAND2_X4 inst_7575 ( .A2(net_19216), .ZN(net_3122), .A1(net_1312) );
NOR2_X2 inst_4628 ( .A1(net_9478), .ZN(net_5067), .A2(net_2128) );
CLKBUF_X2 inst_21943 ( .A(net_21814), .Z(net_21815) );
INV_X4 inst_16452 ( .ZN(net_3451), .A(net_1363) );
NOR2_X2 inst_3794 ( .ZN(net_10029), .A2(net_6761), .A1(net_5782) );
NAND2_X2 inst_9648 ( .ZN(net_10369), .A1(net_10368), .A2(net_10367) );
INV_X2 inst_18904 ( .ZN(net_20592), .A(net_6058) );
INV_X2 inst_18704 ( .ZN(net_8282), .A(net_8281) );
INV_X4 inst_14463 ( .ZN(net_7881), .A(net_4935) );
INV_X4 inst_16317 ( .ZN(net_2960), .A(net_1320) );
NAND2_X2 inst_9608 ( .ZN(net_10725), .A1(net_8543), .A2(net_8470) );
NAND2_X2 inst_7730 ( .A1(net_20296), .ZN(net_18820), .A2(net_17809) );
INV_X4 inst_13945 ( .A(net_11598), .ZN(net_8631) );
NOR2_X2 inst_3652 ( .ZN(net_11669), .A2(net_11096), .A1(net_8102) );
CLKBUF_X2 inst_21747 ( .A(net_21618), .Z(net_21619) );
INV_X8 inst_12428 ( .A(net_20932), .ZN(net_1848) );
INV_X2 inst_19621 ( .A(net_20975), .ZN(net_37) );
INV_X4 inst_18185 ( .A(net_20968), .ZN(net_16385) );
INV_X4 inst_14513 ( .ZN(net_7854), .A(net_4816) );
NOR2_X2 inst_5043 ( .A2(net_1970), .ZN(net_1088), .A1(net_86) );
INV_X4 inst_17635 ( .A(net_1435), .ZN(net_731) );
INV_X4 inst_18266 ( .A(net_19444), .ZN(net_19441) );
INV_X4 inst_13751 ( .ZN(net_9869), .A(net_7621) );
NAND2_X4 inst_6907 ( .A2(net_18889), .A1(net_18888), .ZN(net_17914) );
NAND2_X2 inst_9331 ( .ZN(net_14215), .A1(net_10819), .A2(net_9141) );
XNOR2_X2 inst_602 ( .B(net_16842), .ZN(net_16097), .A(net_631) );
INV_X2 inst_18945 ( .ZN(net_5680), .A(net_5679) );
XNOR2_X2 inst_135 ( .B(net_21220), .ZN(net_18290), .A(net_18166) );
NAND2_X2 inst_10091 ( .ZN(net_13278), .A1(net_11468), .A2(net_8622) );
NAND2_X2 inst_11711 ( .ZN(net_2982), .A2(net_2278), .A1(net_1547) );
NAND2_X4 inst_7673 ( .ZN(net_1225), .A1(net_879), .A2(net_841) );
INV_X4 inst_17705 ( .ZN(net_846), .A(net_214) );
DFF_X1 inst_19858 ( .D(net_17263), .CK(net_22368), .Q(x687) );
AND3_X2 inst_21151 ( .A2(net_8097), .ZN(net_3352), .A3(net_3351), .A1(net_2779) );
NAND2_X2 inst_10037 ( .ZN(net_10166), .A1(net_8722), .A2(net_6822) );
INV_X4 inst_18241 ( .A(net_21238), .ZN(net_2673) );
NAND2_X2 inst_9321 ( .ZN(net_12331), .A1(net_12330), .A2(net_9068) );
NOR2_X4 inst_3117 ( .ZN(net_5005), .A1(net_3984), .A2(net_1905) );
INV_X4 inst_16763 ( .ZN(net_6089), .A(net_154) );
NAND3_X2 inst_6072 ( .ZN(net_20307), .A3(net_19350), .A1(net_19349), .A2(net_5699) );
NOR2_X2 inst_3770 ( .A2(net_11627), .ZN(net_11620), .A1(net_10290) );
NAND2_X2 inst_8157 ( .ZN(net_17992), .A1(net_17941), .A2(net_17892) );
INV_X4 inst_13863 ( .ZN(net_9126), .A(net_7458) );
INV_X4 inst_16260 ( .ZN(net_1643), .A(net_1353) );
NOR3_X2 inst_2709 ( .ZN(net_13719), .A1(net_13718), .A3(net_12707), .A2(net_5027) );
XNOR2_X2 inst_224 ( .ZN(net_17505), .A(net_17089), .B(net_501) );
INV_X4 inst_14756 ( .A(net_9282), .ZN(net_7740) );
INV_X4 inst_14003 ( .A(net_8587), .ZN(net_6356) );
NAND2_X2 inst_9661 ( .ZN(net_19542), .A2(net_12038), .A1(net_11874) );
NOR2_X2 inst_3635 ( .ZN(net_12188), .A1(net_10276), .A2(net_8729) );
INV_X4 inst_16481 ( .ZN(net_9450), .A(net_7153) );
NAND4_X2 inst_5399 ( .A3(net_15413), .ZN(net_14781), .A1(net_14619), .A2(net_13387), .A4(net_10272) );
NOR2_X2 inst_5058 ( .ZN(net_1008), .A1(net_987), .A2(net_380) );
DFF_X2 inst_19768 ( .QN(net_20860), .D(net_18861), .CK(net_22054) );
INV_X4 inst_14297 ( .A(net_9055), .ZN(net_6858) );
OAI211_X2 inst_2406 ( .ZN(net_15728), .B(net_15074), .A(net_14711), .C1(net_13873), .C2(net_12871) );
NAND2_X2 inst_8796 ( .ZN(net_19310), .A2(net_15212), .A1(net_13867) );
INV_X4 inst_17994 ( .A(net_21178), .ZN(net_643) );
SDFF_X2 inst_801 ( .Q(net_20850), .SE(net_18847), .SI(net_17965), .D(net_720), .CK(net_21267) );
NAND2_X2 inst_10617 ( .ZN(net_13107), .A1(net_6587), .A2(net_6561) );
INV_X4 inst_16873 ( .A(net_1330), .ZN(net_1048) );
SDFF_X2 inst_870 ( .Q(net_21207), .SI(net_17088), .SE(net_125), .CK(net_22437), .D(x5903) );
INV_X4 inst_12544 ( .ZN(net_18399), .A(net_18337) );
NAND2_X2 inst_9660 ( .ZN(net_13103), .A1(net_13026), .A2(net_8340) );
XOR2_X2 inst_11 ( .A(net_21126), .Z(net_17067), .B(net_17066) );
INV_X4 inst_15537 ( .A(net_7968), .ZN(net_3251) );
INV_X4 inst_13468 ( .A(net_10343), .ZN(net_9670) );
AOI21_X2 inst_20568 ( .ZN(net_14167), .A(net_14166), .B1(net_12215), .B2(net_10727) );
NAND2_X4 inst_7688 ( .ZN(net_705), .A1(net_264), .A2(net_234) );
OAI21_X2 inst_2276 ( .A(net_8543), .ZN(net_7132), .B1(net_5574), .B2(net_3015) );
NAND2_X2 inst_8892 ( .ZN(net_15114), .A1(net_15113), .A2(net_13961) );
AOI21_X2 inst_20843 ( .ZN(net_9264), .A(net_9263), .B2(net_4595), .B1(net_2157) );
OAI21_X2 inst_2301 ( .ZN(net_20177), .A(net_8682), .B2(net_5644), .B1(net_2850) );
INV_X2 inst_18404 ( .A(net_16774), .ZN(net_16412) );
NAND2_X2 inst_8202 ( .ZN(net_17938), .A2(net_17749), .A1(net_17654) );
XNOR2_X2 inst_557 ( .B(net_17534), .A(net_17426), .ZN(net_6372) );
INV_X4 inst_13639 ( .A(net_13728), .ZN(net_12069) );
INV_X4 inst_14300 ( .ZN(net_5732), .A(net_5536) );
NAND2_X2 inst_11154 ( .ZN(net_4197), .A2(net_2717), .A1(net_1683) );
NOR2_X4 inst_3279 ( .A1(net_19222), .ZN(net_2668), .A2(net_318) );
SDFF_X2 inst_823 ( .Q(net_21143), .SI(net_17609), .SE(net_125), .CK(net_21668), .D(x3521) );
OAI21_X4 inst_1461 ( .ZN(net_15244), .B2(net_14119), .B1(net_10366), .A(net_2528) );
NAND2_X2 inst_8809 ( .ZN(net_15619), .A2(net_14885), .A1(net_10683) );
NOR2_X2 inst_3773 ( .A2(net_10720), .ZN(net_10257), .A1(net_8622) );
CLKBUF_X2 inst_21444 ( .A(net_21315), .Z(net_21316) );
NOR2_X2 inst_4767 ( .ZN(net_4429), .A2(net_3019), .A1(net_2976) );
NAND2_X2 inst_10608 ( .A2(net_20782), .ZN(net_13054), .A1(net_6861) );
INV_X2 inst_19014 ( .ZN(net_5000), .A(net_4999) );
INV_X4 inst_13154 ( .ZN(net_20000), .A(net_14335) );
INV_X2 inst_19230 ( .A(net_3686), .ZN(net_3377) );
NAND3_X4 inst_5620 ( .ZN(net_11467), .A1(net_11466), .A2(net_11465), .A3(net_11464) );
NAND2_X2 inst_11409 ( .ZN(net_7714), .A2(net_2051), .A1(net_90) );
NAND2_X4 inst_7104 ( .ZN(net_13560), .A1(net_10705), .A2(net_9917) );
NAND2_X2 inst_7746 ( .ZN(net_18784), .A1(net_18783), .A2(net_18782) );
NAND2_X2 inst_9976 ( .ZN(net_8875), .A1(net_8874), .A2(net_6515) );
NAND2_X2 inst_8342 ( .A1(net_17763), .ZN(net_17489), .A2(net_17488) );
AOI21_X2 inst_20682 ( .ZN(net_12300), .B2(net_10757), .B1(net_6316), .A(net_2248) );
INV_X4 inst_18121 ( .A(net_20882), .ZN(net_761) );
INV_X4 inst_14084 ( .ZN(net_11357), .A(net_6215) );
INV_X4 inst_16544 ( .ZN(net_11062), .A(net_7298) );
OAI21_X4 inst_1413 ( .A(net_20888), .B2(net_19579), .B1(net_19578), .ZN(net_16172) );
CLKBUF_X2 inst_22502 ( .A(net_22373), .Z(net_22374) );
INV_X4 inst_13320 ( .ZN(net_11521), .A(net_11520) );
NOR2_X2 inst_3993 ( .ZN(net_8272), .A1(net_8221), .A2(net_4570) );
NAND2_X4 inst_6926 ( .A2(net_19018), .A1(net_19017), .ZN(net_17742) );
NAND2_X2 inst_11140 ( .A1(net_8179), .ZN(net_4245), .A2(net_4244) );
CLKBUF_X2 inst_22577 ( .A(net_21898), .Z(net_22449) );
AOI22_X2 inst_20024 ( .ZN(net_10511), .B1(net_10134), .A1(net_8533), .A2(net_6519), .B2(net_5956) );
INV_X4 inst_17615 ( .ZN(net_6599), .A(net_3745) );
INV_X4 inst_13272 ( .ZN(net_12499), .A(net_11265) );
INV_X4 inst_16161 ( .ZN(net_15356), .A(net_1449) );
OAI21_X2 inst_2169 ( .A(net_9972), .ZN(net_8929), .B2(net_6146), .B1(net_1180) );
AOI21_X2 inst_20625 ( .B1(net_13709), .ZN(net_13447), .B2(net_8946), .A(net_8212) );
NAND2_X2 inst_11903 ( .ZN(net_2056), .A1(net_1568), .A2(net_1567) );
INV_X4 inst_15258 ( .ZN(net_3693), .A(net_2782) );
OAI221_X4 inst_1326 ( .C1(net_21228), .ZN(net_16479), .B1(net_16281), .A(net_16264), .B2(net_15813), .C2(net_15722) );
INV_X4 inst_18065 ( .A(net_20953), .ZN(net_1470) );
NAND2_X2 inst_8960 ( .ZN(net_14708), .A2(net_13283), .A1(net_4154) );
INV_X4 inst_16473 ( .ZN(net_1962), .A(net_1786) );
INV_X4 inst_14938 ( .ZN(net_3536), .A(net_3535) );
NAND2_X2 inst_8191 ( .ZN(net_19300), .A2(net_17785), .A1(net_17269) );
NAND2_X2 inst_11920 ( .A2(net_1583), .ZN(net_1540), .A1(net_703) );
NOR2_X2 inst_4238 ( .A1(net_7193), .ZN(net_6567), .A2(net_4730) );
NAND2_X2 inst_9496 ( .A1(net_14743), .ZN(net_12593), .A2(net_11478) );
NAND4_X2 inst_5275 ( .A4(net_20306), .A1(net_20305), .ZN(net_19504), .A2(net_15502), .A3(net_14704) );
INV_X4 inst_18029 ( .A(net_21013), .ZN(net_799) );
INV_X2 inst_18800 ( .ZN(net_7419), .A(net_7418) );
INV_X4 inst_14791 ( .ZN(net_4008), .A(net_4007) );
INV_X2 inst_19237 ( .ZN(net_3325), .A(net_3324) );
INV_X4 inst_14887 ( .A(net_3665), .ZN(net_3664) );
INV_X4 inst_16374 ( .ZN(net_10962), .A(net_703) );
NAND2_X2 inst_9197 ( .ZN(net_13090), .A1(net_13089), .A2(net_11362) );
NAND3_X2 inst_6127 ( .ZN(net_13743), .A3(net_13742), .A1(net_12040), .A2(net_3103) );
INV_X4 inst_14867 ( .ZN(net_4700), .A(net_3754) );
OAI21_X2 inst_2154 ( .A(net_13213), .ZN(net_9279), .B2(net_9278), .B1(net_3239) );
CLKBUF_X2 inst_22218 ( .A(net_22089), .Z(net_22090) );
INV_X4 inst_16487 ( .A(net_9254), .ZN(net_5712) );
NOR2_X2 inst_4602 ( .ZN(net_5011), .A1(net_3760), .A2(net_1544) );
NOR3_X4 inst_2602 ( .ZN(net_18612), .A1(net_18603), .A3(net_15805), .A2(net_15271) );
XNOR2_X2 inst_109 ( .ZN(net_18518), .A(net_18401), .B(net_17761) );
OR2_X2 inst_1182 ( .ZN(net_7829), .A1(net_4750), .A2(net_4749) );
NAND2_X4 inst_6875 ( .ZN(net_18310), .A2(net_18151), .A1(net_18127) );
NOR2_X2 inst_3983 ( .ZN(net_8350), .A2(net_8081), .A1(net_3518) );
INV_X4 inst_15066 ( .ZN(net_4672), .A(net_3295) );
INV_X4 inst_17311 ( .ZN(net_15300), .A(net_15108) );
INV_X8 inst_12275 ( .ZN(net_2745), .A(net_1191) );
NAND2_X2 inst_11019 ( .ZN(net_6978), .A2(net_6953), .A1(net_3750) );
AOI211_X2 inst_21050 ( .ZN(net_12421), .C2(net_8450), .A(net_4832), .B(net_4761), .C1(net_1864) );
NAND3_X2 inst_5984 ( .ZN(net_14543), .A2(net_14542), .A1(net_13341), .A3(net_12970) );
OAI21_X4 inst_1444 ( .B2(net_20725), .B1(net_20724), .ZN(net_18876), .A(net_1868) );
NAND2_X2 inst_11993 ( .A1(net_1645), .ZN(net_1210), .A2(net_369) );
NAND4_X2 inst_5490 ( .ZN(net_12250), .A4(net_12249), .A3(net_9915), .A1(net_7956), .A2(net_7266) );
CLKBUF_X2 inst_22187 ( .A(net_22058), .Z(net_22059) );
INV_X4 inst_17226 ( .ZN(net_1114), .A(net_173) );
OR2_X2 inst_1231 ( .ZN(net_6439), .A2(net_2240), .A1(net_222) );
AOI21_X2 inst_20419 ( .A(net_15366), .ZN(net_15250), .B2(net_14120), .B1(net_4748) );
CLKBUF_X2 inst_21771 ( .A(net_21642), .Z(net_21643) );
INV_X2 inst_19680 ( .A(net_20515), .ZN(net_20514) );
INV_X4 inst_15557 ( .ZN(net_2323), .A(net_2111) );
SDFF_X2 inst_904 ( .Q(net_21168), .D(net_16851), .SE(net_263), .CK(net_22426), .SI(x4980) );
AOI221_X4 inst_20073 ( .B2(net_19715), .B1(net_19714), .ZN(net_18916), .C2(net_15563), .A(net_13923), .C1(net_7318) );
CLKBUF_X2 inst_21546 ( .A(net_21417), .Z(net_21418) );
NAND2_X2 inst_12100 ( .A2(net_20875), .ZN(net_1998), .A1(net_493) );
NAND2_X2 inst_10628 ( .A1(net_13534), .ZN(net_6554), .A2(net_6553) );
INV_X4 inst_13147 ( .ZN(net_19513), .A(net_14532) );
OAI21_X2 inst_2159 ( .B2(net_9698), .ZN(net_9249), .A(net_3345), .B1(net_2345) );
INV_X4 inst_18012 ( .A(net_21086), .ZN(net_681) );
NAND2_X4 inst_7051 ( .A2(net_19899), .A1(net_19898), .ZN(net_19449) );
NAND3_X2 inst_6266 ( .ZN(net_12969), .A2(net_12968), .A3(net_11644), .A1(net_6826) );
NOR2_X2 inst_3923 ( .A1(net_11186), .ZN(net_8781), .A2(net_8780) );
INV_X4 inst_16042 ( .ZN(net_1612), .A(net_1611) );
NOR2_X2 inst_4831 ( .ZN(net_2414), .A2(net_1886), .A1(net_1185) );
SDFF_X2 inst_757 ( .Q(net_20872), .SE(net_18837), .SI(net_18527), .D(net_451), .CK(net_21861) );
CLKBUF_X2 inst_22899 ( .A(net_21804), .Z(net_22771) );
OAI21_X2 inst_1627 ( .ZN(net_20448), .B2(net_15444), .A(net_15104), .B1(net_14081) );
INV_X2 inst_18629 ( .ZN(net_9481), .A(net_9480) );
INV_X4 inst_12670 ( .ZN(net_17783), .A(net_17782) );
INV_X4 inst_17857 ( .ZN(net_311), .A(net_109) );
CLKBUF_X2 inst_22010 ( .A(net_21425), .Z(net_21882) );
INV_X4 inst_13557 ( .A(net_10873), .ZN(net_10726) );
INV_X4 inst_12994 ( .ZN(net_16792), .A(net_16643) );
NOR2_X2 inst_3817 ( .A2(net_11388), .ZN(net_9802), .A1(net_9801) );
INV_X4 inst_15201 ( .A(net_4677), .ZN(net_2912) );
INV_X4 inst_15458 ( .ZN(net_2717), .A(net_2481) );
NOR2_X2 inst_5065 ( .ZN(net_963), .A1(net_930), .A2(net_106) );
OAI22_X2 inst_1256 ( .ZN(net_17634), .B1(net_17633), .A2(net_17576), .B2(net_17299), .A1(net_17204) );
INV_X4 inst_17204 ( .ZN(net_2456), .A(net_1645) );
INV_X4 inst_15710 ( .ZN(net_12504), .A(net_1986) );
CLKBUF_X2 inst_21898 ( .A(net_21769), .Z(net_21770) );
AND3_X2 inst_21149 ( .A3(net_13512), .A1(net_7033), .ZN(net_5321), .A2(net_588) );
NAND2_X2 inst_9549 ( .ZN(net_11031), .A2(net_10919), .A1(net_652) );
INV_X4 inst_15752 ( .ZN(net_4508), .A(net_3703) );
AND2_X2 inst_21334 ( .ZN(net_4346), .A1(net_4345), .A2(net_2982) );
OAI21_X2 inst_1903 ( .B1(net_20150), .ZN(net_13269), .A(net_10260), .B2(net_7450) );
INV_X4 inst_14254 ( .ZN(net_13194), .A(net_5755) );
INV_X2 inst_19550 ( .A(net_3002), .ZN(net_905) );
NAND2_X2 inst_9503 ( .ZN(net_11341), .A2(net_11340), .A1(net_8269) );
NAND2_X2 inst_11230 ( .ZN(net_3950), .A2(net_3949), .A1(net_1790) );
INV_X4 inst_13716 ( .ZN(net_14442), .A(net_7827) );
OAI211_X2 inst_2554 ( .A(net_12063), .ZN(net_10476), .B(net_10475), .C1(net_7394), .C2(net_4560) );
INV_X4 inst_16993 ( .ZN(net_3617), .A(net_1798) );
NAND2_X2 inst_9423 ( .A2(net_11632), .ZN(net_11630), .A1(net_11629) );
INV_X4 inst_14422 ( .A(net_5051), .ZN(net_5050) );
INV_X4 inst_15295 ( .ZN(net_3788), .A(net_2461) );
NOR3_X4 inst_2604 ( .ZN(net_19846), .A1(net_16028), .A3(net_15905), .A2(net_15395) );
INV_X2 inst_18684 ( .ZN(net_14747), .A(net_7254) );
INV_X4 inst_16159 ( .ZN(net_3906), .A(net_1452) );
AND4_X2 inst_21101 ( .A1(net_14314), .A3(net_13621), .ZN(net_12750), .A2(net_11801), .A4(net_11800) );
INV_X4 inst_17776 ( .ZN(net_801), .A(net_550) );
INV_X4 inst_15019 ( .A(net_8981), .ZN(net_5166) );
NOR2_X4 inst_3248 ( .ZN(net_4303), .A1(net_2246), .A2(net_1578) );
CLKBUF_X2 inst_21952 ( .A(net_21308), .Z(net_21824) );
AOI211_X2 inst_21073 ( .B(net_8559), .ZN(net_7683), .C2(net_4610), .C1(net_3389), .A(net_3321) );
AOI21_X2 inst_20549 ( .ZN(net_19261), .B1(net_14367), .B2(net_12476), .A(net_9687) );
INV_X4 inst_16961 ( .ZN(net_902), .A(net_449) );
INV_X4 inst_18303 ( .A(net_20487), .ZN(net_20486) );
INV_X8 inst_12329 ( .A(net_1697), .ZN(net_950) );
OAI21_X2 inst_2110 ( .A(net_10864), .ZN(net_10044), .B2(net_5320), .B1(net_2412) );
INV_X4 inst_16702 ( .ZN(net_3991), .A(net_1395) );
NAND2_X2 inst_9774 ( .A1(net_14075), .ZN(net_9792), .A2(net_9791) );
INV_X4 inst_13896 ( .ZN(net_9169), .A(net_7202) );
NAND2_X4 inst_7463 ( .ZN(net_5652), .A2(net_2430), .A1(net_2094) );
CLKBUF_X2 inst_21817 ( .A(net_21334), .Z(net_21689) );
INV_X4 inst_15051 ( .A(net_3321), .ZN(net_3319) );
INV_X2 inst_18492 ( .A(net_13676), .ZN(net_12333) );
INV_X4 inst_12914 ( .ZN(net_17025), .A(net_16670) );
OAI21_X2 inst_2057 ( .ZN(net_10704), .B2(net_6904), .B1(net_5513), .A(net_630) );
CLKBUF_X2 inst_22131 ( .A(net_21842), .Z(net_22003) );
INV_X4 inst_15217 ( .ZN(net_4371), .A(net_2882) );
INV_X4 inst_13408 ( .ZN(net_13132), .A(net_10350) );
SDFF_X2 inst_843 ( .Q(net_21149), .SI(net_17317), .SE(net_125), .CK(net_22313), .D(x5723) );
NAND2_X2 inst_10710 ( .ZN(net_9467), .A2(net_5933), .A1(net_1186) );
INV_X2 inst_19290 ( .ZN(net_2871), .A(net_2870) );
NOR2_X1 inst_5146 ( .ZN(net_17688), .A1(net_17651), .A2(net_17644) );
CLKBUF_X2 inst_21512 ( .A(net_21383), .Z(net_21384) );
INV_X4 inst_14974 ( .A(net_9989), .ZN(net_4477) );
SDFF_X2 inst_916 ( .Q(net_21212), .D(net_16651), .SE(net_263), .CK(net_22204), .SI(x7607) );
OAI21_X2 inst_1722 ( .ZN(net_15097), .B2(net_12973), .B1(net_9790), .A(net_3383) );
NAND3_X4 inst_5570 ( .A2(net_19024), .A1(net_19023), .ZN(net_15873), .A3(net_15103) );
INV_X4 inst_13799 ( .ZN(net_11086), .A(net_7558) );
AOI21_X2 inst_20921 ( .ZN(net_7217), .B1(net_7025), .B2(net_3855), .A(net_1000) );
NAND2_X2 inst_8754 ( .A1(net_16259), .ZN(net_15913), .A2(net_15496) );
NAND2_X4 inst_7300 ( .ZN(net_9061), .A2(net_5551), .A1(net_5550) );
NAND3_X2 inst_6409 ( .A1(net_13147), .ZN(net_11960), .A3(net_11959), .A2(net_5968) );
NOR2_X2 inst_3665 ( .A1(net_13734), .ZN(net_11559), .A2(net_11558) );
INV_X4 inst_17433 ( .ZN(net_1574), .A(net_809) );
AOI21_X2 inst_20503 ( .ZN(net_14646), .B1(net_12658), .B2(net_12089), .A(net_5266) );
INV_X4 inst_16680 ( .ZN(net_7427), .A(net_1634) );
INV_X4 inst_16111 ( .ZN(net_2581), .A(net_2241) );
OAI211_X2 inst_2525 ( .ZN(net_11787), .C1(net_11786), .A(net_11721), .B(net_10267), .C2(net_9626) );
NOR2_X4 inst_2968 ( .ZN(net_7690), .A1(net_4567), .A2(net_874) );
INV_X4 inst_12875 ( .A(net_16946), .ZN(net_16945) );
NAND2_X2 inst_7916 ( .ZN(net_18457), .A1(net_18399), .A2(net_18343) );
NOR2_X4 inst_2964 ( .ZN(net_7859), .A1(net_6606), .A2(net_4842) );
NAND2_X2 inst_11760 ( .A1(net_5173), .ZN(net_2092), .A2(net_1152) );
NOR2_X2 inst_3721 ( .ZN(net_10969), .A1(net_10968), .A2(net_10409) );
OAI21_X2 inst_2349 ( .ZN(net_3724), .B1(net_2998), .B2(net_2305), .A(net_373) );
NAND2_X2 inst_8855 ( .ZN(net_15363), .A1(net_15362), .A2(net_14369) );
XNOR2_X2 inst_646 ( .B(net_17113), .ZN(net_390), .A(net_389) );
NOR2_X2 inst_5076 ( .ZN(net_10175), .A2(net_1231), .A1(net_30) );
NAND3_X2 inst_6667 ( .A2(net_10114), .ZN(net_8290), .A3(net_6182), .A1(net_761) );
NOR2_X2 inst_4032 ( .ZN(net_7970), .A2(net_6213), .A1(net_4054) );
INV_X4 inst_14310 ( .A(net_8976), .ZN(net_6805) );
NOR2_X4 inst_3169 ( .ZN(net_7168), .A2(net_5595), .A1(net_3784) );
INV_X4 inst_13278 ( .ZN(net_12450), .A(net_11173) );
NAND2_X2 inst_9841 ( .ZN(net_9551), .A1(net_9550), .A2(net_6163) );
NAND4_X2 inst_5344 ( .ZN(net_15441), .A2(net_14498), .A3(net_14301), .A1(net_12654), .A4(net_10331) );
NAND2_X2 inst_11119 ( .ZN(net_10575), .A2(net_4303), .A1(net_409) );
INV_X4 inst_14248 ( .A(net_10709), .ZN(net_9764) );
NAND2_X2 inst_9799 ( .ZN(net_11070), .A2(net_9776), .A1(net_8707) );
NOR3_X2 inst_2788 ( .ZN(net_5369), .A1(net_2502), .A3(net_1908), .A2(net_1037) );
NAND3_X2 inst_6015 ( .ZN(net_14404), .A3(net_14330), .A1(net_11332), .A2(net_9756) );
NAND2_X2 inst_11891 ( .ZN(net_19258), .A1(net_3293), .A2(net_1595) );
INV_X2 inst_19191 ( .ZN(net_3663), .A(net_3662) );
NAND3_X2 inst_6565 ( .A2(net_11168), .ZN(net_10481), .A3(net_10480), .A1(net_4777) );
NAND2_X2 inst_10415 ( .ZN(net_12226), .A1(net_7244), .A2(net_6795) );
NAND2_X2 inst_10194 ( .A1(net_10550), .ZN(net_10280), .A2(net_8006) );
XNOR2_X2 inst_168 ( .ZN(net_17828), .A(net_17827), .B(net_10801) );
CLKBUF_X2 inst_22253 ( .A(net_22124), .Z(net_22125) );
NAND2_X2 inst_9139 ( .ZN(net_13438), .A1(net_13437), .A2(net_13399) );
INV_X4 inst_16173 ( .ZN(net_5635), .A(net_2627) );
CLKBUF_X2 inst_22614 ( .A(net_22241), .Z(net_22486) );
DFF_X1 inst_19917 ( .D(net_16620), .CK(net_21573), .Q(x622) );
NAND2_X2 inst_8688 ( .ZN(net_16417), .A1(net_16393), .A2(net_16339) );
SDFF_X2 inst_991 ( .QN(net_21050), .D(net_413), .SE(net_263), .CK(net_22502), .SI(x2186) );
NAND2_X2 inst_10642 ( .A1(net_13848), .ZN(net_6370), .A2(net_6369) );
XNOR2_X2 inst_170 ( .A(net_17827), .ZN(net_17825), .B(net_10802) );
NAND2_X2 inst_9160 ( .ZN(net_13381), .A2(net_10603), .A1(net_6934) );
DFF_X1 inst_19836 ( .D(net_17523), .CK(net_21360), .Q(x311) );
NOR2_X2 inst_3691 ( .ZN(net_11325), .A1(net_11324), .A2(net_8142) );
INV_X4 inst_17371 ( .A(net_3780), .ZN(net_3108) );
INV_X4 inst_13159 ( .ZN(net_14841), .A(net_14257) );
DFF_X1 inst_19803 ( .D(net_18181), .CK(net_22823), .Q(x1121) );
NAND2_X2 inst_7823 ( .A2(net_18648), .ZN(net_18647), .A1(net_17010) );
OAI21_X2 inst_1857 ( .ZN(net_13942), .A(net_13941), .B1(net_13940), .B2(net_11193) );
NAND2_X2 inst_11536 ( .ZN(net_20717), .A1(net_6867), .A2(net_2925) );
XNOR2_X2 inst_468 ( .B(net_16267), .ZN(net_13298), .A(net_7353) );
OR2_X4 inst_1099 ( .A1(net_20543), .ZN(net_5348), .A2(net_3241) );
INV_X2 inst_19064 ( .ZN(net_4648), .A(net_4647) );
NAND3_X2 inst_6611 ( .A3(net_12126), .A2(net_12025), .ZN(net_9079), .A1(net_7781) );
INV_X4 inst_17973 ( .A(net_20997), .ZN(net_1883) );
NOR2_X2 inst_4428 ( .A2(net_20803), .ZN(net_6062), .A1(net_624) );
CLKBUF_X2 inst_21876 ( .A(net_21747), .Z(net_21748) );
INV_X4 inst_16805 ( .ZN(net_2400), .A(net_1004) );
INV_X4 inst_14762 ( .ZN(net_9921), .A(net_4058) );
NOR2_X2 inst_4889 ( .ZN(net_2100), .A2(net_2099), .A1(net_1999) );
OAI21_X2 inst_2190 ( .ZN(net_8719), .B1(net_7068), .B2(net_4806), .A(net_816) );
XNOR2_X2 inst_429 ( .B(net_21115), .ZN(net_16952), .A(net_16479) );
NAND2_X2 inst_10298 ( .ZN(net_9434), .A2(net_5102), .A1(net_1916) );
INV_X4 inst_18343 ( .A(net_20768), .ZN(net_20767) );
INV_X4 inst_17255 ( .ZN(net_7487), .A(net_1231) );
NAND2_X2 inst_7808 ( .ZN(net_18685), .A1(net_18684), .A2(net_18678) );
INV_X2 inst_18774 ( .ZN(net_7556), .A(net_7555) );
NAND3_X2 inst_5995 ( .ZN(net_14443), .A1(net_14442), .A3(net_14441), .A2(net_14262) );
INV_X4 inst_13824 ( .ZN(net_11004), .A(net_9633) );
INV_X4 inst_13567 ( .A(net_14214), .ZN(net_9136) );
INV_X4 inst_18079 ( .A(net_20987), .ZN(net_2313) );
NOR2_X2 inst_3467 ( .ZN(net_14599), .A2(net_13256), .A1(net_7213) );
INV_X2 inst_19717 ( .A(net_20773), .ZN(net_20772) );
NOR2_X4 inst_3064 ( .ZN(net_8081), .A1(net_4268), .A2(net_3131) );
NOR2_X2 inst_3676 ( .ZN(net_15278), .A2(net_11555), .A1(net_11441) );
CLKBUF_X2 inst_21506 ( .A(net_21377), .Z(net_21378) );
AOI21_X2 inst_20278 ( .B2(net_19291), .B1(net_19290), .A(net_16390), .ZN(net_16315) );
INV_X4 inst_15480 ( .ZN(net_12401), .A(net_2903) );
NAND2_X2 inst_7948 ( .ZN(net_18404), .A2(net_18279), .A1(net_18238) );
NOR2_X2 inst_4033 ( .ZN(net_7967), .A1(net_6253), .A2(net_4589) );
INV_X2 inst_18807 ( .ZN(net_7376), .A(net_7134) );
INV_X2 inst_18528 ( .ZN(net_11100), .A(net_11099) );
INV_X4 inst_14210 ( .ZN(net_13226), .A(net_5917) );
NAND2_X2 inst_8538 ( .ZN(net_16998), .A2(net_16518), .A1(net_16432) );
NOR2_X2 inst_5044 ( .A2(net_2671), .ZN(net_1087), .A1(net_1086) );
NOR2_X4 inst_2899 ( .ZN(net_10871), .A1(net_9322), .A2(net_9321) );
AOI222_X1 inst_20067 ( .ZN(net_15961), .B2(net_15950), .B1(net_15524), .A1(net_15312), .A2(net_14922), .C1(net_12609), .C2(net_8322) );
INV_X4 inst_15510 ( .ZN(net_7097), .A(net_4820) );
CLKBUF_X2 inst_22546 ( .A(net_21263), .Z(net_22418) );
INV_X4 inst_14222 ( .ZN(net_7559), .A(net_6198) );
NOR2_X2 inst_4096 ( .ZN(net_20049), .A2(net_7235), .A1(net_5475) );
CLKBUF_X2 inst_22137 ( .A(net_22008), .Z(net_22009) );
NAND2_X2 inst_10927 ( .A1(net_9571), .ZN(net_6344), .A2(net_5215) );
NAND3_X2 inst_6808 ( .ZN(net_3809), .A3(net_2950), .A2(net_874), .A1(net_120) );
INV_X4 inst_15323 ( .ZN(net_15889), .A(net_15818) );
INV_X4 inst_12508 ( .A(net_18608), .ZN(net_18607) );
XNOR2_X1 inst_689 ( .A(net_16848), .ZN(net_16837), .B(net_16836) );
NOR2_X2 inst_4453 ( .ZN(net_6193), .A2(net_5445), .A1(net_874) );
NOR3_X2 inst_2689 ( .ZN(net_14353), .A2(net_13568), .A3(net_10329), .A1(net_7190) );
INV_X2 inst_19306 ( .A(net_3756), .ZN(net_2729) );
DFF_X1 inst_19863 ( .D(net_17098), .CK(net_22364), .Q(x839) );
INV_X4 inst_16306 ( .ZN(net_1728), .A(net_1644) );
INV_X4 inst_16123 ( .ZN(net_12100), .A(net_1124) );
NAND2_X2 inst_9622 ( .ZN(net_10671), .A2(net_8545), .A1(net_4343) );
INV_X4 inst_12630 ( .ZN(net_17967), .A(net_17938) );
INV_X2 inst_18499 ( .ZN(net_12272), .A(net_10811) );
NAND3_X2 inst_6272 ( .ZN(net_12946), .A2(net_12945), .A3(net_12944), .A1(net_4513) );
INV_X4 inst_17532 ( .ZN(net_1491), .A(net_391) );
INV_X4 inst_13587 ( .A(net_10732), .ZN(net_8910) );
NAND2_X2 inst_8685 ( .ZN(net_16434), .A1(net_16385), .A2(net_16370) );
OAI21_X2 inst_1615 ( .A(net_20872), .B2(net_20312), .B1(net_20311), .ZN(net_16088) );
INV_X4 inst_16718 ( .A(net_7886), .ZN(net_1903) );
NAND2_X2 inst_9148 ( .ZN(net_13403), .A1(net_10875), .A2(net_10650) );
NAND2_X2 inst_11434 ( .ZN(net_6432), .A1(net_3332), .A2(net_3331) );
NAND2_X4 inst_7503 ( .ZN(net_2281), .A2(net_2168), .A1(net_1711) );
INV_X8 inst_12406 ( .ZN(net_179), .A(net_132) );
INV_X4 inst_13760 ( .A(net_9642), .ZN(net_9220) );
NAND2_X2 inst_8313 ( .A2(net_20507), .ZN(net_17582), .A1(net_17335) );
OAI21_X2 inst_2145 ( .ZN(net_20171), .B2(net_13673), .B1(net_11562), .A(net_6602) );
CLKBUF_X2 inst_21949 ( .A(net_21271), .Z(net_21821) );
INV_X4 inst_17890 ( .ZN(net_69), .A(net_68) );
SDFF_X2 inst_709 ( .Q(net_20926), .SE(net_18856), .SI(net_18815), .D(net_510), .CK(net_22030) );
OAI211_X4 inst_2375 ( .C2(net_19267), .C1(net_19266), .ZN(net_16228), .A(net_15314), .B(net_15255) );
NAND3_X2 inst_5725 ( .ZN(net_16124), .A3(net_15715), .A2(net_15351), .A1(net_10961) );
INV_X2 inst_18431 ( .ZN(net_14806), .A(net_14213) );
INV_X4 inst_13400 ( .ZN(net_19778), .A(net_8986) );
NAND2_X2 inst_12080 ( .A1(net_949), .A2(net_937), .ZN(net_778) );
NAND2_X2 inst_9956 ( .ZN(net_8920), .A1(net_8919), .A2(net_7309) );
INV_X2 inst_19434 ( .A(net_2118), .ZN(net_1742) );
INV_X4 inst_12517 ( .A(net_20936), .ZN(net_18601) );
INV_X8 inst_12331 ( .A(net_928), .ZN(net_821) );
NAND2_X2 inst_12106 ( .A2(net_21219), .ZN(net_397), .A1(net_396) );
NAND2_X4 inst_7389 ( .ZN(net_4978), .A1(net_2285), .A2(net_955) );
NOR2_X2 inst_4610 ( .ZN(net_4696), .A1(net_3729), .A2(net_2804) );
INV_X4 inst_13350 ( .ZN(net_12674), .A(net_11707) );
NOR2_X2 inst_4403 ( .ZN(net_19252), .A1(net_5129), .A2(net_4075) );
INV_X2 inst_19076 ( .ZN(net_4601), .A(net_4600) );
CLKBUF_X2 inst_22820 ( .A(net_22691), .Z(net_22692) );
CLKBUF_X2 inst_21643 ( .A(net_21514), .Z(net_21515) );
INV_X4 inst_14589 ( .ZN(net_4471), .A(net_4470) );
NAND2_X2 inst_11432 ( .ZN(net_4555), .A2(net_2032), .A1(net_252) );
NAND2_X2 inst_9885 ( .ZN(net_9424), .A2(net_6106), .A1(net_2649) );
CLKBUF_X2 inst_22446 ( .A(net_22317), .Z(net_22318) );
NOR2_X4 inst_2935 ( .ZN(net_7324), .A2(net_5304), .A1(net_5228) );
CLKBUF_X2 inst_21804 ( .A(net_21646), .Z(net_21676) );
NAND2_X4 inst_7653 ( .A2(net_20800), .ZN(net_1556), .A1(net_973) );
CLKBUF_X2 inst_22788 ( .A(net_21731), .Z(net_22660) );
NOR2_X2 inst_3369 ( .A1(net_21192), .A2(net_16994), .ZN(net_16827) );
INV_X4 inst_13612 ( .ZN(net_18899), .A(net_7061) );
INV_X4 inst_17545 ( .ZN(net_2965), .A(net_167) );
INV_X4 inst_16507 ( .ZN(net_9894), .A(net_6696) );
NAND2_X2 inst_10924 ( .ZN(net_5231), .A2(net_5230), .A1(net_3854) );
INV_X4 inst_14444 ( .A(net_6665), .ZN(net_6140) );
NAND2_X2 inst_9202 ( .ZN(net_13079), .A2(net_13078), .A1(net_10304) );
NAND2_X2 inst_10179 ( .A1(net_11439), .ZN(net_8194), .A2(net_8086) );
CLKBUF_X2 inst_21585 ( .A(net_21345), .Z(net_21457) );
XNOR2_X2 inst_415 ( .B(net_21159), .ZN(net_17451), .A(net_16762) );
AOI21_X2 inst_20481 ( .ZN(net_20823), .B1(net_20240), .B2(net_14430), .A(net_7442) );
NAND2_X2 inst_10592 ( .A1(net_6896), .ZN(net_6642), .A2(net_6641) );
INV_X4 inst_17508 ( .ZN(net_5449), .A(net_1740) );
NAND2_X2 inst_12005 ( .A1(net_3426), .ZN(net_2681), .A2(net_285) );
NAND2_X2 inst_7866 ( .ZN(net_18555), .A1(net_18512), .A2(net_18486) );
NAND2_X4 inst_7652 ( .ZN(net_984), .A1(net_336), .A2(net_331) );
NAND2_X4 inst_7291 ( .A2(net_7151), .ZN(net_6970), .A1(net_4952) );
INV_X4 inst_17348 ( .ZN(net_3187), .A(net_193) );
INV_X4 inst_15772 ( .A(net_11007), .ZN(net_6934) );
NAND2_X2 inst_9074 ( .A1(net_20897), .ZN(net_13838), .A2(net_12510) );
NAND3_X2 inst_6278 ( .ZN(net_12904), .A3(net_12744), .A1(net_8607), .A2(net_7971) );
INV_X4 inst_16601 ( .ZN(net_4194), .A(net_167) );
CLKBUF_X2 inst_22898 ( .A(net_22769), .Z(net_22770) );
INV_X4 inst_15494 ( .ZN(net_2429), .A(net_2428) );
NAND2_X2 inst_10869 ( .ZN(net_6703), .A1(net_5448), .A2(net_3982) );
INV_X4 inst_14185 ( .ZN(net_12757), .A(net_7877) );
NAND2_X2 inst_10408 ( .ZN(net_10715), .A2(net_10465), .A1(net_4760) );
OAI21_X2 inst_1561 ( .B1(net_18003), .ZN(net_17264), .B2(net_16763), .A(net_2440) );
OAI21_X2 inst_2104 ( .A(net_11651), .ZN(net_10060), .B1(net_8402), .B2(net_6290) );
INV_X8 inst_12190 ( .A(net_16594), .ZN(net_16588) );
INV_X8 inst_12437 ( .ZN(net_20462), .A(net_20461) );
NAND2_X2 inst_9530 ( .A1(net_12487), .ZN(net_11110), .A2(net_9113) );
OAI211_X2 inst_2573 ( .C1(net_11366), .A(net_11245), .ZN(net_8966), .B(net_8965), .C2(net_2279) );
INV_X4 inst_16701 ( .A(net_5673), .ZN(net_2271) );
NAND2_X2 inst_8762 ( .A1(net_16359), .ZN(net_15884), .A2(net_15643) );
NAND2_X2 inst_7733 ( .ZN(net_18816), .A2(net_18785), .A1(net_17704) );
NAND3_X2 inst_6233 ( .ZN(net_13218), .A1(net_10410), .A3(net_10033), .A2(net_5457) );
INV_X4 inst_14760 ( .A(net_5587), .ZN(net_4061) );
CLKBUF_X2 inst_22285 ( .A(net_21318), .Z(net_22157) );
INV_X2 inst_19405 ( .A(net_2753), .ZN(net_1989) );
INV_X4 inst_14564 ( .A(net_7711), .ZN(net_7581) );
OAI21_X2 inst_2096 ( .ZN(net_10092), .A(net_10091), .B1(net_5803), .B2(net_5709) );
NAND2_X2 inst_10169 ( .ZN(net_14235), .A1(net_13076), .A2(net_4997) );
XNOR2_X2 inst_552 ( .B(net_16648), .A(net_16607), .ZN(net_713) );
NOR2_X2 inst_4793 ( .ZN(net_7348), .A1(net_2773), .A2(net_1678) );
AOI21_X4 inst_20145 ( .B1(net_20829), .ZN(net_15851), .B2(net_15694), .A(net_13142) );
INV_X2 inst_18394 ( .A(net_16874), .ZN(net_16521) );
NOR2_X2 inst_4997 ( .A2(net_5673), .A1(net_2872), .ZN(net_1368) );
INV_X4 inst_12483 ( .ZN(net_18701), .A(net_18683) );
OAI21_X2 inst_1564 ( .ZN(net_20086), .B2(net_16996), .A(net_16660), .B1(net_16659) );
NAND2_X4 inst_6985 ( .A1(net_20708), .A2(net_19455), .ZN(net_17183) );
NAND2_X2 inst_10995 ( .ZN(net_8478), .A1(net_8190), .A2(net_4920) );
AND3_X2 inst_21131 ( .ZN(net_14894), .A2(net_14893), .A3(net_14866), .A1(net_12544) );
INV_X4 inst_18256 ( .A(net_20957), .ZN(net_123) );
AOI21_X4 inst_20114 ( .B2(net_20960), .B1(net_20828), .ZN(net_20331), .A(net_15948) );
INV_X2 inst_19618 ( .A(net_21229), .ZN(net_40) );
NAND3_X2 inst_6477 ( .ZN(net_11277), .A3(net_11276), .A1(net_7783), .A2(net_7772) );
NAND2_X2 inst_8064 ( .ZN(net_18188), .A2(net_18187), .A1(net_17762) );
INV_X4 inst_15260 ( .ZN(net_5503), .A(net_2791) );
NAND2_X2 inst_9492 ( .ZN(net_15598), .A1(net_12295), .A2(net_9436) );
XNOR2_X2 inst_356 ( .ZN(net_16891), .A(net_16885), .B(net_14915) );
NAND2_X2 inst_9311 ( .ZN(net_12358), .A1(net_11897), .A2(net_9338) );
INV_X4 inst_17627 ( .ZN(net_1165), .A(net_294) );
NAND3_X4 inst_5587 ( .ZN(net_19125), .A3(net_13639), .A1(net_10387), .A2(net_10090) );
NAND2_X2 inst_10735 ( .ZN(net_7330), .A2(net_5770), .A1(net_5229) );
INV_X4 inst_16696 ( .ZN(net_1069), .A(net_1068) );
AOI211_X2 inst_21028 ( .C1(net_15481), .ZN(net_14565), .C2(net_12015), .B(net_9084), .A(net_8215) );
NAND2_X4 inst_6884 ( .A2(net_19207), .A1(net_19206), .ZN(net_18226) );
NAND2_X2 inst_9267 ( .ZN(net_14866), .A1(net_12609), .A2(net_12324) );
NAND2_X2 inst_9105 ( .A1(net_13922), .ZN(net_13731), .A2(net_11711) );
NOR2_X2 inst_4286 ( .A1(net_7465), .ZN(net_6050), .A2(net_3388) );
INV_X4 inst_16004 ( .ZN(net_3334), .A(net_1659) );
OAI21_X2 inst_1935 ( .ZN(net_18902), .B1(net_12930), .B2(net_9253), .A(net_3466) );
NAND3_X2 inst_6032 ( .ZN(net_14360), .A3(net_14359), .A2(net_11607), .A1(net_8623) );
NAND2_X2 inst_9332 ( .A1(net_13032), .ZN(net_12301), .A2(net_9063) );
INV_X4 inst_14949 ( .ZN(net_5874), .A(net_3512) );
NAND2_X2 inst_8678 ( .A2(net_16774), .A1(net_16469), .ZN(net_16455) );
INV_X2 inst_19133 ( .ZN(net_4182), .A(net_4181) );
NAND2_X2 inst_8235 ( .A2(net_17876), .ZN(net_17753), .A1(net_17752) );
INV_X4 inst_15927 ( .ZN(net_2516), .A(net_1734) );
INV_X4 inst_13884 ( .ZN(net_11882), .A(net_7341) );
OAI21_X2 inst_2140 ( .ZN(net_13209), .A(net_9972), .B2(net_9971), .B1(net_7159) );
INV_X4 inst_14501 ( .ZN(net_7790), .A(net_3851) );
NAND2_X2 inst_9641 ( .ZN(net_10390), .A1(net_10389), .A2(net_7764) );
NAND2_X2 inst_11386 ( .ZN(net_9650), .A2(net_3673), .A1(net_3530) );
NAND2_X2 inst_9499 ( .A1(net_14684), .ZN(net_11410), .A2(net_9830) );
AND2_X4 inst_21200 ( .A2(net_12041), .ZN(net_8794), .A1(net_8793) );
INV_X4 inst_15648 ( .ZN(net_2112), .A(net_1224) );
AOI21_X2 inst_20610 ( .ZN(net_13701), .A(net_13700), .B1(net_11061), .B2(net_10446) );
INV_X4 inst_13120 ( .ZN(net_19128), .A(net_15220) );
INV_X2 inst_19130 ( .ZN(net_4258), .A(net_4257) );
OAI21_X2 inst_1559 ( .ZN(net_17623), .B1(net_17445), .A(net_17179), .B2(net_17178) );
NAND2_X2 inst_8830 ( .ZN(net_19474), .A1(net_15831), .A2(net_15133) );
NAND3_X2 inst_6752 ( .A2(net_10536), .ZN(net_5721), .A1(net_5674), .A3(net_3430) );
SDFF_X2 inst_927 ( .Q(net_21132), .SE(net_17277), .D(net_16508), .CK(net_21634), .SI(x3910) );
CLKBUF_X2 inst_22359 ( .A(net_21667), .Z(net_22231) );
INV_X4 inst_13304 ( .ZN(net_12242), .A(net_12241) );
NAND2_X4 inst_7420 ( .ZN(net_5659), .A2(net_2058), .A1(net_1160) );
INV_X4 inst_13258 ( .ZN(net_19036), .A(net_11641) );
XNOR2_X2 inst_73 ( .ZN(net_18758), .A(net_18677), .B(net_16832) );
OAI21_X4 inst_1488 ( .B1(net_19369), .ZN(net_13396), .A(net_12522), .B2(net_6792) );
OAI21_X2 inst_1719 ( .ZN(net_19711), .A(net_14678), .B2(net_13931), .B1(net_9651) );
CLKBUF_X2 inst_22426 ( .A(net_21760), .Z(net_22298) );
NOR2_X2 inst_4690 ( .ZN(net_8345), .A2(net_3113), .A1(net_1776) );
NAND2_X2 inst_9236 ( .ZN(net_12711), .A2(net_12710), .A1(net_5064) );
SDFF_X2 inst_890 ( .Q(net_21223), .SI(net_16888), .SE(net_125), .CK(net_22220), .D(x7268) );
INV_X4 inst_12510 ( .A(net_18620), .ZN(net_18609) );
INV_X8 inst_12352 ( .ZN(net_722), .A(net_264) );
OAI21_X2 inst_1851 ( .ZN(net_14007), .A(net_14006), .B1(net_11142), .B2(net_9986) );
NAND3_X2 inst_5911 ( .ZN(net_15015), .A3(net_12822), .A1(net_9760), .A2(net_8743) );
INV_X4 inst_12896 ( .ZN(net_20632), .A(net_16864) );
NOR2_X2 inst_4514 ( .A2(net_6407), .A1(net_4194), .ZN(net_4185) );
INV_X2 inst_18842 ( .ZN(net_6691), .A(net_6690) );
NAND2_X4 inst_6903 ( .A2(net_19120), .A1(net_19119), .ZN(net_17924) );
OR2_X2 inst_1168 ( .ZN(net_6991), .A1(net_6990), .A2(net_6989) );
INV_X4 inst_12963 ( .ZN(net_16670), .A(net_16579) );
NAND2_X4 inst_7681 ( .ZN(net_1057), .A1(net_314), .A2(net_163) );
INV_X4 inst_17808 ( .ZN(net_934), .A(net_119) );
INV_X4 inst_15395 ( .ZN(net_4791), .A(net_2543) );
INV_X4 inst_15092 ( .ZN(net_3250), .A(net_3249) );
NOR2_X2 inst_4363 ( .ZN(net_5504), .A1(net_5503), .A2(net_4270) );
OR2_X2 inst_1161 ( .ZN(net_12185), .A2(net_10477), .A1(net_2212) );
NOR2_X2 inst_3362 ( .A1(net_17415), .ZN(net_17279), .A2(net_12872) );
INV_X4 inst_17743 ( .ZN(net_535), .A(net_152) );
INV_X4 inst_17308 ( .ZN(net_986), .A(net_601) );
INV_X4 inst_17177 ( .ZN(net_901), .A(net_856) );
INV_X4 inst_15667 ( .A(net_3278), .ZN(net_3039) );
INV_X4 inst_17521 ( .ZN(net_7230), .A(net_401) );
INV_X4 inst_17897 ( .ZN(net_1404), .A(net_955) );
INV_X4 inst_14096 ( .ZN(net_6186), .A(net_6185) );
INV_X4 inst_18062 ( .A(net_21203), .ZN(net_9712) );
INV_X4 inst_16739 ( .ZN(net_1380), .A(net_1048) );
AOI21_X2 inst_20815 ( .ZN(net_10075), .A(net_10074), .B2(net_4743), .B1(net_2898) );
NAND2_X2 inst_10703 ( .ZN(net_6033), .A1(net_4815), .A2(net_3477) );
OAI211_X2 inst_2388 ( .ZN(net_16273), .C2(net_15829), .A(net_15811), .B(net_14292), .C1(net_4436) );
DFF_X2 inst_19770 ( .QN(net_20868), .D(net_18586), .CK(net_22192) );
AOI21_X2 inst_20363 ( .ZN(net_15640), .B2(net_14434), .A(net_11868), .B1(net_1850) );
INV_X4 inst_15984 ( .ZN(net_12546), .A(net_9914) );
NAND3_X2 inst_5633 ( .ZN(net_18751), .A2(net_18738), .A1(net_18737), .A3(net_18663) );
NOR2_X2 inst_4309 ( .ZN(net_7415), .A1(net_6358), .A2(net_5908) );
NAND2_X2 inst_11642 ( .ZN(net_3966), .A2(net_2319), .A1(net_2193) );
NOR3_X4 inst_2634 ( .A3(net_20334), .ZN(net_19144), .A1(net_5024), .A2(net_4473) );
NOR2_X2 inst_3711 ( .ZN(net_11003), .A1(net_11002), .A2(net_11001) );
INV_X4 inst_16812 ( .ZN(net_14195), .A(net_238) );
INV_X4 inst_16408 ( .ZN(net_6733), .A(net_5785) );
INV_X4 inst_17178 ( .ZN(net_4403), .A(net_731) );
NAND2_X4 inst_7568 ( .A1(net_19150), .ZN(net_3075), .A2(net_1581) );
XNOR2_X2 inst_650 ( .B(net_634), .ZN(net_379), .A(net_378) );
XNOR2_X2 inst_289 ( .A(net_17166), .ZN(net_17149), .B(net_16462) );
CLKBUF_X2 inst_22103 ( .A(net_21260), .Z(net_21975) );
NAND2_X2 inst_8674 ( .A1(net_20791), .A2(net_16594), .ZN(net_16460) );
INV_X4 inst_12467 ( .ZN(net_18788), .A(net_18787) );
NAND2_X2 inst_8701 ( .A1(net_21220), .ZN(net_16314), .A2(net_16134) );
NAND2_X2 inst_8643 ( .A1(net_20068), .ZN(net_16572), .A2(net_16571) );
XNOR2_X1 inst_679 ( .B(net_21160), .ZN(net_18627), .A(net_18626) );
INV_X4 inst_17472 ( .ZN(net_999), .A(net_110) );
NAND3_X4 inst_5627 ( .ZN(net_9111), .A1(net_7436), .A2(net_7395), .A3(net_2058) );
INV_X4 inst_16666 ( .ZN(net_1474), .A(net_1127) );
INV_X4 inst_12532 ( .ZN(net_18386), .A(net_18385) );
NAND2_X4 inst_7689 ( .ZN(net_752), .A1(net_684), .A2(net_211) );
NOR2_X2 inst_3364 ( .ZN(net_17159), .A1(net_16868), .A2(net_16693) );
OAI21_X4 inst_1351 ( .B2(net_19510), .B1(net_19509), .A(net_18601), .ZN(net_18596) );
NAND2_X2 inst_10443 ( .A2(net_11984), .ZN(net_7185), .A1(net_6603) );
XOR2_X2 inst_44 ( .A(net_21181), .Z(net_534), .B(net_533) );
NOR2_X2 inst_4433 ( .ZN(net_19627), .A1(net_7153), .A2(net_4784) );
CLKBUF_X2 inst_21988 ( .A(net_21422), .Z(net_21860) );
INV_X4 inst_16501 ( .ZN(net_15411), .A(net_14490) );
INV_X4 inst_13994 ( .ZN(net_6414), .A(net_5273) );
CLKBUF_X2 inst_21437 ( .A(net_21283), .Z(net_21309) );
INV_X4 inst_12805 ( .ZN(net_17323), .A(net_17214) );
XNOR2_X2 inst_435 ( .ZN(net_16266), .A(net_16265), .B(net_15958) );
NAND2_X2 inst_11563 ( .ZN(net_2812), .A1(net_1949), .A2(net_1466) );
NAND2_X2 inst_10791 ( .ZN(net_10306), .A2(net_5590), .A1(net_952) );
NAND2_X2 inst_10305 ( .ZN(net_11839), .A1(net_7867), .A2(net_7866) );
AOI21_X2 inst_20600 ( .B2(net_20717), .B1(net_20716), .ZN(net_13837), .A(net_442) );
INV_X2 inst_19470 ( .A(net_3592), .ZN(net_3214) );
INV_X4 inst_13474 ( .ZN(net_9629), .A(net_9628) );
NOR2_X2 inst_3787 ( .ZN(net_10090), .A1(net_10089), .A2(net_7728) );
NOR2_X2 inst_4982 ( .A1(net_7858), .ZN(net_3711), .A2(net_2773) );
INV_X4 inst_13633 ( .ZN(net_10245), .A(net_6891) );
OAI21_X2 inst_1923 ( .A(net_14472), .ZN(net_13022), .B2(net_11489), .B1(net_6331) );
NOR3_X2 inst_2748 ( .A2(net_12530), .ZN(net_12466), .A3(net_10950), .A1(net_9312) );
NOR2_X4 inst_3013 ( .ZN(net_7317), .A1(net_5605), .A2(net_5572) );
NAND2_X2 inst_9201 ( .A1(net_13093), .ZN(net_13084), .A2(net_10296) );
NOR2_X2 inst_4744 ( .ZN(net_5545), .A2(net_3196), .A1(net_1376) );
DFF_X1 inst_19828 ( .D(net_17664), .CK(net_22551), .Q(x8) );
CLKBUF_X2 inst_22372 ( .A(net_22243), .Z(net_22244) );
NOR2_X2 inst_5087 ( .A1(net_20851), .A2(net_3861), .ZN(net_1201) );
NAND2_X2 inst_9130 ( .A1(net_15104), .ZN(net_13528), .A2(net_10789) );
NAND2_X4 inst_7563 ( .ZN(net_2391), .A2(net_770), .A1(net_295) );
INV_X4 inst_14656 ( .A(net_15369), .ZN(net_4364) );
NAND2_X2 inst_11127 ( .ZN(net_12994), .A1(net_7890), .A2(net_4279) );
INV_X4 inst_13931 ( .ZN(net_8176), .A(net_5541) );
NOR3_X2 inst_2734 ( .ZN(net_12822), .A1(net_10125), .A3(net_8753), .A2(net_7351) );
NOR2_X2 inst_4920 ( .A2(net_6538), .ZN(net_4209), .A1(net_170) );
INV_X4 inst_14956 ( .ZN(net_19998), .A(net_3499) );
INV_X2 inst_18959 ( .ZN(net_5447), .A(net_5446) );
NAND2_X2 inst_11608 ( .ZN(net_4495), .A2(net_4293), .A1(net_1381) );
NAND3_X2 inst_6518 ( .A1(net_11243), .ZN(net_10650), .A3(net_7869), .A2(net_6962) );
SDFF_X2 inst_855 ( .Q(net_21200), .SI(net_17211), .SE(net_125), .CK(net_21657), .D(x6089) );
DFF_X1 inst_19867 ( .D(net_17067), .CK(net_21337), .Q(x256) );
OAI21_X2 inst_2039 ( .ZN(net_11299), .A(net_11263), .B1(net_9728), .B2(net_9625) );
INV_X4 inst_15241 ( .ZN(net_2820), .A(net_2819) );
NOR2_X4 inst_3233 ( .ZN(net_4330), .A1(net_2532), .A2(net_1622) );
CLKBUF_X2 inst_22043 ( .A(net_21914), .Z(net_21915) );
INV_X4 inst_15226 ( .A(net_3767), .ZN(net_2858) );
NAND3_X2 inst_5866 ( .A3(net_20740), .A1(net_20739), .ZN(net_20289), .A2(net_5690) );
CLKBUF_X2 inst_21604 ( .A(net_21475), .Z(net_21476) );
NAND4_X2 inst_5466 ( .A1(net_19215), .ZN(net_19133), .A2(net_11272), .A3(net_10630), .A4(net_8987) );
NAND2_X4 inst_7588 ( .A1(net_20676), .ZN(net_1834), .A2(net_1333) );
NAND2_X2 inst_10160 ( .ZN(net_9730), .A1(net_8260), .A2(net_6185) );
NOR2_X2 inst_4295 ( .A1(net_6321), .ZN(net_5973), .A2(net_5972) );
XNOR2_X2 inst_518 ( .ZN(net_5237), .A(net_5236), .B(net_1897) );
INV_X2 inst_19196 ( .ZN(net_4596), .A(net_3627) );
NAND3_X2 inst_5894 ( .A3(net_20423), .A2(net_20422), .ZN(net_20126), .A1(net_13326) );
NAND2_X2 inst_8242 ( .ZN(net_17805), .A1(net_17556), .A2(net_17468) );
NOR2_X2 inst_3863 ( .ZN(net_9389), .A2(net_9388), .A1(net_3822) );
CLKBUF_X2 inst_22081 ( .A(net_21656), .Z(net_21953) );
OAI21_X2 inst_2345 ( .ZN(net_4359), .A(net_4358), .B2(net_4357), .B1(net_3216) );
INV_X16 inst_19742 ( .ZN(net_981), .A(net_915) );
NAND2_X1 inst_12157 ( .A1(net_7295), .ZN(net_6747), .A2(net_5498) );
INV_X4 inst_18081 ( .A(net_21150), .ZN(net_481) );
NAND3_X2 inst_6538 ( .A3(net_12782), .ZN(net_10577), .A1(net_7421), .A2(net_6254) );
NOR2_X2 inst_3602 ( .ZN(net_12533), .A1(net_12532), .A2(net_11479) );
NAND2_X2 inst_9614 ( .ZN(net_10710), .A1(net_10709), .A2(net_10708) );
INV_X4 inst_15967 ( .ZN(net_3351), .A(net_3205) );
INV_X4 inst_14291 ( .A(net_10435), .ZN(net_6949) );
NAND2_X4 inst_7582 ( .ZN(net_3068), .A2(net_1625), .A1(net_756) );
NAND4_X2 inst_5260 ( .A4(net_19781), .A1(net_19780), .ZN(net_16231), .A2(net_15266), .A3(net_13793) );
INV_X4 inst_12637 ( .ZN(net_20107), .A(net_17914) );
NAND2_X2 inst_11815 ( .A2(net_9090), .ZN(net_6476), .A1(net_1828) );
INV_X4 inst_17291 ( .ZN(net_3332), .A(net_225) );
INV_X8 inst_12336 ( .ZN(net_1014), .A(net_987) );
NAND4_X4 inst_5190 ( .A3(net_18914), .A1(net_18913), .ZN(net_16517), .A4(net_16232), .A2(net_14355) );
OAI21_X4 inst_1354 ( .ZN(net_18357), .B2(net_18299), .A(net_18216), .B1(net_17820) );
SDFF_X2 inst_970 ( .QN(net_21094), .D(net_746), .SE(net_263), .CK(net_21772), .SI(x1483) );
INV_X4 inst_18088 ( .A(net_21242), .ZN(net_103) );
NAND3_X2 inst_6731 ( .ZN(net_20408), .A2(net_6484), .A1(net_3763), .A3(net_2821) );
OAI22_X2 inst_1278 ( .ZN(net_16155), .B1(net_16051), .A1(net_16050), .A2(net_15776), .B2(net_14539) );
NOR2_X2 inst_3763 ( .ZN(net_10305), .A2(net_8678), .A1(net_7642) );
AOI21_X2 inst_20534 ( .ZN(net_20363), .B1(net_20229), .A(net_12925), .B2(net_11910) );
NAND2_X2 inst_10136 ( .ZN(net_8329), .A1(net_8328), .A2(net_6277) );
SDFF_X2 inst_749 ( .Q(net_20975), .SE(net_18581), .SI(net_18542), .D(net_11047), .CK(net_21910) );
INV_X4 inst_15159 ( .ZN(net_3430), .A(net_3039) );
NAND2_X2 inst_11975 ( .ZN(net_2279), .A1(net_1329), .A2(net_1328) );
SDFF_X2 inst_1030 ( .QN(net_20997), .D(net_1883), .SE(net_263), .CK(net_21828), .SI(x3079) );
AOI21_X2 inst_20902 ( .ZN(net_7717), .A(net_5479), .B2(net_4182), .B1(net_3966) );
NOR3_X2 inst_2649 ( .A3(net_19564), .A1(net_19563), .ZN(net_18890), .A2(net_5321) );
CLKBUF_X2 inst_21940 ( .A(net_21358), .Z(net_21812) );
NAND2_X2 inst_11441 ( .ZN(net_3474), .A2(net_3301), .A1(net_2727) );
CLKBUF_X2 inst_21700 ( .A(net_21571), .Z(net_21572) );
NOR2_X2 inst_3828 ( .ZN(net_11673), .A1(net_8874), .A2(net_6147) );
AND2_X4 inst_21261 ( .ZN(net_9031), .A2(net_4770), .A1(net_3842) );
NAND3_X2 inst_5841 ( .ZN(net_15484), .A3(net_14680), .A1(net_12136), .A2(net_8183) );
NAND2_X4 inst_6898 ( .A2(net_19301), .A1(net_19300), .ZN(net_17997) );
CLKBUF_X2 inst_22875 ( .A(net_22531), .Z(net_22747) );
INV_X4 inst_17006 ( .ZN(net_13343), .A(net_866) );
SDFF_X2 inst_1006 ( .QN(net_21026), .D(net_688), .SE(net_263), .CK(net_21955), .SI(x2554) );
OAI21_X2 inst_1985 ( .B2(net_12762), .ZN(net_12059), .A(net_10049), .B1(net_855) );
NAND2_X4 inst_7311 ( .ZN(net_6779), .A2(net_5875), .A1(net_4369) );
INV_X4 inst_17981 ( .A(net_21003), .ZN(net_1874) );
INV_X4 inst_14878 ( .ZN(net_6315), .A(net_3681) );
INV_X4 inst_13519 ( .A(net_9380), .ZN(net_9379) );
NAND2_X2 inst_10473 ( .A1(net_11245), .ZN(net_6985), .A2(net_6983) );
NAND2_X2 inst_9817 ( .A2(net_13880), .ZN(net_9653), .A1(net_9652) );
AOI21_X2 inst_20839 ( .A(net_9647), .B1(net_9569), .ZN(net_9275), .B2(net_3280) );
NOR2_X2 inst_5134 ( .A1(net_230), .ZN(net_187), .A2(net_54) );
NAND2_X4 inst_7180 ( .ZN(net_10876), .A1(net_9349), .A2(net_9348) );
NAND2_X2 inst_8691 ( .ZN(net_19338), .A1(net_16402), .A2(net_16270) );
NOR2_X2 inst_4753 ( .ZN(net_4224), .A1(net_3075), .A2(net_115) );
NAND2_X2 inst_10960 ( .ZN(net_6827), .A1(net_5077), .A2(net_5076) );
CLKBUF_X2 inst_21681 ( .A(net_21552), .Z(net_21553) );
INV_X4 inst_16168 ( .A(net_8128), .ZN(net_2528) );
NAND2_X2 inst_11885 ( .ZN(net_5295), .A1(net_1608), .A2(net_1359) );
NAND2_X2 inst_10082 ( .ZN(net_8636), .A2(net_8635), .A1(net_1505) );
AOI21_X2 inst_20881 ( .ZN(net_8279), .A(net_8278), .B1(net_6264), .B2(net_2848) );
NAND2_X2 inst_11957 ( .ZN(net_1879), .A2(net_1394), .A1(net_225) );
NOR2_X2 inst_4947 ( .ZN(net_1673), .A2(net_1672), .A1(net_61) );
AOI21_X2 inst_20747 ( .ZN(net_11381), .A(net_11380), .B2(net_11379), .B1(net_7113) );
NAND2_X2 inst_8915 ( .ZN(net_14964), .A1(net_14465), .A2(net_13646) );
NAND2_X2 inst_11671 ( .ZN(net_8714), .A2(net_2519), .A1(net_2375) );
AOI211_X2 inst_21015 ( .ZN(net_15556), .B(net_14741), .C1(net_10947), .A(net_10161), .C2(net_9022) );
INV_X4 inst_15986 ( .A(net_13999), .ZN(net_2520) );
INV_X2 inst_18456 ( .ZN(net_13379), .A(net_13378) );
INV_X4 inst_18208 ( .A(net_21190), .ZN(net_11888) );
NAND3_X2 inst_5783 ( .A1(net_19649), .ZN(net_19099), .A3(net_12911), .A2(net_6355) );
INV_X4 inst_16413 ( .ZN(net_2300), .A(net_1258) );
INV_X4 inst_15701 ( .ZN(net_2648), .A(net_2005) );
NAND3_X2 inst_6457 ( .ZN(net_11537), .A2(net_11536), .A3(net_11535), .A1(net_9330) );
INV_X2 inst_19211 ( .A(net_6432), .ZN(net_3507) );
NAND2_X2 inst_9898 ( .ZN(net_13102), .A1(net_9366), .A2(net_4822) );
AOI21_X2 inst_20761 ( .A(net_14014), .ZN(net_11129), .B1(net_6308), .B2(net_2383) );
NOR2_X2 inst_4184 ( .ZN(net_8062), .A1(net_6207), .A2(net_3837) );
AOI21_X2 inst_20853 ( .B1(net_9611), .ZN(net_9070), .A(net_8076), .B2(net_5301) );
NAND3_X2 inst_6531 ( .A1(net_11374), .ZN(net_10599), .A2(net_10598), .A3(net_10597) );
NAND2_X2 inst_11517 ( .ZN(net_5013), .A1(net_2739), .A2(net_1366) );
NOR2_X4 inst_3238 ( .ZN(net_4400), .A1(net_3244), .A2(net_2006) );
NOR2_X4 inst_2854 ( .A2(net_13012), .ZN(net_12724), .A1(net_1927) );
NOR2_X4 inst_3030 ( .ZN(net_6146), .A2(net_3929), .A1(net_3567) );
NAND2_X2 inst_7717 ( .ZN(net_18845), .A2(net_18803), .A1(net_17565) );
OAI21_X2 inst_2230 ( .ZN(net_8193), .A(net_7538), .B1(net_4333), .B2(net_3610) );
NAND3_X4 inst_5630 ( .ZN(net_4787), .A3(net_3805), .A2(net_3804), .A1(net_1331) );
INV_X4 inst_13028 ( .A(net_16465), .ZN(net_16414) );
INV_X2 inst_18621 ( .ZN(net_9577), .A(net_9576) );
INV_X4 inst_17512 ( .ZN(net_1345), .A(net_143) );
NAND2_X2 inst_10511 ( .ZN(net_8826), .A1(net_6884), .A2(net_6883) );
CLKBUF_X2 inst_21776 ( .A(net_21643), .Z(net_21648) );
CLKBUF_X2 inst_21564 ( .A(net_21435), .Z(net_21436) );
INV_X4 inst_13820 ( .A(net_12738), .ZN(net_7513) );
NAND2_X2 inst_10481 ( .ZN(net_10597), .A1(net_7975), .A2(net_6960) );
INV_X4 inst_14964 ( .ZN(net_6357), .A(net_2667) );
AOI21_X2 inst_20318 ( .A(net_20960), .B2(net_20255), .B1(net_20254), .ZN(net_15948) );
INV_X4 inst_18153 ( .A(net_21099), .ZN(net_431) );
INV_X4 inst_14174 ( .A(net_12447), .ZN(net_5995) );
NOR2_X2 inst_4477 ( .ZN(net_5651), .A1(net_4288), .A2(net_4091) );
OAI211_X2 inst_2391 ( .ZN(net_16165), .C1(net_15991), .A(net_15911), .B(net_15637), .C2(net_14803) );
NAND2_X4 inst_7606 ( .ZN(net_2561), .A2(net_1669), .A1(net_621) );
AOI21_X4 inst_20234 ( .ZN(net_12437), .B1(net_12436), .B2(net_8376), .A(net_7490) );
INV_X4 inst_17588 ( .ZN(net_709), .A(net_336) );
INV_X4 inst_14837 ( .ZN(net_11258), .A(net_3863) );
OAI21_X2 inst_2239 ( .ZN(net_20736), .A(net_8328), .B1(net_7653), .B2(net_6071) );
INV_X4 inst_15601 ( .ZN(net_12852), .A(net_2368) );
NAND2_X2 inst_10027 ( .A2(net_10625), .ZN(net_8752), .A1(net_3396) );
AOI21_X2 inst_20509 ( .ZN(net_14631), .B1(net_14630), .B2(net_11954), .A(net_10642) );
NAND3_X2 inst_6335 ( .A2(net_13412), .ZN(net_12445), .A3(net_12444), .A1(net_4885) );
OAI21_X2 inst_1639 ( .ZN(net_15951), .B1(net_15950), .A(net_15372), .B2(net_15227) );
INV_X4 inst_13645 ( .ZN(net_9672), .A(net_6847) );
NAND2_X2 inst_11468 ( .ZN(net_3157), .A1(net_3156), .A2(net_3155) );
NAND2_X2 inst_10717 ( .A1(net_6736), .ZN(net_5911), .A2(net_5910) );
INV_X4 inst_15443 ( .ZN(net_2882), .A(net_2500) );
INV_X4 inst_14743 ( .ZN(net_6808), .A(net_5571) );
NOR2_X1 inst_5155 ( .A1(net_14990), .A2(net_10475), .ZN(net_8814) );
AND3_X2 inst_21136 ( .ZN(net_13207), .A1(net_13206), .A3(net_13205), .A2(net_12928) );
DFF_X2 inst_19779 ( .D(net_5512), .Q(net_25), .CK(net_21512) );
NAND2_X2 inst_10365 ( .ZN(net_9102), .A2(net_4568), .A1(net_154) );
NAND2_X2 inst_11071 ( .ZN(net_4484), .A2(net_4196), .A1(net_703) );
CLKBUF_X2 inst_21857 ( .A(net_21431), .Z(net_21729) );
NAND2_X2 inst_9756 ( .ZN(net_10009), .A1(net_10008), .A2(net_6882) );
NAND2_X4 inst_7403 ( .ZN(net_4479), .A2(net_4326), .A1(net_3311) );
XNOR2_X2 inst_155 ( .ZN(net_17960), .A(net_17865), .B(net_17331) );
AOI21_X4 inst_20197 ( .ZN(net_20725), .B2(net_19181), .B1(net_19180), .A(net_13576) );
NOR2_X2 inst_4858 ( .ZN(net_5681), .A1(net_2422), .A2(net_2273) );
NAND2_X2 inst_10170 ( .ZN(net_9703), .A1(net_8224), .A2(net_4947) );
NAND3_X2 inst_6043 ( .ZN(net_14263), .A3(net_14262), .A2(net_12072), .A1(net_9652) );
NAND4_X2 inst_5309 ( .ZN(net_20604), .A4(net_14786), .A1(net_12145), .A3(net_10674), .A2(net_9928) );
XOR2_X1 inst_55 ( .A(net_21122), .B(net_16846), .Z(net_16831) );
OAI21_X2 inst_2280 ( .A(net_13274), .ZN(net_6880), .B1(net_6457), .B2(net_2780) );
NAND2_X2 inst_9872 ( .ZN(net_9470), .A1(net_9461), .A2(net_7409) );
NAND2_X4 inst_7097 ( .A1(net_18943), .ZN(net_14052), .A2(net_14051) );
NOR2_X2 inst_4127 ( .ZN(net_6965), .A2(net_6482), .A1(net_3625) );
INV_X4 inst_17786 ( .A(net_6078), .ZN(net_138) );
INV_X4 inst_17440 ( .ZN(net_7173), .A(net_475) );
NAND2_X2 inst_11634 ( .ZN(net_2622), .A2(net_783), .A1(net_222) );
DFF_X1 inst_19839 ( .D(net_17325), .CK(net_21608), .Q(x643) );
XNOR2_X2 inst_323 ( .B(net_17247), .A(net_17040), .ZN(net_17034) );
OAI21_X4 inst_1494 ( .ZN(net_13780), .B1(net_12525), .B2(net_4724), .A(net_749) );
AOI211_X2 inst_21005 ( .ZN(net_15890), .C1(net_15889), .C2(net_15176), .A(net_13186), .B(net_13183) );
INV_X4 inst_17792 ( .A(net_3745), .ZN(net_134) );
NOR2_X2 inst_3525 ( .ZN(net_19761), .A1(net_11576), .A2(net_8749) );
INV_X4 inst_12734 ( .A(net_17586), .ZN(net_17550) );
NAND2_X2 inst_10479 ( .A2(net_10629), .ZN(net_6975), .A1(net_3245) );
CLKBUF_X2 inst_21542 ( .A(net_21380), .Z(net_21414) );
NOR2_X2 inst_3449 ( .ZN(net_14935), .A2(net_13775), .A1(net_11787) );
INV_X16 inst_19733 ( .ZN(net_3915), .A(net_765) );
INV_X4 inst_18236 ( .A(net_21218), .ZN(net_396) );
INV_X4 inst_17748 ( .ZN(net_1002), .A(net_169) );
INV_X4 inst_17332 ( .ZN(net_2314), .A(net_129) );
OAI221_X2 inst_1340 ( .ZN(net_14228), .C1(net_14227), .C2(net_14226), .B2(net_13746), .A(net_12812), .B1(net_11460) );
OAI21_X4 inst_1481 ( .B2(net_20002), .B1(net_20001), .ZN(net_14481), .A(net_14153) );
INV_X4 inst_14275 ( .ZN(net_17366), .A(net_15537) );
INV_X4 inst_18326 ( .A(net_20923), .ZN(net_20541) );
INV_X2 inst_18563 ( .ZN(net_10780), .A(net_10779) );
INV_X4 inst_14785 ( .ZN(net_4543), .A(net_4023) );
INV_X4 inst_13194 ( .ZN(net_14125), .A(net_13464) );
NAND2_X2 inst_10191 ( .ZN(net_8156), .A1(net_7173), .A2(net_4461) );
NAND2_X2 inst_7794 ( .ZN(net_18783), .A2(net_18703), .A1(net_17064) );
INV_X4 inst_13349 ( .ZN(net_11028), .A(net_11027) );
AOI21_X2 inst_20576 ( .ZN(net_14105), .B1(net_14104), .B2(net_10574), .A(net_8595) );
INV_X4 inst_17164 ( .ZN(net_1784), .A(net_930) );
NAND2_X2 inst_9355 ( .ZN(net_18898), .A2(net_9893), .A1(net_884) );
NAND2_X2 inst_8788 ( .ZN(net_20093), .A1(net_15636), .A2(net_15163) );
INV_X4 inst_16968 ( .ZN(net_1764), .A(net_898) );
NAND2_X2 inst_10128 ( .ZN(net_8352), .A2(net_8351), .A1(net_6010) );
NAND2_X2 inst_7707 ( .ZN(net_18868), .A2(net_18857), .A1(net_18855) );
NAND2_X2 inst_10204 ( .A2(net_8867), .ZN(net_8119), .A1(net_4995) );
NOR2_X4 inst_3217 ( .ZN(net_4462), .A2(net_2483), .A1(net_1955) );
NAND2_X2 inst_9556 ( .ZN(net_11008), .A1(net_11007), .A2(net_11006) );
NAND3_X2 inst_6440 ( .ZN(net_11812), .A2(net_11811), .A3(net_9599), .A1(net_5953) );
INV_X4 inst_14506 ( .A(net_11212), .ZN(net_4825) );
NOR2_X2 inst_4376 ( .A1(net_5754), .ZN(net_5389), .A2(net_3740) );
AOI21_X2 inst_20452 ( .ZN(net_15063), .B1(net_13493), .B2(net_11789), .A(net_1275) );
NAND2_X2 inst_11778 ( .ZN(net_2029), .A2(net_253), .A1(x6071) );
NAND3_X2 inst_6023 ( .ZN(net_14381), .A3(net_11619), .A2(net_9306), .A1(net_7839) );
INV_X4 inst_17845 ( .A(net_790), .ZN(net_99) );
INV_X2 inst_18547 ( .A(net_12791), .ZN(net_10944) );
NOR2_X4 inst_3044 ( .A1(net_19213), .ZN(net_6213), .A2(net_3402) );
NAND4_X2 inst_5443 ( .ZN(net_13884), .A3(net_13883), .A4(net_11329), .A1(net_9867), .A2(net_8876) );
CLKBUF_X2 inst_22701 ( .A(net_22572), .Z(net_22573) );
INV_X4 inst_14493 ( .ZN(net_9932), .A(net_4845) );
NAND2_X2 inst_11914 ( .A2(net_4516), .ZN(net_3221), .A1(net_168) );
CLKBUF_X2 inst_21388 ( .A(net_21256), .Z(net_21260) );
INV_X8 inst_12324 ( .ZN(net_4711), .A(net_2339) );
OR2_X4 inst_1072 ( .ZN(net_8754), .A1(net_8753), .A2(net_8703) );
CLKBUF_X2 inst_22653 ( .A(net_22524), .Z(net_22525) );
OAI21_X2 inst_1993 ( .ZN(net_19514), .A(net_15077), .B1(net_10927), .B2(net_6756) );
CLKBUF_X2 inst_22884 ( .A(net_21942), .Z(net_22756) );
INV_X4 inst_15744 ( .A(net_16076), .ZN(net_1947) );
INV_X4 inst_14193 ( .ZN(net_12968), .A(net_5976) );
NAND2_X2 inst_9791 ( .A1(net_10539), .ZN(net_9720), .A2(net_9719) );
INV_X4 inst_15439 ( .A(net_9301), .ZN(net_3067) );
NAND3_X2 inst_6671 ( .ZN(net_7762), .A2(net_7751), .A3(net_5893), .A1(net_5082) );
INV_X4 inst_17326 ( .ZN(net_3737), .A(net_1740) );
INV_X4 inst_15580 ( .ZN(net_2270), .A(net_2269) );
CLKBUF_X2 inst_22940 ( .A(net_22811), .Z(net_22812) );
NAND3_X2 inst_6470 ( .ZN(net_11294), .A2(net_11293), .A3(net_11292), .A1(net_2784) );
NOR2_X2 inst_3617 ( .ZN(net_12371), .A1(net_12370), .A2(net_5879) );
NAND2_X2 inst_10893 ( .A1(net_20562), .ZN(net_8975), .A2(net_5400) );
OAI21_X4 inst_1377 ( .B1(net_19930), .ZN(net_19423), .B2(net_16357), .A(net_16223) );
INV_X4 inst_15513 ( .A(net_10292), .ZN(net_2407) );
AND2_X4 inst_21249 ( .ZN(net_4343), .A1(net_1165), .A2(net_955) );
INV_X4 inst_14828 ( .ZN(net_6588), .A(net_5393) );
OAI21_X2 inst_2201 ( .ZN(net_8561), .A(net_8560), .B1(net_8559), .B2(net_5367) );
NAND2_X2 inst_10581 ( .ZN(net_6677), .A2(net_6676), .A1(net_4385) );
AND2_X4 inst_21227 ( .ZN(net_7947), .A2(net_2867), .A1(net_837) );
INV_X4 inst_14144 ( .ZN(net_20019), .A(net_6061) );
INV_X4 inst_15835 ( .ZN(net_3367), .A(net_3082) );
NAND3_X2 inst_5671 ( .A3(net_19569), .A1(net_19568), .ZN(net_16374), .A2(net_12755) );
INV_X4 inst_17084 ( .ZN(net_3707), .A(net_3185) );
INV_X4 inst_15990 ( .ZN(net_1910), .A(net_573) );
NOR2_X2 inst_4911 ( .A2(net_2681), .ZN(net_1926), .A1(net_1925) );
NOR2_X2 inst_4525 ( .ZN(net_7000), .A1(net_3970), .A2(net_131) );
NOR2_X2 inst_4115 ( .ZN(net_20625), .A2(net_12952), .A1(net_7058) );
INV_X4 inst_13264 ( .ZN(net_12661), .A(net_12660) );
NAND2_X2 inst_8174 ( .A2(net_20774), .ZN(net_17941), .A1(net_17882) );
NAND2_X2 inst_8417 ( .ZN(net_17326), .A1(net_16927), .A2(net_16753) );
NAND3_X4 inst_5591 ( .ZN(net_15144), .A2(net_13317), .A3(net_13288), .A1(net_6673) );
OAI21_X2 inst_1687 ( .B1(net_15553), .ZN(net_15397), .A(net_14558), .B2(net_12263) );
INV_X4 inst_14983 ( .A(net_4807), .ZN(net_3412) );
OAI21_X2 inst_1970 ( .ZN(net_12228), .A(net_9142), .B2(net_6411), .B1(net_5415) );
NAND2_X4 inst_7137 ( .A1(net_19773), .ZN(net_10083), .A2(net_7887) );
INV_X8 inst_12211 ( .ZN(net_9635), .A(net_6247) );
NAND3_X2 inst_6790 ( .ZN(net_9798), .A1(net_7010), .A2(net_4108), .A3(net_2831) );
INV_X4 inst_14100 ( .ZN(net_9373), .A(net_6178) );
NAND2_X2 inst_10256 ( .ZN(net_7997), .A2(net_6079), .A1(net_5020) );
CLKBUF_X2 inst_21385 ( .A(net_21256), .Z(net_21257) );
NAND2_X4 inst_7417 ( .A1(net_19529), .ZN(net_5322), .A2(net_131) );
CLKBUF_X2 inst_22807 ( .A(net_22678), .Z(net_22679) );
INV_X4 inst_12576 ( .A(net_18210), .ZN(net_18176) );
CLKBUF_X2 inst_22086 ( .A(net_21957), .Z(net_21958) );
NOR2_X2 inst_4842 ( .A1(net_3456), .ZN(net_2364), .A2(net_1367) );
NOR3_X2 inst_2663 ( .ZN(net_20246), .A3(net_12990), .A1(net_12297), .A2(net_8883) );
NOR2_X4 inst_3289 ( .A2(net_20495), .ZN(net_3121), .A1(net_1204) );
AOI21_X2 inst_20381 ( .A(net_21220), .ZN(net_15543), .B2(net_14594), .B1(net_13115) );
NAND2_X4 inst_7477 ( .ZN(net_3476), .A1(net_2585), .A2(net_2584) );
INV_X4 inst_15911 ( .ZN(net_10383), .A(net_8741) );
INV_X4 inst_15597 ( .ZN(net_2897), .A(net_2225) );
NAND2_X2 inst_7930 ( .ZN(net_18441), .A1(net_18414), .A2(net_17822) );
INV_X4 inst_12650 ( .ZN(net_17869), .A(net_17868) );
NAND2_X2 inst_12116 ( .ZN(net_1164), .A2(net_279), .A1(net_222) );
NAND2_X2 inst_10508 ( .A1(net_11461), .ZN(net_10242), .A2(net_3987) );
INV_X2 inst_19453 ( .A(net_2532), .ZN(net_1539) );
NAND2_X2 inst_12087 ( .A2(net_2495), .A1(net_1596), .ZN(net_1053) );
XNOR2_X2 inst_401 ( .A(net_19449), .ZN(net_16681), .B(net_16680) );
NAND2_X2 inst_8086 ( .ZN(net_18139), .A2(net_18116), .A1(net_16643) );
NOR2_X4 inst_3210 ( .ZN(net_5370), .A1(net_3065), .A2(net_61) );
CLKBUF_X2 inst_22904 ( .A(net_22775), .Z(net_22776) );
NAND4_X4 inst_5200 ( .ZN(net_16902), .A4(net_16326), .A1(net_16084), .A3(net_15888), .A2(net_10822) );
NAND3_X2 inst_6145 ( .ZN(net_13685), .A2(net_12866), .A1(net_12463), .A3(net_7804) );
NOR2_X2 inst_4653 ( .ZN(net_3465), .A2(net_3326), .A1(net_2357) );
NAND3_X2 inst_6087 ( .ZN(net_13953), .A1(net_12438), .A2(net_11116), .A3(net_8523) );
NAND2_X2 inst_12028 ( .ZN(net_1005), .A1(net_311), .A2(net_193) );
INV_X4 inst_17466 ( .ZN(net_995), .A(net_141) );
INV_X4 inst_14823 ( .ZN(net_4911), .A(net_3909) );
INV_X2 inst_18630 ( .ZN(net_9449), .A(net_9448) );
NOR2_X2 inst_4465 ( .ZN(net_4514), .A2(net_3908), .A1(net_2625) );
INV_X4 inst_13107 ( .ZN(net_15735), .A(net_15529) );
INV_X8 inst_12281 ( .ZN(net_9109), .A(net_3682) );
NOR2_X2 inst_4865 ( .ZN(net_12142), .A2(net_2886), .A1(net_2242) );
CLKBUF_X2 inst_21880 ( .A(net_21751), .Z(net_21752) );
INV_X4 inst_13479 ( .ZN(net_12907), .A(net_10300) );
NAND2_X2 inst_8548 ( .ZN(net_16796), .A2(net_16789), .A1(net_580) );
SDFF_X2 inst_930 ( .QN(net_21020), .D(net_714), .SE(net_263), .CK(net_21974), .SI(x2666) );
NAND2_X4 inst_7634 ( .A1(net_2388), .ZN(net_1467), .A2(net_938) );
NAND2_X2 inst_11908 ( .ZN(net_2269), .A1(net_1955), .A2(net_1625) );
NAND3_X2 inst_6801 ( .A2(net_21238), .ZN(net_10444), .A1(net_1887), .A3(net_170) );
INV_X4 inst_15248 ( .ZN(net_4864), .A(net_3820) );
NAND2_X2 inst_8494 ( .A2(net_17107), .A1(net_17099), .ZN(net_16944) );
CLKBUF_X2 inst_22273 ( .A(net_22144), .Z(net_22145) );
CLKBUF_X2 inst_22824 ( .A(net_22695), .Z(net_22696) );
NAND2_X2 inst_10453 ( .ZN(net_7038), .A2(net_7037), .A1(net_6533) );
NAND3_X2 inst_6622 ( .A2(net_14334), .A3(net_11766), .ZN(net_9054), .A1(net_9053) );
INV_X2 inst_18931 ( .ZN(net_5851), .A(net_5850) );
AOI21_X2 inst_20638 ( .ZN(net_13275), .B1(net_13274), .A(net_12069), .B2(net_9886) );
INV_X4 inst_13650 ( .ZN(net_14897), .A(net_8154) );
NOR2_X2 inst_3874 ( .ZN(net_9362), .A2(net_9361), .A1(net_5492) );
NAND2_X2 inst_9168 ( .A1(net_13362), .ZN(net_13361), .A2(net_10526) );
OAI22_X2 inst_1251 ( .ZN(net_18494), .A1(net_18493), .A2(net_18409), .B2(net_18408), .B1(net_17243) );
INV_X8 inst_12245 ( .ZN(net_3438), .A(net_2794) );
CLKBUF_X2 inst_21521 ( .A(net_21392), .Z(net_21393) );
NAND2_X4 inst_7360 ( .A1(net_20807), .ZN(net_7596), .A2(net_847) );
CLKBUF_X2 inst_22054 ( .A(net_21925), .Z(net_21926) );
INV_X4 inst_12488 ( .ZN(net_18683), .A(net_18669) );
CLKBUF_X2 inst_22038 ( .A(net_21909), .Z(net_21910) );
NAND2_X2 inst_10300 ( .A1(net_7885), .ZN(net_7884), .A2(net_4847) );
NAND2_X2 inst_10270 ( .ZN(net_19795), .A1(net_12675), .A2(net_8101) );
NAND2_X4 inst_7433 ( .ZN(net_4537), .A2(net_3300), .A1(net_1842) );
NAND2_X2 inst_9937 ( .ZN(net_9145), .A2(net_7101), .A1(net_5727) );
INV_X2 inst_18412 ( .ZN(net_16115), .A(net_16027) );
INV_X4 inst_15411 ( .ZN(net_14179), .A(net_2528) );
CLKBUF_X2 inst_22125 ( .A(net_21996), .Z(net_21997) );
NAND2_X4 inst_7369 ( .ZN(net_8696), .A1(net_4323), .A2(net_4322) );
OAI21_X2 inst_2172 ( .ZN(net_8925), .A(net_8924), .B2(net_8284), .B1(net_2205) );
NAND2_X2 inst_8005 ( .A2(net_18312), .ZN(net_18304), .A1(net_17300) );
XNOR2_X2 inst_667 ( .A(net_21160), .B(net_21128), .ZN(net_14414) );
CLKBUF_X2 inst_21903 ( .A(net_21774), .Z(net_21775) );
CLKBUF_X2 inst_22950 ( .A(net_22821), .Z(net_22822) );
INV_X4 inst_15885 ( .ZN(net_12295), .A(net_5509) );
INV_X4 inst_12646 ( .ZN(net_17880), .A(net_17879) );
NAND2_X2 inst_8870 ( .ZN(net_15299), .A2(net_14245), .A1(net_4892) );
NOR2_X4 inst_2896 ( .ZN(net_10906), .A1(net_7478), .A2(net_6201) );
INV_X4 inst_17477 ( .ZN(net_1513), .A(net_123) );
NAND2_X2 inst_8732 ( .ZN(net_16057), .A1(net_15691), .A2(net_15559) );
NOR3_X2 inst_2691 ( .ZN(net_14339), .A3(net_11449), .A2(net_7462), .A1(net_7228) );
INV_X2 inst_19254 ( .ZN(net_3213), .A(net_3212) );
INV_X4 inst_14401 ( .ZN(net_6252), .A(net_5113) );
NAND3_X2 inst_6311 ( .ZN(net_12748), .A2(net_12644), .A1(net_10997), .A3(net_6735) );
OAI21_X2 inst_1511 ( .B2(net_20471), .ZN(net_18767), .A(net_18716), .B1(net_18715) );
NAND2_X4 inst_7543 ( .A1(net_5169), .ZN(net_2541), .A2(net_2291) );
NAND2_X2 inst_10777 ( .ZN(net_10525), .A1(net_6856), .A2(net_5613) );
INV_X4 inst_17839 ( .ZN(net_2123), .A(net_1339) );
CLKBUF_X2 inst_22772 ( .A(net_21255), .Z(net_22644) );
NAND2_X2 inst_8977 ( .ZN(net_14512), .A1(net_14511), .A2(net_12845) );
NAND3_X2 inst_6645 ( .A2(net_20571), .ZN(net_13591), .A1(net_8748), .A3(net_6218) );
NOR2_X2 inst_4243 ( .ZN(net_6540), .A2(net_4992), .A1(net_2220) );
INV_X4 inst_18126 ( .A(net_20914), .ZN(net_109) );
AOI21_X4 inst_20144 ( .ZN(net_15852), .B1(net_15690), .B2(net_15306), .A(net_14306) );
INV_X4 inst_14344 ( .A(net_15869), .ZN(net_9006) );
INV_X4 inst_13659 ( .ZN(net_9616), .A(net_8114) );
OAI21_X4 inst_1504 ( .ZN(net_10057), .A(net_10056), .B1(net_7583), .B2(net_6132) );
INV_X4 inst_17730 ( .ZN(net_570), .A(net_74) );
NOR2_X2 inst_3403 ( .ZN(net_15815), .A2(net_15329), .A1(net_13454) );
INV_X2 inst_18878 ( .ZN(net_6196), .A(net_6195) );
NAND3_X2 inst_5830 ( .ZN(net_15531), .A2(net_14728), .A3(net_14717), .A1(net_12942) );
NAND2_X2 inst_9802 ( .ZN(net_11697), .A1(net_11148), .A2(net_7584) );
INV_X2 inst_19088 ( .ZN(net_7392), .A(net_4569) );
INV_X2 inst_18961 ( .ZN(net_5426), .A(net_5168) );
NAND2_X2 inst_9006 ( .ZN(net_14280), .A1(net_14279), .A2(net_13550) );
NAND2_X4 inst_7518 ( .ZN(net_3847), .A2(net_2094), .A1(net_1375) );
NAND2_X4 inst_7242 ( .ZN(net_12038), .A2(net_6996), .A1(net_896) );
NOR2_X2 inst_3807 ( .ZN(net_9837), .A2(net_7430), .A1(net_4122) );
INV_X4 inst_17825 ( .ZN(net_4073), .A(net_1733) );
OR2_X4 inst_1069 ( .A1(net_14622), .ZN(net_11117), .A2(net_11116) );
INV_X4 inst_12719 ( .ZN(net_17542), .A(net_17541) );
CLKBUF_X2 inst_22648 ( .A(net_22519), .Z(net_22520) );
NAND2_X2 inst_11327 ( .ZN(net_3746), .A1(net_3745), .A2(net_3247) );
INV_X2 inst_18954 ( .A(net_11766), .ZN(net_5540) );
INV_X4 inst_14153 ( .ZN(net_7485), .A(net_6026) );
INV_X4 inst_13083 ( .ZN(net_18944), .A(net_15986) );
NAND2_X2 inst_10326 ( .ZN(net_12742), .A2(net_7790), .A1(net_7676) );
NOR2_X2 inst_3541 ( .A1(net_14463), .ZN(net_14201), .A2(net_13371) );
CLKBUF_X2 inst_21624 ( .A(net_21465), .Z(net_21496) );
NAND2_X2 inst_11503 ( .A1(net_4073), .ZN(net_3934), .A2(net_2506) );
INV_X4 inst_13825 ( .ZN(net_11001), .A(net_10431) );
INV_X4 inst_17744 ( .ZN(net_172), .A(net_171) );
NAND4_X4 inst_5167 ( .ZN(net_18147), .A2(net_18054), .A1(net_18045), .A4(net_15651), .A3(net_15437) );
NOR2_X2 inst_3850 ( .A1(net_20077), .ZN(net_9535), .A2(net_9359) );
INV_X4 inst_16678 ( .A(net_7679), .ZN(net_5372) );
INV_X4 inst_16533 ( .A(net_10759), .ZN(net_8462) );
INV_X4 inst_12582 ( .ZN(net_19956), .A(net_18183) );
CLKBUF_X2 inst_21581 ( .A(net_21365), .Z(net_21453) );
INV_X4 inst_14368 ( .ZN(net_8254), .A(net_5199) );
NAND2_X2 inst_10972 ( .A1(net_9785), .ZN(net_4972), .A2(net_3570) );
OAI21_X2 inst_1786 ( .A(net_14949), .ZN(net_14650), .B1(net_12485), .B2(net_10478) );
INV_X4 inst_15271 ( .ZN(net_5081), .A(net_2762) );
INV_X4 inst_15688 ( .ZN(net_2032), .A(net_2031) );
XNOR2_X2 inst_496 ( .A(net_9194), .ZN(net_9005), .B(net_1856) );
NAND2_X2 inst_10639 ( .ZN(net_6420), .A2(net_4290), .A1(net_3580) );
NAND2_X4 inst_7174 ( .ZN(net_19465), .A1(net_7364), .A2(net_7010) );
CLKBUF_X2 inst_22550 ( .A(net_22421), .Z(net_22422) );
INV_X8 inst_12356 ( .ZN(net_10714), .A(net_251) );
NAND2_X2 inst_10304 ( .ZN(net_11824), .A2(net_5847), .A1(net_5459) );
NAND4_X2 inst_5369 ( .ZN(net_15237), .A4(net_14016), .A3(net_11734), .A1(net_9073), .A2(net_8656) );
INV_X4 inst_16889 ( .ZN(net_1154), .A(net_222) );
DFF_X1 inst_19823 ( .D(net_17776), .CK(net_22118), .Q(x462) );
NAND2_X2 inst_9011 ( .ZN(net_14260), .A2(net_12715), .A1(net_12581) );
NAND3_X2 inst_5733 ( .ZN(net_16080), .A1(net_15788), .A2(net_15632), .A3(net_15258) );
NAND2_X4 inst_6867 ( .ZN(net_18390), .A2(net_18212), .A1(net_18184) );
NOR2_X2 inst_3749 ( .ZN(net_10461), .A2(net_7287), .A1(net_6729) );
NOR3_X4 inst_2620 ( .A3(net_18987), .A1(net_18986), .ZN(net_15476), .A2(net_12678) );
INV_X4 inst_17115 ( .A(net_8190), .ZN(net_5984) );
OAI21_X2 inst_1633 ( .ZN(net_16017), .B2(net_15441), .B1(net_5190), .A(net_828) );
INV_X8 inst_12425 ( .A(net_20899), .ZN(net_2274) );
OAI22_X2 inst_1262 ( .B1(net_21125), .ZN(net_17274), .B2(net_16950), .A2(net_16787), .A1(net_738) );
NAND4_X2 inst_5303 ( .ZN(net_15871), .A4(net_15298), .A2(net_13762), .A1(net_13404), .A3(net_8809) );
NAND2_X2 inst_9364 ( .ZN(net_12132), .A2(net_12131), .A1(net_12011) );
NAND2_X2 inst_8048 ( .ZN(net_18228), .A2(net_18198), .A1(net_17845) );
INV_X4 inst_16882 ( .ZN(net_1519), .A(net_996) );
NAND3_X2 inst_6799 ( .A2(net_5727), .ZN(net_3447), .A3(net_3446), .A1(net_899) );
NOR2_X2 inst_3856 ( .ZN(net_9475), .A1(net_9474), .A2(net_4983) );
INV_X8 inst_12453 ( .A(net_20923), .ZN(net_20568) );
CLKBUF_X2 inst_22929 ( .A(net_22800), .Z(net_22801) );
AOI22_X2 inst_19997 ( .ZN(net_14364), .A1(net_14363), .A2(net_12473), .B1(net_10756), .B2(net_9089) );
NOR2_X2 inst_5091 ( .A1(net_2329), .ZN(net_1156), .A2(net_257) );
INV_X4 inst_14169 ( .ZN(net_7474), .A(net_6006) );
NAND2_X2 inst_11650 ( .ZN(net_8554), .A2(net_1587), .A1(net_1545) );
INV_X4 inst_12577 ( .ZN(net_18175), .A(net_18174) );
NAND2_X2 inst_11482 ( .ZN(net_7104), .A1(net_2125), .A2(net_896) );
NAND3_X2 inst_6432 ( .ZN(net_11879), .A3(net_11878), .A2(net_6976), .A1(net_5231) );
AOI21_X2 inst_20847 ( .ZN(net_9117), .B2(net_5619), .B1(net_5338), .A(net_320) );
INV_X4 inst_16891 ( .ZN(net_4299), .A(net_952) );
NAND2_X2 inst_10716 ( .ZN(net_12813), .A2(net_5933), .A1(net_4876) );
INV_X4 inst_16615 ( .ZN(net_8720), .A(net_4270) );
OR2_X4 inst_1077 ( .A1(net_11296), .A2(net_11029), .ZN(net_7933) );
AOI21_X2 inst_20537 ( .ZN(net_14492), .B1(net_12425), .B2(net_11471), .A(net_8568) );
INV_X4 inst_15495 ( .ZN(net_5674), .A(net_1582) );
NAND3_X2 inst_6461 ( .ZN(net_11378), .A2(net_11290), .A1(net_5983), .A3(net_5110) );
NOR3_X2 inst_2757 ( .ZN(net_20300), .A2(net_20020), .A1(net_20019), .A3(net_9973) );
OAI21_X2 inst_1932 ( .A(net_14612), .ZN(net_12936), .B1(net_12935), .B2(net_12934) );
CLKBUF_X2 inst_22108 ( .A(net_21979), .Z(net_21980) );
NAND2_X2 inst_10822 ( .ZN(net_12782), .A2(net_5743), .A1(net_5204) );
NAND2_X2 inst_9733 ( .ZN(net_10109), .A1(net_10108), .A2(net_7664) );
NAND2_X2 inst_7884 ( .ZN(net_18516), .A1(net_18467), .A2(net_17759) );
NOR2_X2 inst_3704 ( .ZN(net_11093), .A2(net_7376), .A1(net_1663) );
INV_X4 inst_13903 ( .ZN(net_7085), .A(net_7084) );
NAND2_X2 inst_11828 ( .ZN(net_3007), .A1(net_2292), .A2(net_1644) );
INV_X2 inst_18792 ( .ZN(net_7447), .A(net_7446) );
INV_X4 inst_17129 ( .ZN(net_1789), .A(net_660) );
SDFF_X2 inst_1052 ( .QN(net_21021), .D(net_443), .SE(net_263), .CK(net_21942), .SI(x2659) );
OAI22_X2 inst_1280 ( .ZN(net_15389), .A2(net_13963), .B1(net_11485), .A1(net_10292), .B2(net_3712) );
AOI21_X2 inst_20913 ( .B2(net_10638), .A(net_10386), .ZN(net_7340), .B1(net_2262) );
AOI21_X4 inst_20181 ( .ZN(net_20192), .B2(net_19249), .B1(net_19248), .A(net_11562) );
INV_X4 inst_12740 ( .ZN(net_17440), .A(net_17439) );
NAND3_X2 inst_6435 ( .ZN(net_11831), .A2(net_11830), .A1(net_9778), .A3(net_9010) );
NAND4_X2 inst_5362 ( .ZN(net_15308), .A4(net_13597), .A3(net_11527), .A1(net_11122), .A2(net_8776) );
INV_X4 inst_13904 ( .ZN(net_7064), .A(net_5640) );
NAND2_X2 inst_9578 ( .ZN(net_10931), .A1(net_10930), .A2(net_10929) );
NAND3_X2 inst_6112 ( .ZN(net_13887), .A3(net_12526), .A1(net_8291), .A2(net_5069) );
NAND3_X2 inst_6200 ( .ZN(net_13308), .A2(net_13307), .A3(net_13306), .A1(net_8552) );
CLKBUF_X2 inst_22070 ( .A(net_21388), .Z(net_21942) );
AND2_X2 inst_21369 ( .ZN(net_2121), .A2(net_154), .A1(net_48) );
AOI21_X4 inst_20111 ( .B2(net_20904), .ZN(net_20198), .B1(net_19102), .A(net_15763) );
INV_X4 inst_14975 ( .ZN(net_4444), .A(net_3433) );
INV_X4 inst_16513 ( .ZN(net_3458), .A(net_807) );
XNOR2_X2 inst_134 ( .B(net_20297), .ZN(net_18244), .A(net_17115) );
OAI211_X2 inst_2409 ( .ZN(net_15526), .C1(net_15506), .B(net_14165), .C2(net_13895), .A(net_10537) );
NOR2_X4 inst_3322 ( .ZN(net_1687), .A2(net_814), .A1(net_776) );
NOR2_X2 inst_3425 ( .ZN(net_20700), .A2(net_14983), .A1(net_10380) );
OAI21_X2 inst_2328 ( .ZN(net_5290), .B1(net_5289), .B2(net_5288), .A(net_4355) );
NAND2_X2 inst_8060 ( .ZN(net_19392), .A2(net_18198), .A1(net_18171) );
NAND3_X2 inst_5779 ( .ZN(net_15846), .A3(net_15357), .A1(net_13570), .A2(net_9456) );
INV_X4 inst_14890 ( .A(net_4645), .ZN(net_3660) );
INV_X4 inst_18285 ( .ZN(net_20751), .A(net_20205) );
INV_X4 inst_13541 ( .ZN(net_12962), .A(net_9200) );
NOR2_X4 inst_2912 ( .ZN(net_9771), .A1(net_8316), .A2(net_6150) );
SDFF_X2 inst_762 ( .Q(net_20934), .SE(net_18856), .SI(net_18518), .D(net_695), .CK(net_21430) );
NOR2_X4 inst_3025 ( .ZN(net_6560), .A1(net_3531), .A2(net_3297) );
INV_X4 inst_15472 ( .ZN(net_19348), .A(net_2033) );
INV_X4 inst_15600 ( .ZN(net_4279), .A(net_2213) );
NAND2_X4 inst_7530 ( .ZN(net_3820), .A1(net_2117), .A2(net_954) );
INV_X4 inst_16649 ( .ZN(net_2660), .A(net_143) );
NAND2_X2 inst_10434 ( .ZN(net_7205), .A1(net_7204), .A2(net_7203) );
INV_X4 inst_16171 ( .ZN(net_15375), .A(net_6415) );
NOR2_X2 inst_4530 ( .ZN(net_6960), .A2(net_4010), .A1(net_1200) );
NAND2_X2 inst_11882 ( .ZN(net_6487), .A1(net_1617), .A2(net_247) );
AOI21_X2 inst_20425 ( .ZN(net_19241), .B1(net_14171), .B2(net_14117), .A(net_12104) );
INV_X4 inst_14607 ( .ZN(net_13588), .A(net_7346) );
AOI211_X2 inst_21034 ( .ZN(net_14349), .C1(net_14348), .C2(net_12312), .A(net_11560), .B(net_10303) );
INV_X4 inst_13843 ( .ZN(net_7479), .A(net_7478) );
OAI21_X2 inst_1956 ( .ZN(net_12535), .B1(net_9223), .B2(net_6942), .A(net_5725) );
NAND2_X2 inst_8378 ( .ZN(net_17351), .A2(net_17350), .A1(net_13949) );
NAND2_X2 inst_10687 ( .ZN(net_7517), .A1(net_6097), .A2(net_3795) );
NAND2_X2 inst_10935 ( .ZN(net_9094), .A1(net_4288), .A2(net_3669) );
SDFF_X2 inst_751 ( .Q(net_20928), .SE(net_18863), .SI(net_18533), .D(net_393), .CK(net_21440) );
DFF_X1 inst_19871 ( .D(net_17028), .CK(net_21599), .Q(x733) );
INV_X2 inst_19195 ( .ZN(net_3637), .A(net_3636) );
NOR2_X2 inst_4283 ( .A2(net_6172), .ZN(net_6084), .A1(net_6083) );
OAI211_X2 inst_2471 ( .A(net_14545), .ZN(net_13847), .B(net_13846), .C1(net_13781), .C2(net_12907) );
NOR2_X4 inst_3244 ( .ZN(net_3080), .A1(net_2712), .A2(net_2532) );
NOR2_X2 inst_3821 ( .ZN(net_9780), .A2(net_9779), .A1(net_4002) );
NAND2_X4 inst_7443 ( .ZN(net_4310), .A2(net_3187), .A1(net_2404) );
NAND3_X2 inst_5981 ( .ZN(net_14571), .A1(net_12709), .A3(net_11761), .A2(net_8484) );
INV_X4 inst_14554 ( .ZN(net_6210), .A(net_4589) );
INV_X4 inst_12675 ( .ZN(net_17739), .A(net_17738) );
INV_X4 inst_13330 ( .ZN(net_11157), .A(net_9868) );
NOR2_X2 inst_4623 ( .ZN(net_3608), .A1(net_2439), .A2(net_2170) );
NOR2_X2 inst_3835 ( .ZN(net_11543), .A1(net_10151), .A2(net_9690) );
CLKBUF_X2 inst_22483 ( .A(net_21630), .Z(net_22355) );
AOI21_X2 inst_20415 ( .B1(net_20677), .ZN(net_20160), .A(net_8275), .B2(net_6580) );
OAI21_X2 inst_2117 ( .B2(net_20211), .ZN(net_20099), .A(net_11297), .B1(net_8287) );
NOR2_X4 inst_3140 ( .ZN(net_4724), .A1(net_2647), .A2(net_640) );
INV_X4 inst_13812 ( .ZN(net_12992), .A(net_7536) );
NAND2_X2 inst_12035 ( .ZN(net_1637), .A2(net_1596), .A1(net_965) );
CLKBUF_X2 inst_22259 ( .A(net_22130), .Z(net_22131) );
INV_X4 inst_17775 ( .ZN(net_14600), .A(net_293) );
INV_X4 inst_14600 ( .A(net_7849), .ZN(net_6798) );
NAND2_X2 inst_11941 ( .A1(net_20889), .A2(net_10714), .ZN(net_8107) );
INV_X8 inst_12308 ( .ZN(net_2384), .A(net_476) );
NAND2_X2 inst_11200 ( .A1(net_8341), .ZN(net_5142), .A2(net_3295) );
NOR2_X2 inst_4642 ( .ZN(net_3394), .A2(net_3393), .A1(net_2085) );
NAND2_X4 inst_7340 ( .ZN(net_4866), .A1(net_4865), .A2(net_4864) );
NOR2_X4 inst_3316 ( .ZN(net_1064), .A2(net_684), .A1(net_211) );
INV_X2 inst_19051 ( .A(net_7031), .ZN(net_4738) );
NAND2_X2 inst_9385 ( .ZN(net_19941), .A2(net_8923), .A1(net_7916) );
NOR2_X2 inst_4411 ( .A1(net_6812), .ZN(net_6189), .A2(net_5054) );
CLKBUF_X2 inst_21649 ( .A(net_21296), .Z(net_21521) );
NAND2_X2 inst_11471 ( .ZN(net_4257), .A2(net_1575), .A1(net_1525) );
CLKBUF_X2 inst_22026 ( .A(net_21897), .Z(net_21898) );
NAND2_X2 inst_7772 ( .ZN(net_18740), .A2(net_18689), .A1(net_18674) );
NOR2_X2 inst_4014 ( .ZN(net_10300), .A1(net_8037), .A2(net_8002) );
INV_X4 inst_17087 ( .ZN(net_1091), .A(net_547) );
NOR2_X2 inst_3694 ( .ZN(net_20041), .A1(net_8125), .A2(net_7997) );
INV_X4 inst_16272 ( .ZN(net_20201), .A(net_1346) );
CLKBUF_X2 inst_21987 ( .A(net_21858), .Z(net_21859) );
INV_X4 inst_15204 ( .ZN(net_5194), .A(net_2906) );
NOR2_X2 inst_4882 ( .ZN(net_2173), .A1(net_2118), .A2(net_345) );
AOI21_X2 inst_20958 ( .B1(net_8836), .ZN(net_5334), .A(net_4167), .B2(net_2088) );
NOR3_X2 inst_2698 ( .ZN(net_14094), .A3(net_10485), .A1(net_8864), .A2(net_3650) );
NAND2_X2 inst_9908 ( .ZN(net_9334), .A1(net_7822), .A2(net_4823) );
OAI211_X2 inst_2518 ( .ZN(net_11896), .A(net_11895), .B(net_11894), .C1(net_11893), .C2(net_3200) );
NOR2_X2 inst_3460 ( .A1(net_16127), .ZN(net_14692), .A2(net_13160) );
NOR2_X1 inst_5152 ( .ZN(net_20055), .A1(net_7921), .A2(net_7065) );
CLKBUF_X2 inst_22326 ( .A(net_21648), .Z(net_22198) );
NAND3_X4 inst_5544 ( .A3(net_19556), .A1(net_19555), .ZN(net_16885), .A2(net_13188) );
INV_X2 inst_19342 ( .ZN(net_19122), .A(net_2448) );
AOI221_X2 inst_20085 ( .C1(net_16214), .ZN(net_15939), .C2(net_14777), .A(net_13806), .B2(net_13738), .B1(net_10175) );
OAI21_X2 inst_2075 ( .ZN(net_10588), .B1(net_10587), .A(net_9126), .B2(net_6458) );
OAI21_X2 inst_1911 ( .ZN(net_13077), .A(net_13076), .B1(net_9622), .B2(net_7100) );
AOI21_X2 inst_20663 ( .ZN(net_12938), .A(net_12937), .B2(net_12262), .B1(net_4154) );
NAND3_X2 inst_5689 ( .ZN(net_16289), .A1(net_16107), .A2(net_15961), .A3(net_15786) );
NAND2_X2 inst_10841 ( .ZN(net_6765), .A2(net_5559), .A1(net_5205) );
INV_X4 inst_15528 ( .A(net_10031), .ZN(net_7295) );
XNOR2_X2 inst_585 ( .ZN(net_582), .A(net_581), .B(net_580) );
INV_X4 inst_15846 ( .A(net_7663), .ZN(net_3525) );
NAND2_X2 inst_8816 ( .ZN(net_15580), .A1(net_15573), .A2(net_14843) );
NAND4_X2 inst_5435 ( .ZN(net_13957), .A1(net_13956), .A2(net_13955), .A4(net_11153), .A3(net_7711) );
NOR2_X2 inst_5107 ( .ZN(net_4615), .A1(net_1848), .A2(net_262) );
CLKBUF_X2 inst_21417 ( .A(net_21288), .Z(net_21289) );
NAND3_X2 inst_5763 ( .ZN(net_15932), .A3(net_15244), .A1(net_14590), .A2(net_14205) );
NAND2_X2 inst_11171 ( .A1(net_20551), .ZN(net_9008), .A2(net_2459) );
INV_X2 inst_18428 ( .ZN(net_14876), .A(net_14338) );
NAND2_X1 inst_12137 ( .ZN(net_17475), .A1(net_17474), .A2(net_17358) );
NAND3_X2 inst_6453 ( .ZN(net_11723), .A2(net_10202), .A1(net_8077), .A3(net_5452) );
OAI211_X2 inst_2428 ( .ZN(net_15162), .B(net_13937), .A(net_11162), .C2(net_10837), .C1(net_9289) );
NOR2_X2 inst_5115 ( .A2(net_20860), .A1(net_20859), .ZN(net_446) );
INV_X4 inst_14382 ( .ZN(net_8372), .A(net_5168) );
CLKBUF_X2 inst_22458 ( .A(net_22329), .Z(net_22330) );
NAND2_X4 inst_7553 ( .ZN(net_2970), .A2(net_1755), .A1(net_1754) );
INV_X2 inst_18966 ( .ZN(net_5320), .A(net_5319) );
INV_X4 inst_17264 ( .ZN(net_2569), .A(net_193) );
OR2_X4 inst_1124 ( .ZN(net_6524), .A2(net_1376), .A1(net_31) );
NOR2_X2 inst_4086 ( .ZN(net_19787), .A1(net_7125), .A2(net_6857) );
NAND2_X2 inst_11091 ( .ZN(net_5972), .A2(net_4361), .A1(net_3244) );
AOI21_X4 inst_20156 ( .B1(net_19827), .B2(net_15753), .ZN(net_15714), .A(net_12572) );
OAI211_X2 inst_2555 ( .B(net_16009), .ZN(net_10432), .A(net_10431), .C2(net_4556), .C1(net_4252) );
INV_X4 inst_13922 ( .ZN(net_9329), .A(net_7873) );
NAND2_X4 inst_6966 ( .A2(net_20064), .A1(net_20063), .ZN(net_18704) );
INV_X2 inst_18526 ( .A(net_11632), .ZN(net_11109) );
INV_X4 inst_13447 ( .ZN(net_14405), .A(net_9758) );
NAND4_X4 inst_5240 ( .ZN(net_19879), .A4(net_19075), .A1(net_19074), .A3(net_9491), .A2(net_8926) );
INV_X8 inst_12450 ( .A(net_20557), .ZN(net_20555) );
NAND4_X2 inst_5343 ( .ZN(net_20759), .A3(net_15457), .A1(net_14747), .A2(net_14467), .A4(net_12702) );
AOI21_X4 inst_20173 ( .B2(net_19571), .B1(net_19570), .ZN(net_15548), .A(net_14994) );
NOR2_X2 inst_3714 ( .A2(net_13324), .ZN(net_10990), .A1(net_10989) );
INV_X8 inst_12317 ( .ZN(net_1741), .A(net_211) );
INV_X8 inst_12269 ( .ZN(net_2697), .A(net_1268) );
NAND4_X2 inst_5285 ( .ZN(net_20272), .A4(net_19242), .A1(net_19241), .A2(net_13068), .A3(net_12482) );
INV_X4 inst_17972 ( .A(net_21116), .ZN(net_16648) );
CLKBUF_X2 inst_22082 ( .A(net_21953), .Z(net_21954) );
AOI21_X2 inst_20705 ( .ZN(net_12113), .B1(net_9320), .B2(net_8346), .A(net_5748) );
NAND3_X2 inst_6658 ( .A3(net_8507), .ZN(net_8465), .A1(net_4925), .A2(net_3083) );
NAND3_X4 inst_5611 ( .ZN(net_19543), .A2(net_9689), .A1(net_7987), .A3(net_7324) );
OAI22_X2 inst_1304 ( .A1(net_13544), .B1(net_13504), .A2(net_11556), .ZN(net_10494), .B2(net_4097) );
NAND2_X2 inst_9027 ( .ZN(net_14084), .A1(net_13752), .A2(net_11913) );
NAND3_X2 inst_6815 ( .ZN(net_5588), .A1(net_4526), .A2(net_3134), .A3(net_2348) );
NOR2_X4 inst_3292 ( .ZN(net_2296), .A2(net_1261), .A1(net_74) );
NAND2_X2 inst_8575 ( .A1(net_17115), .ZN(net_16730), .A2(net_16729) );
NAND2_X2 inst_7751 ( .ZN(net_18775), .A2(net_18739), .A1(net_18680) );
NOR2_X2 inst_5024 ( .A1(net_20859), .ZN(net_1177), .A2(net_867) );
INV_X2 inst_19458 ( .A(net_2097), .ZN(net_1977) );
AOI21_X2 inst_20927 ( .ZN(net_7098), .A(net_7097), .B2(net_7096), .B1(net_3315) );
SDFF_X2 inst_919 ( .Q(net_21124), .D(net_16500), .SE(net_253), .CK(net_21521), .SI(x4261) );
NAND2_X2 inst_10530 ( .ZN(net_18907), .A1(net_6826), .A2(net_6825) );
INV_X4 inst_12772 ( .A(net_17334), .ZN(net_17333) );
OAI21_X2 inst_1916 ( .ZN(net_13048), .B2(net_9538), .A(net_9364), .B1(net_2988) );
NAND2_X2 inst_9705 ( .A1(net_11784), .ZN(net_10203), .A2(net_10202) );
INV_X4 inst_14057 ( .ZN(net_9642), .A(net_8022) );
INV_X8 inst_12403 ( .A(net_766), .ZN(net_82) );
OAI21_X2 inst_1797 ( .ZN(net_14504), .B2(net_11630), .B1(net_11002), .A(net_10309) );
INV_X4 inst_17447 ( .ZN(net_4876), .A(net_81) );
NOR2_X2 inst_4408 ( .A1(net_9396), .ZN(net_8312), .A2(net_5081) );
NOR3_X2 inst_2708 ( .ZN(net_13903), .A1(net_11947), .A3(net_9700), .A2(net_8312) );
NAND3_X2 inst_6197 ( .ZN(net_13312), .A3(net_9872), .A1(net_9369), .A2(net_2760) );
INV_X4 inst_14694 ( .ZN(net_13156), .A(net_5371) );
NAND2_X2 inst_9866 ( .ZN(net_11528), .A2(net_7827), .A1(net_1790) );
NOR2_X2 inst_3530 ( .ZN(net_13572), .A1(net_13571), .A2(net_10506) );
NOR2_X2 inst_5009 ( .ZN(net_2097), .A1(net_1289), .A2(net_236) );
NOR2_X2 inst_4785 ( .A2(net_5859), .A1(net_4259), .ZN(net_2854) );
INV_X4 inst_13552 ( .ZN(net_12310), .A(net_9165) );
NAND2_X2 inst_7785 ( .ZN(net_18725), .A2(net_18713), .A1(net_17069) );
OAI211_X2 inst_2592 ( .ZN(net_5281), .B(net_5280), .C2(net_3777), .A(net_3267), .C1(net_1704) );
INV_X4 inst_18297 ( .A(net_20469), .ZN(net_20468) );
CLKBUF_X2 inst_22817 ( .A(net_22688), .Z(net_22689) );
INV_X4 inst_12752 ( .ZN(net_17412), .A(net_17411) );
NAND2_X4 inst_7331 ( .A2(net_6394), .ZN(net_4943), .A1(net_4942) );
NOR2_X4 inst_3116 ( .ZN(net_6908), .A1(net_3991), .A2(net_3937) );
INV_X4 inst_17106 ( .A(net_14945), .ZN(net_1062) );
INV_X4 inst_15624 ( .ZN(net_2154), .A(net_2153) );
NOR2_X2 inst_4378 ( .A1(net_9926), .ZN(net_5365), .A2(net_5364) );
INV_X4 inst_14682 ( .ZN(net_11808), .A(net_4297) );
NAND2_X2 inst_9682 ( .ZN(net_10259), .A2(net_7757), .A1(net_7325) );
AOI21_X2 inst_20793 ( .ZN(net_20035), .B1(net_10659), .B2(net_10493), .A(net_4338) );
INV_X4 inst_15824 ( .ZN(net_19875), .A(net_1052) );
INV_X4 inst_15589 ( .A(net_3178), .ZN(net_2254) );
INV_X4 inst_15552 ( .A(net_13383), .ZN(net_11505) );
XNOR2_X2 inst_114 ( .ZN(net_18507), .A(net_18416), .B(net_17510) );
NAND2_X2 inst_11767 ( .ZN(net_2693), .A2(net_2093), .A1(net_2074) );
NAND2_X4 inst_7116 ( .ZN(net_13742), .A2(net_11050), .A1(net_11017) );
OAI21_X2 inst_2278 ( .ZN(net_7130), .A(net_7129), .B2(net_7128), .B1(net_2404) );
NOR2_X2 inst_4866 ( .ZN(net_4084), .A2(net_1427), .A1(net_222) );
NAND2_X2 inst_11415 ( .ZN(net_3403), .A2(net_3402), .A1(net_3181) );
NAND2_X2 inst_7924 ( .ZN(net_18449), .A1(net_18333), .A2(net_18281) );
NAND2_X2 inst_7800 ( .ZN(net_20811), .A2(net_20210), .A1(net_18653) );
NOR2_X2 inst_4150 ( .A1(net_8199), .ZN(net_6904), .A2(net_4493) );
NAND2_X2 inst_9630 ( .ZN(net_10519), .A1(net_7936), .A2(net_5767) );
INV_X8 inst_12371 ( .A(net_336), .ZN(net_136) );
XNOR2_X2 inst_534 ( .ZN(net_1677), .B(net_1676), .A(net_408) );
INV_X8 inst_12422 ( .A(net_20916), .ZN(net_1697) );
CLKBUF_X2 inst_22710 ( .A(net_21505), .Z(net_22582) );
INV_X4 inst_16879 ( .A(net_7917), .ZN(net_7129) );
NAND2_X2 inst_8636 ( .A1(net_17177), .A2(net_16596), .ZN(net_16583) );
INV_X4 inst_17268 ( .ZN(net_6604), .A(net_2585) );
INV_X4 inst_13816 ( .ZN(net_7523), .A(net_7522) );
INV_X2 inst_18679 ( .ZN(net_8809), .A(net_8808) );
INV_X2 inst_19203 ( .ZN(net_3551), .A(net_3550) );
NAND2_X2 inst_9033 ( .ZN(net_14068), .A1(net_13922), .A2(net_11870) );
INV_X4 inst_16476 ( .A(net_2862), .ZN(net_1406) );
NAND2_X2 inst_10682 ( .ZN(net_6136), .A1(net_6135), .A2(net_6040) );
NAND3_X4 inst_5618 ( .ZN(net_11952), .A3(net_11720), .A2(net_7969), .A1(net_7179) );
CLKBUF_X2 inst_22917 ( .A(net_22404), .Z(net_22789) );
INV_X2 inst_18632 ( .ZN(net_9442), .A(net_9441) );
INV_X4 inst_15318 ( .ZN(net_3606), .A(net_2002) );
NAND4_X4 inst_5193 ( .A4(net_18937), .A1(net_18936), .ZN(net_18214), .A3(net_16310), .A2(net_15968) );
NOR2_X4 inst_2836 ( .ZN(net_15310), .A2(net_14406), .A1(net_13137) );
NOR2_X2 inst_4336 ( .ZN(net_9463), .A2(net_5698), .A1(net_809) );
INV_X4 inst_17350 ( .ZN(net_1101), .A(net_316) );
INV_X4 inst_16448 ( .ZN(net_18965), .A(net_1225) );
INV_X4 inst_18227 ( .A(net_21232), .ZN(net_1376) );
NAND2_X2 inst_10424 ( .A1(net_10765), .ZN(net_7223), .A2(net_6805) );
NOR3_X2 inst_2770 ( .ZN(net_8640), .A2(net_8639), .A1(net_8326), .A3(net_6017) );
NAND2_X2 inst_11735 ( .ZN(net_5367), .A2(net_3281), .A1(net_170) );
NAND2_X2 inst_9184 ( .ZN(net_13139), .A1(net_13138), .A2(net_10401) );
INV_X4 inst_14542 ( .A(net_6255), .ZN(net_4642) );
INV_X2 inst_19444 ( .A(net_9894), .ZN(net_1627) );
INV_X4 inst_15010 ( .A(net_15936), .ZN(net_15897) );
NOR2_X2 inst_4573 ( .ZN(net_4846), .A2(net_3260), .A1(net_1759) );
CLKBUF_X2 inst_22478 ( .A(net_21996), .Z(net_22350) );
NOR2_X2 inst_3444 ( .ZN(net_14965), .A1(net_14837), .A2(net_13649) );
NAND2_X4 inst_7284 ( .A1(net_19482), .ZN(net_5728), .A2(net_117) );
NAND2_X2 inst_10848 ( .ZN(net_7252), .A1(net_6812), .A2(net_4013) );
NAND2_X2 inst_9295 ( .ZN(net_19737), .A1(net_12401), .A2(net_9168) );
INV_X4 inst_14926 ( .A(net_4914), .ZN(net_3557) );
NOR2_X2 inst_4732 ( .A1(net_20489), .ZN(net_3969), .A2(net_3075) );
INV_X4 inst_17655 ( .A(net_20851), .ZN(net_2828) );
OAI21_X2 inst_2348 ( .ZN(net_3726), .A(net_3725), .B1(net_2844), .B2(net_2235) );
NOR2_X2 inst_4021 ( .ZN(net_9565), .A2(net_8022), .A1(net_5877) );
NAND2_X2 inst_11059 ( .ZN(net_8189), .A2(net_3693), .A1(net_1161) );
AOI21_X2 inst_20823 ( .ZN(net_19588), .B1(net_19515), .B2(net_8924), .A(net_4244) );
NAND2_X2 inst_9827 ( .A1(net_9658), .ZN(net_9624), .A2(net_9623) );
INV_X2 inst_18421 ( .ZN(net_15402), .A(net_15145) );
NAND2_X2 inst_8290 ( .A2(net_20461), .ZN(net_18889), .A1(net_17492) );
AOI21_X2 inst_20300 ( .ZN(net_16121), .B1(net_15995), .B2(net_15727), .A(net_14032) );
NAND2_X2 inst_11114 ( .A2(net_20579), .ZN(net_9055), .A1(net_7661) );
NAND2_X2 inst_7713 ( .ZN(net_18852), .A2(net_18835), .A1(net_18821) );
NOR2_X2 inst_5080 ( .ZN(net_871), .A1(net_709), .A2(net_106) );
NOR2_X2 inst_4666 ( .ZN(net_8803), .A2(net_3253), .A1(net_154) );
INV_X4 inst_16104 ( .ZN(net_14493), .A(net_9727) );
INV_X4 inst_14115 ( .ZN(net_6149), .A(net_6148) );
OAI21_X4 inst_1465 ( .B1(net_15697), .ZN(net_15164), .A(net_14250), .B2(net_13933) );
NAND4_X2 inst_5265 ( .ZN(net_16186), .A1(net_15828), .A4(net_15363), .A2(net_10766), .A3(net_9045) );
INV_X4 inst_13009 ( .A(net_16590), .ZN(net_16537) );
INV_X2 inst_19469 ( .A(net_1449), .ZN(net_1447) );
NAND3_X2 inst_6550 ( .A3(net_13728), .ZN(net_10532), .A1(net_6381), .A2(net_4969) );
INV_X4 inst_17205 ( .ZN(net_3988), .A(net_90) );
INV_X4 inst_15069 ( .ZN(net_5872), .A(net_3275) );
INV_X4 inst_18334 ( .A(net_20571), .ZN(net_20570) );
NOR2_X2 inst_4215 ( .ZN(net_8688), .A1(net_6636), .A2(net_5520) );
INV_X4 inst_15259 ( .ZN(net_2778), .A(net_2777) );
SDFF_X2 inst_999 ( .QN(net_21000), .SE(net_2426), .D(net_450), .CK(net_21839), .SI(x3021) );
NAND2_X2 inst_7805 ( .ZN(net_18689), .A2(net_18656), .A1(net_17394) );
INV_X8 inst_12378 ( .ZN(net_334), .A(net_121) );
INV_X2 inst_19105 ( .A(net_6225), .ZN(net_4497) );
NAND2_X2 inst_8083 ( .ZN(net_18150), .A1(net_18097), .A2(net_18083) );
CLKBUF_X2 inst_21547 ( .A(net_21418), .Z(net_21419) );
OAI21_X2 inst_1846 ( .ZN(net_14017), .A(net_11407), .B2(net_11305), .B1(net_11141) );
INV_X2 inst_19389 ( .A(net_4214), .ZN(net_2084) );
OAI21_X2 inst_2139 ( .ZN(net_13169), .B1(net_9974), .B2(net_9973), .A(net_4990) );
INV_X4 inst_17565 ( .ZN(net_10699), .A(net_6838) );
NOR2_X2 inst_4278 ( .ZN(net_6113), .A1(net_6112), .A2(net_4598) );
NAND2_X2 inst_10236 ( .ZN(net_8042), .A1(net_8041), .A2(net_6121) );
XNOR2_X2 inst_186 ( .ZN(net_17761), .B(net_17760), .A(net_17457) );
NOR2_X2 inst_4271 ( .ZN(net_7540), .A1(net_6131), .A2(net_4544) );
INV_X4 inst_16066 ( .A(net_2278), .ZN(net_1573) );
NAND2_X2 inst_10756 ( .ZN(net_6248), .A2(net_4373), .A1(net_2214) );
NAND2_X2 inst_9820 ( .A1(net_10098), .ZN(net_9644), .A2(net_5720) );
NOR2_X4 inst_3071 ( .ZN(net_5778), .A2(net_3682), .A1(net_2514) );
AOI21_X4 inst_20100 ( .B2(net_20848), .B1(net_19165), .ZN(net_18879), .A(net_15872) );
NAND2_X2 inst_10395 ( .A1(net_9072), .ZN(net_7291), .A2(net_6967) );
NAND2_X2 inst_11963 ( .ZN(net_4963), .A1(net_167), .A2(net_86) );
INV_X4 inst_13536 ( .ZN(net_12417), .A(net_9209) );
NAND2_X2 inst_8283 ( .A1(net_20524), .ZN(net_17624), .A2(net_17623) );
SDFF_X2 inst_863 ( .Q(net_21221), .SI(net_17167), .SE(net_125), .CK(net_21472), .D(x7336) );
INV_X2 inst_19484 ( .A(net_4516), .ZN(net_1337) );
INV_X4 inst_16821 ( .ZN(net_1112), .A(net_995) );
NAND2_X2 inst_8669 ( .ZN(net_16471), .A1(net_16470), .A2(net_16469) );
NAND3_X2 inst_6315 ( .ZN(net_12576), .A3(net_12508), .A2(net_12501), .A1(net_5163) );
OAI21_X4 inst_1385 ( .A(net_20888), .B2(net_19364), .B1(net_19363), .ZN(net_16325) );
INV_X4 inst_15288 ( .A(net_3940), .ZN(net_3532) );
NAND3_X2 inst_6513 ( .A2(net_12283), .A3(net_12282), .ZN(net_10753), .A1(net_3724) );
NAND3_X2 inst_5921 ( .ZN(net_14983), .A3(net_13110), .A2(net_10523), .A1(net_6686) );
AOI21_X2 inst_20758 ( .ZN(net_11202), .B2(net_9504), .B1(net_4872), .A(net_3880) );
NAND3_X2 inst_5770 ( .ZN(net_20395), .A2(net_15403), .A3(net_15120), .A1(net_14202) );
OAI21_X2 inst_1573 ( .A(net_16385), .ZN(net_16348), .B1(net_16102), .B2(net_14827) );
NAND3_X4 inst_5521 ( .A3(net_19058), .A1(net_19057), .ZN(net_18649), .A2(net_15683) );
NAND2_X2 inst_8394 ( .ZN(net_19351), .A1(net_17278), .A2(net_17162) );
OAI21_X4 inst_1390 ( .A(net_20856), .B2(net_20053), .B1(net_20052), .ZN(net_19317) );
INV_X2 inst_18738 ( .ZN(net_10135), .A(net_7920) );
XNOR2_X2 inst_229 ( .B(net_21183), .ZN(net_17497), .A(net_17198) );
NAND2_X2 inst_9124 ( .A1(net_14346), .ZN(net_13537), .A2(net_11030) );
INV_X2 inst_19008 ( .ZN(net_5019), .A(net_5018) );
INV_X4 inst_12920 ( .ZN(net_16821), .A(net_16663) );
NAND2_X2 inst_9596 ( .ZN(net_10841), .A1(net_10840), .A2(net_7451) );
NOR2_X2 inst_4992 ( .A1(net_4299), .ZN(net_3155), .A2(net_1397) );
AND2_X2 inst_21283 ( .ZN(net_13111), .A2(net_11620), .A1(net_9043) );
NOR2_X2 inst_4689 ( .A2(net_11845), .ZN(net_7122), .A1(net_165) );
INV_X4 inst_17063 ( .ZN(net_2953), .A(net_819) );
NAND2_X2 inst_11719 ( .ZN(net_3304), .A1(net_2431), .A2(net_2260) );
NAND3_X2 inst_6151 ( .ZN(net_13677), .A2(net_13676), .A1(net_11205), .A3(net_8941) );
NAND2_X2 inst_9187 ( .ZN(net_13130), .A1(net_13129), .A2(net_11690) );
OAI21_X2 inst_2131 ( .ZN(net_9995), .A(net_9994), .B2(net_9993), .B1(net_8122) );
NAND2_X2 inst_12007 ( .A1(net_2563), .ZN(net_1566), .A2(net_1165) );
NAND2_X2 inst_9949 ( .ZN(net_10424), .A2(net_8941), .A1(net_6356) );
NAND2_X4 inst_7297 ( .ZN(net_11587), .A2(net_5572), .A1(net_5571) );
NAND2_X2 inst_8804 ( .ZN(net_19386), .A2(net_15355), .A1(net_14439) );
CLKBUF_X2 inst_22869 ( .A(net_22740), .Z(net_22741) );
NAND2_X2 inst_9453 ( .ZN(net_11512), .A1(net_11511), .A2(net_9645) );
XNOR2_X2 inst_421 ( .B(net_21132), .ZN(net_16508), .A(net_16506) );
NAND2_X2 inst_11263 ( .ZN(net_9887), .A1(net_3900), .A2(net_3819) );
NAND2_X4 inst_7016 ( .ZN(net_17237), .A1(net_16603), .A2(net_16468) );
SDFF_X2 inst_816 ( .Q(net_21161), .SI(net_17772), .SE(net_125), .CK(net_21484), .D(x5290) );
NAND2_X2 inst_11000 ( .ZN(net_6048), .A2(net_3498), .A1(net_703) );
INV_X4 inst_16824 ( .ZN(net_15156), .A(net_449) );
INV_X4 inst_12911 ( .A(net_16909), .ZN(net_16685) );
NOR3_X2 inst_2798 ( .ZN(net_2675), .A1(net_2674), .A2(net_2673), .A3(net_170) );
CLKBUF_X2 inst_21899 ( .A(net_21770), .Z(net_21771) );
INV_X4 inst_12903 ( .ZN(net_17101), .A(net_17099) );
INV_X4 inst_12692 ( .ZN(net_17645), .A(net_17644) );
INV_X4 inst_13694 ( .ZN(net_11399), .A(net_7929) );
NAND2_X4 inst_7596 ( .ZN(net_3138), .A1(net_1583), .A2(net_958) );
AOI21_X2 inst_20884 ( .A(net_7915), .ZN(net_7824), .B2(net_6336), .B1(net_2692) );
OR2_X4 inst_1108 ( .ZN(net_2448), .A1(net_1503), .A2(net_1355) );
INV_X2 inst_19013 ( .ZN(net_5002), .A(net_5001) );
NOR2_X1 inst_5148 ( .A1(net_10952), .ZN(net_10951), .A2(net_10950) );
INV_X2 inst_19519 ( .A(net_1633), .ZN(net_1121) );
NOR2_X2 inst_4534 ( .A1(net_7886), .A2(net_4229), .ZN(net_4040) );
CLKBUF_X2 inst_21405 ( .A(net_21249), .Z(net_21277) );
NAND2_X2 inst_8286 ( .A2(net_20584), .ZN(net_17622), .A1(net_17324) );
INV_X4 inst_15901 ( .ZN(net_9247), .A(net_1745) );
NAND2_X2 inst_11422 ( .ZN(net_6927), .A1(net_3368), .A2(net_3367) );
INV_X4 inst_16288 ( .ZN(net_6613), .A(net_896) );
NAND2_X2 inst_8604 ( .A2(net_20765), .ZN(net_18971), .A1(net_3434) );
CLKBUF_X2 inst_22134 ( .A(net_21536), .Z(net_22006) );
NAND2_X2 inst_9718 ( .ZN(net_10163), .A1(net_10162), .A2(net_7713) );
AOI21_X2 inst_20307 ( .B2(net_19036), .B1(net_19035), .ZN(net_16066), .A(net_15753) );
OAI21_X2 inst_1543 ( .B1(net_18003), .ZN(net_17836), .B2(net_17608), .A(net_2526) );
INV_X4 inst_16954 ( .ZN(net_14764), .A(net_1000) );
INV_X4 inst_16214 ( .A(net_15366), .ZN(net_1915) );
CLKBUF_X2 inst_22960 ( .A(net_22831), .Z(net_22832) );
INV_X4 inst_13892 ( .ZN(net_11876), .A(net_4453) );
NAND2_X4 inst_7290 ( .A2(net_20211), .ZN(net_12035), .A1(net_5595) );
OR2_X4 inst_1118 ( .ZN(net_6433), .A1(net_602), .A2(net_151) );
INV_X4 inst_15341 ( .ZN(net_5789), .A(net_2596) );
NAND2_X4 inst_6978 ( .ZN(net_17490), .A2(net_16904), .A1(net_16714) );
NAND3_X2 inst_6109 ( .ZN(net_13893), .A3(net_13049), .A1(net_11412), .A2(net_9660) );
DFF_X1 inst_19901 ( .D(net_16987), .CK(net_21583), .Q(x659) );
INV_X4 inst_17768 ( .A(net_20851), .ZN(net_8304) );
NAND2_X2 inst_10948 ( .ZN(net_8333), .A1(net_5120), .A2(net_4967) );
XNOR2_X2 inst_473 ( .A(net_13655), .ZN(net_11889), .B(net_11888) );
AOI21_X2 inst_20275 ( .B1(net_21220), .ZN(net_20260), .B2(net_16082), .A(net_15543) );
INV_X4 inst_15114 ( .ZN(net_3489), .A(net_2382) );
NAND2_X2 inst_10140 ( .ZN(net_19551), .A1(net_13922), .A2(net_6956) );
INV_X4 inst_16258 ( .ZN(net_2099), .A(net_1364) );
INV_X4 inst_17303 ( .ZN(net_4874), .A(net_86) );
OAI21_X2 inst_2211 ( .A(net_14751), .ZN(net_8530), .B2(net_8529), .B1(net_6853) );
NOR2_X4 inst_3083 ( .ZN(net_5696), .A1(net_4383), .A2(net_4226) );
NAND2_X2 inst_9170 ( .ZN(net_13356), .A1(net_13355), .A2(net_10541) );
CLKBUF_X2 inst_22175 ( .A(net_21667), .Z(net_22047) );
INV_X4 inst_12609 ( .ZN(net_18085), .A(net_18080) );
INV_X4 inst_15336 ( .ZN(net_13984), .A(net_11380) );
NAND2_X2 inst_9917 ( .A2(net_10540), .ZN(net_9299), .A1(net_3633) );
INV_X4 inst_12942 ( .ZN(net_17123), .A(net_16789) );
AOI21_X2 inst_20553 ( .B1(net_19086), .ZN(net_14300), .A(net_11426), .B2(net_11258) );
INV_X2 inst_18821 ( .ZN(net_8335), .A(net_7302) );
INV_X4 inst_15371 ( .A(net_3829), .ZN(net_2570) );
NAND2_X2 inst_11034 ( .A1(net_8021), .ZN(net_5924), .A2(net_2570) );
OAI21_X4 inst_1404 ( .B2(net_19085), .B1(net_19084), .ZN(net_18925), .A(net_16368) );
NOR2_X4 inst_2989 ( .ZN(net_7477), .A1(net_5598), .A2(net_2563) );
NAND3_X2 inst_5880 ( .ZN(net_15282), .A3(net_14140), .A1(net_12318), .A2(net_2320) );
NOR2_X2 inst_3479 ( .ZN(net_14380), .A1(net_12998), .A2(net_12047) );
NOR2_X2 inst_4704 ( .A2(net_4150), .ZN(net_4126), .A1(net_3760) );
NOR2_X2 inst_3575 ( .ZN(net_12716), .A2(net_12328), .A1(net_11131) );
NAND2_X2 inst_9238 ( .ZN(net_12706), .A2(net_12705), .A1(net_3840) );
NOR2_X2 inst_4493 ( .A1(net_10714), .ZN(net_6618), .A2(net_2857) );
INV_X2 inst_19368 ( .ZN(net_2216), .A(net_1230) );
NAND2_X2 inst_8484 ( .ZN(net_16975), .A2(net_16974), .A1(net_16639) );
NAND2_X2 inst_10180 ( .ZN(net_13941), .A2(net_8191), .A1(net_5448) );
NAND2_X4 inst_7251 ( .ZN(net_10026), .A1(net_5121), .A2(net_3297) );
NAND3_X2 inst_5669 ( .ZN(net_16377), .A3(net_16180), .A2(net_15881), .A1(net_7668) );
INV_X4 inst_16556 ( .ZN(net_2380), .A(net_1057) );
NAND2_X2 inst_10941 ( .ZN(net_6284), .A2(net_5170), .A1(net_165) );
OAI21_X4 inst_1395 ( .A(net_16394), .ZN(net_16278), .B1(net_15989), .B2(net_15733) );
OAI211_X2 inst_2477 ( .ZN(net_13513), .C1(net_13512), .C2(net_12523), .A(net_10706), .B(net_1053) );
AOI21_X2 inst_20492 ( .ZN(net_14754), .B2(net_12288), .A(net_11089), .B1(net_2341) );
INV_X4 inst_14660 ( .ZN(net_18584), .A(net_18025) );
NAND4_X2 inst_5460 ( .A1(net_13490), .ZN(net_13332), .A2(net_13007), .A4(net_11638), .A3(net_8939) );
INV_X4 inst_17316 ( .A(net_3842), .ZN(net_1253) );
NAND2_X2 inst_11424 ( .ZN(net_8963), .A2(net_3819), .A1(net_3737) );
NAND2_X2 inst_8322 ( .A2(net_20583), .ZN(net_17559), .A1(net_17323) );
NOR2_X2 inst_4838 ( .ZN(net_2372), .A2(net_2371), .A1(net_1953) );
AOI22_X2 inst_19974 ( .ZN(net_15626), .A1(net_14709), .A2(net_14443), .B2(net_5676), .B1(net_60) );
OAI21_X2 inst_1875 ( .ZN(net_13694), .A(net_13693), .B2(net_10773), .B1(net_10292) );
NAND2_X2 inst_10005 ( .A1(net_13177), .ZN(net_8812), .A2(net_8811) );
NOR2_X4 inst_3190 ( .ZN(net_4448), .A2(net_2442), .A1(net_555) );
NAND2_X2 inst_8459 ( .ZN(net_17055), .A1(net_16824), .A2(net_16605) );
NAND2_X2 inst_10873 ( .A2(net_6437), .ZN(net_5428), .A1(net_2659) );
NOR2_X2 inst_3397 ( .ZN(net_19525), .A2(net_15491), .A1(net_15225) );
INV_X4 inst_13286 ( .ZN(net_12415), .A(net_12414) );
NAND4_X2 inst_5484 ( .A4(net_12992), .ZN(net_12472), .A2(net_12471), .A3(net_11757), .A1(net_7157) );
NAND2_X2 inst_11544 ( .A2(net_7397), .ZN(net_6484), .A1(net_1494) );
NOR2_X2 inst_4421 ( .ZN(net_6129), .A1(net_5205), .A2(net_3539) );
AOI21_X2 inst_20599 ( .ZN(net_19986), .B1(net_13703), .B2(net_13101), .A(net_7808) );
NAND2_X2 inst_8448 ( .A2(net_17330), .ZN(net_17102), .A1(net_17101) );
NOR2_X2 inst_4233 ( .ZN(net_6582), .A2(net_6581), .A1(net_5494) );
NAND2_X4 inst_7128 ( .ZN(net_12972), .A2(net_10319), .A1(net_9758) );
NAND3_X2 inst_5905 ( .ZN(net_15126), .A3(net_13390), .A2(net_10149), .A1(net_8289) );
NOR2_X2 inst_3968 ( .A1(net_10709), .ZN(net_8414), .A2(net_8413) );
INV_X4 inst_16535 ( .A(net_8067), .ZN(net_5576) );
NAND2_X2 inst_8208 ( .ZN(net_17862), .A2(net_17707), .A1(net_17612) );
INV_X2 inst_19023 ( .ZN(net_4938), .A(net_4937) );
INV_X4 inst_13010 ( .A(net_16590), .ZN(net_16436) );
NOR2_X2 inst_4633 ( .ZN(net_3527), .A1(net_2417), .A2(net_1256) );
INV_X4 inst_16349 ( .ZN(net_1398), .A(net_908) );
CLKBUF_X2 inst_21489 ( .A(net_21254), .Z(net_21361) );
NAND2_X2 inst_8113 ( .ZN(net_18103), .A2(net_18099), .A1(net_17487) );
INV_X4 inst_15845 ( .ZN(net_3933), .A(net_1835) );
INV_X4 inst_14871 ( .ZN(net_4654), .A(net_3693) );
NAND3_X2 inst_6660 ( .ZN(net_8452), .A2(net_7727), .A1(net_4888), .A3(net_4360) );
NAND2_X2 inst_10915 ( .ZN(net_5345), .A2(net_3874), .A1(net_86) );
NAND2_X2 inst_8027 ( .ZN(net_18268), .A2(net_18180), .A1(net_17281) );
NAND3_X2 inst_6411 ( .ZN(net_11955), .A2(net_9398), .A1(net_7086), .A3(net_6562) );
AOI21_X2 inst_20269 ( .A(net_20880), .B2(net_20326), .B1(net_20325), .ZN(net_18051) );
NAND2_X2 inst_9525 ( .A1(net_11612), .ZN(net_11123), .A2(net_7630) );
NAND2_X2 inst_8769 ( .ZN(net_15866), .A2(net_15641), .A1(net_15605) );
XNOR2_X2 inst_618 ( .B(net_17774), .ZN(net_484), .A(net_483) );
OAI211_X2 inst_2444 ( .ZN(net_14763), .C1(net_14600), .A(net_14402), .C2(net_11814), .B(net_8621) );
NAND2_X2 inst_11980 ( .ZN(net_1315), .A1(net_771), .A2(net_259) );
NOR2_X4 inst_3057 ( .ZN(net_8284), .A2(net_3627), .A1(net_2264) );
OAI211_X2 inst_2462 ( .C1(net_20550), .B(net_14331), .ZN(net_14148), .C2(net_9198), .A(net_7481) );
NAND3_X2 inst_6706 ( .ZN(net_12217), .A1(net_7455), .A3(net_4388), .A2(net_1058) );
XNOR2_X2 inst_474 ( .ZN(net_11885), .A(net_11884), .B(net_2432) );
INV_X2 inst_18865 ( .ZN(net_11234), .A(net_8867) );
NAND3_X4 inst_5561 ( .ZN(net_19101), .A2(net_15446), .A1(net_15310), .A3(net_14834) );
CLKBUF_X2 inst_22215 ( .A(net_22086), .Z(net_22087) );
AOI21_X2 inst_20657 ( .ZN(net_13033), .B1(net_13032), .A(net_12641), .B2(net_6543) );
XNOR2_X2 inst_626 ( .B(net_15585), .ZN(net_462), .A(net_461) );
CLKBUF_X2 inst_22169 ( .A(net_21990), .Z(net_22041) );
INV_X4 inst_15955 ( .ZN(net_15058), .A(net_10151) );
INV_X4 inst_15560 ( .ZN(net_15099), .A(net_8983) );
INV_X4 inst_14497 ( .ZN(net_6007), .A(net_4842) );
NAND2_X2 inst_11539 ( .A1(net_7968), .ZN(net_2920), .A2(net_2919) );
NAND2_X2 inst_9879 ( .ZN(net_9451), .A1(net_9450), .A2(net_7406) );
NAND2_X4 inst_7476 ( .ZN(net_4438), .A1(net_2697), .A2(net_1981) );
INV_X4 inst_18143 ( .A(net_21146), .ZN(net_16982) );
INV_X4 inst_16568 ( .A(net_5591), .ZN(net_4056) );
NAND2_X2 inst_10247 ( .ZN(net_13582), .A1(net_8014), .A2(net_1670) );
NAND2_X2 inst_8880 ( .ZN(net_15187), .A1(net_15186), .A2(net_14656) );
NAND2_X2 inst_11457 ( .ZN(net_12495), .A1(net_6617), .A2(net_3224) );
INV_X4 inst_12641 ( .ZN(net_17905), .A(net_17904) );
SDFF_X2 inst_798 ( .Q(net_20916), .SE(net_18577), .SI(net_17986), .D(net_528), .CK(net_21273) );
INV_X4 inst_12648 ( .ZN(net_17873), .A(net_17872) );
CLKBUF_X2 inst_22091 ( .A(net_21962), .Z(net_21963) );
INV_X4 inst_16382 ( .ZN(net_6041), .A(net_2264) );
INV_X4 inst_18215 ( .A(net_21231), .ZN(net_1790) );
INV_X4 inst_16838 ( .ZN(net_9310), .A(net_567) );
NOR2_X2 inst_4340 ( .ZN(net_5688), .A1(net_5687), .A2(net_4294) );
OAI21_X4 inst_1434 ( .B2(net_20685), .B1(net_20684), .A(net_16210), .ZN(net_15945) );
INV_X4 inst_12727 ( .ZN(net_20318), .A(net_17504) );
OAI21_X2 inst_1886 ( .ZN(net_13516), .B2(net_13515), .A(net_11060), .B1(net_1379) );
INV_X2 inst_18357 ( .ZN(net_18447), .A(net_18446) );
NAND2_X2 inst_10211 ( .ZN(net_12091), .A2(net_6278), .A1(net_1790) );
INV_X4 inst_16435 ( .ZN(net_12320), .A(net_10590) );
INV_X4 inst_12889 ( .A(net_16870), .ZN(net_16811) );
NAND2_X2 inst_8831 ( .ZN(net_15538), .A1(net_15537), .A2(net_15117) );
AOI21_X2 inst_20589 ( .ZN(net_13939), .A(net_13596), .B2(net_11288), .B1(net_3099) );
NAND2_X2 inst_8778 ( .ZN(net_15814), .A2(net_15358), .A1(net_14060) );
NOR2_X2 inst_4349 ( .ZN(net_5620), .A1(net_3845), .A2(net_2564) );
OAI21_X4 inst_1457 ( .B2(net_20171), .B1(net_20170), .ZN(net_15290), .A(net_15289) );
NAND2_X2 inst_8627 ( .A1(net_21157), .A2(net_16605), .ZN(net_16598) );
NAND2_X2 inst_10552 ( .ZN(net_8027), .A1(net_5950), .A2(net_4956) );
INV_X4 inst_16635 ( .ZN(net_6635), .A(net_86) );
AOI22_X2 inst_20016 ( .ZN(net_11335), .A1(net_8205), .A2(net_7619), .B1(net_5701), .B2(net_4117) );
INV_X4 inst_13244 ( .ZN(net_13191), .A(net_12227) );
NAND2_X2 inst_8209 ( .A2(net_19772), .A1(net_19771), .ZN(net_17861) );
NAND2_X2 inst_11254 ( .ZN(net_10429), .A2(net_4084), .A1(net_573) );
CLKBUF_X2 inst_22009 ( .A(net_21880), .Z(net_21881) );
NOR2_X2 inst_3662 ( .ZN(net_11583), .A1(net_11582), .A2(net_9787) );
INV_X4 inst_18117 ( .A(net_21225), .ZN(net_279) );
NOR3_X2 inst_2670 ( .ZN(net_14828), .A3(net_13471), .A2(net_5913), .A1(net_4168) );
INV_X4 inst_15726 ( .ZN(net_2761), .A(net_1459) );
NAND2_X2 inst_10983 ( .A2(net_5136), .ZN(net_4955), .A1(net_4481) );
NAND2_X2 inst_8380 ( .ZN(net_17345), .A2(net_17344), .A1(net_17059) );
NOR2_X4 inst_2974 ( .ZN(net_9465), .A1(net_5754), .A2(net_5698) );
INV_X4 inst_16965 ( .ZN(net_9994), .A(net_6631) );
OAI21_X2 inst_1895 ( .ZN(net_13363), .A(net_13362), .B2(net_9970), .B1(net_8433) );
NAND2_X2 inst_8476 ( .ZN(net_17012), .A2(net_17008), .A1(net_16788) );
NOR3_X2 inst_2730 ( .ZN(net_13185), .A2(net_13184), .A3(net_13183), .A1(net_7216) );
INV_X2 inst_19159 ( .ZN(net_3973), .A(net_3972) );
SDFF_X2 inst_737 ( .Q(net_20899), .SE(net_18856), .SI(net_18553), .D(net_649), .CK(net_22261) );
AOI21_X2 inst_20486 ( .ZN(net_20722), .B1(net_15362), .B2(net_13434), .A(net_10978) );
INV_X2 inst_19667 ( .ZN(net_20480), .A(net_20478) );
NAND2_X2 inst_11725 ( .ZN(net_2233), .A2(net_2232), .A1(net_1289) );
INV_X2 inst_19504 ( .ZN(net_1247), .A(net_1246) );
NAND2_X2 inst_11178 ( .ZN(net_8495), .A2(net_4112), .A1(net_2660) );
AOI21_X2 inst_20780 ( .B1(net_13310), .ZN(net_10560), .A(net_8524), .B2(net_6401) );
INV_X4 inst_16373 ( .A(net_4042), .ZN(net_1622) );
NAND2_X2 inst_8990 ( .ZN(net_14466), .A1(net_14465), .A2(net_12948) );
CLKBUF_X2 inst_22024 ( .A(net_21895), .Z(net_21896) );
XNOR2_X2 inst_545 ( .ZN(net_740), .A(net_739), .B(net_738) );
INV_X4 inst_16905 ( .ZN(net_1254), .A(net_420) );
INV_X4 inst_15819 ( .A(net_10386), .ZN(net_8338) );
NAND2_X2 inst_8373 ( .ZN(net_19395), .A1(net_17359), .A2(net_17358) );
DFF_X1 inst_19832 ( .D(net_17447), .CK(net_22546), .Q(x0) );
NAND2_X2 inst_10189 ( .ZN(net_8165), .A1(net_8164), .A2(net_8163) );
NAND2_X2 inst_8132 ( .ZN(net_18041), .A2(net_18029), .A1(net_18022) );
INV_X4 inst_17733 ( .ZN(net_4915), .A(net_4478) );
NAND2_X4 inst_6854 ( .A2(net_19947), .A1(net_19946), .ZN(net_18473) );
CLKBUF_X2 inst_21475 ( .A(net_21346), .Z(net_21347) );
INV_X4 inst_14475 ( .ZN(net_5764), .A(net_3403) );
INV_X8 inst_12188 ( .ZN(net_16727), .A(net_16439) );
NAND3_X2 inst_6682 ( .A2(net_7755), .ZN(net_7733), .A1(net_6429), .A3(net_3470) );
INV_X4 inst_13595 ( .ZN(net_8775), .A(net_7276) );
CLKBUF_X2 inst_21499 ( .A(net_21370), .Z(net_21371) );
NAND2_X2 inst_7832 ( .ZN(net_18636), .A2(net_18609), .A1(net_16775) );
NAND2_X2 inst_8624 ( .A1(net_19422), .ZN(net_16601), .A2(net_16415) );
NAND3_X2 inst_5878 ( .ZN(net_15284), .A1(net_14232), .A3(net_12502), .A2(net_6747) );
INV_X4 inst_14383 ( .A(net_10638), .ZN(net_5167) );
AOI21_X4 inst_20194 ( .ZN(net_19916), .B1(net_15088), .B2(net_13221), .A(net_13052) );
NAND2_X2 inst_8910 ( .ZN(net_14973), .A1(net_14972), .A2(net_13664) );
INV_X4 inst_13356 ( .ZN(net_10973), .A(net_10972) );
CLKBUF_X2 inst_21979 ( .A(net_21850), .Z(net_21851) );
NAND3_X2 inst_6573 ( .ZN(net_10463), .A2(net_10462), .A1(net_8038), .A3(net_7305) );
INV_X4 inst_13067 ( .ZN(net_16299), .A(net_16227) );
INV_X8 inst_12347 ( .ZN(net_928), .A(net_334) );
NAND2_X2 inst_10559 ( .A2(net_10950), .ZN(net_8670), .A1(net_6598) );
INV_X4 inst_13879 ( .ZN(net_10873), .A(net_7364) );
NOR2_X2 inst_4415 ( .A1(net_8007), .ZN(net_5036), .A2(net_5035) );
NOR2_X2 inst_4209 ( .A1(net_15374), .A2(net_13147), .ZN(net_6649) );
NAND2_X2 inst_10266 ( .A1(net_12440), .ZN(net_10192), .A2(net_6245) );
NAND3_X2 inst_6635 ( .ZN(net_8977), .A2(net_8976), .A3(net_8975), .A1(net_6941) );
CLKBUF_X2 inst_21957 ( .A(net_21454), .Z(net_21829) );
INV_X4 inst_15932 ( .ZN(net_2013), .A(net_1727) );
NAND2_X2 inst_10275 ( .ZN(net_7961), .A2(net_7960), .A1(net_6631) );
INV_X2 inst_18746 ( .ZN(net_7889), .A(net_7888) );
NAND2_X2 inst_8561 ( .A1(net_21189), .A2(net_20501), .ZN(net_16747) );
NAND2_X2 inst_8972 ( .ZN(net_14518), .A2(net_12865), .A1(net_11476) );
INV_X4 inst_16781 ( .ZN(net_9518), .A(net_238) );
DFF_X2 inst_19782 ( .QN(net_21105), .D(net_2455), .CK(net_21681) );
NAND2_X2 inst_12072 ( .ZN(net_1572), .A2(net_834), .A1(net_85) );
NAND3_X2 inst_5828 ( .ZN(net_15534), .A1(net_15124), .A3(net_14102), .A2(net_8835) );
NOR2_X2 inst_4260 ( .ZN(net_6244), .A2(net_6243), .A1(net_1091) );
NAND2_X2 inst_10218 ( .ZN(net_20269), .A2(net_8085), .A1(net_2448) );
NAND2_X2 inst_8072 ( .A2(net_18192), .ZN(net_18164), .A1(net_16867) );
NOR2_X2 inst_3484 ( .ZN(net_19869), .A1(net_12634), .A2(net_10004) );
INV_X4 inst_13868 ( .A(net_9476), .ZN(net_9118) );
SDFF_X2 inst_942 ( .QN(net_21010), .D(net_686), .SE(net_253), .CK(net_21902), .SI(x2881) );
NAND2_X2 inst_7755 ( .ZN(net_18790), .A2(net_18748), .A1(net_18727) );
NAND2_X2 inst_12077 ( .A2(net_1848), .ZN(net_1118), .A1(net_791) );
NAND2_X2 inst_8269 ( .A2(net_17683), .A1(net_17660), .ZN(net_17655) );
INV_X4 inst_13174 ( .ZN(net_14389), .A(net_13929) );
NAND3_X2 inst_6603 ( .A3(net_13320), .ZN(net_9880), .A2(net_7832), .A1(net_4929) );
AOI22_X2 inst_19967 ( .ZN(net_15850), .A2(net_15322), .B1(net_14865), .B2(net_12573), .A1(net_449) );
AOI21_X2 inst_20430 ( .ZN(net_15184), .B2(net_13902), .B1(net_11377), .A(net_3309) );
NAND2_X4 inst_7338 ( .ZN(net_4878), .A2(net_4396), .A1(net_663) );
NAND2_X4 inst_7353 ( .ZN(net_7873), .A2(net_5333), .A1(net_2744) );
NOR2_X2 inst_4501 ( .ZN(net_4254), .A1(net_4253), .A2(net_3231) );
INV_X2 inst_19225 ( .A(net_10444), .ZN(net_3440) );
NAND2_X4 inst_7144 ( .ZN(net_13307), .A2(net_9754), .A1(net_7591) );
NOR2_X2 inst_4252 ( .ZN(net_6359), .A1(net_6127), .A2(net_2620) );
NAND2_X2 inst_11758 ( .ZN(net_2849), .A2(net_2096), .A1(net_1380) );
AOI21_X2 inst_20951 ( .ZN(net_5749), .B1(net_5748), .A(net_4334), .B2(net_3161) );
NAND3_X2 inst_6356 ( .ZN(net_12092), .A3(net_12091), .A2(net_11805), .A1(net_11647) );
CLKBUF_X2 inst_22170 ( .A(net_21393), .Z(net_22042) );
NAND2_X2 inst_8258 ( .ZN(net_17694), .A1(net_17589), .A2(net_17408) );
INV_X2 inst_18728 ( .ZN(net_8065), .A(net_8064) );
NAND4_X2 inst_5451 ( .A2(net_20757), .A1(net_20756), .ZN(net_19694), .A4(net_7566), .A3(net_5657) );
AOI22_X2 inst_20034 ( .A1(net_10386), .ZN(net_8463), .B1(net_8462), .A2(net_6997), .B2(net_4670) );
INV_X4 inst_16929 ( .ZN(net_8836), .A(net_7260) );
INV_X4 inst_16124 ( .A(net_2846), .ZN(net_1484) );
NAND3_X2 inst_6393 ( .ZN(net_19521), .A2(net_11718), .A1(net_11276), .A3(net_9522) );
XNOR2_X2 inst_418 ( .A(net_16677), .ZN(net_16533), .B(net_14414) );
INV_X4 inst_17368 ( .ZN(net_14027), .A(net_60) );
NOR2_X2 inst_3961 ( .ZN(net_8591), .A2(net_6479), .A1(net_4287) );
INV_X2 inst_19155 ( .A(net_7093), .ZN(net_3994) );
CLKBUF_X2 inst_22851 ( .A(net_22722), .Z(net_22723) );
CLKBUF_X2 inst_22194 ( .A(net_21836), .Z(net_22066) );
NAND2_X2 inst_9526 ( .A1(net_11236), .ZN(net_11122), .A2(net_7626) );
NAND2_X2 inst_11851 ( .A2(net_9310), .A1(net_2348), .ZN(net_1694) );
NAND3_X2 inst_5871 ( .A2(net_20696), .A1(net_20695), .ZN(net_20112), .A3(net_12828) );
NAND2_X2 inst_10016 ( .ZN(net_13335), .A2(net_8154), .A1(net_6867) );
AOI21_X2 inst_20666 ( .B1(net_13375), .ZN(net_12921), .A(net_11315), .B2(net_9270) );
INV_X4 inst_16241 ( .ZN(net_4088), .A(net_1826) );
INV_X4 inst_13957 ( .ZN(net_8060), .A(net_5473) );
OR2_X2 inst_1177 ( .A1(net_15375), .ZN(net_5377), .A2(net_5376) );
OAI211_X2 inst_2548 ( .ZN(net_10821), .A(net_5648), .C2(net_4639), .B(net_3270), .C1(net_2174) );
NAND2_X2 inst_11494 ( .ZN(net_11363), .A2(net_3087), .A1(net_90) );
NOR2_X2 inst_5127 ( .ZN(net_266), .A2(net_265), .A1(net_74) );
NAND2_X2 inst_8022 ( .ZN(net_19949), .A1(net_18405), .A2(net_18260) );
INV_X4 inst_12587 ( .A(net_18166), .ZN(net_18134) );
NAND2_X2 inst_9051 ( .A1(net_19859), .ZN(net_14013), .A2(net_10031) );
OAI21_X2 inst_1666 ( .B1(net_19580), .ZN(net_19140), .B2(net_15690), .A(net_12192) );
INV_X4 inst_17916 ( .ZN(net_14714), .A(net_10216) );
SDFF_X2 inst_735 ( .Q(net_20942), .SE(net_18581), .SI(net_18558), .D(net_3755), .CK(net_22757) );
CLKBUF_X2 inst_22796 ( .A(net_22667), .Z(net_22668) );
OAI21_X2 inst_1529 ( .ZN(net_18005), .B2(net_17899), .A(net_1281), .B1(net_253) );
INV_X2 inst_18992 ( .A(net_6842), .ZN(net_5085) );
INV_X4 inst_16798 ( .ZN(net_15468), .A(net_11032) );
INV_X8 inst_12445 ( .ZN(net_20508), .A(net_17110) );
NAND2_X2 inst_10426 ( .ZN(net_12932), .A2(net_7221), .A1(net_2344) );
NAND2_X2 inst_7890 ( .ZN(net_18506), .A2(net_18444), .A1(net_18397) );
OAI21_X2 inst_1653 ( .B2(net_20193), .B1(net_20192), .ZN(net_18880), .A(net_9656) );
CLKBUF_X2 inst_22141 ( .A(net_22012), .Z(net_22013) );
INV_X4 inst_17230 ( .ZN(net_19537), .A(net_699) );
AOI21_X2 inst_20647 ( .ZN(net_13071), .B1(net_13070), .B2(net_12870), .A(net_11107) );
INV_X2 inst_18777 ( .ZN(net_10639), .A(net_7690) );
INV_X4 inst_13376 ( .ZN(net_10877), .A(net_10876) );
NAND2_X4 inst_7220 ( .ZN(net_9104), .A1(net_7393), .A2(net_6314) );
AOI21_X2 inst_20739 ( .A(net_12401), .ZN(net_11436), .B2(net_11435), .B1(net_4414) );
INV_X4 inst_18052 ( .A(net_20961), .ZN(net_862) );
NAND2_X2 inst_11627 ( .ZN(net_3031), .A1(net_2557), .A2(net_2519) );
NOR2_X4 inst_2984 ( .A2(net_20859), .ZN(net_9743), .A1(net_4583) );
NOR2_X4 inst_3258 ( .ZN(net_4157), .A2(net_2241), .A1(net_1645) );
INV_X4 inst_13002 ( .ZN(net_17048), .A(net_16902) );
NAND2_X1 inst_12150 ( .A1(net_13192), .ZN(net_10612), .A2(net_7257) );
INV_X2 inst_19250 ( .A(net_4024), .ZN(net_3257) );
OAI21_X2 inst_1805 ( .A(net_15156), .ZN(net_14475), .B2(net_11648), .B1(net_8562) );
NOR2_X2 inst_3563 ( .ZN(net_12918), .A2(net_11156), .A1(net_4488) );
INV_X4 inst_18339 ( .ZN(net_20708), .A(net_16485) );
INV_X4 inst_16628 ( .ZN(net_8854), .A(net_1111) );
NAND2_X2 inst_9675 ( .ZN(net_14296), .A1(net_13023), .A2(net_8174) );
INV_X4 inst_16088 ( .ZN(net_2739), .A(net_1467) );
NAND2_X2 inst_8231 ( .ZN(net_17791), .A2(net_17666), .A1(net_17398) );
NAND2_X2 inst_8936 ( .ZN(net_14849), .A2(net_14182), .A1(net_4690) );
NOR3_X2 inst_2752 ( .A3(net_15280), .ZN(net_11988), .A2(net_8602), .A1(net_3445) );
NAND2_X2 inst_10095 ( .ZN(net_13179), .A1(net_8616), .A2(net_7879) );
INV_X4 inst_16140 ( .ZN(net_2522), .A(net_1104) );
OAI22_X2 inst_1281 ( .ZN(net_15368), .A2(net_13909), .B2(net_12806), .A1(net_4452), .B1(net_4384) );
INV_X2 inst_19032 ( .ZN(net_4882), .A(net_4881) );
OAI21_X2 inst_1509 ( .ZN(net_18861), .B2(net_18843), .B1(net_18025), .A(net_7390) );
NOR2_X4 inst_3088 ( .ZN(net_6616), .A2(net_4027), .A1(net_1255) );
NAND2_X2 inst_10386 ( .A1(net_15224), .ZN(net_10746), .A2(net_5610) );
NAND2_X2 inst_9000 ( .ZN(net_14288), .A2(net_13482), .A1(net_11384) );
INV_X4 inst_15858 ( .ZN(net_14055), .A(net_11572) );
NOR2_X2 inst_3782 ( .ZN(net_10125), .A2(net_7974), .A1(net_5414) );
INV_X4 inst_15754 ( .A(net_8485), .ZN(net_5149) );
NAND2_X4 inst_7486 ( .A2(net_19418), .ZN(net_2461), .A1(net_218) );
INV_X4 inst_15101 ( .ZN(net_12419), .A(net_10231) );
INV_X4 inst_15466 ( .ZN(net_3344), .A(net_3110) );
NAND3_X2 inst_6630 ( .A3(net_19858), .ZN(net_19720), .A1(net_8758), .A2(net_6926) );
INV_X4 inst_15378 ( .ZN(net_14337), .A(net_2565) );
CLKBUF_X2 inst_22293 ( .A(net_22101), .Z(net_22165) );
NAND2_X2 inst_8054 ( .A1(net_19956), .ZN(net_18212), .A2(net_18211) );
NAND3_X2 inst_5809 ( .ZN(net_15655), .A3(net_14870), .A2(net_9233), .A1(net_8582) );
OR2_X2 inst_1140 ( .ZN(net_19362), .A2(net_11479), .A1(net_9180) );
AOI211_X2 inst_21036 ( .ZN(net_14144), .C2(net_10772), .C1(net_8473), .B(net_7128), .A(net_6022) );
INV_X4 inst_15637 ( .ZN(net_2806), .A(net_2546) );
INV_X2 inst_19696 ( .A(net_20551), .ZN(net_20550) );
AOI21_X2 inst_20559 ( .ZN(net_14267), .B2(net_12416), .B1(net_7700), .A(net_2371) );
NAND2_X2 inst_9251 ( .A1(net_13659), .ZN(net_12664), .A2(net_7895) );
NAND3_X2 inst_6140 ( .A3(net_19632), .ZN(net_13715), .A2(net_13472), .A1(net_12636) );
OAI21_X2 inst_1800 ( .ZN(net_14484), .A(net_14483), .B2(net_12521), .B1(net_8428) );
NOR2_X2 inst_4773 ( .ZN(net_3690), .A1(net_1772), .A2(net_1703) );
NAND2_X2 inst_8463 ( .A2(net_20498), .ZN(net_17050), .A1(net_16820) );
NAND2_X2 inst_11087 ( .ZN(net_4395), .A1(net_4394), .A2(net_2168) );
XNOR2_X2 inst_448 ( .ZN(net_14911), .B(net_14910), .A(net_12874) );
AOI21_X2 inst_20374 ( .ZN(net_15603), .B1(net_15602), .B2(net_14256), .A(net_4238) );
NAND3_X2 inst_5966 ( .ZN(net_14777), .A3(net_13419), .A2(net_13354), .A1(net_12699) );
NAND3_X2 inst_5680 ( .A3(net_19791), .A1(net_19790), .ZN(net_16331), .A2(net_12756) );
DFF_X1 inst_19813 ( .QN(net_21201), .D(net_17976), .CK(net_21444) );
NAND2_X2 inst_10253 ( .ZN(net_8001), .A2(net_6085), .A1(net_5017) );
NAND3_X2 inst_6056 ( .ZN(net_14224), .A2(net_14211), .A3(net_13610), .A1(net_13432) );
NOR2_X2 inst_4921 ( .ZN(net_3548), .A1(net_2493), .A2(net_1933) );
INV_X4 inst_14367 ( .ZN(net_6305), .A(net_5202) );
CLKBUF_X2 inst_21631 ( .A(net_21319), .Z(net_21503) );
AND2_X4 inst_21175 ( .ZN(net_20326), .A1(net_12194), .A2(net_12193) );
NAND2_X2 inst_9374 ( .ZN(net_12014), .A2(net_12013), .A1(net_4714) );
CLKBUF_X2 inst_21498 ( .A(net_21369), .Z(net_21370) );
NAND2_X2 inst_10862 ( .ZN(net_11819), .A1(net_11472), .A2(net_5437) );
NAND2_X2 inst_10053 ( .A1(net_13418), .ZN(net_8691), .A2(net_6819) );
INV_X4 inst_16072 ( .ZN(net_2975), .A(net_2278) );
INV_X2 inst_18624 ( .ZN(net_9561), .A(net_9560) );
INV_X4 inst_13017 ( .ZN(net_16492), .A(net_16425) );
NAND2_X2 inst_8212 ( .ZN(net_19301), .A2(net_17784), .A1(net_17268) );
OAI221_X2 inst_1343 ( .ZN(net_13459), .C2(net_13458), .C1(net_13198), .A(net_7362), .B1(net_5415), .B2(net_5307) );
NAND2_X2 inst_9068 ( .ZN(net_13979), .A2(net_12201), .A1(net_10073) );
NAND2_X2 inst_8050 ( .ZN(net_18261), .A1(net_18159), .A2(net_18133) );
CLKBUF_X2 inst_21737 ( .A(net_21250), .Z(net_21609) );
AOI21_X2 inst_20909 ( .B1(net_11702), .B2(net_10246), .A(net_8959), .ZN(net_7375) );
INV_X4 inst_16133 ( .ZN(net_15026), .A(net_1046) );
NAND2_X4 inst_7536 ( .ZN(net_1945), .A1(net_817), .A2(net_106) );
NOR2_X2 inst_4054 ( .ZN(net_10218), .A2(net_6566), .A1(net_6207) );
NAND2_X2 inst_7813 ( .ZN(net_18713), .A1(net_18641), .A2(net_18630) );
NAND3_X2 inst_6713 ( .ZN(net_7101), .A2(net_4214), .A3(net_4063), .A1(net_3893) );
OR2_X2 inst_1246 ( .ZN(net_8556), .A1(net_2673), .A2(net_119) );
NOR2_X4 inst_3185 ( .ZN(net_5590), .A1(net_2836), .A2(net_222) );
INV_X4 inst_17419 ( .ZN(net_3284), .A(net_143) );
NOR2_X2 inst_4679 ( .ZN(net_5384), .A2(net_3013), .A1(net_1376) );
CLKBUF_X2 inst_22467 ( .A(net_21373), .Z(net_22339) );
AOI21_X2 inst_20783 ( .B1(net_20406), .ZN(net_10555), .B2(net_9324), .A(net_5661) );
NAND2_X2 inst_11699 ( .ZN(net_3884), .A2(net_2073), .A1(net_1376) );
NAND2_X2 inst_11269 ( .ZN(net_3892), .A2(net_2106), .A1(net_955) );
CLKBUF_X2 inst_22895 ( .A(net_22766), .Z(net_22767) );
CLKBUF_X2 inst_22666 ( .A(net_22537), .Z(net_22538) );
INV_X4 inst_13163 ( .ZN(net_14811), .A(net_14230) );
CLKBUF_X2 inst_22183 ( .A(net_21863), .Z(net_22055) );
INV_X4 inst_15881 ( .ZN(net_2687), .A(net_1781) );
NAND3_X2 inst_5647 ( .A3(net_20357), .A1(net_20356), .ZN(net_16895), .A2(net_16362) );
CLKBUF_X2 inst_22225 ( .A(net_22096), .Z(net_22097) );
NAND2_X2 inst_10623 ( .A1(net_9666), .ZN(net_6565), .A2(net_6564) );
NAND3_X4 inst_5580 ( .A3(net_19728), .A1(net_19727), .ZN(net_19637), .A2(net_15598) );
INV_X8 inst_12180 ( .ZN(net_19982), .A(net_16553) );
INV_X4 inst_16351 ( .ZN(net_1295), .A(net_1288) );
NAND2_X2 inst_8568 ( .ZN(net_16740), .A2(net_16588), .A1(net_16516) );
OAI21_X2 inst_2029 ( .ZN(net_11313), .A(net_8455), .B2(net_7608), .B1(net_5480) );
INV_X4 inst_17298 ( .A(net_4288), .ZN(net_4253) );
NAND2_X2 inst_10632 ( .ZN(net_8113), .A2(net_6443), .A1(net_2828) );
INV_X4 inst_12812 ( .ZN(net_17205), .A(net_17204) );
NAND2_X2 inst_8779 ( .ZN(net_15809), .A2(net_15282), .A1(net_1411) );
NOR2_X2 inst_4936 ( .ZN(net_2200), .A2(net_1226), .A1(net_170) );
INV_X4 inst_15037 ( .A(net_3353), .ZN(net_3346) );
CLKBUF_X2 inst_21781 ( .A(net_21381), .Z(net_21653) );
INV_X4 inst_16528 ( .A(net_6924), .ZN(net_6092) );
AOI21_X2 inst_20858 ( .A(net_11443), .ZN(net_8902), .B2(net_8901), .B1(net_4622) );
CLKBUF_X2 inst_21694 ( .A(net_21565), .Z(net_21566) );
INV_X2 inst_18784 ( .A(net_9532), .ZN(net_7502) );
OAI21_X2 inst_1965 ( .A(net_14593), .ZN(net_12302), .B1(net_8564), .B2(net_7306) );
INV_X4 inst_16033 ( .ZN(net_2295), .A(net_1795) );
NOR2_X2 inst_3915 ( .A2(net_14544), .ZN(net_10303), .A1(net_3170) );
NAND4_X2 inst_5419 ( .ZN(net_14426), .A4(net_12437), .A1(net_11393), .A2(net_9410), .A3(net_2619) );
NAND2_X2 inst_8144 ( .A2(net_20129), .A1(net_20128), .ZN(net_18021) );
NAND3_X2 inst_5743 ( .A3(net_20160), .A1(net_20159), .A2(net_19231), .ZN(net_18930) );
INV_X2 inst_19127 ( .ZN(net_4298), .A(net_4297) );
NAND4_X2 inst_5422 ( .ZN(net_14244), .A4(net_13600), .A2(net_7829), .A3(net_6627), .A1(net_4131) );
INV_X2 inst_18913 ( .A(net_9954), .ZN(net_6016) );
CLKBUF_X2 inst_21916 ( .A(net_21509), .Z(net_21788) );
INV_X4 inst_15785 ( .ZN(net_12763), .A(net_12708) );
NOR2_X4 inst_3285 ( .A2(net_1981), .ZN(net_1557), .A1(net_1556) );
AND2_X4 inst_21216 ( .A2(net_11255), .A1(net_10389), .ZN(net_6296) );
NAND2_X4 inst_6948 ( .ZN(net_20464), .A1(net_17182), .A2(net_17056) );
NAND3_X2 inst_6492 ( .ZN(net_11163), .A2(net_11162), .A3(net_11161), .A1(net_5807) );
INV_X2 inst_19234 ( .ZN(net_3354), .A(net_3353) );
INV_X4 inst_14091 ( .ZN(net_7560), .A(net_4633) );
INV_X4 inst_14934 ( .ZN(net_5933), .A(net_4849) );
NAND2_X2 inst_11931 ( .A1(net_20875), .ZN(net_2474), .A2(net_1487) );
NAND2_X2 inst_11790 ( .A1(net_4030), .A2(net_2066), .ZN(net_1967) );
NAND2_X2 inst_11568 ( .A1(net_4511), .ZN(net_2790), .A2(net_2735) );
NOR2_X2 inst_4460 ( .ZN(net_4618), .A2(net_4529), .A1(net_2587) );
INV_X4 inst_18046 ( .A(net_21053), .ZN(net_616) );
NAND2_X2 inst_8336 ( .ZN(net_17514), .A1(net_17513), .A2(net_17512) );
INV_X4 inst_12559 ( .ZN(net_18360), .A(net_18273) );
NAND2_X2 inst_11681 ( .A2(net_5285), .ZN(net_4347), .A1(net_2344) );
NAND2_X4 inst_7002 ( .ZN(net_17374), .A1(net_16713), .A2(net_16712) );
NOR2_X4 inst_2804 ( .ZN(net_18247), .A1(net_18149), .A2(net_18148) );
NOR2_X2 inst_5131 ( .A2(net_396), .ZN(net_224), .A1(net_221) );
CLKBUF_X2 inst_22245 ( .A(net_22116), .Z(net_22117) );
AOI211_X2 inst_21079 ( .ZN(net_6396), .B(net_4747), .A(net_3413), .C1(net_1985), .C2(net_1905) );
SDFF_X2 inst_772 ( .Q(net_20962), .SE(net_18576), .SI(net_18487), .D(net_687), .CK(net_21246) );
NAND3_X2 inst_6738 ( .A3(net_10837), .ZN(net_6465), .A1(net_6464), .A2(net_4870) );
NOR2_X2 inst_3682 ( .ZN(net_11423), .A1(net_11422), .A2(net_10124) );
NOR2_X2 inst_4940 ( .ZN(net_2967), .A1(net_2221), .A2(net_1535) );
NOR2_X2 inst_4583 ( .ZN(net_6572), .A1(net_3823), .A2(net_168) );
INV_X4 inst_13282 ( .ZN(net_12435), .A(net_11163) );
INV_X4 inst_15141 ( .ZN(net_5451), .A(net_3114) );
NAND2_X2 inst_10525 ( .ZN(net_8937), .A2(net_6846), .A1(net_1103) );
INV_X4 inst_14396 ( .ZN(net_12640), .A(net_5121) );
NOR2_X2 inst_4870 ( .ZN(net_2906), .A1(net_1500), .A2(net_546) );
NAND4_X2 inst_5454 ( .ZN(net_13455), .A3(net_10644), .A4(net_8801), .A1(net_8177), .A2(net_6576) );
INV_X4 inst_17047 ( .ZN(net_1160), .A(net_131) );
NAND3_X2 inst_6224 ( .ZN(net_13237), .A3(net_13129), .A1(net_8425), .A2(net_6638) );
AND2_X4 inst_21194 ( .ZN(net_10380), .A1(net_10379), .A2(net_7762) );
NAND3_X2 inst_6761 ( .ZN(net_10364), .A1(net_9146), .A3(net_5579), .A2(net_1033) );
XNOR2_X2 inst_606 ( .B(net_16599), .ZN(net_519), .A(net_518) );
NOR2_X4 inst_2942 ( .A2(net_20548), .ZN(net_8303), .A1(net_6926) );
NAND2_X2 inst_9929 ( .ZN(net_9184), .A1(net_9183), .A2(net_5841) );
INV_X4 inst_16496 ( .ZN(net_3244), .A(net_2007) );
INV_X4 inst_13875 ( .ZN(net_19617), .A(net_9838) );
NAND2_X2 inst_10287 ( .ZN(net_7934), .A2(net_5897), .A1(net_1478) );
NAND2_X2 inst_8167 ( .ZN(net_17963), .A1(net_17962), .A2(net_17961) );
XNOR2_X2 inst_139 ( .A(net_20505), .ZN(net_18181), .B(net_9194) );
INV_X4 inst_13767 ( .A(net_12612), .ZN(net_7605) );
INV_X4 inst_15813 ( .ZN(net_12669), .A(net_10765) );
NAND2_X2 inst_10856 ( .ZN(net_7272), .A1(net_5454), .A2(net_4263) );
NAND2_X2 inst_8903 ( .ZN(net_15061), .A2(net_13987), .A1(net_10832) );
INV_X4 inst_12548 ( .ZN(net_18286), .A(net_18285) );
OAI22_X2 inst_1316 ( .B1(net_8138), .ZN(net_5777), .A1(net_5776), .B2(net_5775), .A2(net_3508) );
CLKBUF_X2 inst_22020 ( .A(net_21891), .Z(net_21892) );
CLKBUF_X2 inst_21396 ( .A(net_21252), .Z(net_21268) );
NAND2_X2 inst_8400 ( .ZN(net_17388), .A2(net_16958), .A1(net_16796) );
NOR2_X2 inst_3551 ( .ZN(net_13083), .A1(net_13082), .A2(net_13081) );
NAND3_X4 inst_5528 ( .A3(net_20669), .A1(net_20668), .ZN(net_17777), .A2(net_16126) );
INV_X2 inst_18504 ( .ZN(net_11991), .A(net_10566) );
NAND3_X2 inst_6521 ( .ZN(net_19533), .A1(net_10636), .A2(net_10635), .A3(net_10634) );
AOI21_X2 inst_20984 ( .A(net_664), .ZN(net_455), .B2(net_26), .B1(net_25) );
XNOR2_X2 inst_191 ( .B(net_21137), .ZN(net_17682), .A(net_17681) );
INV_X4 inst_16552 ( .ZN(net_9681), .A(net_1209) );
NAND2_X2 inst_8908 ( .ZN(net_19799), .A2(net_13670), .A1(net_11786) );
NAND2_X2 inst_9328 ( .A1(net_14496), .ZN(net_12304), .A2(net_10661) );
INV_X4 inst_13485 ( .ZN(net_19524), .A(net_11849) );
NOR2_X2 inst_4538 ( .A2(net_4066), .ZN(net_4021), .A1(net_4020) );
NAND4_X4 inst_5212 ( .ZN(net_16425), .A4(net_16206), .A2(net_16146), .A1(net_16074), .A3(net_15791) );
INV_X4 inst_13988 ( .ZN(net_7798), .A(net_5345) );
AND3_X2 inst_21145 ( .ZN(net_7735), .A3(net_5853), .A2(net_5292), .A1(net_2987) );
CLKBUF_X2 inst_22787 ( .A(net_22658), .Z(net_22659) );
INV_X4 inst_18279 ( .ZN(net_20071), .A(net_20069) );
NAND2_X4 inst_6892 ( .A2(net_18070), .ZN(net_18060), .A1(net_16013) );
AOI21_X4 inst_20208 ( .B1(net_20839), .ZN(net_14574), .A(net_12589), .B2(net_278) );
NOR2_X2 inst_3879 ( .ZN(net_10869), .A2(net_9320), .A1(net_731) );
NAND4_X2 inst_5269 ( .A4(net_18962), .A1(net_18961), .ZN(net_16139), .A3(net_15192), .A2(net_14329) );
AND4_X2 inst_21098 ( .ZN(net_13461), .A1(net_13460), .A4(net_13150), .A3(net_12787), .A2(net_8536) );
CLKBUF_X2 inst_22634 ( .A(net_22505), .Z(net_22506) );
AND2_X4 inst_21237 ( .ZN(net_8800), .A2(net_5284), .A1(net_4715) );
INV_X2 inst_19143 ( .ZN(net_4103), .A(net_4102) );
NAND3_X2 inst_6544 ( .A3(net_12126), .A2(net_11964), .ZN(net_10564), .A1(net_5796) );
INV_X8 inst_12201 ( .ZN(net_11504), .A(net_9593) );
OAI21_X2 inst_2184 ( .A(net_11389), .ZN(net_8834), .B2(net_4960), .B1(net_4087) );
INV_X4 inst_13296 ( .ZN(net_12349), .A(net_12348) );
INV_X2 inst_19723 ( .A(net_20790), .ZN(net_20789) );
NOR3_X2 inst_2665 ( .ZN(net_14988), .A3(net_12811), .A1(net_11633), .A2(net_11211) );
OR2_X2 inst_1132 ( .ZN(net_14290), .A1(net_14289), .A2(net_12619) );
INV_X4 inst_14415 ( .A(net_13472), .ZN(net_6211) );
INV_X4 inst_17619 ( .ZN(net_445), .A(net_129) );
SDFF_X2 inst_968 ( .QN(net_21007), .D(net_2403), .SE(net_263), .CK(net_21846), .SI(x2957) );
NOR2_X2 inst_4700 ( .ZN(net_4141), .A2(net_3172), .A1(net_1020) );
INV_X4 inst_13531 ( .ZN(net_11532), .A(net_9222) );
NOR2_X2 inst_4441 ( .ZN(net_4808), .A2(net_4807), .A1(net_961) );
INV_X2 inst_19213 ( .A(net_4798), .ZN(net_3488) );
INV_X4 inst_15024 ( .A(net_4989), .ZN(net_4584) );
AOI221_X2 inst_20075 ( .ZN(net_19339), .B1(net_16281), .C1(net_16054), .C2(net_15802), .B2(net_13698), .A(net_5316) );
INV_X2 inst_19512 ( .A(net_1921), .ZN(net_1183) );
NOR2_X4 inst_3153 ( .ZN(net_4051), .A1(net_3311), .A2(net_1230) );
NAND3_X2 inst_6076 ( .ZN(net_20059), .A2(net_14092), .A3(net_12972), .A1(net_12294) );
INV_X4 inst_14357 ( .ZN(net_5998), .A(net_5254) );
NAND2_X2 inst_11990 ( .ZN(net_2309), .A2(net_1329), .A1(net_1044) );
NOR2_X2 inst_4004 ( .ZN(net_8110), .A2(net_8109), .A1(net_3874) );
INV_X4 inst_12708 ( .ZN(net_17568), .A(net_17567) );
CLKBUF_X2 inst_21690 ( .A(net_21561), .Z(net_21562) );
INV_X4 inst_15352 ( .A(net_14472), .ZN(net_14465) );
INV_X2 inst_18513 ( .A(net_14542), .ZN(net_11578) );
INV_X4 inst_17312 ( .ZN(net_7260), .A(net_1020) );
NAND2_X2 inst_11838 ( .A1(net_10183), .A2(net_2744), .ZN(net_1739) );
NAND2_X2 inst_8887 ( .ZN(net_15145), .A2(net_14097), .A1(net_5736) );
NOR2_X2 inst_3798 ( .ZN(net_9882), .A1(net_6868), .A2(net_6605) );
INV_X4 inst_18137 ( .A(net_21132), .ZN(net_16794) );
NAND4_X4 inst_5232 ( .A4(net_19265), .A1(net_19264), .ZN(net_18901), .A3(net_13757), .A2(net_11228) );
NOR2_X2 inst_4109 ( .ZN(net_7089), .A2(net_6641), .A1(net_4130) );
INV_X2 inst_19449 ( .ZN(net_2166), .A(net_1189) );
NOR2_X2 inst_4192 ( .ZN(net_8008), .A2(net_6725), .A1(net_154) );
NAND2_X2 inst_10048 ( .ZN(net_8698), .A1(net_8697), .A2(net_8696) );
NOR2_X4 inst_3004 ( .A1(net_9692), .ZN(net_7876), .A2(net_3187) );
INV_X8 inst_12396 ( .A(net_220), .ZN(net_160) );
NOR2_X2 inst_4672 ( .ZN(net_5371), .A2(net_3947), .A1(net_3019) );
INV_X4 inst_14438 ( .ZN(net_6159), .A(net_4998) );
INV_X8 inst_12363 ( .ZN(net_2094), .A(net_195) );
INV_X4 inst_17355 ( .ZN(net_3063), .A(net_115) );
INV_X4 inst_17024 ( .ZN(net_11511), .A(net_904) );
OAI211_X2 inst_2456 ( .ZN(net_14317), .B(net_14316), .C1(net_14315), .C2(net_14314), .A(net_13621) );
NOR2_X4 inst_2887 ( .A1(net_20100), .ZN(net_11038), .A2(net_9667) );
NAND2_X1 inst_12162 ( .A1(net_6207), .A2(net_3836), .ZN(net_2362) );
NAND2_X2 inst_11120 ( .A1(net_20574), .ZN(net_8976), .A2(net_4302) );
INV_X2 inst_18655 ( .A(net_11020), .ZN(net_9214) );
INV_X4 inst_16972 ( .ZN(net_6712), .A(net_3748) );
NAND2_X2 inst_8805 ( .ZN(net_19085), .A1(net_15567), .A2(net_15354) );
OAI21_X4 inst_1473 ( .B2(net_19544), .B1(net_19543), .ZN(net_18929), .A(net_14308) );
CLKBUF_X2 inst_22157 ( .A(net_22028), .Z(net_22029) );
NAND4_X2 inst_5334 ( .A2(net_19587), .A1(net_19586), .ZN(net_15535), .A4(net_14698), .A3(net_13056) );
INV_X4 inst_12793 ( .ZN(net_17273), .A(net_17272) );
NAND2_X2 inst_9306 ( .ZN(net_12375), .A1(net_10920), .A2(net_9116) );
INV_X4 inst_16248 ( .ZN(net_4457), .A(net_2994) );
INV_X4 inst_18099 ( .A(net_20869), .ZN(net_938) );
XNOR2_X2 inst_632 ( .B(net_16833), .ZN(net_7648), .A(net_634) );
INV_X2 inst_18435 ( .ZN(net_19704), .A(net_13906) );
XOR2_X2 inst_0 ( .B(net_21157), .Z(net_18676), .A(net_18628) );
INV_X4 inst_13934 ( .ZN(net_12902), .A(net_6844) );
AND2_X4 inst_21203 ( .ZN(net_11560), .A2(net_8044), .A1(net_7950) );
INV_X4 inst_17242 ( .A(net_2183), .ZN(net_1547) );
INV_X2 inst_19582 ( .ZN(net_964), .A(net_183) );
NAND2_X2 inst_11405 ( .ZN(net_6231), .A1(net_4221), .A2(net_1073) );
INV_X4 inst_14582 ( .A(net_6509), .ZN(net_4499) );
NAND2_X2 inst_11199 ( .ZN(net_5155), .A2(net_4862), .A1(net_4075) );
AOI211_X2 inst_20996 ( .C1(net_21220), .ZN(net_16255), .C2(net_15943), .B(net_10316), .A(net_6593) );
INV_X8 inst_12266 ( .ZN(net_2810), .A(net_1457) );
NAND2_X2 inst_8994 ( .ZN(net_14447), .A2(net_13136), .A1(net_7165) );
AOI21_X4 inst_20099 ( .B1(net_20694), .ZN(net_18927), .B2(net_16390), .A(net_16251) );
INV_X4 inst_13520 ( .ZN(net_9352), .A(net_9351) );
OAI21_X2 inst_1983 ( .ZN(net_12071), .A(net_12070), .B2(net_12069), .B1(net_5182) );
INV_X4 inst_13748 ( .ZN(net_10208), .A(net_9578) );
NAND2_X4 inst_7323 ( .A2(net_20554), .ZN(net_6247), .A1(net_4371) );
CLKBUF_X2 inst_21430 ( .A(net_21301), .Z(net_21302) );
AOI21_X2 inst_20342 ( .B1(net_16127), .ZN(net_15764), .B2(net_14775), .A(net_13108) );
INV_X4 inst_17343 ( .ZN(net_1016), .A(net_937) );
OAI21_X2 inst_1948 ( .A(net_12638), .ZN(net_12581), .B2(net_12525), .B1(net_2238) );
NAND2_X4 inst_7158 ( .A1(net_11465), .ZN(net_10972), .A2(net_9540) );
NAND2_X2 inst_8409 ( .ZN(net_19044), .A2(net_17235), .A1(net_16688) );
INV_X2 inst_19346 ( .A(net_2674), .ZN(net_2427) );
INV_X4 inst_15148 ( .ZN(net_9493), .A(net_3077) );
NAND2_X2 inst_8266 ( .A2(net_17683), .ZN(net_17659), .A1(net_17658) );
XNOR2_X2 inst_422 ( .ZN(net_16507), .A(net_16506), .B(net_1516) );
INV_X4 inst_16281 ( .A(net_9324), .ZN(net_8865) );
AOI21_X2 inst_20621 ( .A(net_15166), .ZN(net_13489), .B2(net_9012), .B1(net_7855) );
OAI21_X2 inst_2243 ( .ZN(net_7377), .B1(net_5797), .A(net_4546), .B2(net_2787) );
CLKBUF_X2 inst_22095 ( .A(net_21842), .Z(net_21967) );
OAI21_X4 inst_1426 ( .ZN(net_19274), .B1(net_16030), .A(net_15629), .B2(net_15476) );
NAND2_X2 inst_9021 ( .A1(net_15064), .ZN(net_14165), .A2(net_12230) );
NOR2_X2 inst_4812 ( .A2(net_6945), .ZN(net_4580), .A1(net_3351) );
NOR2_X4 inst_3090 ( .ZN(net_5474), .A2(net_4293), .A1(net_2582) );
INV_X4 inst_14466 ( .ZN(net_7871), .A(net_4921) );
INV_X4 inst_17050 ( .ZN(net_4792), .A(net_952) );
INV_X4 inst_14635 ( .A(net_14837), .ZN(net_4384) );
NAND2_X2 inst_10012 ( .ZN(net_8786), .A1(net_8785), .A2(net_8176) );
CLKBUF_X2 inst_22540 ( .A(net_22411), .Z(net_22412) );
INV_X4 inst_17751 ( .A(net_14029), .ZN(net_442) );
INV_X4 inst_14624 ( .ZN(net_4623), .A(net_4398) );
NAND2_X2 inst_8355 ( .A2(net_17488), .ZN(net_17462), .A1(net_17077) );
NOR2_X2 inst_4879 ( .A1(net_4259), .ZN(net_2188), .A2(net_2187) );
NOR2_X2 inst_4695 ( .ZN(net_4148), .A1(net_3915), .A2(net_2189) );
NOR2_X2 inst_4142 ( .ZN(net_8883), .A1(net_7260), .A2(net_3975) );
INV_X4 inst_17871 ( .A(net_227), .ZN(net_84) );
NAND2_X2 inst_12125 ( .ZN(net_352), .A2(net_199), .A1(net_63) );
NAND2_X2 inst_8513 ( .ZN(net_19680), .A1(net_16538), .A2(net_16523) );
INV_X4 inst_17591 ( .ZN(net_609), .A(net_333) );
NAND2_X2 inst_11260 ( .ZN(net_3910), .A2(net_2468), .A1(net_1163) );
NAND2_X2 inst_9097 ( .ZN(net_20382), .A2(net_13780), .A1(net_13673) );
INV_X4 inst_12680 ( .ZN(net_17729), .A(net_17728) );
INV_X8 inst_12206 ( .ZN(net_12436), .A(net_9751) );
INV_X4 inst_15267 ( .ZN(net_4405), .A(net_3834) );
INV_X4 inst_14774 ( .ZN(net_5108), .A(net_4047) );
NOR2_X4 inst_2859 ( .ZN(net_13819), .A1(net_11688), .A2(net_4995) );
INV_X4 inst_18036 ( .A(net_21173), .ZN(net_618) );
XNOR2_X2 inst_397 ( .B(net_21150), .A(net_20525), .ZN(net_16756) );
XNOR2_X2 inst_504 ( .ZN(net_8993), .B(net_5737), .A(net_2403) );
NAND2_X2 inst_8601 ( .A2(net_21118), .ZN(net_19667), .A1(net_16675) );
INV_X4 inst_14240 ( .ZN(net_11230), .A(net_5794) );
OAI22_X2 inst_1297 ( .ZN(net_11835), .A2(net_11834), .A1(net_10292), .B2(net_5125), .B1(net_2302) );
AOI211_X2 inst_21070 ( .ZN(net_7698), .B(net_5565), .C1(net_3514), .C2(net_3333), .A(net_3264) );
NOR2_X4 inst_3194 ( .A2(net_3984), .ZN(net_3863), .A1(net_3083) );
NOR2_X2 inst_3884 ( .ZN(net_9293), .A2(net_6266), .A1(net_4741) );
INV_X4 inst_13831 ( .A(net_9696), .ZN(net_7498) );
INV_X4 inst_16937 ( .A(net_1981), .ZN(net_924) );
NAND3_X2 inst_6296 ( .ZN(net_12818), .A2(net_10878), .A1(net_5508), .A3(net_5410) );
OR2_X2 inst_1173 ( .ZN(net_6003), .A1(net_6002), .A2(net_6001) );
AND2_X2 inst_21279 ( .A1(net_15026), .ZN(net_13585), .A2(net_13584) );
NAND2_X2 inst_9708 ( .ZN(net_10196), .A1(net_10195), .A2(net_10194) );
NOR2_X4 inst_2908 ( .ZN(net_8589), .A1(net_8588), .A2(net_6477) );
AOI21_X2 inst_20925 ( .B2(net_8938), .ZN(net_7171), .A(net_7170), .B1(net_3448) );
NOR2_X2 inst_5019 ( .A2(net_2490), .ZN(net_1232), .A1(net_1231) );
NAND2_X2 inst_9507 ( .ZN(net_11331), .A2(net_8153), .A1(net_5415) );
INV_X4 inst_17438 ( .ZN(net_11032), .A(net_10688) );
AOI21_X2 inst_20262 ( .ZN(net_18071), .B2(net_18070), .B1(net_15904), .A(net_13097) );
NOR2_X2 inst_4893 ( .A1(net_6599), .ZN(net_6457), .A2(net_3027) );
NAND3_X2 inst_5875 ( .A3(net_19906), .A1(net_19905), .ZN(net_15303), .A2(net_11316) );
AOI22_X2 inst_20003 ( .A1(net_14346), .ZN(net_13429), .B1(net_10298), .A2(net_9079), .B2(net_7754) );
NAND2_X2 inst_11318 ( .A1(net_20551), .ZN(net_8505), .A2(net_2770) );
NAND2_X2 inst_8514 ( .A1(net_17445), .ZN(net_16916), .A2(net_16911) );
NAND3_X2 inst_6717 ( .ZN(net_6777), .A2(net_6776), .A3(net_2830), .A1(net_1536) );
INV_X4 inst_17070 ( .ZN(net_1103), .A(net_955) );
NAND2_X2 inst_9807 ( .A1(net_14700), .ZN(net_9684), .A2(net_9683) );
NAND2_X2 inst_9089 ( .ZN(net_13795), .A2(net_12459), .A1(net_11389) );
INV_X4 inst_13684 ( .ZN(net_7974), .A(net_7973) );
NAND2_X2 inst_9302 ( .A1(net_15270), .ZN(net_12376), .A2(net_9119) );
INV_X4 inst_12995 ( .ZN(net_16630), .A(net_16488) );
NAND3_X2 inst_6283 ( .ZN(net_12892), .A3(net_12891), .A1(net_7055), .A2(net_2353) );
NAND2_X4 inst_7380 ( .A1(net_20566), .ZN(net_9046), .A2(net_4302) );
CLKBUF_X2 inst_22164 ( .A(net_22035), .Z(net_22036) );
NAND2_X4 inst_7387 ( .A2(net_20842), .ZN(net_7727), .A1(net_2139) );
NAND3_X2 inst_5857 ( .ZN(net_15400), .A1(net_14599), .A3(net_13140), .A2(net_12243) );
NAND2_X2 inst_9463 ( .ZN(net_11488), .A2(net_11487), .A1(net_10709) );
OAI21_X2 inst_1774 ( .ZN(net_14686), .B2(net_11945), .B1(net_11696), .A(net_11407) );
NAND2_X2 inst_8032 ( .ZN(net_18330), .A2(net_18188), .A1(net_18163) );
INV_X4 inst_12596 ( .ZN(net_18140), .A(net_18118) );
SDFF_X2 inst_985 ( .QN(net_21052), .D(net_736), .SE(net_263), .CK(net_22516), .SI(x2160) );
INV_X4 inst_12473 ( .ZN(net_18759), .A(net_18758) );
CLKBUF_X2 inst_21835 ( .A(net_21706), .Z(net_21707) );
NAND2_X4 inst_6943 ( .ZN(net_19017), .A2(net_17487), .A1(net_17307) );
INV_X4 inst_16202 ( .ZN(net_13576), .A(net_1663) );
INV_X2 inst_19300 ( .ZN(net_6406), .A(net_2776) );
INV_X4 inst_12985 ( .A(net_16843), .ZN(net_16642) );
NAND2_X2 inst_10627 ( .ZN(net_7804), .A1(net_7253), .A2(net_6555) );
INV_X4 inst_17408 ( .ZN(net_9325), .A(net_7268) );
INV_X2 inst_19286 ( .A(net_3883), .ZN(net_2880) );
INV_X4 inst_14208 ( .ZN(net_5925), .A(net_5924) );
INV_X4 inst_12563 ( .ZN(net_18224), .A(net_18223) );
NAND3_X2 inst_5918 ( .A3(net_20460), .A1(net_20459), .ZN(net_15007), .A2(net_11319) );
AOI21_X2 inst_20787 ( .B2(net_13146), .ZN(net_10548), .B1(net_5029), .A(net_855) );
INV_X4 inst_12969 ( .ZN(net_16688), .A(net_16517) );
CLKBUF_X2 inst_22152 ( .A(net_22023), .Z(net_22024) );
OAI21_X2 inst_2007 ( .ZN(net_11408), .A(net_11407), .B2(net_11406), .B1(net_2677) );
NOR2_X2 inst_3644 ( .ZN(net_12017), .A2(net_8810), .A1(net_5080) );
NAND2_X2 inst_10965 ( .A2(net_5165), .ZN(net_5058), .A1(net_4025) );
AND2_X2 inst_21354 ( .A1(net_20859), .ZN(net_2776), .A2(net_1216) );
SDFF_X2 inst_805 ( .Q(net_20946), .SE(net_18576), .SI(net_17959), .D(net_672), .CK(net_21264) );
NAND2_X2 inst_9991 ( .A1(net_12401), .ZN(net_12166), .A2(net_8845) );
NAND3_X2 inst_6005 ( .ZN(net_14425), .A3(net_12441), .A1(net_9371), .A2(net_3534) );
INV_X4 inst_17822 ( .ZN(net_337), .A(net_230) );
INV_X8 inst_12387 ( .ZN(net_195), .A(net_110) );
AOI211_X2 inst_21062 ( .ZN(net_9906), .A(net_9905), .C1(net_5250), .B(net_4487), .C2(net_1464) );
INV_X4 inst_12664 ( .ZN(net_17806), .A(net_17805) );
CLKBUF_X2 inst_22677 ( .A(net_22548), .Z(net_22549) );
INV_X4 inst_13735 ( .ZN(net_7657), .A(net_7656) );
NAND3_X4 inst_5603 ( .ZN(net_19359), .A3(net_12540), .A1(net_12434), .A2(net_9215) );
INV_X4 inst_14257 ( .A(net_8411), .ZN(net_5750) );
NAND3_X2 inst_6569 ( .ZN(net_10468), .A2(net_10467), .A3(net_9055), .A1(net_4709) );
XNOR2_X2 inst_373 ( .B(net_21200), .A(net_17517), .ZN(net_16841) );
INV_X4 inst_17801 ( .A(net_152), .ZN(net_124) );
DFF_X1 inst_19910 ( .D(net_16758), .CK(net_22788), .Q(x1238) );
OAI21_X2 inst_1868 ( .ZN(net_13733), .B2(net_12673), .A(net_9263), .B1(net_7645) );
INV_X4 inst_13672 ( .ZN(net_9576), .A(net_8029) );
NAND2_X2 inst_11428 ( .ZN(net_4415), .A2(net_3268), .A1(net_143) );
NAND2_X2 inst_9537 ( .A1(net_11764), .ZN(net_11066), .A2(net_11065) );
XOR2_X2 inst_22 ( .B(net_21118), .A(net_16764), .Z(net_16755) );
INV_X2 inst_19139 ( .ZN(net_4131), .A(net_4130) );
INV_X4 inst_13914 ( .A(net_13588), .ZN(net_6955) );
NOR2_X4 inst_3099 ( .ZN(net_5233), .A2(net_2620), .A1(net_502) );
INV_X4 inst_13289 ( .ZN(net_13440), .A(net_11051) );
NAND2_X4 inst_7034 ( .A1(net_19433), .ZN(net_16739), .A2(net_16414) );
SDFF_X2 inst_767 ( .Q(net_20972), .SE(net_18864), .SI(net_18507), .D(net_9259), .CK(net_22745) );
NAND2_X4 inst_7657 ( .ZN(net_1109), .A2(net_928), .A1(net_58) );
INV_X4 inst_14065 ( .ZN(net_9553), .A(net_8006) );
NOR2_X2 inst_3356 ( .ZN(net_17685), .A2(net_17638), .A1(net_17120) );
NAND2_X2 inst_10405 ( .A1(net_8976), .ZN(net_7271), .A2(net_7270) );
CLKBUF_X2 inst_21549 ( .A(net_21420), .Z(net_21421) );
INV_X2 inst_19429 ( .ZN(net_20836), .A(net_2422) );
CLKBUF_X2 inst_22855 ( .A(net_22726), .Z(net_22727) );
INV_X4 inst_18270 ( .A(net_19452), .ZN(net_19450) );
NAND2_X2 inst_7914 ( .ZN(net_18459), .A2(net_18348), .A1(net_18293) );
INV_X4 inst_15374 ( .ZN(net_18025), .A(net_29) );
CLKBUF_X2 inst_21658 ( .A(net_21529), .Z(net_21530) );
NOR2_X2 inst_4310 ( .ZN(net_8632), .A1(net_5940), .A2(net_5900) );
NAND2_X2 inst_8943 ( .ZN(net_19328), .A1(net_14731), .A2(net_13237) );
XNOR2_X2 inst_526 ( .A(net_21201), .B(net_5616), .ZN(net_3437) );
OR2_X2 inst_1178 ( .A1(net_13095), .ZN(net_5363), .A2(net_5362) );
NOR2_X4 inst_3104 ( .ZN(net_10034), .A1(net_4066), .A2(net_2746) );
NAND2_X2 inst_9174 ( .ZN(net_13346), .A2(net_10451), .A1(net_7968) );
OAI21_X4 inst_1450 ( .B2(net_19309), .B1(net_19308), .ZN(net_15448), .A(net_333) );
NAND2_X2 inst_8423 ( .ZN(net_20098), .A1(net_19455), .A2(net_16810) );
NAND3_X2 inst_6689 ( .A2(net_12474), .ZN(net_7707), .A1(net_2951), .A3(net_2772) );
NAND4_X2 inst_5511 ( .A1(net_11845), .ZN(net_10800), .A2(net_8980), .A3(net_8565), .A4(net_7079) );
NOR2_X4 inst_3123 ( .ZN(net_4940), .A2(net_4020), .A1(net_3977) );
NAND2_X2 inst_11592 ( .ZN(net_2691), .A2(net_2518), .A1(net_1064) );
NAND2_X2 inst_11149 ( .A1(net_8991), .ZN(net_7011), .A2(net_4209) );
NAND2_X2 inst_10645 ( .ZN(net_7644), .A2(net_6362), .A1(net_5900) );
INV_X4 inst_16098 ( .ZN(net_2642), .A(net_1331) );
NOR2_X2 inst_3725 ( .ZN(net_13629), .A1(net_9171), .A2(net_8246) );
NAND4_X2 inst_5400 ( .ZN(net_14780), .A3(net_12932), .A1(net_12632), .A4(net_12007), .A2(net_10890) );
CLKBUF_X2 inst_22845 ( .A(net_22716), .Z(net_22717) );
OAI21_X2 inst_1592 ( .A(net_16260), .ZN(net_16243), .B2(net_15898), .B1(net_9318) );
OAI21_X2 inst_1770 ( .ZN(net_14695), .A(net_14694), .B2(net_11952), .B1(net_11533) );
CLKBUF_X2 inst_22947 ( .A(net_22818), .Z(net_22819) );
NOR2_X2 inst_3413 ( .ZN(net_15641), .A2(net_14992), .A1(net_13519) );
NAND3_X2 inst_6095 ( .A3(net_14678), .A2(net_14617), .ZN(net_13925), .A1(net_12023) );
NOR2_X2 inst_4483 ( .ZN(net_4705), .A1(net_4329), .A2(net_4328) );
INV_X4 inst_12857 ( .ZN(net_19530), .A(net_16898) );
CLKBUF_X2 inst_21786 ( .A(net_21292), .Z(net_21658) );
CLKBUF_X2 inst_21400 ( .A(net_21267), .Z(net_21272) );
INV_X4 inst_15617 ( .ZN(net_4009), .A(net_2165) );
NAND2_X2 inst_11109 ( .A1(net_20548), .ZN(net_4327), .A2(net_4326) );
INV_X4 inst_14132 ( .ZN(net_7927), .A(net_5411) );
INV_X4 inst_16776 ( .ZN(net_19108), .A(net_802) );
INV_X2 inst_18734 ( .A(net_8736), .ZN(net_7983) );
OAI21_X4 inst_1419 ( .B2(net_19496), .B1(net_19495), .ZN(net_19485), .A(net_16394) );
INV_X4 inst_14544 ( .ZN(net_9698), .A(net_4623) );
OAI211_X2 inst_2501 ( .ZN(net_12814), .A(net_12813), .B(net_12812), .C2(net_11225), .C1(net_5415) );
INV_X2 inst_18665 ( .A(net_12475), .ZN(net_9177) );
CLKBUF_X2 inst_21983 ( .A(net_21726), .Z(net_21855) );
INV_X4 inst_14164 ( .ZN(net_7478), .A(net_6014) );
INV_X4 inst_16233 ( .A(net_9542), .ZN(net_7903) );
INV_X2 inst_18796 ( .ZN(net_7431), .A(net_7430) );
INV_X4 inst_16657 ( .ZN(net_6617), .A(net_5220) );
AND2_X2 inst_21371 ( .ZN(net_3482), .A2(net_143), .A1(net_112) );
INV_X4 inst_13314 ( .ZN(net_11624), .A(net_11623) );
OAI211_X4 inst_2378 ( .B(net_20738), .A(net_20737), .C1(net_19032), .ZN(net_16061), .C2(net_15039) );
INV_X4 inst_15942 ( .ZN(net_2486), .A(net_2114) );
NAND3_X2 inst_6302 ( .ZN(net_12803), .A2(net_12802), .A1(net_9433), .A3(net_8788) );
INV_X4 inst_14137 ( .ZN(net_9416), .A(net_6086) );
NAND2_X2 inst_9996 ( .ZN(net_10317), .A1(net_8836), .A2(net_8303) );
CLKBUF_X2 inst_21740 ( .A(net_21611), .Z(net_21612) );
AOI21_X2 inst_20421 ( .B1(net_15248), .ZN(net_15222), .B2(net_14090), .A(net_8259) );
AOI21_X2 inst_20428 ( .ZN(net_15200), .B2(net_13982), .B1(net_13338), .A(net_1052) );
INV_X4 inst_14392 ( .ZN(net_9152), .A(net_8901) );
INV_X4 inst_13874 ( .ZN(net_7412), .A(net_7411) );
INV_X4 inst_13164 ( .ZN(net_14809), .A(net_14224) );
CLKBUF_X2 inst_22838 ( .A(net_22709), .Z(net_22710) );
INV_X4 inst_16472 ( .A(net_11511), .ZN(net_11088) );
NAND2_X2 inst_12079 ( .A1(net_1682), .ZN(net_1323), .A2(net_896) );
INV_X4 inst_15237 ( .ZN(net_6492), .A(net_2151) );
NAND2_X2 inst_10072 ( .A1(net_10515), .ZN(net_8654), .A2(net_6704) );
INV_X4 inst_17482 ( .A(net_10714), .ZN(net_8021) );
NAND2_X2 inst_11153 ( .ZN(net_4202), .A2(net_2117), .A1(net_768) );
INV_X4 inst_16885 ( .A(net_7173), .ZN(net_1292) );
INV_X4 inst_16018 ( .ZN(net_13416), .A(net_10917) );
INV_X4 inst_15569 ( .ZN(net_3010), .A(net_2562) );
NAND2_X2 inst_12031 ( .ZN(net_1336), .A2(net_459), .A1(net_223) );
INV_X4 inst_14560 ( .ZN(net_6191), .A(net_4567) );
NAND3_X2 inst_6740 ( .ZN(net_6456), .A2(net_6455), .A3(net_5675), .A1(net_2986) );
NAND2_X2 inst_10501 ( .A1(net_10714), .ZN(net_10367), .A2(net_6920) );
NAND2_X2 inst_10796 ( .ZN(net_8973), .A2(net_3936), .A1(net_624) );
NAND2_X2 inst_8847 ( .ZN(net_15398), .A2(net_14562), .A1(net_13526) );
INV_X4 inst_16616 ( .ZN(net_1500), .A(net_1119) );
NOR2_X2 inst_3801 ( .ZN(net_9857), .A2(net_9476), .A1(net_5625) );
NOR2_X2 inst_4177 ( .ZN(net_8136), .A2(net_6725), .A1(net_4403) );
NAND2_X2 inst_9350 ( .ZN(net_12182), .A2(net_9902), .A1(net_731) );
INV_X4 inst_17187 ( .ZN(net_5458), .A(net_721) );
NAND3_X2 inst_6491 ( .ZN(net_11166), .A2(net_11165), .A3(net_11164), .A1(net_7491) );
INV_X4 inst_15870 ( .ZN(net_13709), .A(net_7210) );
INV_X4 inst_13133 ( .ZN(net_15263), .A(net_14860) );
NAND2_X2 inst_9193 ( .ZN(net_13113), .A1(net_13112), .A2(net_10350) );
OAI21_X2 inst_2155 ( .A(net_11929), .ZN(net_9277), .B2(net_9276), .B1(net_2759) );
INV_X4 inst_12927 ( .A(net_17233), .ZN(net_16657) );
NAND3_X2 inst_6352 ( .ZN(net_12159), .A3(net_11763), .A1(net_9913), .A2(net_7288) );
XNOR2_X2 inst_464 ( .B(net_16334), .ZN(net_13282), .A(net_9007) );
INV_X4 inst_13428 ( .ZN(net_9896), .A(net_8465) );
NAND4_X2 inst_5360 ( .ZN(net_15318), .A2(net_13727), .A3(net_12399), .A1(net_11491), .A4(net_10062) );
INV_X4 inst_13392 ( .ZN(net_12157), .A(net_7475) );
XNOR2_X2 inst_341 ( .B(net_21140), .ZN(net_16963), .A(net_16487) );
INV_X4 inst_15194 ( .A(net_4188), .ZN(net_2929) );
INV_X8 inst_12313 ( .ZN(net_1787), .A(net_372) );
INV_X4 inst_14961 ( .ZN(net_3479), .A(net_3478) );
INV_X4 inst_13090 ( .ZN(net_15979), .A(net_15862) );
INV_X4 inst_14006 ( .ZN(net_6343), .A(net_6342) );
NAND2_X2 inst_11095 ( .A1(net_5342), .ZN(net_4354), .A2(net_2186) );
OAI21_X2 inst_2359 ( .ZN(net_1098), .B1(net_1097), .A(net_978), .B2(net_664) );
NOR2_X2 inst_3702 ( .ZN(net_11101), .A2(net_7570), .A1(net_7144) );
NAND2_X2 inst_11229 ( .ZN(net_3952), .A2(net_2762), .A1(net_2585) );
AOI21_X2 inst_20372 ( .B1(net_20351), .ZN(net_15608), .B2(net_15607), .A(net_9101) );
NAND2_X2 inst_8526 ( .ZN(net_16900), .A2(net_16899), .A1(net_7771) );
INV_X4 inst_17090 ( .ZN(net_1403), .A(net_803) );
INV_X4 inst_13913 ( .ZN(net_8845), .A(net_6966) );
INV_X4 inst_13031 ( .A(net_16718), .ZN(net_16437) );
NAND2_X2 inst_8505 ( .A2(net_20502), .ZN(net_16926), .A1(net_9255) );
NAND3_X4 inst_5556 ( .ZN(net_19609), .A2(net_15860), .A3(net_15472), .A1(net_6554) );
NAND3_X1 inst_6826 ( .ZN(net_6463), .A3(net_4837), .A2(net_3101), .A1(net_2713) );
CLKBUF_X2 inst_22698 ( .A(net_22569), .Z(net_22570) );
NAND2_X2 inst_10226 ( .A2(net_11192), .ZN(net_8063), .A1(net_60) );
INV_X2 inst_19160 ( .A(net_5543), .ZN(net_4969) );
NAND2_X2 inst_8840 ( .ZN(net_15456), .A2(net_14976), .A1(net_14628) );
NOR2_X2 inst_4968 ( .ZN(net_6451), .A1(net_1588), .A2(net_1300) );
INV_X4 inst_14319 ( .ZN(net_5461), .A(net_5460) );
CLKBUF_X2 inst_21550 ( .A(net_21421), .Z(net_21422) );
NAND2_X2 inst_10122 ( .A2(net_9832), .ZN(net_8373), .A1(net_4526) );
NOR2_X2 inst_4162 ( .A1(net_9083), .ZN(net_8215), .A2(net_6521) );
INV_X2 inst_19572 ( .ZN(net_1196), .A(net_658) );
CLKBUF_X2 inst_21575 ( .A(net_21244), .Z(net_21447) );
AOI21_X2 inst_20650 ( .ZN(net_13057), .B2(net_9837), .B1(net_7788), .A(net_652) );
NAND4_X4 inst_5171 ( .A3(net_19339), .A1(net_19338), .ZN(net_16870), .A4(net_16304), .A2(net_14882) );
INV_X4 inst_12936 ( .A(net_17126), .ZN(net_16639) );
INV_X2 inst_18600 ( .ZN(net_9919), .A(net_8489) );
INV_X4 inst_17812 ( .A(net_20897), .ZN(net_278) );
INV_X4 inst_14363 ( .ZN(net_5219), .A(net_5218) );
NOR2_X4 inst_3201 ( .ZN(net_3515), .A1(net_3054), .A2(net_2017) );
INV_X4 inst_17554 ( .A(net_4945), .ZN(net_4323) );
INV_X4 inst_17930 ( .A(net_21104), .ZN(net_55) );
INV_X4 inst_14532 ( .ZN(net_12457), .A(net_4700) );
INV_X4 inst_16080 ( .ZN(net_3084), .A(net_1548) );
XNOR2_X2 inst_251 ( .ZN(net_17311), .A(net_17310), .B(net_13289) );
NAND2_X2 inst_10651 ( .A1(net_13504), .ZN(net_6350), .A2(net_6349) );
OAI21_X2 inst_1552 ( .ZN(net_17703), .A(net_17452), .B1(net_17451), .B2(net_17450) );
OAI21_X2 inst_1524 ( .B2(net_19386), .B1(net_19385), .ZN(net_18896), .A(net_18067) );
INV_X4 inst_18171 ( .A(net_20973), .ZN(net_74) );
INV_X4 inst_13983 ( .ZN(net_13460), .A(net_6578) );
NAND2_X2 inst_9369 ( .ZN(net_12110), .A1(net_12109), .A2(net_9936) );
NOR2_X2 inst_4789 ( .A2(net_7663), .ZN(net_2793), .A1(net_1146) );
NOR2_X2 inst_4977 ( .ZN(net_6444), .A2(net_1542), .A1(net_417) );
INV_X4 inst_15481 ( .ZN(net_5579), .A(net_3102) );
NAND2_X2 inst_9892 ( .ZN(net_12842), .A2(net_9384), .A1(net_5246) );
NAND2_X2 inst_7781 ( .ZN(net_18727), .A2(net_18723), .A1(net_18645) );
INV_X2 inst_18522 ( .ZN(net_11336), .A(net_10027) );
INV_X4 inst_15734 ( .ZN(net_2602), .A(net_2140) );
INV_X4 inst_13628 ( .A(net_10452), .ZN(net_9772) );
SDFF_X2 inst_898 ( .Q(net_21123), .D(net_16773), .SE(net_263), .CK(net_21532), .SI(x4285) );
OAI21_X2 inst_1977 ( .A(net_13058), .ZN(net_12146), .B1(net_8721), .B2(net_8227) );
OAI21_X2 inst_1793 ( .A(net_15677), .ZN(net_14598), .B2(net_11723), .B1(net_9265) );
NAND2_X2 inst_8012 ( .ZN(net_18294), .A2(net_18244), .A1(net_17261) );
NAND2_X2 inst_9223 ( .ZN(net_12951), .A2(net_12950), .A1(net_4719) );
NAND2_X2 inst_9747 ( .ZN(net_19904), .A1(net_10082), .A2(net_8383) );
NAND2_X2 inst_11804 ( .ZN(net_4162), .A2(net_3648), .A1(net_3493) );
NAND4_X2 inst_5299 ( .ZN(net_15904), .A2(net_15291), .A4(net_14691), .A1(net_14364), .A3(net_13028) );
NAND2_X2 inst_10805 ( .ZN(net_8982), .A1(net_7975), .A2(net_5543) );
NAND3_X2 inst_5697 ( .A3(net_20302), .A1(net_20301), .ZN(net_19387), .A2(net_14854) );
OAI21_X2 inst_2291 ( .ZN(net_6515), .A(net_5181), .B2(net_2899), .B1(net_2841) );
NAND2_X2 inst_8230 ( .ZN(net_17792), .A1(net_17669), .A2(net_17524) );
NOR2_X2 inst_4822 ( .ZN(net_12954), .A2(net_3182), .A1(net_143) );
NOR2_X4 inst_3132 ( .A1(net_19008), .ZN(net_4823), .A2(net_3830) );
INV_X4 inst_16572 ( .ZN(net_6538), .A(net_827) );
INV_X4 inst_13835 ( .ZN(net_11251), .A(net_7492) );
INV_X2 inst_18768 ( .ZN(net_7593), .A(net_7592) );
INV_X4 inst_16419 ( .ZN(net_3385), .A(net_168) );
NAND2_X4 inst_7395 ( .ZN(net_5199), .A1(net_2966), .A2(net_809) );
NOR2_X2 inst_4999 ( .ZN(net_1365), .A2(net_1364), .A1(net_493) );
NAND3_X2 inst_6071 ( .ZN(net_14123), .A3(net_10551), .A1(net_8875), .A2(net_5702) );
AOI21_X2 inst_20444 ( .B1(net_20889), .ZN(net_15120), .B2(net_13219), .A(net_12128) );
NAND3_X2 inst_5819 ( .ZN(net_15594), .A1(net_14890), .A2(net_13494), .A3(net_13146) );
NOR2_X2 inst_3910 ( .A1(net_11366), .A2(net_10606), .ZN(net_10339) );
AOI21_X4 inst_20258 ( .ZN(net_4225), .A(net_3297), .B1(net_2166), .B2(net_2101) );
CLKBUF_X2 inst_22907 ( .A(net_22778), .Z(net_22779) );
INV_X2 inst_18540 ( .ZN(net_11011), .A(net_11010) );
OAI221_X2 inst_1332 ( .C1(net_15858), .ZN(net_15551), .A(net_15143), .C2(net_13309), .B1(net_10947), .B2(net_9021) );
OAI21_X2 inst_1841 ( .A(net_15334), .ZN(net_14025), .B2(net_10271), .B1(net_3738) );
NOR2_X2 inst_3345 ( .A2(net_18147), .ZN(net_18087), .A1(net_12455) );
AND2_X4 inst_21211 ( .ZN(net_11906), .A1(net_8639), .A2(net_6670) );
NOR2_X4 inst_3264 ( .ZN(net_2716), .A1(net_1462), .A2(net_168) );
INV_X4 inst_16802 ( .ZN(net_15191), .A(net_1012) );
OAI21_X2 inst_2332 ( .ZN(net_4691), .A(net_4690), .B2(net_3648), .B1(net_3554) );
INV_X4 inst_13415 ( .A(net_12875), .ZN(net_11623) );
NAND2_X2 inst_9082 ( .ZN(net_13817), .A2(net_12567), .A1(net_652) );
INV_X4 inst_13431 ( .ZN(net_9874), .A(net_8439) );
CLKBUF_X2 inst_22539 ( .A(net_22410), .Z(net_22411) );
INV_X2 inst_18538 ( .ZN(net_13669), .A(net_11038) );
INV_X4 inst_17455 ( .ZN(net_1175), .A(net_186) );
INV_X4 inst_16019 ( .ZN(net_2779), .A(net_1647) );
NAND3_X2 inst_5946 ( .ZN(net_14891), .A1(net_13721), .A3(net_9552), .A2(net_3000) );
OAI21_X2 inst_2310 ( .A(net_8179), .ZN(net_5745), .B2(net_4304), .B1(net_2854) );
CLKBUF_X2 inst_22755 ( .A(net_21800), .Z(net_22627) );
INV_X4 inst_14327 ( .ZN(net_7958), .A(net_4276) );
NOR2_X2 inst_5017 ( .ZN(net_7399), .A2(net_951), .A1(net_112) );
AOI21_X2 inst_20545 ( .B1(net_19738), .ZN(net_14398), .B2(net_11186), .A(net_9563) );
OAI22_X2 inst_1290 ( .ZN(net_12879), .A2(net_12878), .B1(net_12877), .A1(net_11681), .B2(net_7041) );
INV_X4 inst_16461 ( .ZN(net_5157), .A(net_809) );
NAND2_X2 inst_7939 ( .ZN(net_18425), .A1(net_18367), .A2(net_18307) );
NAND2_X2 inst_11451 ( .ZN(net_4307), .A2(net_2405), .A1(net_2361) );
NAND3_X2 inst_6342 ( .A3(net_14643), .ZN(net_12252), .A1(net_9052), .A2(net_3370) );
NAND3_X2 inst_5845 ( .ZN(net_15443), .A3(net_14398), .A2(net_8463), .A1(net_7899) );
NOR2_X2 inst_5038 ( .A1(net_1699), .ZN(net_1490), .A2(net_133) );
CLKBUF_X2 inst_21535 ( .A(net_21406), .Z(net_21407) );
INV_X4 inst_18090 ( .A(net_20927), .ZN(net_513) );
INV_X4 inst_13399 ( .ZN(net_10492), .A(net_8989) );
NOR2_X2 inst_5142 ( .A1(net_1271), .A2(net_386), .ZN(net_141) );
NAND3_X2 inst_5757 ( .ZN(net_19994), .A1(net_15701), .A3(net_15139), .A2(net_8532) );
CLKBUF_X2 inst_21714 ( .A(net_21585), .Z(net_21586) );
NOR2_X2 inst_4899 ( .ZN(net_2000), .A1(net_1999), .A2(net_1998) );
INV_X4 inst_15865 ( .ZN(net_1960), .A(net_1804) );
CLKBUF_X2 inst_21909 ( .A(net_21780), .Z(net_21781) );
INV_X4 inst_12604 ( .ZN(net_18142), .A(net_18084) );
NOR2_X2 inst_5079 ( .ZN(net_7237), .A2(net_884), .A1(net_68) );
NAND3_X2 inst_6429 ( .ZN(net_11916), .A3(net_11915), .A1(net_9846), .A2(net_3932) );
NOR2_X2 inst_3861 ( .A1(net_20569), .A2(net_13497), .ZN(net_11478) );
CLKBUF_X2 inst_21559 ( .A(net_21392), .Z(net_21431) );
INV_X4 inst_15809 ( .ZN(net_3384), .A(net_1390) );
NOR2_X2 inst_4399 ( .A2(net_9295), .ZN(net_8360), .A1(net_5173) );
NAND2_X2 inst_11547 ( .A1(net_3133), .ZN(net_2885), .A2(net_2884) );
NAND2_X2 inst_9847 ( .ZN(net_9538), .A1(net_7576), .A2(net_7099) );
NAND2_X2 inst_9840 ( .ZN(net_9562), .A2(net_8019), .A1(net_7613) );
INV_X4 inst_16864 ( .A(net_14657), .ZN(net_14159) );
NOR2_X2 inst_4196 ( .ZN(net_19922), .A2(net_13840), .A1(net_13093) );
CLKBUF_X2 inst_22296 ( .A(net_21851), .Z(net_22168) );
CLKBUF_X2 inst_21458 ( .A(net_21329), .Z(net_21330) );
NAND2_X2 inst_10672 ( .ZN(net_9766), .A1(net_6981), .A2(net_6166) );
SDFF_X2 inst_1014 ( .QN(net_21082), .D(net_473), .SE(net_263), .CK(net_22573), .SI(x1686) );
OAI211_X2 inst_2531 ( .C1(net_13926), .ZN(net_11745), .A(net_11744), .C2(net_11743), .B(net_9583) );
NAND2_X2 inst_10009 ( .A1(net_12504), .A2(net_11627), .ZN(net_10293) );
NAND3_X2 inst_6781 ( .ZN(net_4294), .A2(net_2247), .A3(net_1576), .A1(net_1534) );
INV_X2 inst_19480 ( .A(net_2337), .ZN(net_1386) );
INV_X4 inst_14918 ( .ZN(net_19022), .A(net_4826) );
NAND2_X2 inst_11879 ( .A1(net_20798), .A2(net_5259), .ZN(net_1621) );
CLKBUF_X2 inst_22720 ( .A(net_22591), .Z(net_22592) );
INV_X4 inst_16597 ( .A(net_3713), .ZN(net_1137) );
INV_X2 inst_18363 ( .A(net_18112), .ZN(net_18106) );
INV_X8 inst_12299 ( .ZN(net_9571), .A(net_6849) );
INV_X4 inst_16479 ( .ZN(net_1206), .A(net_1205) );
OAI21_X2 inst_1680 ( .ZN(net_20223), .B2(net_14450), .B1(net_9093), .A(net_238) );
INV_X4 inst_15221 ( .ZN(net_5032), .A(net_2868) );
OAI21_X2 inst_1626 ( .B1(net_19128), .ZN(net_16029), .B2(net_14643), .A(net_13665) );
INV_X4 inst_12834 ( .ZN(net_17278), .A(net_17125) );
INV_X4 inst_16323 ( .ZN(net_1313), .A(net_1110) );
CLKBUF_X2 inst_21947 ( .A(net_21818), .Z(net_21819) );
INV_X8 inst_12271 ( .ZN(net_2430), .A(net_1179) );
AND2_X2 inst_21359 ( .A2(net_4615), .A1(net_1583), .ZN(net_1483) );
NAND3_X2 inst_6528 ( .A2(net_11245), .ZN(net_10607), .A3(net_10606), .A1(net_6832) );
NAND2_X2 inst_9789 ( .ZN(net_9742), .A2(net_9741), .A1(net_8744) );
NAND2_X2 inst_9117 ( .A1(net_15573), .ZN(net_13567), .A2(net_13566) );
NOR2_X2 inst_3894 ( .ZN(net_9182), .A2(net_9181), .A1(net_4156) );
NAND2_X2 inst_8037 ( .ZN(net_18255), .A1(net_18237), .A2(net_18169) );
AOI21_X2 inst_20580 ( .ZN(net_14080), .A(net_13375), .B2(net_10305), .B1(net_3649) );
NAND2_X2 inst_10132 ( .ZN(net_12031), .A2(net_9832), .A1(net_8341) );
NAND4_X2 inst_5385 ( .ZN(net_19476), .A3(net_15018), .A4(net_13171), .A1(net_13124), .A2(net_12547) );
OR2_X4 inst_1087 ( .ZN(net_4976), .A1(net_4975), .A2(net_4791) );
INV_X4 inst_17055 ( .A(net_2179), .ZN(net_1689) );
AOI21_X2 inst_20355 ( .ZN(net_15695), .B1(net_15694), .B2(net_15016), .A(net_13977) );
INV_X4 inst_13701 ( .ZN(net_12079), .A(net_7882) );
INV_X4 inst_14453 ( .ZN(net_19515), .A(net_9623) );
NAND2_X2 inst_10061 ( .A1(net_13999), .ZN(net_8680), .A2(net_8635) );
OAI21_X4 inst_1375 ( .B1(net_20649), .ZN(net_16424), .B2(net_16368), .A(net_16291) );
INV_X8 inst_12199 ( .ZN(net_15860), .A(net_15711) );
INV_X4 inst_15693 ( .A(net_2757), .ZN(net_2022) );
NAND2_X2 inst_7966 ( .ZN(net_18367), .A2(net_18288), .A1(net_18205) );
INV_X2 inst_19097 ( .A(net_5952), .ZN(net_4541) );
INV_X2 inst_19373 ( .A(net_3217), .ZN(net_2186) );
NOR2_X2 inst_4564 ( .ZN(net_4431), .A2(net_3903), .A1(net_454) );
INV_X4 inst_15134 ( .ZN(net_3983), .A(net_2234) );
NAND2_X2 inst_9290 ( .ZN(net_12461), .A2(net_9402), .A1(net_8182) );
NAND4_X2 inst_5258 ( .A2(net_20117), .A1(net_20116), .A4(net_20096), .ZN(net_16328), .A3(net_15793) );
INV_X8 inst_12235 ( .ZN(net_5909), .A(net_3562) );
NAND2_X2 inst_11209 ( .ZN(net_4501), .A1(net_4042), .A2(net_3439) );
OAI211_X2 inst_2564 ( .A(net_12813), .ZN(net_9868), .B(net_9867), .C2(net_4474), .C1(net_81) );
CLKBUF_X2 inst_22504 ( .A(net_22375), .Z(net_22376) );
INV_X4 inst_15173 ( .A(net_4355), .ZN(net_3011) );
OR2_X4 inst_1082 ( .ZN(net_5892), .A2(net_5891), .A1(net_948) );
INV_X4 inst_15185 ( .ZN(net_3667), .A(net_2966) );
NOR3_X2 inst_2677 ( .ZN(net_20251), .A3(net_19809), .A1(net_19808), .A2(net_10457) );
NAND2_X2 inst_10068 ( .A1(net_11747), .A2(net_11324), .ZN(net_10126) );
XNOR2_X2 inst_105 ( .ZN(net_18527), .A(net_18460), .B(net_18360) );
INV_X2 inst_18529 ( .ZN(net_11097), .A(net_11096) );
NOR2_X2 inst_3518 ( .A1(net_14151), .ZN(net_13771), .A2(net_12515) );
INV_X2 inst_18888 ( .ZN(net_9702), .A(net_6132) );
OAI21_X2 inst_2161 ( .ZN(net_9142), .B2(net_5368), .B1(net_3744), .A(net_934) );
NAND2_X2 inst_8294 ( .ZN(net_17612), .A2(net_17611), .A1(net_17197) );
XNOR2_X2 inst_625 ( .B(net_15294), .ZN(net_464), .A(net_463) );
AOI21_X2 inst_20944 ( .ZN(net_6397), .B1(net_4672), .B2(net_3883), .A(net_2877) );
DFF_X1 inst_19802 ( .D(net_18172), .CK(net_22395), .Q(x797) );
INV_X4 inst_16855 ( .ZN(net_10286), .A(net_4403) );
NAND3_X2 inst_6747 ( .ZN(net_5800), .A2(net_5799), .A3(net_2871), .A1(net_1817) );
INV_X4 inst_14041 ( .ZN(net_10728), .A(net_6262) );
NAND2_X2 inst_8119 ( .A1(net_20073), .ZN(net_19342), .A2(net_18079) );
AND2_X2 inst_21338 ( .A2(net_4687), .ZN(net_3166), .A1(net_3165) );
INV_X2 inst_19269 ( .A(net_3262), .ZN(net_3062) );
XNOR2_X2 inst_181 ( .ZN(net_17768), .B(net_17767), .A(net_17334) );
INV_X4 inst_17460 ( .ZN(net_14720), .A(net_14563) );
INV_X4 inst_13212 ( .ZN(net_20176), .A(net_12834) );
NAND2_X2 inst_8964 ( .ZN(net_14679), .A1(net_14678), .A2(net_13312) );
NAND2_X2 inst_8329 ( .ZN(net_17545), .A2(net_17544), .A1(net_13299) );
NAND4_X4 inst_5215 ( .A4(net_19366), .A1(net_19365), .ZN(net_16778), .A3(net_16208), .A2(net_14041) );
AOI21_X2 inst_20937 ( .ZN(net_6469), .A(net_6468), .B1(net_5260), .B2(net_2475) );
INV_X2 inst_19674 ( .A(net_20497), .ZN(net_20496) );
INV_X4 inst_17470 ( .ZN(net_12398), .A(net_442) );
INV_X4 inst_17479 ( .ZN(net_1142), .A(net_191) );
CLKBUF_X2 inst_21484 ( .A(net_21338), .Z(net_21356) );
NAND2_X2 inst_10885 ( .ZN(net_5411), .A2(net_5291), .A1(net_3682) );
INV_X4 inst_16723 ( .ZN(net_2241), .A(net_820) );
AOI21_X4 inst_20165 ( .B1(net_19973), .ZN(net_15635), .B2(net_15499), .A(net_13660) );
INV_X2 inst_18568 ( .A(net_12962), .ZN(net_10771) );
NAND2_X2 inst_9738 ( .ZN(net_13046), .A1(net_12306), .A2(net_9391) );
SDFF_X2 inst_713 ( .Q(net_20952), .SE(net_18865), .SI(net_18809), .D(net_611), .CK(net_21499) );
NAND2_X2 inst_10125 ( .ZN(net_8362), .A1(net_8361), .A2(net_8360) );
CLKBUF_X2 inst_22957 ( .A(net_22828), .Z(net_22829) );
INV_X4 inst_16548 ( .A(net_2953), .ZN(net_2733) );
NAND2_X4 inst_6918 ( .ZN(net_18208), .A1(net_17582), .A2(net_17516) );
CLKBUF_X2 inst_22682 ( .A(net_22553), .Z(net_22554) );
INV_X2 inst_19176 ( .ZN(net_3803), .A(net_3802) );
INV_X4 inst_17578 ( .A(net_10714), .ZN(net_8707) );
NAND2_X2 inst_11508 ( .A2(net_3861), .ZN(net_3531), .A1(net_2143) );
INV_X4 inst_16492 ( .ZN(net_6911), .A(net_117) );
INV_X4 inst_15256 ( .ZN(net_5127), .A(net_2786) );
NAND2_X2 inst_7768 ( .ZN(net_18746), .A2(net_18745), .A1(net_17732) );
INV_X4 inst_17036 ( .A(net_1547), .ZN(net_840) );
INV_X4 inst_14062 ( .ZN(net_9610), .A(net_6246) );
NOR2_X4 inst_3208 ( .ZN(net_5521), .A2(net_3026), .A1(net_3025) );
NAND2_X4 inst_7410 ( .ZN(net_6629), .A2(net_3861), .A1(net_2791) );
NOR2_X2 inst_4134 ( .ZN(net_6954), .A1(net_6953), .A2(net_6952) );
NOR2_X2 inst_3507 ( .ZN(net_13973), .A2(net_12003), .A1(net_8845) );
XNOR2_X2 inst_271 ( .B(net_21171), .ZN(net_17217), .A(net_17216) );
AND2_X2 inst_21304 ( .ZN(net_9752), .A2(net_9751), .A1(net_8539) );
NAND2_X2 inst_11918 ( .A2(net_20581), .ZN(net_1546), .A1(net_1545) );
NAND3_X2 inst_6705 ( .A3(net_10042), .A2(net_8467), .ZN(net_7345), .A1(net_3833) );
OR2_X2 inst_1230 ( .ZN(net_5302), .A1(net_2329), .A2(net_2107) );
INV_X4 inst_16979 ( .ZN(net_10819), .A(net_487) );
NAND2_X2 inst_10844 ( .ZN(net_11340), .A2(net_4356), .A1(net_535) );
NAND2_X4 inst_7262 ( .ZN(net_10643), .A2(net_9478), .A1(net_6579) );
NOR2_X2 inst_3535 ( .A1(net_14395), .ZN(net_13454), .A2(net_10780) );
INV_X4 inst_17880 ( .ZN(net_550), .A(net_386) );
NAND2_X2 inst_9344 ( .A1(net_16046), .ZN(net_12207), .A2(net_8911) );
INV_X4 inst_14685 ( .A(net_11860), .ZN(net_7849) );
NOR2_X2 inst_3497 ( .ZN(net_14087), .A1(net_12412), .A2(net_10632) );
INV_X4 inst_17752 ( .ZN(net_710), .A(net_166) );
OR3_X2 inst_1064 ( .A3(net_2744), .ZN(net_2678), .A1(net_2476), .A2(net_761) );
NAND4_X2 inst_5416 ( .ZN(net_14581), .A2(net_11561), .A3(net_11495), .A4(net_10301), .A1(net_9763) );
INV_X4 inst_17193 ( .ZN(net_712), .A(net_711) );
INV_X4 inst_14875 ( .ZN(net_3687), .A(net_3686) );
AOI21_X2 inst_20631 ( .ZN(net_13393), .B1(net_12184), .B2(net_8752), .A(net_1051) );
INV_X2 inst_19605 ( .A(net_21223), .ZN(net_98) );
NAND2_X2 inst_11110 ( .A2(net_6942), .ZN(net_5554), .A1(net_1830) );
NOR2_X2 inst_3599 ( .ZN(net_12553), .A2(net_9595), .A1(net_6912) );
CLKBUF_X2 inst_22623 ( .A(net_22050), .Z(net_22495) );
INV_X4 inst_14335 ( .ZN(net_8344), .A(net_5391) );
INV_X4 inst_14539 ( .A(net_6357), .ZN(net_4651) );
CLKBUF_X2 inst_21607 ( .A(net_21478), .Z(net_21479) );
INV_X4 inst_17490 ( .ZN(net_1415), .A(net_459) );
INV_X4 inst_13727 ( .A(net_7798), .ZN(net_7797) );
INV_X4 inst_17737 ( .ZN(net_2329), .A(net_304) );
NAND2_X2 inst_12124 ( .ZN(net_734), .A1(net_279), .A2(net_189) );
NAND4_X4 inst_5208 ( .ZN(net_20766), .A1(net_16238), .A4(net_16060), .A2(net_15885), .A3(net_5261) );
NOR2_X2 inst_3581 ( .ZN(net_12684), .A2(net_10982), .A1(net_8111) );
NAND2_X2 inst_9930 ( .ZN(net_9159), .A2(net_7114), .A1(net_112) );
AOI21_X2 inst_20304 ( .ZN(net_20657), .B1(net_19552), .B2(net_15804), .A(net_14947) );
NOR2_X2 inst_4833 ( .ZN(net_2379), .A2(net_1844), .A1(net_1707) );
OAI21_X2 inst_2065 ( .ZN(net_10675), .A(net_9968), .B1(net_9348), .B2(net_5586) );
NAND2_X2 inst_10765 ( .ZN(net_5640), .A2(net_5639), .A1(net_5623) );
OAI21_X2 inst_2251 ( .A(net_14617), .ZN(net_7297), .B2(net_5525), .B1(net_3612) );
NOR2_X2 inst_3987 ( .A1(net_15224), .ZN(net_8320), .A2(net_7280) );
INV_X4 inst_18008 ( .A(net_20964), .ZN(net_85) );
AOI21_X2 inst_20593 ( .ZN(net_13932), .B2(net_11284), .B1(net_9367), .A(net_6739) );
INV_X4 inst_12825 ( .ZN(net_17157), .A(net_17156) );
INV_X4 inst_13720 ( .ZN(net_12809), .A(net_7814) );
NOR2_X2 inst_5124 ( .ZN(net_276), .A2(net_51), .A1(net_38) );
INV_X2 inst_18797 ( .ZN(net_7426), .A(net_7425) );
INV_X4 inst_13226 ( .ZN(net_19371), .A(net_13595) );
OAI21_X2 inst_1899 ( .ZN(net_13352), .A(net_10108), .B2(net_9957), .B1(net_6644) );
NAND2_X4 inst_7200 ( .A1(net_19210), .ZN(net_10221), .A2(net_7941) );
NAND2_X2 inst_9349 ( .ZN(net_12186), .A1(net_12185), .A2(net_12184) );
OAI211_X2 inst_2569 ( .C2(net_11245), .ZN(net_9025), .A(net_9024), .C1(net_9023), .B(net_3207) );
NAND2_X2 inst_10573 ( .A2(net_7258), .ZN(net_6694), .A1(net_4820) );
AOI21_X2 inst_20804 ( .ZN(net_10346), .A(net_10345), .B2(net_6167), .B1(net_2781) );
NAND2_X2 inst_10197 ( .A2(net_9999), .ZN(net_8135), .A1(net_8041) );
NAND2_X2 inst_9048 ( .ZN(net_14041), .A2(net_12081), .A1(net_10569) );
INV_X2 inst_19113 ( .ZN(net_4456), .A(net_4455) );
NOR3_X2 inst_2716 ( .ZN(net_13466), .A1(net_10342), .A3(net_9036), .A2(net_8620) );
INV_X4 inst_17529 ( .ZN(net_1176), .A(net_412) );
NOR2_X4 inst_3228 ( .ZN(net_7146), .A1(net_2546), .A2(net_1485) );
NAND2_X2 inst_9212 ( .ZN(net_13043), .A2(net_11287), .A1(net_9360) );
OAI21_X2 inst_2124 ( .A(net_12546), .ZN(net_10014), .B1(net_6855), .B2(net_4523) );
AND3_X4 inst_21122 ( .ZN(net_12570), .A3(net_12569), .A2(net_11348), .A1(net_3664) );
INV_X4 inst_13268 ( .ZN(net_12594), .A(net_12593) );
INV_X4 inst_17095 ( .ZN(net_9342), .A(net_6028) );
OAI21_X4 inst_1435 ( .B2(net_19929), .B1(net_19928), .ZN(net_15928), .A(net_15633) );
NAND2_X2 inst_11582 ( .A1(net_3904), .ZN(net_2725), .A2(net_2042) );
NOR2_X2 inst_3746 ( .ZN(net_10549), .A2(net_8672), .A1(net_7940) );
INV_X4 inst_15610 ( .ZN(net_13556), .A(net_10383) );
INV_X8 inst_12288 ( .ZN(net_1836), .A(net_845) );
NAND2_X2 inst_10810 ( .ZN(net_5528), .A2(net_5527), .A1(net_538) );
NOR2_X2 inst_4121 ( .ZN(net_7036), .A1(net_7035), .A2(net_4767) );
NOR3_X2 inst_2640 ( .A3(net_20102), .A1(net_20101), .ZN(net_18957), .A2(net_13921) );
CLKBUF_X2 inst_21468 ( .A(net_21294), .Z(net_21340) );
INV_X4 inst_16588 ( .A(net_5358), .ZN(net_1146) );
INV_X4 inst_12732 ( .ZN(net_17683), .A(net_17662) );
NAND2_X2 inst_8162 ( .ZN(net_17972), .A1(net_17925), .A2(net_17406) );
INV_X4 inst_18184 ( .A(net_21161), .ZN(net_615) );
NAND2_X2 inst_7908 ( .ZN(net_18469), .A2(net_18389), .A1(net_18327) );
NOR2_X2 inst_4448 ( .A1(net_5435), .A2(net_5232), .ZN(net_4775) );
INV_X4 inst_17042 ( .ZN(net_1085), .A(net_1011) );
CLKBUF_X2 inst_22130 ( .A(net_22001), .Z(net_22002) );
INV_X4 inst_17642 ( .ZN(net_1545), .A(net_284) );
INV_X2 inst_18941 ( .ZN(net_5802), .A(net_5801) );
NOR2_X2 inst_4784 ( .ZN(net_3881), .A2(net_2130), .A1(net_222) );
DFF_X1 inst_19927 ( .QN(net_21108), .D(net_10154), .CK(net_22465) );
INV_X4 inst_17998 ( .A(net_21201), .ZN(net_89) );
INV_X4 inst_15155 ( .ZN(net_14511), .A(net_12784) );
INV_X2 inst_19625 ( .A(net_21237), .ZN(net_119) );
NAND2_X4 inst_7207 ( .ZN(net_12945), .A1(net_8083), .A2(net_5008) );
INV_X8 inst_12256 ( .ZN(net_3797), .A(net_2522) );
AOI211_X2 inst_21054 ( .ZN(net_11782), .A(net_11781), .B(net_10284), .C1(net_9762), .C2(net_4402) );
INV_X4 inst_14716 ( .ZN(net_6436), .A(net_4196) );
NOR2_X4 inst_3321 ( .ZN(net_1042), .A1(net_507), .A2(net_129) );
INV_X4 inst_16464 ( .ZN(net_6091), .A(net_5459) );
XNOR2_X2 inst_333 ( .B(net_21184), .ZN(net_16995), .A(net_16994) );
NAND2_X4 inst_7684 ( .ZN(net_1131), .A1(net_330), .A2(net_136) );
NAND3_X2 inst_5988 ( .ZN(net_19203), .A2(net_14536), .A1(net_13344), .A3(net_12950) );
NAND2_X2 inst_8368 ( .A1(net_20585), .ZN(net_19048), .A2(net_17370) );
INV_X4 inst_18069 ( .A(net_21216), .ZN(net_168) );
NAND4_X2 inst_5279 ( .ZN(net_20828), .A2(net_20183), .A1(net_20182), .A4(net_14570), .A3(net_7297) );
NAND2_X2 inst_11934 ( .A1(net_2246), .ZN(net_1884), .A2(net_1119) );
NAND2_X2 inst_11394 ( .A1(net_6089), .ZN(net_4857), .A2(net_3497) );
NAND2_X2 inst_9335 ( .ZN(net_12294), .A1(net_10956), .A2(net_8956) );
NAND2_X2 inst_10953 ( .ZN(net_5093), .A2(net_3415), .A1(net_2533) );
DFF_X1 inst_19898 ( .D(net_16875), .CK(net_21588), .Q(x480) );
NAND2_X2 inst_10897 ( .ZN(net_5394), .A2(net_5393), .A1(net_955) );
NOR3_X2 inst_2764 ( .ZN(net_10458), .A1(net_6722), .A3(net_6467), .A2(net_5132) );
NAND3_X2 inst_6246 ( .ZN(net_13151), .A2(net_13150), .A3(net_13149), .A1(net_5425) );
INV_X4 inst_13755 ( .ZN(net_7617), .A(net_7616) );
INV_X4 inst_17722 ( .A(net_965), .ZN(net_190) );
NAND2_X2 inst_11065 ( .A2(net_5872), .ZN(net_4524), .A1(net_1988) );
NAND3_X2 inst_6155 ( .ZN(net_13670), .A3(net_13669), .A1(net_8420), .A2(net_3547) );
NAND3_X2 inst_5774 ( .ZN(net_15892), .A1(net_15412), .A3(net_15171), .A2(net_13866) );
CLKBUF_X2 inst_22766 ( .A(net_22637), .Z(net_22638) );
AOI21_X2 inst_20757 ( .B1(net_20486), .ZN(net_11206), .B2(net_9512), .A(net_4897) );
NAND2_X2 inst_9664 ( .ZN(net_10322), .A1(net_8117), .A2(net_7742) );
NAND2_X2 inst_8719 ( .A1(net_21220), .ZN(net_16179), .A2(net_15956) );
NAND2_X2 inst_11610 ( .A2(net_2727), .ZN(net_2612), .A1(net_1329) );
INV_X2 inst_19579 ( .A(net_2964), .ZN(net_494) );
CLKBUF_X2 inst_21394 ( .A(net_21248), .Z(net_21266) );
NOR2_X4 inst_3178 ( .ZN(net_4277), .A1(net_2208), .A2(net_703) );
NOR2_X2 inst_4203 ( .ZN(net_14881), .A2(net_6683), .A1(net_1790) );
NAND2_X2 inst_9972 ( .ZN(net_8887), .A1(net_8886), .A2(net_8885) );
NOR2_X4 inst_2840 ( .ZN(net_14768), .A2(net_14135), .A1(net_7889) );
AND2_X2 inst_21327 ( .ZN(net_5624), .A1(net_5623), .A2(net_5362) );
INV_X4 inst_16313 ( .ZN(net_3725), .A(net_1323) );
INV_X4 inst_12521 ( .ZN(net_18504), .A(net_18503) );
NAND2_X2 inst_10939 ( .A1(net_12070), .ZN(net_5185), .A2(net_5184) );
AOI21_X4 inst_20129 ( .B2(net_19940), .B1(net_19939), .A(net_16210), .ZN(net_16143) );
INV_X4 inst_14214 ( .ZN(net_19379), .A(net_8398) );
NOR3_X2 inst_2781 ( .A2(net_14151), .A1(net_8399), .ZN(net_6529), .A3(net_6528) );
NAND2_X2 inst_9544 ( .A1(net_11678), .ZN(net_11052), .A2(net_9222) );
INV_X4 inst_13190 ( .ZN(net_20048), .A(net_13533) );
CLKBUF_X2 inst_22098 ( .A(net_21909), .Z(net_21970) );
CLKBUF_X2 inst_22618 ( .A(net_22489), .Z(net_22490) );
NAND2_X2 inst_11043 ( .ZN(net_9963), .A1(net_9131), .A2(net_4722) );
INV_X4 inst_18262 ( .ZN(net_19636), .A(net_19432) );
INV_X4 inst_12780 ( .ZN(net_18420), .A(net_17307) );
OAI211_X2 inst_2402 ( .ZN(net_15870), .C1(net_15869), .B(net_15341), .C2(net_14240), .A(net_6978) );
INV_X4 inst_18245 ( .A(net_21118), .ZN(net_670) );
NAND2_X2 inst_8877 ( .ZN(net_19559), .A1(net_15245), .A2(net_14750) );
NOR3_X4 inst_2616 ( .A3(net_19271), .A1(net_19270), .ZN(net_19013), .A2(net_5323) );
INV_X4 inst_17701 ( .ZN(net_1740), .A(net_307) );
INV_X4 inst_14627 ( .A(net_5590), .ZN(net_4397) );
NAND2_X2 inst_8095 ( .ZN(net_18126), .A1(net_18098), .A2(net_18082) );
AOI21_X2 inst_20977 ( .A(net_4840), .ZN(net_4215), .B2(net_4214), .B1(net_1392) );
DFF_X1 inst_19854 ( .D(net_17153), .CK(net_21600), .Q(x708) );
OAI21_X2 inst_2113 ( .ZN(net_10036), .B2(net_5613), .B1(net_4988), .A(net_948) );
NAND4_X4 inst_5249 ( .ZN(net_20715), .A4(net_8825), .A2(net_8787), .A1(net_8329), .A3(net_5710) );
OAI21_X2 inst_1820 ( .A(net_14687), .ZN(net_14158), .B2(net_10528), .B1(net_8908) );
INV_X4 inst_15674 ( .ZN(net_19805), .A(net_3246) );
NAND2_X2 inst_8253 ( .ZN(net_17709), .A2(net_17708), .A1(net_17201) );
NAND2_X4 inst_6998 ( .ZN(net_17344), .A1(net_16728), .A2(net_16573) );
NAND3_X2 inst_6065 ( .ZN(net_20252), .A3(net_19831), .A1(net_19830), .A2(net_7967) );
NOR2_X2 inst_4729 ( .ZN(net_5434), .A1(net_3131), .A2(net_3026) );
OAI21_X2 inst_2271 ( .A(net_14458), .ZN(net_7141), .B2(net_7140), .B1(net_5560) );
NAND3_X2 inst_6209 ( .ZN(net_13277), .A3(net_13173), .A2(net_10608), .A1(net_10020) );
NAND2_X2 inst_7793 ( .ZN(net_18710), .A2(net_18666), .A1(net_17075) );
INV_X4 inst_16119 ( .ZN(net_3546), .A(net_1490) );
NAND2_X2 inst_10314 ( .ZN(net_9375), .A1(net_7975), .A2(net_7846) );
NOR2_X2 inst_3779 ( .A2(net_11979), .ZN(net_11520), .A1(net_10141) );
AOI21_X4 inst_20157 ( .ZN(net_15710), .B2(net_14979), .A(net_11103), .B1(net_1915) );
AOI21_X2 inst_20609 ( .ZN(net_13717), .B2(net_10848), .B1(net_9313), .A(net_7777) );
NAND2_X2 inst_11644 ( .ZN(net_2615), .A2(net_1058), .A1(net_86) );
SDFF_X2 inst_697 ( .Q(net_20923), .SI(net_18848), .SE(net_18847), .D(net_351), .CK(net_21298) );
NAND2_X2 inst_11150 ( .A2(net_7395), .ZN(net_4600), .A1(net_2195) );
INV_X4 inst_14035 ( .ZN(net_7475), .A(net_5134) );
NAND4_X4 inst_5159 ( .A4(net_18916), .A1(net_18915), .ZN(net_18617), .A3(net_15578), .A2(net_13801) );
INV_X1 inst_19761 ( .A(net_3136), .ZN(net_2086) );
NAND2_X2 inst_10350 ( .ZN(net_12236), .A2(net_7494), .A1(net_532) );
INV_X2 inst_18756 ( .A(net_10754), .ZN(net_7645) );
NAND2_X4 inst_7527 ( .ZN(net_2901), .A1(net_2252), .A2(net_2012) );
INV_X4 inst_13941 ( .ZN(net_6818), .A(net_6817) );
NAND2_X2 inst_11512 ( .ZN(net_3003), .A1(net_3002), .A2(net_1899) );
AOI21_X2 inst_20879 ( .B1(net_9579), .B2(net_9558), .ZN(net_8435), .A(net_5379) );
CLKBUF_X2 inst_22258 ( .A(net_22129), .Z(net_22130) );
AND2_X2 inst_21274 ( .ZN(net_20228), .A1(net_14509), .A2(net_11901) );
INV_X8 inst_12307 ( .ZN(net_11297), .A(net_4874) );
INV_X2 inst_19547 ( .ZN(net_1668), .A(net_920) );
INV_X2 inst_19200 ( .ZN(net_20023), .A(net_2514) );
NAND2_X2 inst_8758 ( .A1(net_16743), .ZN(net_15908), .A2(net_15515) );
INV_X4 inst_12975 ( .ZN(net_16655), .A(net_16510) );
INV_X4 inst_17252 ( .ZN(net_10667), .A(net_117) );
INV_X4 inst_14853 ( .ZN(net_3825), .A(net_3824) );
INV_X4 inst_13972 ( .ZN(net_7942), .A(net_6664) );
INV_X4 inst_16279 ( .ZN(net_1342), .A(net_732) );
INV_X4 inst_15165 ( .ZN(net_11860), .A(net_4348) );
INV_X4 inst_14198 ( .ZN(net_5969), .A(net_5968) );
INV_X4 inst_16656 ( .ZN(net_9421), .A(net_6856) );
OAI21_X2 inst_2004 ( .ZN(net_20822), .A(net_10667), .B2(net_7471), .B1(net_4192) );
INV_X4 inst_15894 ( .ZN(net_2617), .A(net_1775) );
XNOR2_X2 inst_220 ( .B(net_21132), .A(net_19442), .ZN(net_17511) );
AOI22_X2 inst_20008 ( .ZN(net_12853), .A1(net_12852), .A2(net_12851), .B2(net_6952), .B1(net_1986) );
XNOR2_X2 inst_245 ( .B(net_21114), .ZN(net_17318), .A(net_16984) );
NAND2_X4 inst_6991 ( .A2(net_19866), .A1(net_19865), .ZN(net_17513) );
NAND2_X2 inst_9779 ( .A1(net_11440), .ZN(net_9770), .A2(net_7592) );
CLKBUF_X2 inst_22858 ( .A(net_21972), .Z(net_22730) );
INV_X4 inst_15584 ( .A(net_16035), .ZN(net_2266) );
NOR2_X2 inst_4111 ( .ZN(net_19589), .A2(net_7068), .A1(net_5646) );
CLKBUF_X2 inst_22888 ( .A(net_22759), .Z(net_22760) );
INV_X2 inst_19728 ( .A(net_20800), .ZN(net_20799) );
INV_X2 inst_19146 ( .ZN(net_4097), .A(net_4096) );
NAND2_X2 inst_8388 ( .ZN(net_19158), .A2(net_17415), .A1(net_16596) );
INV_X4 inst_18164 ( .A(net_21068), .ZN(net_415) );
INV_X4 inst_16867 ( .ZN(net_6930), .A(net_4211) );
NAND2_X2 inst_8768 ( .ZN(net_20750), .A1(net_15876), .A2(net_15622) );
AOI21_X2 inst_20772 ( .A(net_10947), .ZN(net_10642), .B1(net_10641), .B2(net_6869) );
XNOR2_X2 inst_147 ( .ZN(net_18040), .A(net_18010), .B(net_17276) );
XNOR2_X2 inst_313 ( .B(net_20526), .ZN(net_17081), .A(net_16681) );
OAI21_X2 inst_1676 ( .A(net_16743), .ZN(net_15544), .B2(net_14595), .B1(net_13113) );
NOR2_X2 inst_4170 ( .A1(net_20537), .ZN(net_8159), .A2(net_4479) );
NAND2_X2 inst_8480 ( .A1(net_20516), .A2(net_17007), .ZN(net_17005) );
SDFF_X2 inst_1041 ( .QN(net_21034), .D(net_518), .SE(net_263), .CK(net_21950), .SI(x2420) );
OAI21_X2 inst_2086 ( .ZN(net_10399), .A(net_10398), .B2(net_7085), .B1(net_2580) );
INV_X4 inst_17964 ( .A(net_21230), .ZN(net_3867) );
INV_X4 inst_12918 ( .ZN(net_16919), .A(net_16665) );
NAND2_X2 inst_8743 ( .ZN(net_19988), .A1(net_15744), .A2(net_15653) );
NAND2_X2 inst_8570 ( .ZN(net_16737), .A1(net_16436), .A2(net_16416) );
NAND2_X2 inst_8195 ( .A2(net_20775), .ZN(net_17892), .A1(net_17881) );
INV_X4 inst_12789 ( .A(net_17293), .ZN(net_17292) );
AOI21_X2 inst_20572 ( .B1(net_19410), .ZN(net_14133), .B2(net_10031), .A(net_7687) );
XNOR2_X2 inst_553 ( .A(net_21121), .ZN(net_10801), .B(net_742) );
NAND2_X2 inst_9271 ( .ZN(net_15029), .A2(net_10904), .A1(net_7394) );
NOR2_X4 inst_3331 ( .ZN(net_2919), .A1(net_879), .A2(net_234) );
XNOR2_X2 inst_242 ( .ZN(net_17332), .A(net_16880), .B(net_240) );
NAND2_X2 inst_8950 ( .A1(net_15607), .ZN(net_14725), .A2(net_13303) );
INV_X4 inst_16843 ( .ZN(net_15690), .A(net_9656) );
INV_X4 inst_16177 ( .ZN(net_3715), .A(net_1431) );
INV_X4 inst_14592 ( .ZN(net_15995), .A(net_12208) );
CLKBUF_X2 inst_21516 ( .A(net_21387), .Z(net_21388) );
INV_X4 inst_16263 ( .ZN(net_1352), .A(net_1351) );
OR2_X2 inst_1186 ( .ZN(net_4564), .A1(net_4563), .A2(net_2117) );
CLKBUF_X2 inst_22918 ( .A(net_22416), .Z(net_22790) );
NAND2_X2 inst_9513 ( .ZN(net_20002), .A1(net_8198), .A2(net_5399) );
CLKBUF_X2 inst_22414 ( .A(net_22285), .Z(net_22286) );
NAND2_X2 inst_10542 ( .ZN(net_6789), .A1(net_6316), .A2(net_5651) );
OAI21_X2 inst_1739 ( .A(net_15217), .ZN(net_15045), .B2(net_12832), .B1(net_6409) );
INV_X4 inst_13712 ( .ZN(net_15280), .A(net_7848) );
INV_X4 inst_14863 ( .ZN(net_19553), .A(net_3765) );
INV_X8 inst_12430 ( .ZN(net_19418), .A(net_1131) );
NAND4_X2 inst_5446 ( .A2(net_20293), .ZN(net_13680), .A1(net_13679), .A4(net_13678), .A3(net_8829) );
NOR2_X2 inst_4956 ( .A1(net_10714), .ZN(net_1994), .A2(net_1637) );
NOR2_X2 inst_3609 ( .ZN(net_12418), .A2(net_12417), .A1(net_8542) );
INV_X4 inst_17631 ( .A(net_4478), .ZN(net_401) );
NAND2_X2 inst_8619 ( .A1(net_16646), .A2(net_16612), .ZN(net_16609) );
INV_X2 inst_19435 ( .ZN(net_1732), .A(net_1163) );
INV_X2 inst_19101 ( .A(net_6001), .ZN(net_4533) );
NAND3_X2 inst_6649 ( .ZN(net_8555), .A1(net_8554), .A3(net_7104), .A2(net_5339) );
INV_X4 inst_13338 ( .ZN(net_14407), .A(net_11108) );
INV_X2 inst_19189 ( .ZN(net_6332), .A(net_4675) );
INV_X4 inst_16809 ( .ZN(net_2994), .A(net_1617) );
NAND2_X2 inst_8221 ( .ZN(net_17879), .A2(net_17659), .A1(net_17585) );
NOR3_X4 inst_2608 ( .ZN(net_20649), .A3(net_19362), .A1(net_19361), .A2(net_15713) );
NAND3_X2 inst_6008 ( .ZN(net_20621), .A1(net_12716), .A2(net_11613), .A3(net_10028) );
CLKBUF_X2 inst_22334 ( .A(net_22205), .Z(net_22206) );
NAND2_X2 inst_11840 ( .A1(net_20921), .ZN(net_10320), .A2(net_146) );
INV_X4 inst_12659 ( .ZN(net_18237), .A(net_18208) );
INV_X4 inst_15873 ( .ZN(net_19669), .A(net_1795) );
INV_X4 inst_14766 ( .ZN(net_5660), .A(net_4054) );
OAI211_X2 inst_2521 ( .ZN(net_11870), .B(net_11869), .A(net_11234), .C1(net_5865), .C2(net_2922) );
XNOR2_X2 inst_385 ( .B(net_21228), .A(net_16799), .ZN(net_16798) );
CLKBUF_X2 inst_21764 ( .A(net_21635), .Z(net_21636) );
AOI21_X2 inst_20434 ( .ZN(net_15167), .B1(net_15166), .B2(net_13915), .A(net_8837) );
INV_X4 inst_14110 ( .ZN(net_6160), .A(net_6159) );
NOR3_X2 inst_2653 ( .A3(net_20398), .A1(net_20397), .ZN(net_15477), .A2(net_10228) );
NAND2_X2 inst_11062 ( .A2(net_4681), .ZN(net_4534), .A1(net_1984) );
INV_X2 inst_19073 ( .ZN(net_4625), .A(net_4624) );
INV_X4 inst_14827 ( .ZN(net_4895), .A(net_3901) );
AOI22_X2 inst_19988 ( .ZN(net_15136), .A2(net_13321), .A1(net_12852), .B2(net_5854), .B1(net_2368) );
NAND2_X2 inst_11324 ( .A1(net_4770), .ZN(net_3752), .A2(net_3751) );
INV_X4 inst_15799 ( .ZN(net_8639), .A(net_6655) );
CLKBUF_X2 inst_21441 ( .A(net_21312), .Z(net_21313) );
NAND2_X2 inst_10696 ( .ZN(net_6070), .A2(net_4416), .A1(net_4056) );
INV_X4 inst_13150 ( .ZN(net_14899), .A(net_14392) );
CLKBUF_X2 inst_21502 ( .A(net_21373), .Z(net_21374) );
XNOR2_X2 inst_596 ( .B(net_16794), .A(net_552), .ZN(net_551) );
NOR3_X2 inst_2771 ( .ZN(net_8499), .A3(net_6848), .A2(net_6841), .A1(net_3761) );
NAND2_X2 inst_8835 ( .ZN(net_19385), .A2(net_14770), .A1(net_13189) );
NOR2_X2 inst_4687 ( .A1(net_20474), .ZN(net_3849), .A2(net_3075) );
CLKBUF_X2 inst_21967 ( .A(net_21838), .Z(net_21839) );
NAND2_X2 inst_9245 ( .ZN(net_12676), .A1(net_12675), .A2(net_12674) );
OAI21_X2 inst_1705 ( .A(net_15343), .ZN(net_15258), .B2(net_13592), .B1(net_5196) );
NAND2_X2 inst_11286 ( .ZN(net_5375), .A2(net_4092), .A1(net_1376) );
NOR2_X2 inst_4664 ( .ZN(net_8322), .A2(net_6455), .A1(net_3278) );
INV_X4 inst_17388 ( .ZN(net_1216), .A(net_335) );
INV_X4 inst_14601 ( .ZN(net_16546), .A(net_4447) );
NOR2_X2 inst_5003 ( .A1(net_20568), .ZN(net_1391), .A2(net_1354) );
INV_X4 inst_15841 ( .A(net_2731), .ZN(net_1846) );
INV_X8 inst_12215 ( .ZN(net_7549), .A(net_6154) );
INV_X4 inst_15454 ( .ZN(net_2487), .A(net_2486) );
NAND3_X2 inst_5798 ( .ZN(net_15718), .A2(net_15112), .A1(net_14133), .A3(net_14105) );
NOR2_X4 inst_3253 ( .ZN(net_6437), .A1(net_2275), .A2(net_498) );
NAND4_X2 inst_5321 ( .A3(net_19506), .A1(net_19505), .ZN(net_18958), .A2(net_14999), .A4(net_14699) );
INV_X4 inst_16378 ( .A(net_10093), .ZN(net_1688) );
INV_X4 inst_14250 ( .ZN(net_7308), .A(net_4458) );
NOR2_X2 inst_4596 ( .ZN(net_8483), .A2(net_3841), .A1(net_388) );
NAND2_X2 inst_9013 ( .ZN(net_19813), .A1(net_13091), .A2(net_12664) );
NAND2_X2 inst_8427 ( .ZN(net_19159), .A2(net_17416), .A1(net_16721) );
INV_X4 inst_18316 ( .A(net_20520), .ZN(net_20518) );
XNOR2_X2 inst_637 ( .B(net_552), .ZN(net_427), .A(net_426) );
INV_X2 inst_18649 ( .ZN(net_11895), .A(net_9227) );
INV_X4 inst_13572 ( .ZN(net_12315), .A(net_9128) );
INV_X4 inst_17211 ( .ZN(net_6028), .A(net_493) );
INV_X2 inst_18834 ( .ZN(net_6763), .A(net_6762) );
INV_X4 inst_16024 ( .A(net_4039), .ZN(net_1892) );
INV_X4 inst_13148 ( .ZN(net_14907), .A(net_14411) );
NAND2_X4 inst_7033 ( .ZN(net_18326), .A1(net_16449), .A2(net_16417) );
INV_X2 inst_18496 ( .ZN(net_12312), .A(net_12311) );
INV_X4 inst_15787 ( .A(net_3133), .ZN(net_1908) );
NAND2_X2 inst_8152 ( .ZN(net_18009), .A1(net_17955), .A2(net_17930) );
NAND2_X2 inst_10159 ( .ZN(net_9732), .A2(net_5050), .A1(net_154) );
NOR2_X2 inst_4762 ( .ZN(net_7072), .A1(net_6377), .A2(net_2987) );
XNOR2_X2 inst_164 ( .B(net_21113), .ZN(net_17849), .A(net_17676) );
NAND2_X2 inst_8534 ( .ZN(net_16861), .A2(net_16670), .A1(net_16668) );
CLKBUF_X2 inst_21879 ( .A(net_21696), .Z(net_21751) );
NAND2_X2 inst_8467 ( .ZN(net_17047), .A2(net_17046), .A1(net_7774) );
CLKBUF_X2 inst_21448 ( .A(net_21273), .Z(net_21320) );
OAI21_X2 inst_2305 ( .B2(net_6537), .ZN(net_5854), .A(net_5853), .B1(net_5852) );
NAND2_X2 inst_10079 ( .ZN(net_13306), .A2(net_7864), .A1(net_5818) );
OAI21_X2 inst_2150 ( .A(net_9795), .ZN(net_9308), .B2(net_3259), .B1(net_1913) );
NAND2_X2 inst_10930 ( .A1(net_5959), .ZN(net_5216), .A2(net_5215) );
NAND2_X2 inst_9770 ( .A1(net_10539), .ZN(net_9800), .A2(net_6986) );
SDFF_X2 inst_946 ( .QN(net_21091), .D(net_584), .SE(net_253), .CK(net_21796), .SI(x1526) );
OAI21_X2 inst_2260 ( .A(net_8667), .ZN(net_7169), .B2(net_7168), .B1(net_4187) );
INV_X2 inst_18804 ( .ZN(net_7410), .A(net_7409) );
NAND2_X2 inst_8141 ( .A1(net_20234), .ZN(net_18026), .A2(net_17859) );
INV_X4 inst_13276 ( .ZN(net_13469), .A(net_12455) );
INV_X2 inst_19048 ( .ZN(net_5915), .A(net_4744) );
NAND2_X2 inst_11700 ( .ZN(net_2306), .A2(net_2305), .A1(net_61) );
NOR2_X2 inst_4625 ( .ZN(net_3604), .A1(net_2285), .A2(net_439) );
NAND2_X4 inst_6951 ( .ZN(net_17602), .A2(net_17147), .A1(net_17009) );
NOR2_X2 inst_3922 ( .A1(net_13076), .ZN(net_10276), .A2(net_8782) );
OAI21_X2 inst_2053 ( .ZN(net_10843), .A(net_7609), .B2(net_6461), .B1(net_4032) );
INV_X2 inst_19654 ( .A(net_20207), .ZN(net_20206) );
NAND2_X2 inst_10539 ( .ZN(net_8114), .A1(net_5005), .A2(net_1085) );
NAND2_X2 inst_10038 ( .ZN(net_13129), .A2(net_8721), .A1(net_1657) );
OAI222_X2 inst_1325 ( .ZN(net_10507), .C1(net_8676), .A2(net_7656), .C2(net_7091), .B1(net_6520), .A1(net_4502), .B2(net_3546) );
CLKBUF_X2 inst_21894 ( .A(net_21435), .Z(net_21766) );
INV_X2 inst_19018 ( .ZN(net_4979), .A(net_4978) );
NAND2_X2 inst_8859 ( .ZN(net_15347), .A1(net_14793), .A2(net_14427) );
INV_X4 inst_17861 ( .ZN(net_1815), .A(net_910) );
CLKBUF_X2 inst_22747 ( .A(net_21639), .Z(net_22619) );
INV_X4 inst_13503 ( .ZN(net_9423), .A(net_9422) );
INV_X4 inst_16684 ( .ZN(net_10323), .A(net_7436) );
NAND2_X4 inst_6873 ( .A2(net_19138), .A1(net_19137), .ZN(net_18312) );
INV_X4 inst_14087 ( .A(net_6210), .ZN(net_6209) );
NOR2_X4 inst_3312 ( .ZN(net_1194), .A2(net_322), .A1(net_108) );
INV_X4 inst_15432 ( .ZN(net_2505), .A(net_2504) );
NAND2_X2 inst_9207 ( .A1(net_15104), .ZN(net_13056), .A2(net_11275) );
INV_X4 inst_17138 ( .ZN(net_14949), .A(net_11032) );
NAND2_X1 inst_12143 ( .ZN(net_16903), .A1(net_16902), .A2(net_16901) );
OR2_X2 inst_1235 ( .A2(net_7780), .ZN(net_1589), .A1(net_168) );
INV_X4 inst_16948 ( .ZN(net_5727), .A(net_1259) );
INV_X4 inst_16760 ( .ZN(net_2554), .A(net_1036) );
INV_X4 inst_15015 ( .ZN(net_13873), .A(net_3379) );
INV_X4 inst_14107 ( .ZN(net_7555), .A(net_6165) );
INV_X4 inst_13143 ( .ZN(net_15073), .A(net_14651) );
INV_X4 inst_16115 ( .ZN(net_2005), .A(net_1493) );
AOI21_X2 inst_20566 ( .ZN(net_19073), .B2(net_13553), .B1(net_13091), .A(net_7047) );
NOR2_X2 inst_3626 ( .ZN(net_20284), .A2(net_10779), .A1(net_6138) );
NOR2_X2 inst_4036 ( .A1(net_8013), .ZN(net_7938), .A2(net_7937) );
NAND4_X4 inst_5244 ( .A1(net_19891), .ZN(net_14784), .A4(net_14783), .A3(net_14782), .A2(net_14448) );
INV_X2 inst_19068 ( .ZN(net_4635), .A(net_4634) );
INV_X4 inst_14942 ( .ZN(net_6182), .A(net_5490) );
INV_X4 inst_13457 ( .ZN(net_11084), .A(net_9723) );
INV_X2 inst_18572 ( .A(net_12378), .ZN(net_10738) );
CLKBUF_X2 inst_21890 ( .A(net_21692), .Z(net_21762) );
OAI21_X2 inst_1600 ( .A(net_20960), .ZN(net_16178), .B2(net_15780), .B1(net_13118) );
NOR2_X4 inst_2850 ( .A1(net_20752), .ZN(net_14817), .A2(net_12784) );
INV_X4 inst_14884 ( .ZN(net_4659), .A(net_3670) );
INV_X4 inst_14268 ( .A(net_8019), .ZN(net_7599) );
NAND4_X4 inst_5163 ( .ZN(net_18112), .A4(net_18068), .A1(net_18063), .A2(net_15678), .A3(net_12207) );
NAND2_X2 inst_9590 ( .ZN(net_10890), .A2(net_7345), .A1(net_60) );
NAND2_X4 inst_7677 ( .ZN(net_1288), .A2(net_814), .A1(net_258) );
SDFF_X2 inst_849 ( .Q(net_21242), .SI(net_17309), .SE(net_125), .CK(net_21548), .D(x6655) );
NAND2_X4 inst_7393 ( .ZN(net_6914), .A1(net_4125), .A2(net_3356) );
INV_X1 inst_19764 ( .A(net_2144), .ZN(net_1577) );
INV_X4 inst_16998 ( .A(net_1823), .ZN(net_1047) );
CLKBUF_X2 inst_22591 ( .A(net_22462), .Z(net_22463) );
XOR2_X2 inst_3 ( .Z(net_18220), .A(net_18093), .B(net_4439) );
INV_X4 inst_14517 ( .A(net_11808), .ZN(net_4811) );
NOR2_X4 inst_3060 ( .ZN(net_7954), .A1(net_4952), .A2(net_4951) );
AOI21_X2 inst_20416 ( .ZN(net_15274), .B1(net_14689), .B2(net_13899), .A(net_11516) );
NAND3_X2 inst_5812 ( .ZN(net_15645), .A3(net_14373), .A1(net_13821), .A2(net_11486) );
NAND2_X2 inst_10041 ( .A2(net_11374), .A1(net_10207), .ZN(net_8716) );
XNOR2_X2 inst_566 ( .B(net_9255), .ZN(net_651), .A(net_650) );
OAI21_X4 inst_1399 ( .A(net_20896), .B2(net_19520), .B1(net_19519), .ZN(net_16244) );
INV_X2 inst_19180 ( .ZN(net_3786), .A(net_3785) );
INV_X8 inst_12301 ( .ZN(net_5043), .A(net_1176) );
NAND2_X2 inst_10613 ( .ZN(net_7848), .A2(net_6573), .A1(net_1714) );
NOR2_X2 inst_4357 ( .ZN(net_5581), .A2(net_5139), .A1(net_1522) );
INV_X4 inst_16456 ( .ZN(net_8138), .A(net_112) );
NOR2_X2 inst_4327 ( .A1(net_12231), .ZN(net_5809), .A2(net_5808) );
INV_X4 inst_16189 ( .ZN(net_15840), .A(net_15312) );
NAND2_X2 inst_11375 ( .ZN(net_18979), .A2(net_2952), .A1(net_2870) );
CLKBUF_X2 inst_21937 ( .A(net_21808), .Z(net_21809) );
NAND2_X2 inst_10419 ( .A1(net_14755), .ZN(net_13787), .A2(net_5552) );
OAI21_X2 inst_2333 ( .ZN(net_4688), .A(net_4687), .B1(net_3607), .B2(net_1876) );
INV_X4 inst_14844 ( .ZN(net_9072), .A(net_3848) );
CLKBUF_X2 inst_21800 ( .A(net_21302), .Z(net_21672) );
INV_X4 inst_15291 ( .ZN(net_5104), .A(net_2717) );
NAND2_X4 inst_7047 ( .A2(net_19238), .A1(net_19237), .ZN(net_16801) );
INV_X2 inst_19713 ( .A(net_20764), .ZN(net_20763) );
NAND2_X2 inst_11345 ( .A2(net_4029), .ZN(net_3657), .A1(net_1182) );
INV_X2 inst_19596 ( .A(net_798), .ZN(net_201) );
NAND3_X2 inst_5928 ( .ZN(net_14938), .A2(net_12900), .A3(net_12733), .A1(net_7899) );
NOR2_X2 inst_5056 ( .A1(net_20558), .ZN(net_1083), .A2(net_61) );
NAND4_X2 inst_5370 ( .ZN(net_15234), .A1(net_14188), .A4(net_14017), .A2(net_12277), .A3(net_11777) );
OAI21_X2 inst_1732 ( .ZN(net_15076), .B2(net_12896), .B1(net_10222), .A(net_238) );
NAND2_X4 inst_7256 ( .ZN(net_7977), .A1(net_6616), .A2(net_6221) );
INV_X2 inst_18697 ( .ZN(net_8336), .A(net_8335) );
NAND3_X2 inst_6119 ( .A2(net_14711), .ZN(net_13861), .A3(net_13278), .A1(net_11512) );
INV_X4 inst_15461 ( .ZN(net_10119), .A(net_7116) );
CLKBUF_X2 inst_22358 ( .A(net_22229), .Z(net_22230) );
NAND3_X2 inst_6269 ( .ZN(net_12959), .A2(net_12958), .A3(net_12957), .A1(net_6790) );
INV_X4 inst_13247 ( .ZN(net_19490), .A(net_11930) );
NAND2_X2 inst_9481 ( .A1(net_14086), .ZN(net_11455), .A2(net_11454) );
NAND3_X2 inst_5858 ( .ZN(net_15399), .A3(net_13973), .A1(net_12719), .A2(net_7582) );
CLKBUF_X2 inst_21813 ( .A(net_21684), .Z(net_21685) );
NOR2_X4 inst_3069 ( .A1(net_7489), .ZN(net_5948), .A2(net_4389) );
NOR2_X2 inst_3631 ( .ZN(net_20195), .A2(net_13119), .A1(net_8669) );
AOI21_X2 inst_20956 ( .ZN(net_5337), .B2(net_4184), .A(net_4174), .B1(net_112) );
OR2_X4 inst_1101 ( .ZN(net_6497), .A2(net_2149), .A1(net_85) );
NAND2_X2 inst_8596 ( .A2(net_19437), .ZN(net_16687), .A1(net_16569) );
INV_X4 inst_17712 ( .ZN(net_2077), .A(net_218) );
NAND3_X2 inst_6652 ( .A2(net_9072), .ZN(net_8547), .A3(net_8546), .A1(net_8033) );
NOR2_X4 inst_2950 ( .ZN(net_8148), .A2(net_4853), .A1(net_154) );
AOI21_X4 inst_20213 ( .B1(net_19247), .ZN(net_19074), .B2(net_10383), .A(net_9722) );
NAND2_X2 inst_8584 ( .ZN(net_16717), .A2(net_16716), .A1(net_16665) );
INV_X4 inst_15777 ( .A(net_2795), .ZN(net_1914) );
INV_X4 inst_17673 ( .A(net_6692), .ZN(net_243) );
NAND2_X2 inst_12013 ( .ZN(net_2240), .A2(net_1699), .A1(net_133) );
INV_X2 inst_19273 ( .ZN(net_3005), .A(net_3004) );
INV_X4 inst_15572 ( .ZN(net_5677), .A(net_1224) );
OAI211_X2 inst_2451 ( .C1(net_20041), .ZN(net_14575), .C2(net_13619), .B(net_11313), .A(net_10334) );
INV_X4 inst_16326 ( .ZN(net_11148), .A(net_7394) );
OR2_X2 inst_1202 ( .A1(net_10031), .ZN(net_3743), .A2(net_3742) );
CLKBUF_X2 inst_22561 ( .A(net_22432), .Z(net_22433) );
CLKBUF_X2 inst_22474 ( .A(net_22197), .Z(net_22346) );
INV_X4 inst_15106 ( .A(net_15099), .ZN(net_8264) );
AOI21_X2 inst_20590 ( .ZN(net_20422), .B1(net_20283), .B2(net_13938), .A(net_9567) );
NAND2_X4 inst_7020 ( .ZN(net_17245), .A1(net_16568), .A2(net_16453) );
OAI21_X2 inst_2227 ( .ZN(net_8461), .B1(net_8460), .A(net_5093), .B2(net_3128) );
XNOR2_X2 inst_660 ( .B(net_16462), .ZN(net_13294), .A(net_738) );
OAI211_X2 inst_2490 ( .ZN(net_13166), .B(net_13165), .C2(net_13164), .A(net_12800), .C1(net_7903) );
INV_X4 inst_14526 ( .ZN(net_20115), .A(net_4767) );
AND4_X4 inst_21091 ( .ZN(net_13337), .A4(net_11555), .A3(net_8916), .A2(net_8206), .A1(net_5524) );
NAND2_X2 inst_10150 ( .A1(net_11045), .ZN(net_8291), .A2(net_5053) );
OAI21_X2 inst_1576 ( .A(net_20928), .B2(net_19951), .B1(net_19950), .ZN(net_16326) );
AOI21_X4 inst_20120 ( .ZN(net_19168), .B1(net_18993), .A(net_14482), .B2(net_14033) );
INV_X4 inst_16712 ( .ZN(net_1060), .A(net_1059) );
NAND2_X2 inst_11532 ( .A2(net_7538), .ZN(net_2931), .A1(net_2617) );
INV_X2 inst_19535 ( .ZN(net_979), .A(net_978) );
NAND3_X2 inst_5642 ( .ZN(net_17459), .A3(net_17044), .A2(net_16192), .A1(net_13825) );
INV_X4 inst_16397 ( .ZN(net_15747), .A(net_14490) );
NAND2_X4 inst_7459 ( .A1(net_19952), .ZN(net_2818), .A2(net_2314) );
NAND2_X2 inst_11898 ( .ZN(net_2986), .A1(net_1582), .A2(net_1166) );
NAND2_X2 inst_8390 ( .A1(net_20633), .ZN(net_19763), .A2(net_16902) );
INV_X4 inst_17141 ( .ZN(net_1058), .A(net_167) );
NAND3_X2 inst_6659 ( .ZN(net_8453), .A2(net_6426), .A3(net_5584), .A1(net_4484) );
INV_X2 inst_18859 ( .ZN(net_6329), .A(net_6328) );
NAND2_X2 inst_7828 ( .A1(net_21162), .ZN(net_18638), .A2(net_18607) );
NOR2_X2 inst_4368 ( .ZN(net_19888), .A1(net_3901), .A2(net_3521) );
DFF_X1 inst_19822 ( .D(net_17682), .CK(net_21368), .Q(x132) );
NAND2_X2 inst_10331 ( .A2(net_20778), .ZN(net_9230), .A1(net_6951) );
CLKBUF_X2 inst_21752 ( .A(net_21623), .Z(net_21624) );
NAND2_X2 inst_11137 ( .ZN(net_9707), .A2(net_7144), .A1(net_5591) );
INV_X4 inst_17604 ( .ZN(net_374), .A(net_193) );
AOI21_X2 inst_20476 ( .B2(net_19171), .B1(net_19170), .ZN(net_14948), .A(net_12203) );
OR2_X2 inst_1147 ( .ZN(net_20144), .A1(net_13538), .A2(net_11836) );
AOI21_X2 inst_20692 ( .ZN(net_12205), .A(net_10417), .B2(net_8388), .B1(net_4816) );
OAI21_X2 inst_1768 ( .ZN(net_14697), .B2(net_12064), .B1(net_7022), .A(net_6528) );
INV_X4 inst_18308 ( .A(net_20501), .ZN(net_20498) );
NAND3_X2 inst_6410 ( .ZN(net_11957), .A3(net_11956), .A1(net_9881), .A2(net_7868) );
INV_X4 inst_12865 ( .ZN(net_16991), .A(net_16990) );
NOR2_X4 inst_2917 ( .ZN(net_10269), .A1(net_6154), .A2(net_107) );
INV_X2 inst_18953 ( .A(net_8696), .ZN(net_5552) );
OAI21_X4 inst_1408 ( .A(net_20920), .B2(net_20417), .B1(net_20416), .ZN(net_16181) );
AOI211_X2 inst_21083 ( .B(net_6002), .ZN(net_5262), .A(net_3039), .C2(net_2852), .C1(net_2829) );
INV_X4 inst_13563 ( .A(net_13483), .ZN(net_9143) );
OAI21_X2 inst_1889 ( .B2(net_19721), .B1(net_19720), .A(net_13530), .ZN(net_13492) );
AOI21_X2 inst_20447 ( .B2(net_20727), .B1(net_20726), .ZN(net_15096), .A(net_828) );
OAI21_X2 inst_2011 ( .ZN(net_11386), .A(net_10377), .B2(net_7540), .B1(net_5088) );
INV_X4 inst_13495 ( .ZN(net_9456), .A(net_9455) );
OAI21_X2 inst_1761 ( .ZN(net_20034), .A(net_14714), .B2(net_11788), .B1(net_11657) );
INV_X4 inst_16000 ( .ZN(net_15924), .A(net_15790) );
NAND3_X2 inst_6582 ( .ZN(net_10438), .A3(net_10437), .A2(net_9633), .A1(net_6073) );
NAND2_X2 inst_9418 ( .A1(net_12866), .A2(net_12061), .ZN(net_11643) );
NAND4_X2 inst_5474 ( .ZN(net_13181), .A1(net_12444), .A2(net_11558), .A4(net_10032), .A3(net_8355) );
XNOR2_X2 inst_84 ( .ZN(net_18573), .B(net_18521), .A(net_18471) );
NAND3_X2 inst_5974 ( .ZN(net_20145), .A3(net_12291), .A1(net_8884), .A2(net_4033) );
XNOR2_X2 inst_173 ( .ZN(net_17870), .A(net_17539), .B(net_17082) );
NAND2_X4 inst_7660 ( .A2(net_20820), .ZN(net_2110), .A1(net_212) );
NAND3_X4 inst_5568 ( .ZN(net_15933), .A3(net_15246), .A2(net_14792), .A1(net_14591) );
NAND3_X2 inst_5821 ( .ZN(net_15591), .A3(net_14229), .A2(net_11605), .A1(net_11123) );
NAND2_X4 inst_7187 ( .ZN(net_19121), .A2(net_8830), .A1(net_8829) );
NAND3_X2 inst_5713 ( .ZN(net_16164), .A1(net_15914), .A3(net_15784), .A2(net_15635) );
NAND2_X2 inst_10493 ( .A1(net_12100), .ZN(net_8301), .A2(net_5095) );
NAND2_X2 inst_8723 ( .A1(net_16402), .ZN(net_16107), .A2(net_15866) );
INV_X4 inst_13047 ( .A(net_16560), .ZN(net_16497) );
OAI21_X2 inst_1943 ( .ZN(net_12715), .A(net_12714), .B2(net_9228), .B1(net_7438) );
NAND2_X2 inst_7847 ( .ZN(net_18597), .A2(net_18583), .A1(net_12085) );
NAND3_X4 inst_5573 ( .ZN(net_19190), .A1(net_15207), .A3(net_15049), .A2(net_8118) );
INV_X2 inst_18598 ( .ZN(net_9978), .A(net_9977) );
OAI21_X2 inst_1531 ( .ZN(net_18011), .B1(net_17958), .A(net_17934), .B2(net_17933) );
AOI21_X2 inst_20619 ( .ZN(net_13519), .B2(net_9032), .B1(net_8323), .A(net_855) );
NAND2_X4 inst_7640 ( .ZN(net_2275), .A2(net_1134), .A1(net_917) );
NAND2_X4 inst_7083 ( .ZN(net_19594), .A1(net_15269), .A2(net_15076) );
AOI21_X2 inst_20964 ( .B1(net_5852), .A(net_5467), .ZN(net_5307), .B2(net_1108) );
AND3_X2 inst_21142 ( .ZN(net_9051), .A1(net_7448), .A3(net_7214), .A2(net_6140) );
NAND2_X2 inst_11706 ( .ZN(net_4248), .A2(net_2278), .A1(net_1154) );
INV_X4 inst_15075 ( .A(net_15628), .ZN(net_15027) );
NOR2_X4 inst_2922 ( .ZN(net_10720), .A1(net_7902), .A2(net_6797) );
NAND2_X2 inst_11831 ( .ZN(net_1858), .A1(net_1699), .A2(net_1092) );
NAND2_X2 inst_11649 ( .ZN(net_3260), .A1(net_1681), .A2(net_1554) );
NAND2_X2 inst_10410 ( .ZN(net_14538), .A1(net_8751), .A2(net_5535) );
INV_X2 inst_18551 ( .A(net_12844), .ZN(net_10913) );
INV_X2 inst_18682 ( .ZN(net_8784), .A(net_8783) );
INV_X4 inst_16036 ( .ZN(net_2674), .A(net_2053) );
SDFF_X2 inst_1037 ( .QN(net_21101), .SE(net_2426), .D(net_1511), .CK(net_22715), .SI(x1373) );
NAND2_X2 inst_7777 ( .ZN(net_18731), .A2(net_18694), .A1(net_17869) );
NAND2_X2 inst_8652 ( .A2(net_20068), .ZN(net_16558), .A1(net_16491) );
NOR2_X2 inst_3596 ( .ZN(net_12586), .A1(net_9484), .A2(net_4152) );
OAI22_X2 inst_1250 ( .ZN(net_18675), .A2(net_18663), .B2(net_18615), .B1(net_17775), .A1(net_17756) );
NAND2_X4 inst_7071 ( .A1(net_20352), .A2(net_16394), .ZN(net_16111) );
AOI21_X2 inst_20471 ( .ZN(net_20455), .B1(net_14981), .B2(net_12839), .A(net_8628) );
NAND2_X2 inst_10240 ( .A2(net_8429), .ZN(net_8032), .A1(net_8031) );
INV_X2 inst_19028 ( .A(net_6707), .ZN(net_4905) );
AOI21_X2 inst_20640 ( .ZN(net_13268), .A(net_10290), .B2(net_9880), .B1(net_5415) );
OAI21_X2 inst_1979 ( .ZN(net_19712), .B1(net_12144), .A(net_8596), .B2(net_8229) );
XNOR2_X2 inst_364 ( .B(net_17534), .A(net_17006), .ZN(net_16873) );
NAND2_X2 inst_11586 ( .A2(net_3282), .A1(net_2980), .ZN(net_2707) );
NAND2_X2 inst_9253 ( .ZN(net_14619), .A2(net_12659), .A1(net_10229) );
NAND2_X2 inst_9283 ( .ZN(net_12547), .A1(net_12546), .A2(net_9677) );
NOR2_X4 inst_2997 ( .ZN(net_10089), .A2(net_5937), .A1(net_454) );
NOR2_X2 inst_4712 ( .ZN(net_4104), .A1(net_3151), .A2(net_3150) );
XNOR2_X2 inst_411 ( .B(net_17294), .ZN(net_16620), .A(net_16619) );
CLKBUF_X2 inst_21590 ( .A(net_21461), .Z(net_21462) );
NAND2_X2 inst_9055 ( .ZN(net_14002), .A2(net_11980), .A1(net_11979) );
NAND2_X2 inst_10380 ( .A1(net_18025), .ZN(net_7386), .A2(net_377) );
NOR2_X2 inst_4026 ( .A2(net_12908), .A1(net_10298), .ZN(net_9555) );
INV_X4 inst_14722 ( .ZN(net_15481), .A(net_14186) );
INV_X4 inst_14649 ( .ZN(net_4638), .A(net_4371) );
NAND2_X2 inst_9395 ( .A2(net_12835), .ZN(net_11704), .A1(net_8933) );
NAND2_X2 inst_11333 ( .A1(net_11311), .ZN(net_9947), .A2(net_3771) );
NAND2_X2 inst_10668 ( .ZN(net_9759), .A1(net_6706), .A2(net_3626) );
NAND2_X2 inst_11010 ( .ZN(net_4875), .A1(net_4874), .A2(net_2700) );
NOR2_X2 inst_4382 ( .ZN(net_6292), .A2(net_5234), .A1(net_2435) );
NAND2_X2 inst_10908 ( .ZN(net_13078), .A1(net_5372), .A2(net_5371) );
INV_X4 inst_14426 ( .ZN(net_10050), .A(net_5041) );
INV_X4 inst_17391 ( .ZN(net_6668), .A(net_81) );
INV_X2 inst_19708 ( .A(net_20577), .ZN(net_20576) );
INV_X4 inst_13480 ( .ZN(net_9588), .A(net_9587) );
INV_X4 inst_17941 ( .A(net_20967), .ZN(net_116) );
NAND2_X2 inst_8708 ( .A1(net_21212), .ZN(net_16276), .A2(net_16103) );
INV_X4 inst_15400 ( .ZN(net_3340), .A(net_1853) );
INV_X4 inst_13297 ( .A(net_12617), .ZN(net_12341) );
INV_X4 inst_14020 ( .ZN(net_11244), .A(net_6294) );
NAND2_X2 inst_9874 ( .ZN(net_9462), .A1(net_9461), .A2(net_9460) );
NAND3_X4 inst_5538 ( .A3(net_20187), .A1(net_20186), .ZN(net_17416), .A2(net_15438) );
XNOR2_X2 inst_61 ( .ZN(net_18822), .A(net_18766), .B(net_16618) );
XNOR2_X2 inst_203 ( .ZN(net_17609), .A(net_17280), .B(net_16857) );
NAND3_X2 inst_5834 ( .ZN(net_15513), .A2(net_14723), .A1(net_14632), .A3(net_14567) );
INV_X2 inst_19681 ( .A(net_20520), .ZN(net_20519) );
INV_X4 inst_14077 ( .ZN(net_7571), .A(net_6222) );
OR2_X2 inst_1139 ( .A1(net_15202), .ZN(net_11509), .A2(net_11508) );
NAND2_X2 inst_10597 ( .ZN(net_10524), .A2(net_6700), .A1(net_242) );
NAND2_X2 inst_8852 ( .ZN(net_15382), .A2(net_14702), .A1(net_14512) );
NOR2_X2 inst_4507 ( .ZN(net_5268), .A1(net_4211), .A2(net_4210) );
INV_X4 inst_17381 ( .ZN(net_6316), .A(net_895) );
INV_X4 inst_14558 ( .ZN(net_6030), .A(net_4570) );
NAND2_X2 inst_9968 ( .ZN(net_8893), .A1(net_7253), .A2(net_7013) );
CLKBUF_X2 inst_22057 ( .A(net_21928), .Z(net_21929) );
NAND2_X4 inst_7631 ( .ZN(net_2006), .A1(net_1513), .A2(net_1343) );
INV_X4 inst_14669 ( .ZN(net_8035), .A(net_5305) );
NAND3_X2 inst_6607 ( .ZN(net_9296), .A2(net_9295), .A3(net_9294), .A1(net_4269) );
XNOR2_X2 inst_456 ( .A(net_17144), .ZN(net_13661), .B(net_1866) );
SDFF_X2 inst_832 ( .Q(net_21141), .SI(net_17509), .SE(net_125), .CK(net_22443), .D(x3608) );
CLKBUF_X2 inst_22588 ( .A(net_22459), .Z(net_22460) );
NAND2_X2 inst_8102 ( .ZN(net_20282), .A2(net_18118), .A1(net_16965) );
XNOR2_X2 inst_275 ( .B(net_21173), .ZN(net_17190), .A(net_17189) );
NAND2_X2 inst_11492 ( .A1(net_7874), .ZN(net_3995), .A2(net_3089) );
NOR2_X2 inst_3728 ( .ZN(net_10889), .A2(net_10888), .A1(net_8553) );
NAND2_X2 inst_11576 ( .ZN(net_6464), .A2(net_4038), .A1(net_154) );
AOI21_X2 inst_20687 ( .ZN(net_12232), .B1(net_12231), .B2(net_8509), .A(net_4489) );
OAI211_X2 inst_2416 ( .C1(net_20635), .ZN(net_15485), .C2(net_15183), .A(net_10691), .B(net_8185) );
INV_X4 inst_17239 ( .ZN(net_659), .A(net_511) );
NOR2_X2 inst_3812 ( .ZN(net_9833), .A1(net_9832), .A2(net_9618) );
INV_X4 inst_17069 ( .ZN(net_2957), .A(net_1607) );
AND2_X4 inst_21245 ( .ZN(net_7080), .A2(net_2412), .A1(net_2339) );
NAND2_X2 inst_7879 ( .ZN(net_18525), .A1(net_18466), .A2(net_18441) );
NOR2_X2 inst_3959 ( .A1(net_20408), .ZN(net_8593), .A2(net_8592) );
INV_X2 inst_19354 ( .A(net_3070), .ZN(net_2815) );
NAND2_X2 inst_9839 ( .ZN(net_19029), .A2(net_9647), .A1(net_9569) );
NOR2_X2 inst_4518 ( .A1(net_10886), .A2(net_4673), .ZN(net_4152) );
NAND2_X2 inst_11185 ( .ZN(net_11174), .A1(net_4111), .A2(net_3055) );
INV_X4 inst_15415 ( .ZN(net_19960), .A(net_1845) );
NAND2_X2 inst_10348 ( .ZN(net_12480), .A2(net_4577), .A1(net_761) );
NAND2_X2 inst_9726 ( .ZN(net_14533), .A1(net_10134), .A2(net_8005) );
NAND2_X4 inst_6832 ( .ZN(net_18807), .A2(net_18729), .A1(net_18700) );
INV_X4 inst_14234 ( .ZN(net_7566), .A(net_5073) );
AOI21_X2 inst_20451 ( .ZN(net_15070), .B1(net_13544), .B2(net_13011), .A(net_7698) );
CLKBUF_X2 inst_22205 ( .A(net_22076), .Z(net_22077) );
NAND2_X2 inst_7958 ( .ZN(net_18391), .A2(net_18390), .A1(net_17155) );
NAND2_X2 inst_11237 ( .A2(net_7155), .ZN(net_3939), .A1(net_1979) );
NOR2_X4 inst_3166 ( .ZN(net_4100), .A1(net_2175), .A2(net_1821) );
INV_X2 inst_19320 ( .ZN(net_2614), .A(net_2613) );
CLKBUF_X2 inst_21874 ( .A(net_21745), .Z(net_21746) );
INV_X4 inst_18131 ( .A(net_21045), .ZN(net_743) );
INV_X4 inst_14218 ( .ZN(net_20042), .A(net_6870) );
NAND2_X4 inst_7452 ( .ZN(net_3773), .A2(net_2253), .A1(net_2108) );
INV_X4 inst_13807 ( .ZN(net_7543), .A(net_7542) );
NOR2_X2 inst_3656 ( .A2(net_15018), .ZN(net_12701), .A1(net_8842) );
INV_X4 inst_12497 ( .A(net_18645), .ZN(net_18628) );
OAI21_X2 inst_2237 ( .ZN(net_7754), .A(net_7753), .B2(net_1325), .B1(net_1016) );
CLKBUF_X2 inst_21970 ( .A(net_21841), .Z(net_21842) );
NAND2_X2 inst_9155 ( .ZN(net_13388), .A1(net_11907), .A2(net_10607) );
INV_X4 inst_14905 ( .ZN(net_6172), .A(net_3589) );
INV_X4 inst_14570 ( .ZN(net_7511), .A(net_3677) );
NAND2_X4 inst_6834 ( .ZN(net_18787), .A2(net_18744), .A1(net_18719) );
INV_X4 inst_18175 ( .A(net_21062), .ZN(net_541) );
INV_X2 inst_18407 ( .A(net_16602), .ZN(net_16476) );
AOI211_X2 inst_21081 ( .A(net_7097), .ZN(net_5264), .B(net_4805), .C2(net_2532), .C1(net_2485) );
AOI21_X4 inst_20135 ( .ZN(net_19798), .B1(net_15876), .B2(net_15560), .A(net_14948) );
NAND2_X2 inst_10701 ( .A1(net_20553), .ZN(net_8759), .A2(net_6042) );
NOR2_X4 inst_2827 ( .ZN(net_16015), .A1(net_15806), .A2(net_15485) );
NAND2_X2 inst_9062 ( .A1(net_15270), .ZN(net_13991), .A2(net_11989) );
OAI211_X2 inst_2448 ( .ZN(net_14626), .B(net_11985), .C2(net_11530), .C1(net_9638), .A(net_5751) );
CLKBUF_X2 inst_22598 ( .A(net_22469), .Z(net_22470) );
AND2_X4 inst_21253 ( .A1(net_20875), .A2(net_1981), .ZN(net_1833) );
INV_X4 inst_17146 ( .ZN(net_1433), .A(net_774) );
OAI211_X2 inst_2541 ( .ZN(net_10828), .B(net_6563), .C2(net_4625), .C1(net_3331), .A(net_2623) );
AND2_X2 inst_21294 ( .ZN(net_19181), .A1(net_12036), .A2(net_8508) );
INV_X4 inst_17525 ( .ZN(net_4074), .A(net_662) );
OAI21_X2 inst_1693 ( .ZN(net_15358), .B2(net_13723), .B1(net_9800), .A(net_3396) );
INV_X2 inst_19690 ( .A(net_20543), .ZN(net_20542) );
DFF_X1 inst_19799 ( .D(net_18195), .CK(net_22400), .Q(x779) );
AOI21_X4 inst_20162 ( .ZN(net_19999), .B1(net_19775), .B2(net_15026), .A(net_14447) );
NOR2_X4 inst_3306 ( .A2(net_20860), .A1(net_2244), .ZN(net_1157) );
SDFF_X2 inst_1020 ( .QN(net_20992), .D(net_361), .SE(net_263), .CK(net_21833), .SI(x3147) );
CLKBUF_X2 inst_22430 ( .A(net_22301), .Z(net_22302) );
NAND2_X2 inst_11007 ( .ZN(net_4880), .A2(net_4023), .A1(net_107) );
INV_X4 inst_17959 ( .A(net_21071), .ZN(net_489) );
NAND2_X2 inst_7721 ( .ZN(net_18838), .A2(net_18814), .A1(net_18798) );
NAND2_X2 inst_11057 ( .ZN(net_4633), .A2(net_4632), .A1(net_3990) );
INV_X4 inst_13886 ( .ZN(net_12280), .A(net_5769) );
INV_X4 inst_16298 ( .ZN(net_4340), .A(net_1341) );
NOR2_X2 inst_3952 ( .ZN(net_19284), .A2(net_7949), .A1(net_2657) );
NAND2_X2 inst_12084 ( .A1(net_20873), .A2(net_3201), .ZN(net_1266) );
NOR2_X2 inst_3588 ( .ZN(net_12625), .A2(net_12624), .A1(net_11198) );
INV_X2 inst_19566 ( .A(net_14657), .ZN(net_784) );
INV_X4 inst_15120 ( .ZN(net_7106), .A(net_6402) );
NAND3_X4 inst_5559 ( .ZN(net_16131), .A3(net_15746), .A1(net_15613), .A2(net_13106) );
OR2_X4 inst_1096 ( .ZN(net_9100), .A1(net_7892), .A2(net_4677) );
INV_X4 inst_16336 ( .A(net_2855), .ZN(net_1826) );
NOR2_X2 inst_4552 ( .ZN(net_4983), .A2(net_3823), .A1(net_3385) );
NAND2_X2 inst_9260 ( .ZN(net_12639), .A1(net_12638), .A2(net_10833) );
CLKBUF_X2 inst_22498 ( .A(net_22369), .Z(net_22370) );
DFF_X1 inst_19843 ( .D(net_17403), .CK(net_21350), .Q(x296) );
NAND3_X2 inst_5637 ( .ZN(net_20504), .A3(net_18069), .A1(net_16226), .A2(net_10817) );
OAI21_X2 inst_1839 ( .ZN(net_14028), .A(net_14027), .B2(net_10258), .B1(net_5284) );
INV_X4 inst_14708 ( .ZN(net_15869), .A(net_14837) );
AOI22_X2 inst_19958 ( .A1(net_21236), .B1(net_16644), .ZN(net_16283), .B2(net_16010), .A2(net_15893) );
INV_X4 inst_18332 ( .A(net_20565), .ZN(net_20564) );
NAND2_X2 inst_8041 ( .ZN(net_18285), .A1(net_18167), .A2(net_18139) );
INV_X4 inst_13095 ( .ZN(net_18947), .A(net_15739) );
SDFF_X2 inst_725 ( .Q(net_20901), .SE(net_18864), .SI(net_18571), .D(net_854), .CK(net_21498) );
INV_X4 inst_12840 ( .ZN(net_17350), .A(net_17227) );
NAND3_X2 inst_6326 ( .ZN(net_12510), .A2(net_7579), .A3(net_4697), .A1(net_2591) );
OAI221_X2 inst_1337 ( .ZN(net_15173), .A(net_14616), .C1(net_14315), .C2(net_12564), .B2(net_8992), .B1(net_2368) );
INV_X4 inst_18181 ( .A(net_20965), .ZN(net_834) );
NAND4_X2 inst_5375 ( .ZN(net_19541), .A4(net_14053), .A1(net_13351), .A3(net_12677), .A2(net_9648) );
NOR2_X4 inst_3096 ( .ZN(net_4218), .A2(net_2648), .A1(net_154) );
AOI22_X2 inst_20001 ( .B1(net_15360), .A1(net_14078), .ZN(net_13866), .A2(net_11591), .B2(net_9845) );
INV_X4 inst_15532 ( .ZN(net_15119), .A(net_14009) );
NOR2_X4 inst_3015 ( .A2(net_20548), .A1(net_7099), .ZN(net_6845) );
INV_X2 inst_19520 ( .ZN(net_1805), .A(net_848) );
CLKBUF_X2 inst_22342 ( .A(net_22213), .Z(net_22214) );
NAND2_X2 inst_11618 ( .A2(net_2891), .ZN(net_2578), .A1(net_1768) );
OAI211_X2 inst_2441 ( .ZN(net_14824), .C1(net_14551), .B(net_13389), .A(net_10540), .C2(net_2936) );
INV_X4 inst_17288 ( .A(net_1922), .ZN(net_629) );
INV_X4 inst_16264 ( .ZN(net_15248), .A(net_14678) );
NAND2_X2 inst_11945 ( .ZN(net_1439), .A1(net_1438), .A2(net_757) );
AOI21_X4 inst_20128 ( .ZN(net_16156), .B1(net_16127), .B2(net_15777), .A(net_15461) );
NAND2_X2 inst_9714 ( .ZN(net_20831), .A1(net_10174), .A2(net_9593) );
NAND2_X4 inst_7427 ( .ZN(net_5329), .A2(net_3493), .A1(net_2139) );
AOI21_X2 inst_20708 ( .ZN(net_12106), .B2(net_12105), .B1(net_8497), .A(net_253) );
SDFF_X2 inst_878 ( .Q(net_21210), .D(net_16933), .SE(net_253), .CK(net_22435), .SI(x5825) );
INV_X4 inst_17099 ( .ZN(net_9339), .A(net_8041) );
NOR2_X2 inst_4959 ( .ZN(net_1629), .A1(net_243), .A2(net_61) );
INV_X2 inst_18707 ( .ZN(net_8243), .A(net_8242) );
INV_X4 inst_13442 ( .ZN(net_11644), .A(net_9794) );
NAND3_X2 inst_6782 ( .A3(net_4820), .A2(net_4704), .ZN(net_4260), .A1(net_4259) );
INV_X2 inst_19669 ( .A(net_20484), .ZN(net_20483) );
OAI21_X2 inst_1926 ( .A(net_13371), .ZN(net_12980), .B2(net_9293), .B1(net_8107) );
NOR2_X2 inst_4351 ( .ZN(net_5619), .A1(net_5618), .A2(net_2613) );
INV_X4 inst_17683 ( .ZN(net_573), .A(net_508) );
INV_X4 inst_16908 ( .ZN(net_14171), .A(net_7173) );
NAND3_X2 inst_6211 ( .ZN(net_13271), .A1(net_9592), .A3(net_8858), .A2(net_8079) );
INV_X4 inst_12761 ( .ZN(net_17389), .A(net_17388) );
NAND3_X2 inst_6383 ( .A2(net_13486), .ZN(net_12023), .A3(net_10475), .A1(net_8228) );
XNOR2_X2 inst_564 ( .ZN(net_672), .A(net_671), .B(net_670) );
AND3_X4 inst_21115 ( .ZN(net_13963), .A3(net_13962), .A1(net_13460), .A2(net_12056) );
INV_X4 inst_12795 ( .ZN(net_17271), .A(net_17270) );
NAND2_X2 inst_10262 ( .ZN(net_12910), .A1(net_7988), .A2(net_5048) );
INV_X4 inst_16913 ( .ZN(net_1828), .A(net_939) );
NAND2_X2 inst_11210 ( .A1(net_20546), .ZN(net_6902), .A2(net_2806) );
NAND3_X2 inst_6500 ( .ZN(net_10835), .A2(net_10834), .A1(net_8409), .A3(net_7069) );
SDFF_X2 inst_934 ( .QN(net_21062), .D(net_541), .SE(net_263), .CK(net_21744), .SI(x2027) );
SDFF_X2 inst_1000 ( .QN(net_21041), .SE(net_2426), .D(net_496), .CK(net_22002), .SI(x2298) );
INV_X4 inst_17398 ( .ZN(net_1881), .A(net_938) );
INV_X2 inst_18606 ( .A(net_9782), .ZN(net_9781) );
INV_X4 inst_18188 ( .A(net_21119), .ZN(net_17494) );
OAI211_X2 inst_2585 ( .C1(net_9131), .A(net_8963), .ZN(net_7083), .B(net_7082), .C2(net_2645) );
NAND2_X2 inst_12044 ( .ZN(net_1181), .A1(net_824), .A2(net_809) );
OAI21_X1 inst_2364 ( .A(net_12004), .ZN(net_7150), .B2(net_7149), .B1(net_2737) );
NOR2_X2 inst_4299 ( .ZN(net_7446), .A1(net_5951), .A2(net_5889) );
INV_X2 inst_18502 ( .ZN(net_12104), .A(net_10668) );
CLKBUF_X2 inst_21465 ( .A(net_21336), .Z(net_21337) );
NAND2_X2 inst_11281 ( .A2(net_3945), .ZN(net_3857), .A1(net_165) );
OAI21_X2 inst_1882 ( .ZN(net_13545), .A(net_13544), .B2(net_9812), .B1(net_9154) );
AOI21_X2 inst_20869 ( .A(net_10917), .B2(net_9956), .ZN(net_8570), .B1(net_8469) );
INV_X4 inst_14510 ( .A(net_11264), .ZN(net_8025) );
INV_X4 inst_13787 ( .A(net_9437), .ZN(net_9204) );
INV_X4 inst_14482 ( .ZN(net_7248), .A(net_4869) );
NAND2_X2 inst_7812 ( .ZN(net_18674), .A2(net_18655), .A1(net_17395) );
INV_X4 inst_17273 ( .ZN(net_1329), .A(net_647) );
NAND2_X2 inst_8441 ( .ZN(net_19154), .A2(net_17007), .A1(net_634) );
NAND2_X2 inst_8218 ( .ZN(net_17838), .A2(net_17706), .A1(net_17640) );
NAND3_X2 inst_6578 ( .ZN(net_10450), .A2(net_10449), .A3(net_8696), .A1(net_4695) );
INV_X2 inst_19174 ( .ZN(net_3810), .A(net_3809) );
INV_X4 inst_16149 ( .ZN(net_9438), .A(net_4156) );
INV_X4 inst_12849 ( .ZN(net_17069), .A(net_17068) );
INV_X4 inst_17686 ( .ZN(net_4288), .A(net_304) );
NAND3_X4 inst_5531 ( .ZN(net_17662), .A3(net_16896), .A2(net_16128), .A1(net_13141) );
NAND4_X2 inst_5397 ( .ZN(net_19512), .A2(net_12769), .A3(net_10777), .A4(net_10572), .A1(net_8585) );
SDFF_X2 inst_727 ( .Q(net_20865), .SE(net_18577), .SI(net_18568), .D(net_464), .CK(net_22457) );
AOI21_X2 inst_20368 ( .B1(net_20396), .B2(net_15831), .ZN(net_15630), .A(net_13652) );
NAND2_X2 inst_11795 ( .ZN(net_3823), .A2(net_2093), .A1(net_1220) );
NOR2_X2 inst_4804 ( .ZN(net_12939), .A2(net_3013), .A1(net_2709) );
CLKBUF_X2 inst_21730 ( .A(net_21491), .Z(net_21602) );
NAND2_X2 inst_11686 ( .ZN(net_11861), .A1(net_6207), .A2(net_2343) );
NOR2_X4 inst_2874 ( .ZN(net_12303), .A1(net_10015), .A2(net_9164) );
INV_X2 inst_19471 ( .A(net_9109), .ZN(net_1441) );
NAND3_X2 inst_6485 ( .ZN(net_11197), .A2(net_11041), .A1(net_6120), .A3(net_5846) );
NOR2_X2 inst_4607 ( .A2(net_3815), .ZN(net_3744), .A1(net_1452) );
OAI211_X2 inst_2431 ( .ZN(net_15030), .B(net_15029), .A(net_13029), .C2(net_12570), .C1(net_1181) );
NAND2_X2 inst_8861 ( .ZN(net_15344), .A1(net_15343), .A2(net_14428) );
NAND2_X2 inst_12052 ( .ZN(net_906), .A1(net_300), .A2(net_117) );
AND2_X4 inst_21189 ( .A1(net_14538), .ZN(net_10750), .A2(net_10749) );
INV_X2 inst_18713 ( .ZN(net_8216), .A(net_8215) );
NAND2_X2 inst_8274 ( .ZN(net_17646), .A2(net_17473), .A1(net_17349) );
DFF_X1 inst_19790 ( .D(net_18651), .CK(net_22123), .Q(x532) );
INV_X4 inst_16085 ( .ZN(net_14430), .A(net_6886) );
NAND2_X4 inst_7607 ( .A1(net_19287), .ZN(net_3102), .A2(net_1735) );
SDFF_X2 inst_953 ( .QN(net_21064), .D(net_530), .SE(net_263), .CK(net_21739), .SI(x2011) );
INV_X4 inst_16605 ( .ZN(net_14865), .A(net_12609) );
INV_X4 inst_13674 ( .A(net_12109), .ZN(net_8005) );
NAND2_X2 inst_11524 ( .A2(net_3757), .ZN(net_3740), .A1(net_182) );
INV_X2 inst_18989 ( .ZN(net_5102), .A(net_5101) );
INV_X2 inst_18811 ( .ZN(net_7335), .A(net_5772) );
NAND4_X2 inst_5483 ( .ZN(net_12484), .A3(net_12483), .A2(net_8833), .A4(net_7691), .A1(net_5937) );
CLKBUF_X2 inst_21613 ( .A(net_21286), .Z(net_21485) );
NAND3_X2 inst_6694 ( .ZN(net_7686), .A1(net_4774), .A2(net_3290), .A3(net_2901) );
NOR2_X2 inst_3373 ( .A2(net_17517), .ZN(net_16672), .A1(net_11872) );
NAND2_X2 inst_8919 ( .ZN(net_14958), .A2(net_13714), .A1(net_13353) );
NOR2_X2 inst_4902 ( .ZN(net_4402), .A1(net_1980), .A2(net_1799) );
AOI22_X2 inst_20050 ( .A1(net_11270), .ZN(net_3706), .A2(net_2584), .B1(net_2388), .B2(net_1283) );
INV_X1 inst_19755 ( .A(net_8245), .ZN(net_6179) );
NAND2_X4 inst_7613 ( .ZN(net_1905), .A2(net_1347), .A1(net_1216) );
INV_X2 inst_19329 ( .ZN(net_2548), .A(net_2547) );
NAND2_X2 inst_11464 ( .ZN(net_4645), .A2(net_1828), .A1(net_1720) );
INV_X4 inst_18072 ( .A(net_21035), .ZN(net_469) );
NAND2_X4 inst_6956 ( .A2(net_19436), .ZN(net_17478), .A1(net_17362) );
NOR2_X2 inst_4720 ( .A1(net_6692), .ZN(net_3125), .A2(net_2396) );
INV_X4 inst_16750 ( .ZN(net_8246), .A(net_6274) );
NAND2_X2 inst_11488 ( .A1(net_4340), .ZN(net_4004), .A2(net_3093) );
INV_X4 inst_17699 ( .ZN(net_1959), .A(net_270) );
NOR2_X2 inst_4986 ( .ZN(net_12712), .A2(net_1470), .A1(net_112) );
INV_X2 inst_18980 ( .A(net_8039), .ZN(net_5148) );
INV_X2 inst_18695 ( .A(net_8879), .ZN(net_8357) );
NAND3_X2 inst_6378 ( .ZN(net_12037), .A2(net_12036), .A3(net_12035), .A1(net_8088) );
XNOR2_X2 inst_294 ( .B(net_21168), .ZN(net_17130), .A(net_17129) );
CLKBUF_X2 inst_21759 ( .A(net_21421), .Z(net_21631) );
INV_X4 inst_13510 ( .A(net_9407), .ZN(net_9406) );
NAND2_X2 inst_8275 ( .ZN(net_17728), .A2(net_17464), .A1(net_17345) );
NAND2_X2 inst_7842 ( .A2(net_20523), .ZN(net_18619), .A1(net_18618) );
INV_X4 inst_15428 ( .A(net_7988), .ZN(net_7867) );
NOR2_X2 inst_3384 ( .ZN(net_16365), .A2(net_16213), .A1(net_16077) );
AOI21_X2 inst_20320 ( .A(net_20889), .B2(net_19015), .B1(net_19014), .ZN(net_15905) );
NAND2_X2 inst_11202 ( .ZN(net_5116), .A2(net_4272), .A1(net_4052) );
SDFF_X2 inst_810 ( .Q(net_21194), .SI(net_17871), .SE(net_125), .CK(net_21419), .D(x6246) );
INV_X4 inst_16540 ( .A(net_10105), .ZN(net_9313) );
NAND2_X2 inst_8982 ( .ZN(net_14498), .A2(net_12739), .A1(net_7394) );
INV_X4 inst_16043 ( .ZN(net_2672), .A(net_1609) );
NAND2_X2 inst_9511 ( .ZN(net_11238), .A2(net_8350), .A1(net_6873) );
INV_X2 inst_18895 ( .ZN(net_9675), .A(net_6101) );
NAND2_X2 inst_9767 ( .ZN(net_11132), .A2(net_9813), .A1(net_8961) );
NOR2_X4 inst_3035 ( .ZN(net_20773), .A2(net_5162), .A1(net_3634) );
INV_X2 inst_18900 ( .ZN(net_11553), .A(net_8221) );
INV_X4 inst_17694 ( .A(net_20889), .ZN(net_588) );
INV_X4 inst_14855 ( .ZN(net_14545), .A(net_3813) );
NAND2_X2 inst_12063 ( .A2(net_9131), .ZN(net_1066), .A1(net_861) );
INV_X4 inst_18015 ( .A(net_20874), .ZN(net_493) );
NAND2_X2 inst_7836 ( .A1(net_18640), .ZN(net_18631), .A2(net_18620) );
INV_X2 inst_19386 ( .ZN(net_2126), .A(net_2125) );
NAND2_X2 inst_10010 ( .ZN(net_8799), .A1(net_8798), .A2(net_8180) );
INV_X4 inst_14573 ( .ZN(net_5917), .A(net_3772) );
NAND2_X2 inst_11984 ( .ZN(net_1281), .A2(net_253), .A1(x4642) );
XNOR2_X2 inst_481 ( .ZN(net_11047), .B(net_7277), .A(net_1855) );
INV_X4 inst_16076 ( .ZN(net_15969), .A(net_15744) );
NAND3_X2 inst_5992 ( .ZN(net_19802), .A1(net_13395), .A3(net_7335), .A2(net_4683) );
INV_X4 inst_16295 ( .ZN(net_1816), .A(net_954) );
NAND2_X2 inst_8633 ( .A1(net_20790), .ZN(net_16589), .A2(net_16588) );
INV_X4 inst_13699 ( .ZN(net_11869), .A(net_7891) );
NAND3_X2 inst_6208 ( .ZN(net_13280), .A2(net_13279), .A3(net_13278), .A1(net_11351) );
INV_X4 inst_16899 ( .ZN(net_1037), .A(net_117) );
INV_X4 inst_13056 ( .ZN(net_16372), .A(net_16331) );
OAI211_X2 inst_2485 ( .B(net_14545), .ZN(net_13478), .A(net_13201), .C2(net_12561), .C1(net_3397) );
INV_X4 inst_16773 ( .ZN(net_1026), .A(net_752) );
NAND2_X2 inst_9087 ( .ZN(net_13798), .A2(net_12458), .A1(net_10052) );
NAND2_X2 inst_10584 ( .ZN(net_7944), .A1(net_6668), .A2(net_6410) );
INV_X4 inst_13353 ( .ZN(net_12666), .A(net_10986) );
OAI21_X2 inst_2217 ( .B1(net_20487), .B2(net_9041), .ZN(net_8517), .A(net_3825) );
INV_X4 inst_16332 ( .ZN(net_19882), .A(net_2855) );
INV_X4 inst_13707 ( .ZN(net_11894), .A(net_7864) );
INV_X2 inst_19482 ( .ZN(net_2798), .A(net_1949) );
SDFF_X2 inst_850 ( .Q(net_21140), .SI(net_17289), .SE(net_945), .CK(net_22156), .D(x3635) );
INV_X4 inst_17719 ( .ZN(net_5239), .A(net_196) );
NAND2_X4 inst_7612 ( .A1(net_20065), .ZN(net_3095), .A2(net_256) );
NAND2_X2 inst_11175 ( .ZN(net_10502), .A1(net_4156), .A2(net_2251) );
AOI22_X2 inst_20039 ( .A1(net_9083), .ZN(net_7349), .B2(net_7348), .A2(net_5381), .B1(net_573) );
CLKBUF_X2 inst_22295 ( .A(net_22166), .Z(net_22167) );
INV_X4 inst_12642 ( .ZN(net_17903), .A(net_17902) );
INV_X4 inst_16912 ( .ZN(net_1033), .A(net_955) );
AOI21_X2 inst_20672 ( .B1(net_19492), .ZN(net_12589), .B2(net_6478), .A(net_69) );
AOI21_X2 inst_20482 ( .ZN(net_14895), .A(net_13653), .B1(net_13544), .B2(net_9114) );
INV_X4 inst_17444 ( .ZN(net_3148), .A(net_2557) );
INV_X4 inst_14485 ( .ZN(net_8083), .A(net_4853) );
OAI211_X2 inst_2438 ( .ZN(net_14978), .B(net_14384), .C1(net_14227), .C2(net_12466), .A(net_6609) );
AND2_X2 inst_21336 ( .A1(net_4361), .ZN(net_3483), .A2(net_3482) );
INV_X4 inst_15577 ( .ZN(net_4087), .A(net_2272) );
NAND2_X2 inst_10391 ( .A2(net_12011), .ZN(net_7310), .A1(net_7309) );
NAND4_X2 inst_5479 ( .A4(net_13697), .ZN(net_12826), .A2(net_12825), .A3(net_10909), .A1(net_5642) );
XNOR2_X2 inst_237 ( .B(net_21124), .ZN(net_17396), .A(net_16947) );
OAI211_X2 inst_2543 ( .ZN(net_10826), .B(net_7397), .C2(net_4629), .A(net_3373), .C1(net_1989) );
NOR3_X2 inst_2772 ( .A2(net_20023), .ZN(net_19731), .A1(net_6842), .A3(net_5015) );
NAND2_X2 inst_11449 ( .A1(net_3804), .ZN(net_3252), .A2(net_2686) );
NAND2_X2 inst_8836 ( .ZN(net_19478), .A2(net_14796), .A1(net_14280) );
INV_X4 inst_17234 ( .A(net_10319), .ZN(net_6879) );
INV_X4 inst_13178 ( .ZN(net_19225), .A(net_13865) );
NAND2_X2 inst_8056 ( .ZN(net_18207), .A2(net_18174), .A1(net_17852) );
INV_X4 inst_17667 ( .ZN(net_249), .A(net_248) );
XOR2_X2 inst_51 ( .A(net_21164), .Z(net_395), .B(net_394) );
SDFF_X2 inst_813 ( .Q(net_21217), .SI(net_17825), .SE(net_125), .CK(net_22246), .D(x7467) );
CLKBUF_X2 inst_21828 ( .A(net_21511), .Z(net_21700) );
INV_X4 inst_17081 ( .ZN(net_15697), .A(net_12398) );
NAND2_X2 inst_10379 ( .A1(net_18025), .ZN(net_7387), .A2(net_432) );
NAND3_X2 inst_6691 ( .ZN(net_7704), .A2(net_7703), .A3(net_5336), .A1(net_3702) );
INV_X4 inst_14874 ( .ZN(net_19374), .A(net_3690) );
INV_X4 inst_13373 ( .ZN(net_12313), .A(net_10893) );
NAND2_X2 inst_11195 ( .ZN(net_10644), .A1(net_5387), .A2(net_3719) );
OAI21_X2 inst_1837 ( .ZN(net_14035), .B2(net_10103), .B1(net_4720), .A(net_855) );
AOI21_X2 inst_20728 ( .ZN(net_11920), .B1(net_11472), .A(net_9938), .B2(net_8690) );
INV_X2 inst_18527 ( .ZN(net_11107), .A(net_11106) );
INV_X4 inst_13198 ( .ZN(net_13933), .A(net_13272) );
NAND2_X2 inst_9100 ( .ZN(net_13767), .A2(net_13766), .A1(net_10634) );
NAND3_X2 inst_5686 ( .A1(net_20650), .ZN(net_16300), .A3(net_15800), .A2(net_15758) );
NAND2_X2 inst_10944 ( .ZN(net_5146), .A1(net_4794), .A2(net_3686) );
DFF_X1 inst_19905 ( .D(net_16702), .CK(net_22789), .Q(x1176) );
NOR2_X4 inst_3291 ( .A2(net_20495), .ZN(net_1338), .A1(net_995) );
XNOR2_X2 inst_64 ( .ZN(net_18809), .A(net_18762), .B(net_17322) );
INV_X4 inst_15904 ( .A(net_4259), .ZN(net_1766) );
INV_X4 inst_13964 ( .ZN(net_7993), .A(net_6714) );
SDFF_X2 inst_743 ( .Q(net_20974), .SE(net_18576), .SI(net_18550), .D(net_5787), .CK(net_22751) );
OAI21_X2 inst_2106 ( .ZN(net_10053), .A(net_10052), .B1(net_4979), .B2(net_3360) );
NOR2_X2 inst_4051 ( .ZN(net_7855), .A1(net_7854), .A2(net_4933) );
NOR3_X2 inst_2723 ( .ZN(net_13252), .A2(net_11781), .A1(net_10599), .A3(net_6285) );
INV_X2 inst_18825 ( .ZN(net_6859), .A(net_6858) );
NAND2_X2 inst_9141 ( .A1(net_14966), .ZN(net_13421), .A2(net_10784) );
NOR2_X2 inst_4265 ( .ZN(net_7562), .A1(net_6207), .A2(net_4553) );
NAND2_X2 inst_8628 ( .ZN(net_16597), .A2(net_16596), .A1(net_5670) );
AOI211_X2 inst_21053 ( .ZN(net_11789), .B(net_11627), .C1(net_10151), .A(net_7437), .C2(net_4717) );
OAI21_X2 inst_1809 ( .ZN(net_14265), .A(net_14264), .B2(net_13566), .B1(net_9231) );
CLKBUF_X2 inst_21974 ( .A(net_21845), .Z(net_21846) );
NAND3_X2 inst_6664 ( .ZN(net_8445), .A3(net_8444), .A1(net_3857), .A2(net_2693) );
CLKBUF_X2 inst_22790 ( .A(net_22661), .Z(net_22662) );
NAND2_X2 inst_8272 ( .ZN(net_17740), .A1(net_17477), .A2(net_17356) );
INV_X4 inst_14602 ( .ZN(net_9194), .A(net_4444) );
INV_X8 inst_12172 ( .ZN(net_18077), .A(net_18073) );
NAND2_X2 inst_11866 ( .A2(net_2384), .ZN(net_1649), .A1(net_225) );
NOR2_X2 inst_4344 ( .ZN(net_6064), .A2(net_2802), .A1(net_348) );
NAND2_X2 inst_8111 ( .A2(net_20219), .ZN(net_18108), .A1(net_16666) );
NAND2_X2 inst_8541 ( .A2(net_19451), .ZN(net_16825), .A1(net_678) );
INV_X4 inst_15404 ( .A(net_5714), .ZN(net_2533) );
INV_X4 inst_14717 ( .ZN(net_15340), .A(net_2368) );
AOI21_X2 inst_20750 ( .ZN(net_11354), .B1(net_11353), .B2(net_11352), .A(net_10389) );
INV_X4 inst_16794 ( .ZN(net_5595), .A(net_1011) );
NOR2_X2 inst_4011 ( .ZN(net_8074), .A1(net_6059), .A2(net_3801) );
INV_X4 inst_17992 ( .A(net_20895), .ZN(net_137) );
NAND2_X2 inst_11478 ( .ZN(net_4068), .A1(net_2673), .A2(net_2200) );
NAND2_X2 inst_10432 ( .A2(net_7235), .ZN(net_7209), .A1(net_6733) );
INV_X4 inst_15556 ( .ZN(net_7892), .A(net_6135) );
INV_X4 inst_17763 ( .ZN(net_3890), .A(net_284) );
INV_X4 inst_14609 ( .ZN(net_12215), .A(net_6579) );
NAND3_X2 inst_6445 ( .ZN(net_11797), .A2(net_9327), .A1(net_8140), .A3(net_6651) );
INV_X4 inst_17322 ( .ZN(net_4900), .A(net_761) );
AND2_X2 inst_21366 ( .A2(net_20860), .A1(net_1662), .ZN(net_1034) );
NAND2_X2 inst_8045 ( .ZN(net_18233), .A2(net_18232), .A1(net_16697) );
NAND2_X4 inst_7436 ( .ZN(net_10435), .A2(net_3915), .A1(net_3374) );
NAND2_X2 inst_11689 ( .A1(net_4042), .ZN(net_2333), .A2(net_2332) );
NOR2_X4 inst_2980 ( .ZN(net_9779), .A1(net_3308), .A2(net_703) );
NAND4_X4 inst_5197 ( .A2(net_19614), .A1(net_19613), .ZN(net_16428), .A4(net_16075), .A3(net_15949) );
DFF_X1 inst_19785 ( .D(net_18676), .CK(net_22133), .Q(x570) );
INV_X2 inst_18861 ( .ZN(net_6320), .A(net_6319) );
AOI21_X2 inst_20643 ( .ZN(net_13190), .B1(net_11678), .B2(net_8763), .A(net_6567) );
NAND2_X2 inst_10184 ( .ZN(net_11900), .A1(net_7903), .A2(net_6241) );
SDFF_X2 inst_915 ( .Q(net_21148), .D(net_16652), .SE(net_263), .CK(net_22207), .SI(x5754) );
NAND2_X2 inst_9869 ( .A1(net_10592), .ZN(net_9479), .A2(net_7544) );
INV_X2 inst_19396 ( .ZN(net_3497), .A(net_2559) );
NOR2_X2 inst_4416 ( .A1(net_6625), .ZN(net_5014), .A2(net_5013) );
NAND2_X2 inst_10008 ( .ZN(net_8801), .A2(net_6463), .A1(net_6112) );
NAND3_X2 inst_5660 ( .ZN(net_16427), .A2(net_16275), .A3(net_16216), .A1(net_11463) );
INV_X4 inst_16343 ( .ZN(net_15692), .A(net_15104) );
INV_X4 inst_14017 ( .ZN(net_11929), .A(net_8254) );
INV_X4 inst_16096 ( .A(net_1999), .ZN(net_1521) );
NAND2_X2 inst_9552 ( .ZN(net_11022), .A2(net_11021), .A1(net_6049) );
INV_X4 inst_14703 ( .ZN(net_14706), .A(net_9263) );
INV_X4 inst_12591 ( .A(net_18153), .ZN(net_18135) );
NOR2_X2 inst_4807 ( .ZN(net_7138), .A1(net_2750), .A2(net_2681) );
AND3_X2 inst_21132 ( .ZN(net_14403), .A2(net_14402), .A3(net_13846), .A1(net_13537) );
OAI21_X2 inst_1668 ( .ZN(net_15663), .A(net_15616), .B2(net_14892), .B1(net_13443) );
AOI21_X2 inst_20595 ( .B1(net_19653), .ZN(net_13901), .B2(net_11062), .A(net_6244) );
INV_X4 inst_16432 ( .A(net_5959), .ZN(net_1245) );
NAND2_X2 inst_11169 ( .ZN(net_5223), .A1(net_4163), .A2(net_4125) );
NAND2_X2 inst_9987 ( .ZN(net_12172), .A1(net_8870), .A2(net_8847) );
INV_X4 inst_15425 ( .A(net_14038), .ZN(net_8870) );
NOR2_X2 inst_4811 ( .A1(net_5220), .ZN(net_3782), .A2(net_2444) );
INV_X4 inst_15935 ( .ZN(net_9903), .A(net_1725) );
NAND2_X2 inst_11942 ( .ZN(net_2787), .A1(net_1445), .A2(net_1395) );
AND2_X2 inst_21345 ( .ZN(net_7136), .A1(net_2686), .A2(net_2685) );
NAND2_X4 inst_7068 ( .A2(net_20872), .A1(net_20262), .ZN(net_16238) );
INV_X2 inst_19350 ( .ZN(net_2397), .A(net_2396) );
INV_X2 inst_18726 ( .ZN(net_20357), .A(net_8102) );
XNOR2_X2 inst_293 ( .A(net_17820), .ZN(net_17132), .B(net_9258) );
NOR2_X2 inst_4741 ( .A2(net_6426), .ZN(net_3044), .A1(net_242) );
NAND2_X2 inst_11078 ( .A2(net_11382), .ZN(net_4463), .A1(net_1627) );
NOR2_X2 inst_3744 ( .ZN(net_10602), .A2(net_7291), .A1(net_5487) );
INV_X4 inst_15346 ( .A(net_5149), .ZN(net_3364) );
INV_X4 inst_17154 ( .ZN(net_9378), .A(net_5450) );
NAND4_X2 inst_5402 ( .ZN(net_14742), .A1(net_11433), .A4(net_10558), .A3(net_10102), .A2(net_8871) );
INV_X2 inst_18976 ( .ZN(net_5188), .A(net_5187) );
NOR2_X4 inst_2953 ( .ZN(net_8134), .A1(net_5311), .A2(net_3069) );
INV_X4 inst_13000 ( .ZN(net_19803), .A(net_16418) );
INV_X4 inst_17614 ( .ZN(net_1922), .A(net_309) );
NAND2_X2 inst_8219 ( .ZN(net_17837), .A2(net_17799), .A1(net_17438) );
XNOR2_X2 inst_98 ( .ZN(net_18542), .A(net_18433), .B(net_17393) );
INV_X2 inst_19392 ( .ZN(net_2067), .A(net_1541) );
NOR2_X4 inst_3087 ( .A2(net_20536), .ZN(net_6267), .A1(net_2813) );
SDFF_X2 inst_959 ( .QN(net_21089), .D(net_707), .SE(net_253), .CK(net_21785), .SI(x1580) );
NAND2_X2 inst_10102 ( .A1(net_8949), .ZN(net_8579), .A2(net_5214) );
INV_X4 inst_14611 ( .ZN(net_7677), .A(net_4428) );
INV_X2 inst_19478 ( .ZN(net_1401), .A(net_1400) );
INV_X2 inst_18397 ( .A(net_16801), .ZN(net_16486) );
INV_X4 inst_13343 ( .A(net_11499), .ZN(net_11082) );
NAND2_X4 inst_7626 ( .ZN(net_1238), .A1(net_1237), .A2(net_106) );
XNOR2_X2 inst_605 ( .B(net_595), .ZN(net_521), .A(net_520) );
NAND2_X2 inst_9998 ( .ZN(net_8828), .A2(net_8112), .A1(net_6061) );
NAND2_X4 inst_7481 ( .ZN(net_20578), .A2(net_19418), .A1(net_1783) );
NOR3_X1 inst_2799 ( .A2(net_11365), .ZN(net_11256), .A3(net_11255), .A1(net_5356) );
NAND2_X2 inst_10988 ( .A2(net_20577), .A1(net_6177), .ZN(net_4936) );
CLKBUF_X2 inst_22489 ( .A(net_22360), .Z(net_22361) );
OAI21_X2 inst_2048 ( .A(net_13494), .ZN(net_10854), .B1(net_6525), .B2(net_5673) );
NOR2_X4 inst_2948 ( .ZN(net_8180), .A1(net_7872), .A2(net_6862) );
NAND2_X2 inst_7900 ( .ZN(net_18483), .A2(net_18429), .A1(net_18379) );
INV_X2 inst_19310 ( .ZN(net_2714), .A(net_2713) );
INV_X2 inst_19364 ( .A(net_2829), .ZN(net_2245) );
NAND2_X2 inst_10396 ( .A1(net_10567), .ZN(net_7290), .A2(net_7289) );
NAND2_X2 inst_11643 ( .ZN(net_5671), .A1(net_2493), .A2(net_1128) );
INV_X4 inst_13850 ( .A(net_7469), .ZN(net_7468) );
CLKBUF_X2 inst_21597 ( .A(net_21468), .Z(net_21469) );
OAI21_X2 inst_1931 ( .A(net_15372), .ZN(net_12940), .B1(net_12939), .B2(net_9664) );
INV_X2 inst_19684 ( .A(net_20526), .ZN(net_20525) );
NOR2_X2 inst_4735 ( .A1(net_20557), .ZN(net_4265), .A2(net_3065) );
NAND3_X2 inst_6631 ( .A3(net_11830), .ZN(net_9017), .A2(net_8442), .A1(net_2351) );
NAND2_X2 inst_11926 ( .A1(net_3226), .A2(net_1593), .ZN(net_1498) );
NAND2_X2 inst_8402 ( .ZN(net_17384), .A2(net_16957), .A1(net_16791) );
NOR2_X4 inst_3002 ( .A1(net_20446), .ZN(net_7564), .A2(net_90) );
INV_X4 inst_13007 ( .ZN(net_16750), .A(net_16615) );
NOR2_X2 inst_4389 ( .ZN(net_6326), .A2(net_5200), .A1(net_154) );
NAND2_X4 inst_6828 ( .ZN(net_18851), .A2(net_18820), .A1(net_18800) );
INV_X4 inst_15153 ( .A(net_15810), .ZN(net_3552) );
NOR2_X4 inst_2940 ( .A1(net_20024), .ZN(net_9793), .A2(net_1376) );
INV_X4 inst_16391 ( .ZN(net_8205), .A(net_5701) );
NAND2_X2 inst_11855 ( .ZN(net_1678), .A1(net_307), .A2(net_222) );
NAND2_X4 inst_7533 ( .A1(net_19516), .ZN(net_2808), .A2(net_879) );
NAND2_X2 inst_9383 ( .ZN(net_19980), .A1(net_9451), .A2(net_8928) );
NAND3_X2 inst_6606 ( .ZN(net_9297), .A1(net_9295), .A2(net_7695), .A3(net_3536) );
AND4_X4 inst_21088 ( .ZN(net_19064), .A1(net_15081), .A4(net_14139), .A3(net_13689), .A2(net_12253) );
NAND2_X2 inst_11267 ( .A1(net_10667), .ZN(net_3894), .A2(net_2438) );
CLKBUF_X2 inst_22434 ( .A(net_22305), .Z(net_22306) );
AOI21_X2 inst_20662 ( .ZN(net_12964), .A(net_10995), .B1(net_10031), .B2(net_9271) );
INV_X4 inst_15048 ( .ZN(net_5060), .A(net_3371) );
NAND2_X4 inst_7022 ( .ZN(net_17378), .A1(net_16561), .A2(net_16450) );
NOR2_X2 inst_3474 ( .ZN(net_14452), .A2(net_12781), .A1(net_10695) );
INV_X4 inst_16136 ( .ZN(net_2289), .A(net_2275) );
INV_X8 inst_12328 ( .A(net_3919), .ZN(net_2327) );
AOI21_X2 inst_20555 ( .ZN(net_14284), .B1(net_12359), .B2(net_9802), .A(net_8959) );
XNOR2_X2 inst_578 ( .A(net_16921), .B(net_16464), .ZN(net_13286) );
INV_X4 inst_17251 ( .ZN(net_656), .A(net_655) );
INV_X4 inst_17913 ( .ZN(net_1581), .A(net_1271) );
INV_X4 inst_16129 ( .ZN(net_13091), .A(net_6886) );
INV_X4 inst_14197 ( .ZN(net_7452), .A(net_5974) );
INV_X4 inst_13063 ( .ZN(net_19161), .A(net_16294) );
INV_X4 inst_17873 ( .ZN(net_1708), .A(net_834) );
INV_X4 inst_15164 ( .ZN(net_5436), .A(net_4248) );
NAND2_X4 inst_7317 ( .ZN(net_8351), .A1(net_5165), .A2(net_131) );
CLKBUF_X2 inst_22783 ( .A(net_22606), .Z(net_22655) );
INV_X2 inst_18355 ( .ZN(net_18626), .A(net_18604) );
OAI21_X4 inst_1498 ( .ZN(net_20838), .A(net_12004), .B2(net_11735), .B1(net_8231) );
OAI21_X4 inst_1358 ( .ZN(net_18273), .A(net_18152), .B2(net_18086), .B1(net_16539) );
NAND2_X2 inst_8343 ( .ZN(net_19931), .A1(net_17472), .A2(net_17242) );
INV_X4 inst_17853 ( .ZN(net_926), .A(net_766) );
INV_X2 inst_18935 ( .ZN(net_20590), .A(net_5833) );
INV_X8 inst_12456 ( .ZN(net_20775), .A(net_20774) );
NOR2_X2 inst_4775 ( .ZN(net_9931), .A2(net_2732), .A1(net_1175) );
INV_X4 inst_16303 ( .ZN(net_3654), .A(net_1211) );
DFF_X1 inst_19818 ( .D(net_17779), .CK(net_22384), .Q(x848) );
NAND2_X2 inst_10831 ( .A1(net_20573), .ZN(net_6770), .A2(net_4051) );
CLKBUF_X2 inst_21428 ( .A(net_21299), .Z(net_21300) );
NOR2_X2 inst_4450 ( .ZN(net_5746), .A1(net_5217), .A2(net_1877) );
CLKBUF_X2 inst_21843 ( .A(net_21714), .Z(net_21715) );
INV_X4 inst_12817 ( .ZN(net_17512), .A(net_17365) );
INV_X4 inst_17856 ( .A(net_8967), .ZN(net_277) );
INV_X8 inst_12460 ( .ZN(net_20807), .A(net_2637) );
NOR2_X4 inst_3182 ( .ZN(net_4353), .A2(net_3122), .A1(net_193) );
AOI21_X2 inst_20730 ( .ZN(net_11774), .B2(net_9443), .B1(net_7230), .A(net_5045) );
INV_X4 inst_14557 ( .ZN(net_7393), .A(net_5698) );
NOR2_X4 inst_2866 ( .ZN(net_12386), .A1(net_11016), .A2(net_11015) );
NAND3_X2 inst_6805 ( .A3(net_20798), .ZN(net_9799), .A1(net_3185), .A2(net_3184) );
NAND2_X2 inst_11528 ( .ZN(net_2956), .A1(net_2955), .A2(net_2005) );
NAND2_X2 inst_11546 ( .ZN(net_2892), .A1(net_2436), .A2(net_1201) );
NAND4_X2 inst_5379 ( .ZN(net_15160), .A4(net_13784), .A2(net_13412), .A3(net_10248), .A1(net_5876) );
SDFF_X2 inst_838 ( .Q(net_21199), .SI(net_17332), .SE(net_125), .CK(net_22163), .D(x6110) );
CLKBUF_X2 inst_22004 ( .A(net_21875), .Z(net_21876) );
CLKBUF_X2 inst_22901 ( .A(net_22772), .Z(net_22773) );
INV_X4 inst_12905 ( .ZN(net_16705), .A(net_16548) );
OAI21_X4 inst_1405 ( .A(net_20896), .B2(net_18885), .B1(net_18884), .ZN(net_16184) );
NAND3_X2 inst_6811 ( .A3(net_20581), .ZN(net_3004), .A1(net_1682), .A2(net_896) );
NOR2_X2 inst_4058 ( .A1(net_11345), .ZN(net_10181), .A2(net_8187) );
CLKBUF_X2 inst_22037 ( .A(net_21908), .Z(net_21909) );
NAND3_X2 inst_6786 ( .ZN(net_19482), .A1(net_4229), .A3(net_1877), .A2(net_1633) );
NAND2_X2 inst_9172 ( .ZN(net_13349), .A1(net_13348), .A2(net_10568) );
NOR3_X2 inst_2749 ( .A2(net_19627), .ZN(net_12433), .A1(net_9122), .A3(net_3831) );
NAND3_X4 inst_5584 ( .A3(net_20432), .A1(net_20431), .ZN(net_20256), .A2(net_14724) );
NAND2_X4 inst_6963 ( .A2(net_19042), .A1(net_19041), .ZN(net_17428) );
CLKBUF_X2 inst_22622 ( .A(net_22493), .Z(net_22494) );
INV_X2 inst_19065 ( .A(net_6176), .ZN(net_4640) );
NAND2_X2 inst_8823 ( .ZN(net_19552), .A2(net_14830), .A1(net_11856) );
AOI21_X2 inst_20626 ( .ZN(net_13445), .B1(net_13444), .B2(net_8944), .A(net_8210) );
NAND2_X2 inst_11118 ( .A1(net_10119), .ZN(net_4314), .A2(net_4313) );
INV_X4 inst_14647 ( .A(net_5480), .ZN(net_4372) );
NAND3_X4 inst_5567 ( .ZN(net_19690), .A3(net_15216), .A1(net_14340), .A2(net_13817) );
OAI21_X2 inst_2013 ( .ZN(net_11383), .B1(net_11382), .A(net_10335), .B2(net_7690) );
AOI22_X2 inst_20030 ( .B1(net_11858), .ZN(net_9898), .B2(net_9897), .A1(net_8186), .A2(net_4924) );
NOR2_X2 inst_4506 ( .A1(net_6750), .ZN(net_4720), .A2(net_4219) );
NOR3_X2 inst_2756 ( .A2(net_11368), .ZN(net_11254), .A3(net_11253), .A1(net_5365) );
NAND2_X2 inst_10071 ( .A1(net_12339), .ZN(net_8656), .A2(net_8655) );
XNOR2_X2 inst_492 ( .B(net_15294), .ZN(net_9238), .A(net_4449) );
NAND2_X2 inst_8635 ( .A1(net_20769), .ZN(net_16585), .A2(net_16584) );
NAND2_X4 inst_7229 ( .A1(net_20637), .ZN(net_7269), .A2(net_7268) );
NAND4_X2 inst_5414 ( .ZN(net_14583), .A4(net_12155), .A1(net_9964), .A2(net_8480), .A3(net_8437) );
INV_X4 inst_18298 ( .A(net_20473), .ZN(net_20472) );
INV_X4 inst_12589 ( .ZN(net_18187), .A(net_18162) );
INV_X8 inst_12292 ( .ZN(net_1666), .A(net_1071) );
XNOR2_X2 inst_82 ( .ZN(net_18655), .A(net_18640), .B(net_17253) );
NOR2_X2 inst_4335 ( .A1(net_13576), .A2(net_10246), .ZN(net_5723) );
NOR2_X2 inst_4187 ( .ZN(net_8045), .A1(net_6743), .A2(net_6742) );
NOR2_X2 inst_4239 ( .ZN(net_7814), .A2(net_4871), .A1(net_1124) );
INV_X4 inst_15586 ( .ZN(net_2782), .A(net_1373) );
DFF_X1 inst_19806 ( .D(net_18156), .CK(net_22390), .Q(x804) );
NAND2_X4 inst_7335 ( .ZN(net_6056), .A2(net_3438), .A1(net_940) );
AND2_X4 inst_21159 ( .ZN(net_19467), .A1(net_14083), .A2(net_11903) );
INV_X8 inst_12171 ( .ZN(net_18153), .A(net_18128) );
OR2_X4 inst_1121 ( .A1(net_2274), .A2(net_1645), .ZN(net_1148) );
INV_X8 inst_12185 ( .ZN(net_16973), .A(net_16808) );
NAND2_X2 inst_8932 ( .ZN(net_20364), .A1(net_13599), .A2(net_12225) );
NOR2_X4 inst_3187 ( .ZN(net_5433), .A2(net_3110), .A1(net_1523) );
CLKBUF_X2 inst_22407 ( .A(net_22278), .Z(net_22279) );
INV_X4 inst_18213 ( .A(net_21157), .ZN(net_16462) );
NAND2_X2 inst_11053 ( .ZN(net_4695), .A1(net_4694), .A2(net_2933) );
INV_X4 inst_17294 ( .ZN(net_5877), .A(net_673) );
XNOR2_X2 inst_307 ( .ZN(net_17093), .A(net_17092), .B(net_10804) );
NAND2_X2 inst_8411 ( .ZN(net_19396), .A1(net_17233), .A2(net_17232) );
CLKBUF_X2 inst_22078 ( .A(net_21949), .Z(net_21950) );
NAND2_X2 inst_8292 ( .ZN(net_17614), .A1(net_17529), .A2(net_17203) );
INV_X4 inst_12663 ( .ZN(net_17808), .A(net_17807) );
INV_X4 inst_18291 ( .A(net_20219), .ZN(net_20217) );
OAI21_X2 inst_2034 ( .ZN(net_11308), .B1(net_11307), .A(net_10976), .B2(net_9776) );
INV_X4 inst_16354 ( .ZN(net_1837), .A(net_1561) );
SDFF_X2 inst_717 ( .Q(net_20922), .SE(net_18856), .SI(net_18757), .D(net_414), .CK(net_21293) );
OAI21_X4 inst_1505 ( .ZN(net_9979), .A(net_5516), .B1(net_4744), .B2(net_4742) );
INV_X4 inst_15097 ( .ZN(net_4503), .A(net_3233) );
NAND2_X2 inst_10439 ( .ZN(net_7194), .A1(net_7193), .A2(net_7192) );
NAND2_X2 inst_8460 ( .A1(net_20069), .ZN(net_17054), .A2(net_16594) );
NAND2_X2 inst_11557 ( .ZN(net_7748), .A2(net_1762), .A1(net_1345) );
NAND2_X4 inst_7166 ( .ZN(net_12528), .A1(net_9356), .A2(net_7874) );
INV_X2 inst_19037 ( .ZN(net_4832), .A(net_4831) );
INV_X2 inst_19495 ( .ZN(net_2326), .A(net_1284) );
INV_X4 inst_16693 ( .ZN(net_4907), .A(net_3750) );
NAND2_X2 inst_7944 ( .ZN(net_18417), .A1(net_18298), .A2(net_18259) );
NOR2_X2 inst_3686 ( .ZN(net_11415), .A1(net_9574), .A2(net_9288) );
INV_X4 inst_15956 ( .ZN(net_8618), .A(net_5576) );
NOR2_X2 inst_3842 ( .A1(net_10319), .ZN(net_9596), .A2(net_7621) );
INV_X8 inst_12186 ( .ZN(net_17445), .A(net_17052) );
OAI21_X2 inst_1703 ( .ZN(net_15291), .B1(net_14157), .B2(net_12529), .A(net_1171) );
NAND3_X2 inst_5886 ( .A3(net_20045), .A1(net_20044), .ZN(net_19523), .A2(net_11795) );
NAND3_X2 inst_6566 ( .ZN(net_10479), .A3(net_7908), .A2(net_5912), .A1(net_5507) );
DFF_X1 inst_19807 ( .D(net_18155), .CK(net_22386), .Q(x815) );
NAND2_X4 inst_7167 ( .ZN(net_11642), .A2(net_9430), .A1(net_6617) );
INV_X2 inst_19488 ( .ZN(net_2218), .A(net_2096) );
INV_X4 inst_18122 ( .A(net_20981), .ZN(net_2515) );
INV_X4 inst_14894 ( .ZN(net_13871), .A(net_4034) );
INV_X4 inst_14139 ( .ZN(net_7510), .A(net_6080) );
INV_X4 inst_13680 ( .ZN(net_7994), .A(net_7993) );
NAND2_X2 inst_7788 ( .A2(net_18721), .ZN(net_18720), .A1(net_17388) );
INV_X4 inst_16358 ( .ZN(net_11572), .A(net_8286) );
NAND2_X2 inst_8934 ( .ZN(net_14854), .A2(net_14148), .A1(net_10054) );
XNOR2_X2 inst_614 ( .B(net_16836), .ZN(net_492), .A(net_491) );
CLKBUF_X2 inst_22876 ( .A(net_22747), .Z(net_22748) );
NAND2_X2 inst_9080 ( .ZN(net_13829), .A2(net_11687), .A1(net_1890) );
INV_X8 inst_12197 ( .ZN(net_16576), .A(net_16337) );
OAI21_X2 inst_1896 ( .A(net_15366), .ZN(net_13360), .B2(net_10009), .B1(net_8424) );
SDFF_X2 inst_1031 ( .QN(net_21029), .D(net_853), .SE(net_263), .CK(net_21881), .SI(x2508) );
SDFF_X2 inst_945 ( .QN(net_20990), .D(net_2472), .SE(net_263), .CK(net_21854), .SI(x3163) );
INV_X4 inst_17012 ( .ZN(net_2009), .A(net_1114) );
XNOR2_X2 inst_369 ( .ZN(net_16847), .A(net_16846), .B(net_7649) );
OAI21_X2 inst_1900 ( .ZN(net_13351), .A(net_13350), .B1(net_11317), .B2(net_8633) );
INV_X4 inst_15044 ( .ZN(net_4398), .A(net_3329) );
INV_X4 inst_12899 ( .A(net_17129), .ZN(net_16948) );
INV_X4 inst_12850 ( .ZN(net_17355), .A(net_17235) );
NAND3_X2 inst_5695 ( .ZN(net_16256), .A3(net_15951), .A2(net_14475), .A1(net_13614) );
NOR2_X4 inst_2916 ( .ZN(net_9669), .A2(net_8160), .A1(net_6233) );
CLKBUF_X2 inst_22067 ( .A(net_21938), .Z(net_21939) );
AOI21_X2 inst_20842 ( .A(net_12295), .ZN(net_9265), .B2(net_4597), .B1(net_2185) );
OAI22_X2 inst_1286 ( .ZN(net_14243), .A2(net_14242), .B1(net_14241), .B2(net_13955), .A1(net_12546) );
NAND2_X2 inst_8812 ( .ZN(net_15611), .A2(net_14925), .A1(net_14476) );
INV_X2 inst_18599 ( .ZN(net_9976), .A(net_9975) );
XNOR2_X2 inst_77 ( .B(net_21161), .ZN(net_18681), .A(net_18680) );
NAND3_X2 inst_6399 ( .ZN(net_11990), .A3(net_11828), .A1(net_9988), .A2(net_7419) );
NAND2_X2 inst_8224 ( .A2(net_20666), .A1(net_20665), .ZN(net_17863) );
INV_X4 inst_17010 ( .ZN(net_7858), .A(net_4711) );
INV_X4 inst_17435 ( .ZN(net_15048), .A(net_278) );
INV_X4 inst_13328 ( .ZN(net_12455), .A(net_11178) );
NAND2_X2 inst_11710 ( .ZN(net_3307), .A2(net_1680), .A1(net_896) );
NAND2_X4 inst_7086 ( .A1(net_20664), .ZN(net_15583), .A2(net_15582) );
NAND2_X2 inst_9642 ( .ZN(net_10387), .A1(net_10386), .A2(net_9815) );
INV_X2 inst_18483 ( .ZN(net_12486), .A(net_11241) );
AND2_X2 inst_21288 ( .ZN(net_12178), .A2(net_12177), .A1(net_12174) );
DFF_X1 inst_19837 ( .D(net_17407), .CK(net_22115), .Q(x329) );
INV_X4 inst_15713 ( .ZN(net_7667), .A(net_1504) );
NAND2_X2 inst_11881 ( .A2(net_5342), .ZN(net_1618), .A1(net_247) );
INV_X2 inst_19070 ( .ZN(net_4629), .A(net_3970) );
AOI21_X2 inst_20397 ( .ZN(net_15439), .A(net_14500), .B2(net_14445), .B1(net_13034) );
INV_X4 inst_13553 ( .ZN(net_10740), .A(net_9164) );
INV_X4 inst_14691 ( .ZN(net_4816), .A(net_3824) );
NAND2_X2 inst_9637 ( .A1(net_14820), .ZN(net_10397), .A2(net_7763) );
INV_X2 inst_19199 ( .A(net_4951), .ZN(net_3587) );
OR2_X2 inst_1234 ( .A2(net_6520), .ZN(net_4198), .A1(net_1515) );
AOI22_X2 inst_20048 ( .A1(net_4502), .ZN(net_4423), .B2(net_2457), .A2(net_1428), .B1(net_303) );
CLKBUF_X2 inst_22945 ( .A(net_22539), .Z(net_22817) );
NAND2_X2 inst_10040 ( .ZN(net_8718), .A1(net_8717), .A2(net_6408) );
INV_X4 inst_16564 ( .ZN(net_14378), .A(net_5716) );
OAI211_X2 inst_2398 ( .ZN(net_16052), .A(net_15480), .C2(net_15170), .B(net_14403), .C1(net_3296) );
OAI211_X2 inst_2595 ( .ZN(net_5257), .C2(net_5256), .A(net_4950), .B(net_4673), .C1(net_1818) );
NAND3_X4 inst_5614 ( .ZN(net_13281), .A1(net_8775), .A3(net_8767), .A2(net_5715) );
NAND2_X2 inst_11938 ( .A1(net_8304), .ZN(net_1958), .A2(net_1477) );
NAND2_X2 inst_9400 ( .ZN(net_11696), .A2(net_11695), .A1(net_5087) );
OAI211_X4 inst_2371 ( .C2(net_20928), .C1(net_19230), .ZN(net_16709), .B(net_16173), .A(net_11661) );
NOR2_X4 inst_2939 ( .A2(net_19488), .A1(net_19487), .ZN(net_7552) );
NAND3_X2 inst_6818 ( .A1(net_4079), .A2(net_3929), .A3(net_2384), .ZN(net_2059) );
OR2_X2 inst_1223 ( .ZN(net_5299), .A1(net_4037), .A2(net_2485) );
NOR3_X2 inst_2785 ( .ZN(net_12927), .A1(net_5733), .A3(net_4406), .A2(net_2454) );
INV_X4 inst_13636 ( .ZN(net_8212), .A(net_8211) );
NAND3_X2 inst_6574 ( .A3(net_11640), .ZN(net_10456), .A2(net_8085), .A1(net_4936) );
INV_X2 inst_18578 ( .A(net_12196), .ZN(net_10402) );
XNOR2_X1 inst_681 ( .A(net_18147), .ZN(net_18105), .B(net_17144) );
NAND4_X2 inst_5432 ( .A2(net_20414), .A1(net_20413), .A3(net_15844), .ZN(net_14108), .A4(net_13632) );
INV_X4 inst_13785 ( .A(net_7571), .ZN(net_7570) );
NAND2_X4 inst_7665 ( .ZN(net_1040), .A1(net_897), .A2(net_805) );
NOR2_X2 inst_4886 ( .A2(net_10810), .A1(net_2164), .ZN(net_2131) );
INV_X4 inst_15376 ( .ZN(net_14363), .A(net_12881) );
OAI21_X2 inst_2010 ( .ZN(net_11387), .A(net_10381), .B1(net_9252), .B2(net_7536) );
INV_X4 inst_13181 ( .ZN(net_14325), .A(net_13853) );
INV_X4 inst_15604 ( .ZN(net_11909), .A(net_2212) );
NAND2_X2 inst_11575 ( .A2(net_9364), .A1(net_3446), .ZN(net_2743) );
AND2_X4 inst_21176 ( .ZN(net_19100), .A2(net_12124), .A1(net_10643) );
NAND3_X4 inst_5547 ( .A3(net_20199), .A1(net_20198), .ZN(net_16520), .A2(net_10825) );
SDFF_X2 inst_871 ( .Q(net_21222), .SI(net_17087), .SE(net_125), .CK(net_21460), .D(x7296) );
NOR3_X2 inst_2684 ( .ZN(net_14438), .A2(net_14437), .A1(net_12803), .A3(net_11252) );
NAND3_X2 inst_6320 ( .ZN(net_12560), .A3(net_10639), .A2(net_8833), .A1(net_5943) );
NAND2_X4 inst_6842 ( .A2(net_19233), .A1(net_19232), .ZN(net_18690) );
OR2_X2 inst_1171 ( .A2(net_7665), .ZN(net_6322), .A1(net_6321) );
INV_X2 inst_18770 ( .A(net_9618), .ZN(net_7579) );
NAND4_X2 inst_5274 ( .ZN(net_16085), .A4(net_15490), .A2(net_14339), .A3(net_13816), .A1(net_12967) );
NAND4_X2 inst_5493 ( .ZN(net_12237), .A1(net_12236), .A3(net_11594), .A4(net_8544), .A2(net_8363) );
NAND3_X4 inst_5616 ( .ZN(net_19924), .A3(net_12124), .A2(net_7522), .A1(net_5686) );
NAND2_X2 inst_8192 ( .ZN(net_17896), .A1(net_17783), .A2(net_17595) );
NAND3_X2 inst_5766 ( .ZN(net_19590), .A3(net_15387), .A2(net_13349), .A1(net_11586) );
CLKBUF_X2 inst_22063 ( .A(net_21934), .Z(net_21935) );
INV_X4 inst_18026 ( .A(net_21130), .ZN(net_17534) );
OAI211_X2 inst_2594 ( .ZN(net_5261), .A(net_5260), .B(net_5259), .C2(net_1807), .C1(net_1521) );
NOR2_X2 inst_5113 ( .A2(net_20876), .A1(net_20875), .ZN(net_556) );
INV_X4 inst_16474 ( .ZN(net_8202), .A(net_1505) );
AND2_X4 inst_21188 ( .ZN(net_14350), .A2(net_10952), .A1(net_1233) );
CLKBUF_X2 inst_21586 ( .A(net_21457), .Z(net_21458) );
INV_X4 inst_14052 ( .ZN(net_19319), .A(net_6250) );
NOR2_X2 inst_3976 ( .ZN(net_18963), .A2(net_9973), .A1(net_8397) );
CLKBUF_X2 inst_22835 ( .A(net_22416), .Z(net_22707) );
NAND2_X2 inst_11773 ( .A1(net_20495), .ZN(net_4673), .A2(net_2350) );
NAND2_X2 inst_9444 ( .ZN(net_13812), .A2(net_11542), .A1(net_2484) );
CLKBUF_X2 inst_21494 ( .A(net_21365), .Z(net_21366) );
INV_X2 inst_19378 ( .ZN(net_2159), .A(net_2158) );
OR2_X4 inst_1119 ( .ZN(net_2751), .A2(net_1002), .A1(net_896) );
INV_X4 inst_15430 ( .ZN(net_2881), .A(net_2506) );
INV_X4 inst_14748 ( .ZN(net_4078), .A(net_4077) );
NOR2_X2 inst_3699 ( .ZN(net_19249), .A1(net_7453), .A2(net_5188) );
NOR2_X2 inst_5082 ( .A2(net_20495), .A1(net_955), .ZN(net_858) );
NAND2_X2 inst_9684 ( .A2(net_11763), .ZN(net_10256), .A1(net_7434) );
NOR2_X2 inst_5050 ( .ZN(net_2337), .A2(net_1588), .A1(net_170) );
NAND2_X2 inst_10947 ( .ZN(net_8980), .A2(net_5127), .A1(net_2376) );
INV_X4 inst_17310 ( .ZN(net_597), .A(net_596) );
AOI21_X2 inst_20353 ( .B1(net_20586), .ZN(net_15701), .A(net_13144), .B2(net_1774) );
NAND2_X2 inst_9112 ( .ZN(net_13581), .A2(net_13580), .A1(net_13364) );
NOR2_X2 inst_4925 ( .A1(net_3696), .ZN(net_2518), .A2(net_1813) );
CLKBUF_X2 inst_22075 ( .A(net_21946), .Z(net_21947) );
CLKBUF_X2 inst_22639 ( .A(net_22510), .Z(net_22511) );
NAND2_X4 inst_7021 ( .ZN(net_17380), .A1(net_16565), .A2(net_16452) );
NOR2_X2 inst_4457 ( .A1(net_5032), .ZN(net_4662), .A2(net_2152) );
NAND3_X2 inst_6133 ( .ZN(net_13738), .A3(net_12607), .A2(net_11083), .A1(net_8410) );
SDFF_X2 inst_903 ( .Q(net_21122), .D(net_16831), .SE(net_263), .CK(net_22431), .SI(x4319) );
INV_X4 inst_14806 ( .ZN(net_3980), .A(net_3979) );
OAI21_X2 inst_1725 ( .A(net_15974), .ZN(net_15092), .B2(net_13061), .B1(net_11780) );
NAND4_X2 inst_5391 ( .ZN(net_14896), .A2(net_12588), .A1(net_12375), .A4(net_11437), .A3(net_9730) );
NAND2_X4 inst_7238 ( .ZN(net_10604), .A1(net_7009), .A2(net_6604) );
CLKBUF_X2 inst_22891 ( .A(net_21379), .Z(net_22763) );
NAND2_X2 inst_8607 ( .A2(net_16996), .ZN(net_16660), .A1(net_16659) );
NAND2_X2 inst_8602 ( .A2(net_17517), .ZN(net_16673), .A1(net_15588) );
NAND2_X2 inst_9700 ( .ZN(net_10214), .A2(net_10213), .A1(net_7485) );
NOR2_X2 inst_3504 ( .ZN(net_13986), .A2(net_12057), .A1(net_11747) );
NOR2_X2 inst_3924 ( .A1(net_9791), .ZN(net_8776), .A2(net_8126) );
AOI21_X2 inst_20918 ( .A(net_10286), .B2(net_9921), .ZN(net_7311), .B1(net_3618) );
INV_X4 inst_17365 ( .ZN(net_3630), .A(net_546) );
INV_X4 inst_14408 ( .ZN(net_11282), .A(net_5095) );
NOR2_X2 inst_4510 ( .ZN(net_6634), .A2(net_1544), .A1(net_167) );
NAND2_X2 inst_9548 ( .ZN(net_11033), .A1(net_11032), .A2(net_10915) );
NOR2_X2 inst_4572 ( .ZN(net_9993), .A2(net_3149), .A1(net_1215) );
NAND4_X4 inst_5189 ( .A4(net_19577), .A1(net_19576), .A3(net_18890), .ZN(net_16524), .A2(net_15963) );
INV_X4 inst_13053 ( .A(net_16556), .ZN(net_16447) );
INV_X4 inst_17995 ( .A(net_20919), .ZN(net_325) );
INV_X4 inst_17904 ( .A(net_1339), .ZN(net_59) );
NAND2_X2 inst_11203 ( .ZN(net_13840), .A2(net_2888), .A1(net_154) );
NOR2_X2 inst_3464 ( .ZN(net_19279), .A2(net_13308), .A1(net_9196) );
SDFF_X2 inst_1044 ( .QN(net_21063), .D(net_520), .SE(net_263), .CK(net_21701), .SI(x2019) );
NAND2_X2 inst_9233 ( .ZN(net_14302), .A1(net_13093), .A2(net_12720) );
NAND3_X2 inst_6187 ( .ZN(net_19566), .A3(net_9155), .A2(net_7981), .A1(net_7066) );
INV_X2 inst_18907 ( .ZN(net_9680), .A(net_8093) );
NAND2_X2 inst_10309 ( .ZN(net_11855), .A2(net_7851), .A1(net_6647) );
NAND2_X4 inst_7554 ( .ZN(net_3070), .A2(net_2497), .A1(net_1752) );
NAND2_X2 inst_9509 ( .ZN(net_12526), .A1(net_10319), .A2(net_7898) );
INV_X4 inst_16377 ( .ZN(net_7812), .A(net_1279) );
INV_X4 inst_16086 ( .ZN(net_8068), .A(net_399) );
INV_X4 inst_14389 ( .A(net_9558), .ZN(net_5138) );
INV_X4 inst_17191 ( .A(net_4205), .ZN(net_1698) );
NAND2_X2 inst_8327 ( .ZN(net_19920), .A2(net_17504), .A1(net_17195) );
NOR2_X4 inst_3014 ( .ZN(net_5975), .A1(net_3131), .A2(net_2585) );
INV_X4 inst_16396 ( .A(net_4704), .ZN(net_2974) );
INV_X4 inst_15112 ( .ZN(net_5574), .A(net_3191) );
NAND3_X2 inst_6256 ( .ZN(net_13003), .A2(net_13002), .A3(net_13001), .A1(net_6152) );
XNOR2_X2 inst_227 ( .ZN(net_17567), .B(net_17500), .A(net_16844) );
OAI21_X2 inst_1532 ( .B1(net_18003), .ZN(net_17977), .B2(net_17849), .A(net_2036) );
NOR2_X2 inst_4303 ( .ZN(net_5938), .A2(net_5937), .A1(net_120) );
NAND3_X2 inst_5861 ( .ZN(net_15339), .A3(net_13735), .A2(net_13678), .A1(net_11310) );
OAI21_X2 inst_2136 ( .ZN(net_9986), .A(net_9985), .B1(net_9984), .B2(net_9983) );
INV_X4 inst_16872 ( .ZN(net_14643), .A(net_14022) );
NOR2_X4 inst_2891 ( .ZN(net_10954), .A1(net_7476), .A2(net_2828) );
INV_X4 inst_17830 ( .ZN(net_1655), .A(net_268) );
INV_X2 inst_18491 ( .ZN(net_12335), .A(net_12334) );
INV_X4 inst_17260 ( .A(net_2709), .ZN(net_1604) );
NAND2_X4 inst_7557 ( .A1(net_20868), .ZN(net_2111), .A2(net_1074) );
NAND2_X2 inst_8642 ( .A1(net_16801), .A2(net_16774), .ZN(net_16573) );
NAND3_X2 inst_6036 ( .ZN(net_14332), .A2(net_14331), .A3(net_14330), .A1(net_7223) );
INV_X2 inst_18381 ( .ZN(net_16785), .A(net_16784) );
NAND2_X2 inst_9944 ( .A1(net_11366), .ZN(net_9059), .A2(net_8247) );
INV_X4 inst_17539 ( .ZN(net_3704), .A(net_153) );
NOR2_X2 inst_5029 ( .A1(net_1798), .ZN(net_1149), .A2(net_1148) );
NAND2_X2 inst_10200 ( .A1(net_10236), .A2(net_9967), .ZN(net_8125) );
INV_X2 inst_18637 ( .A(net_12056), .ZN(net_9390) );
INV_X4 inst_15457 ( .ZN(net_14700), .A(net_14463) );
XNOR2_X2 inst_581 ( .B(net_16982), .ZN(net_600), .A(net_599) );
OAI211_X2 inst_2551 ( .ZN(net_10813), .B(net_10812), .A(net_6459), .C2(net_4611), .C1(net_2980) );
XOR2_X2 inst_28 ( .B(net_21113), .Z(net_15958), .A(net_15957) );
NOR2_X2 inst_4407 ( .ZN(net_6227), .A1(net_6127), .A2(net_5082) );
INV_X4 inst_17928 ( .A(net_21234), .ZN(net_230) );
CLKBUF_X2 inst_22748 ( .A(net_22619), .Z(net_22620) );
INV_X4 inst_16517 ( .A(net_1599), .ZN(net_1188) );
NAND2_X2 inst_9410 ( .A2(net_12999), .ZN(net_11660), .A1(net_11659) );
AOI21_X2 inst_20497 ( .B1(net_20781), .ZN(net_14713), .B2(net_12190), .A(net_7394) );
INV_X4 inst_12656 ( .A(net_17843), .ZN(net_17829) );
NAND2_X2 inst_9434 ( .A1(net_13007), .ZN(net_11595), .A2(net_11594) );
NAND2_X2 inst_9401 ( .ZN(net_11694), .A2(net_11693), .A1(net_8310) );
NAND2_X4 inst_7440 ( .ZN(net_5232), .A1(net_3276), .A2(net_1468) );
INV_X4 inst_15869 ( .ZN(net_2757), .A(net_1799) );
XNOR2_X2 inst_592 ( .B(net_16743), .ZN(net_561), .A(net_560) );
NAND2_X4 inst_7289 ( .ZN(net_5942), .A2(net_5333), .A1(net_4163) );
INV_X4 inst_13841 ( .ZN(net_10874), .A(net_7482) );
NOR2_X2 inst_5143 ( .A2(net_220), .ZN(net_139), .A1(net_39) );
AOI21_X2 inst_20387 ( .ZN(net_19288), .B1(net_14731), .B2(net_14584), .A(net_14401) );
INV_X4 inst_15118 ( .ZN(net_3585), .A(net_3181) );
INV_X4 inst_16621 ( .ZN(net_1113), .A(net_1112) );
INV_X2 inst_19521 ( .A(net_1844), .ZN(net_1108) );
INV_X4 inst_13504 ( .A(net_11832), .ZN(net_9419) );
NAND2_X2 inst_7858 ( .ZN(net_18571), .A1(net_18556), .A2(net_18545) );
INV_X4 inst_14755 ( .ZN(net_8901), .A(net_5475) );
INV_X4 inst_12876 ( .ZN(net_18405), .A(net_18326) );
NOR2_X2 inst_5096 ( .A2(net_834), .ZN(net_806), .A1(net_805) );
NOR2_X2 inst_3948 ( .ZN(net_8615), .A2(net_7965), .A1(net_3052) );
NAND2_X2 inst_11413 ( .A1(net_9943), .ZN(net_5407), .A2(net_4289) );
NAND4_X4 inst_5227 ( .A2(net_19842), .A1(net_19841), .ZN(net_16274), .A4(net_14752), .A3(net_8530) );
INV_X4 inst_16278 ( .ZN(net_1695), .A(net_1420) );
INV_X4 inst_14157 ( .ZN(net_8590), .A(net_7232) );
NAND2_X2 inst_11808 ( .ZN(net_2868), .A2(net_2089), .A1(net_221) );
CLKBUF_X2 inst_22663 ( .A(net_21889), .Z(net_22535) );
INV_X2 inst_18743 ( .ZN(net_7905), .A(net_7904) );
OAI22_X2 inst_1301 ( .ZN(net_11223), .B2(net_10444), .A2(net_10431), .B1(net_9387), .A1(net_7071) );
INV_X4 inst_14109 ( .ZN(net_7553), .A(net_6161) );
XNOR2_X2 inst_647 ( .A(net_17494), .B(net_17247), .ZN(net_13946) );
NOR2_X4 inst_2830 ( .ZN(net_19003), .A2(net_15504), .A1(net_15349) );
INV_X2 inst_19559 ( .A(net_1328), .ZN(net_838) );
INV_X4 inst_12871 ( .A(net_17658), .ZN(net_16951) );
INV_X2 inst_18736 ( .ZN(net_7926), .A(net_7925) );
NOR2_X2 inst_5137 ( .A2(net_1719), .ZN(net_183), .A1(net_107) );
CLKBUF_X2 inst_21705 ( .A(net_21312), .Z(net_21577) );
NOR2_X4 inst_2985 ( .ZN(net_11034), .A2(net_4608), .A1(net_1050) );
AOI21_X2 inst_20978 ( .ZN(net_3712), .A(net_3711), .B1(net_3710), .B2(net_2180) );
NAND2_X2 inst_9821 ( .A1(net_12326), .ZN(net_9643), .A2(net_9642) );
NAND2_X2 inst_8156 ( .ZN(net_18000), .A2(net_17964), .A1(net_17734) );
AOI22_X2 inst_19979 ( .ZN(net_15480), .B1(net_15099), .A2(net_14607), .B2(net_11378), .A1(net_1277) );
SDFF_X2 inst_833 ( .Q(net_21174), .SI(net_17508), .SE(net_125), .CK(net_22164), .D(x4734) );
NAND2_X2 inst_11968 ( .A2(net_5162), .ZN(net_3238), .A1(net_1363) );
XNOR2_X2 inst_118 ( .ZN(net_18475), .A(net_18359), .B(net_17577) );
NOR2_X2 inst_4924 ( .ZN(net_3216), .A2(net_1823), .A1(net_222) );
INV_X4 inst_12709 ( .ZN(net_17566), .A(net_17565) );
INV_X4 inst_14433 ( .ZN(net_5025), .A(net_5024) );
NAND2_X2 inst_10781 ( .A1(net_20923), .A2(net_7146), .ZN(net_6967) );
NAND3_X2 inst_6591 ( .ZN(net_9962), .A3(net_9961), .A2(net_8378), .A1(net_6542) );
OAI21_X2 inst_2037 ( .B1(net_13554), .ZN(net_11304), .B2(net_9741), .A(net_5346) );
NAND2_X2 inst_8578 ( .ZN(net_16726), .A1(net_16630), .A2(net_16537) );
INV_X4 inst_13532 ( .A(net_11435), .ZN(net_9218) );
NAND2_X4 inst_6930 ( .ZN(net_17604), .A1(net_17603), .A2(net_17602) );
NAND2_X2 inst_9102 ( .ZN(net_13763), .A1(net_13762), .A2(net_13761) );
INV_X4 inst_15343 ( .ZN(net_4855), .A(net_1954) );
INV_X8 inst_12276 ( .ZN(net_2037), .A(net_1398) );
SDFF_X2 inst_883 ( .Q(net_21243), .SI(net_16953), .SE(net_125), .CK(net_21538), .D(x6631) );
CLKBUF_X2 inst_22287 ( .A(net_22158), .Z(net_22159) );
INV_X4 inst_12536 ( .ZN(net_18376), .A(net_18375) );
INV_X4 inst_12710 ( .ZN(net_17564), .A(net_17563) );
SDFF_X2 inst_756 ( .Q(net_20932), .SE(net_18858), .SI(net_18531), .D(net_715), .CK(net_21438) );
CLKBUF_X2 inst_21634 ( .A(net_21505), .Z(net_21506) );
INV_X2 inst_19711 ( .A(net_20711), .ZN(net_20710) );
CLKBUF_X2 inst_21854 ( .A(net_21725), .Z(net_21726) );
INV_X4 inst_13423 ( .ZN(net_10783), .A(net_10080) );
NAND2_X2 inst_9270 ( .ZN(net_14873), .A2(net_10910), .A1(net_10714) );
INV_X4 inst_15628 ( .ZN(net_3787), .A(net_3034) );
NAND2_X4 inst_7150 ( .ZN(net_11707), .A2(net_9532), .A1(net_6655) );
INV_X2 inst_19431 ( .ZN(net_2925), .A(net_2242) );
INV_X4 inst_15500 ( .ZN(net_12714), .A(net_2423) );
NAND2_X2 inst_9873 ( .A1(net_10188), .ZN(net_9464), .A2(net_9463) );
NAND2_X2 inst_9685 ( .ZN(net_13101), .A1(net_10255), .A2(net_10254) );
OR2_X2 inst_1165 ( .ZN(net_11725), .A1(net_7156), .A2(net_6384) );
NAND4_X2 inst_5439 ( .ZN(net_19657), .A3(net_12284), .A4(net_12282), .A1(net_10094), .A2(net_8454) );
NAND2_X2 inst_11029 ( .ZN(net_4774), .A1(net_4773), .A2(net_3515) );
NAND2_X2 inst_8891 ( .ZN(net_15116), .A1(net_15048), .A2(net_13958) );
NOR3_X2 inst_2644 ( .ZN(net_15899), .A1(net_15488), .A3(net_15141), .A2(net_10003) );
NAND2_X4 inst_6922 ( .A1(net_20463), .ZN(net_19771), .A2(net_17278) );
CLKBUF_X2 inst_22605 ( .A(net_22476), .Z(net_22477) );
NOR3_X4 inst_2626 ( .ZN(net_19131), .A2(net_12615), .A3(net_12030), .A1(net_10347) );
NAND2_X2 inst_9314 ( .ZN(net_12352), .A1(net_12326), .A2(net_9017) );
NOR2_X2 inst_4629 ( .ZN(net_3594), .A1(net_2142), .A2(net_1863) );
INV_X4 inst_17307 ( .ZN(net_10048), .A(net_603) );
INV_X4 inst_14140 ( .ZN(net_9388), .A(net_6079) );
NAND3_X2 inst_5983 ( .ZN(net_14546), .A2(net_14545), .A3(net_14544), .A1(net_13401) );
INV_X2 inst_19599 ( .A(net_311), .ZN(net_175) );
NAND2_X2 inst_9056 ( .ZN(net_14001), .A1(net_11983), .A2(net_11981) );
INV_X4 inst_17629 ( .ZN(net_290), .A(net_289) );
INV_X4 inst_16825 ( .ZN(net_10550), .A(net_6316) );
NAND2_X4 inst_6883 ( .A2(net_18192), .ZN(net_18165), .A1(net_16757) );
INV_X4 inst_17107 ( .ZN(net_10914), .A(net_5107) );
SDFF_X2 inst_992 ( .QN(net_21055), .D(net_637), .SE(net_263), .CK(net_22501), .SI(x2127) );
INV_X4 inst_18040 ( .A(net_20949), .ZN(net_63) );
XNOR2_X2 inst_488 ( .ZN(net_9259), .A(net_9258), .B(net_1860) );
INV_X4 inst_14085 ( .A(net_6215), .ZN(net_6214) );
NAND2_X2 inst_7809 ( .A2(net_18696), .ZN(net_18682), .A1(net_488) );
NAND4_X4 inst_5196 ( .A2(net_19849), .A1(net_19848), .ZN(net_16843), .A4(net_16152), .A3(net_16144) );
CLKBUF_X2 inst_22611 ( .A(net_21617), .Z(net_22483) );
INV_X4 inst_18269 ( .A(net_19449), .ZN(net_19447) );
NAND2_X2 inst_8666 ( .A1(net_21123), .A2(net_16718), .ZN(net_16474) );
CLKBUF_X2 inst_22813 ( .A(net_22684), .Z(net_22685) );
NAND2_X4 inst_7308 ( .ZN(net_10773), .A1(net_5436), .A2(net_4792) );
XNOR2_X2 inst_254 ( .A(net_17312), .ZN(net_17295), .B(net_17294) );
NAND3_X2 inst_6053 ( .ZN(net_14233), .A3(net_12387), .A1(net_7897), .A2(net_7797) );
NAND2_X2 inst_9543 ( .ZN(net_20681), .A1(net_11432), .A2(net_11053) );
AOI22_X2 inst_20012 ( .ZN(net_20332), .B1(net_13871), .A2(net_11906), .B2(net_10648), .A1(net_4432) );
CLKBUF_X2 inst_22155 ( .A(net_21820), .Z(net_22027) );
OAI21_X4 inst_1412 ( .A(net_20928), .B2(net_19384), .B1(net_19383), .ZN(net_16173) );
NAND2_X2 inst_9862 ( .ZN(net_9494), .A1(net_9493), .A2(net_8475) );
INV_X4 inst_17066 ( .ZN(net_11466), .A(net_4702) );
NAND2_X2 inst_10957 ( .ZN(net_8310), .A2(net_3535), .A1(net_732) );
INV_X4 inst_15382 ( .ZN(net_5409), .A(net_2558) );
INV_X4 inst_13364 ( .ZN(net_13676), .A(net_10912) );
INV_X4 inst_12774 ( .ZN(net_17327), .A(net_17326) );
AOI21_X2 inst_20673 ( .ZN(net_12578), .B2(net_12487), .A(net_10345), .B1(net_7705) );
XNOR2_X2 inst_661 ( .A(net_21168), .B(net_21136), .ZN(net_13951) );
NAND3_X2 inst_6265 ( .ZN(net_12973), .A1(net_12746), .A2(net_10787), .A3(net_7016) );
NAND2_X4 inst_7416 ( .ZN(net_8938), .A1(net_3656), .A2(net_1033) );
NAND2_X2 inst_10817 ( .A1(net_6879), .A2(net_5571), .ZN(net_5508) );
OAI21_X2 inst_2073 ( .ZN(net_10594), .A(net_10593), .B1(net_10592), .B2(net_6447) );
NAND2_X4 inst_7346 ( .ZN(net_8833), .A1(net_5291), .A2(net_399) );
NAND2_X2 inst_8661 ( .A2(net_16815), .ZN(net_16518), .A1(net_4491) );
NAND2_X2 inst_11418 ( .ZN(net_8764), .A2(net_2894), .A1(net_2003) );
NOR2_X2 inst_3984 ( .ZN(net_8347), .A2(net_8345), .A1(net_4811) );
NOR2_X2 inst_4682 ( .ZN(net_5543), .A1(net_3205), .A2(net_2991) );
INV_X4 inst_17161 ( .A(net_2709), .ZN(net_748) );
NAND2_X2 inst_11310 ( .A1(net_20552), .ZN(net_4754), .A2(net_2715) );
XNOR2_X2 inst_419 ( .ZN(net_16532), .A(net_16530), .B(net_5236) );
NAND2_X4 inst_7488 ( .A2(net_20424), .ZN(net_2441), .A1(net_2380) );
INV_X4 inst_12546 ( .ZN(net_18419), .A(net_18288) );
NAND2_X2 inst_12098 ( .ZN(net_839), .A2(net_525), .A1(net_179) );
NAND3_X2 inst_6495 ( .A2(net_15366), .A3(net_14166), .ZN(net_10858), .A1(net_7639) );
INV_X4 inst_15763 ( .ZN(net_13700), .A(net_81) );
NAND2_X4 inst_6941 ( .A2(net_19244), .A1(net_19243), .ZN(net_17572) );
INV_X4 inst_18201 ( .A(net_21241), .ZN(net_1339) );
NAND2_X2 inst_10629 ( .A1(net_6863), .ZN(net_6551), .A2(net_6550) );
CLKBUF_X2 inst_22784 ( .A(net_22655), .Z(net_22656) );
INV_X4 inst_14298 ( .ZN(net_6857), .A(net_5539) );
INV_X4 inst_14283 ( .ZN(net_8057), .A(net_4064) );
INV_X4 inst_16222 ( .A(net_1499), .ZN(net_1387) );
INV_X8 inst_12377 ( .A(net_972), .ZN(net_181) );
NAND2_X2 inst_7898 ( .ZN(net_19692), .A2(net_18383), .A1(net_17887) );
INV_X4 inst_16848 ( .ZN(net_15044), .A(net_10686) );
INV_X4 inst_12749 ( .A(net_18704), .ZN(net_18684) );
NAND2_X2 inst_11160 ( .ZN(net_4190), .A1(net_1972), .A2(net_1142) );
XOR2_X2 inst_34 ( .A(net_21194), .Z(net_695), .B(net_694) );
NOR2_X2 inst_3717 ( .ZN(net_10978), .A2(net_10977), .A1(net_4032) );
NAND2_X2 inst_9120 ( .ZN(net_20170), .A2(net_13558), .A1(net_11894) );
XOR2_X2 inst_12 ( .Z(net_17037), .B(net_17036), .A(net_16657) );
INV_X4 inst_12690 ( .ZN(net_17666), .A(net_17665) );
NAND2_X2 inst_9823 ( .ZN(net_9637), .A1(net_9636), .A2(net_9635) );
INV_X4 inst_13946 ( .ZN(net_7292), .A(net_6798) );
INV_X2 inst_18520 ( .A(net_14533), .ZN(net_13695) );
INV_X2 inst_18674 ( .ZN(net_9114), .A(net_9113) );
NAND2_X2 inst_9856 ( .ZN(net_9511), .A1(net_9510), .A2(net_9509) );
OAI21_X4 inst_1424 ( .ZN(net_18984), .A(net_16210), .B2(net_15493), .B1(net_15152) );
OAI21_X4 inst_1425 ( .B1(net_20169), .ZN(net_16045), .A(net_15821), .B2(net_1915) );
DFF_X1 inst_19830 ( .D(net_17543), .CK(net_21612), .Q(x697) );
OAI21_X2 inst_2198 ( .ZN(net_8572), .A(net_8571), .B1(net_7679), .B2(net_6391) );
XNOR2_X2 inst_258 ( .B(net_21183), .ZN(net_17284), .A(net_16971) );
CLKBUF_X2 inst_22379 ( .A(net_22250), .Z(net_22251) );
OAI211_X2 inst_2405 ( .ZN(net_15732), .C1(net_15731), .C2(net_14526), .A(net_13925), .B(net_11991) );
INV_X4 inst_13126 ( .ZN(net_15383), .A(net_15134) );
NOR2_X4 inst_3076 ( .ZN(net_9971), .A1(net_4789), .A2(net_4383) );
CLKBUF_X2 inst_21472 ( .A(net_21343), .Z(net_21344) );
NAND2_X2 inst_10964 ( .A1(net_6876), .ZN(net_5061), .A2(net_5060) );
XNOR2_X2 inst_482 ( .ZN(net_10805), .A(net_10804), .B(net_5790) );
NAND2_X2 inst_9804 ( .ZN(net_9694), .A1(net_9693), .A2(net_8448) );
INV_X2 inst_19190 ( .ZN(net_3666), .A(net_3665) );
NOR2_X2 inst_3534 ( .ZN(net_13508), .A2(net_11013), .A1(net_2789) );
NOR2_X4 inst_3276 ( .ZN(net_2405), .A1(net_1645), .A2(net_1217) );
NAND2_X2 inst_10230 ( .ZN(net_10146), .A1(net_7995), .A2(net_5162) );
NOR2_X2 inst_3996 ( .ZN(net_20415), .A1(net_10225), .A2(net_8244) );
NAND2_X4 inst_7059 ( .A2(net_20888), .ZN(net_19847), .A1(net_19618) );
XNOR2_X2 inst_539 ( .B(net_21121), .ZN(net_980), .A(net_798) );
INV_X4 inst_12915 ( .ZN(net_17024), .A(net_16669) );
NAND2_X2 inst_11066 ( .ZN(net_4521), .A2(net_3419), .A1(net_154) );
CLKBUF_X2 inst_22601 ( .A(net_22472), .Z(net_22473) );
SDFF_X2 inst_895 ( .Q(net_21134), .D(net_16761), .SE(net_263), .CK(net_21386), .SI(x3820) );
NAND2_X2 inst_11042 ( .ZN(net_7819), .A1(net_6625), .A2(net_4319) );
NAND2_X2 inst_10054 ( .ZN(net_13159), .A2(net_8690), .A1(net_8224) );
AOI221_X2 inst_20087 ( .ZN(net_15678), .C1(net_15677), .C2(net_14440), .B2(net_7993), .A(net_7911), .B1(net_3378) );
AND2_X4 inst_21250 ( .ZN(net_5269), .A1(net_2183), .A2(net_222) );
NAND3_X2 inst_6583 ( .ZN(net_10436), .A3(net_10435), .A2(net_9631), .A1(net_6070) );
CLKBUF_X2 inst_22497 ( .A(net_22072), .Z(net_22369) );
AOI21_X4 inst_20206 ( .B1(net_18912), .ZN(net_14647), .B2(net_11526), .A(net_7696) );
NAND2_X2 inst_10034 ( .A1(net_11189), .ZN(net_8723), .A2(net_6773) );
OAI21_X2 inst_2341 ( .A(net_12478), .ZN(net_4665), .B2(net_4664), .B1(net_3617) );
NAND3_X4 inst_5526 ( .A2(net_19499), .A1(net_19498), .ZN(net_18089), .A3(net_18060) );
NAND2_X2 inst_10685 ( .ZN(net_20314), .A1(net_6127), .A2(net_6126) );
NAND2_X2 inst_10616 ( .ZN(net_15416), .A2(net_14222), .A1(net_2875) );
NOR2_X2 inst_4122 ( .ZN(net_7034), .A1(net_7033), .A2(net_3807) );
INV_X4 inst_12557 ( .ZN(net_18287), .A(net_18200) );
INV_X4 inst_13184 ( .ZN(net_14234), .A(net_13640) );
NAND2_X2 inst_9901 ( .ZN(net_13098), .A2(net_9329), .A1(net_5959) );
INV_X4 inst_16482 ( .ZN(net_1481), .A(net_1204) );
NAND2_X2 inst_10324 ( .ZN(net_9323), .A2(net_7803), .A1(net_3297) );
INV_X4 inst_16340 ( .ZN(net_7874), .A(net_6177) );
NAND2_X2 inst_9189 ( .ZN(net_19597), .A1(net_13126), .A2(net_13125) );
NOR2_X2 inst_4797 ( .ZN(net_4263), .A2(net_3075), .A1(net_628) );
NAND3_X2 inst_6082 ( .A2(net_20784), .ZN(net_13961), .A3(net_11149), .A1(net_8406) );
NAND2_X2 inst_8482 ( .A2(net_17242), .ZN(net_16978), .A1(net_742) );
SDFF_X2 inst_826 ( .Q(net_21197), .SI(net_17547), .SE(net_125), .CK(net_22327), .D(x6178) );
NAND2_X2 inst_9343 ( .ZN(net_12209), .A1(net_12208), .A2(net_12196) );
INV_X4 inst_16541 ( .A(net_15343), .ZN(net_15245) );
NOR2_X2 inst_4002 ( .A1(net_14006), .ZN(net_8143), .A2(net_7248) );
INV_X4 inst_14009 ( .ZN(net_13442), .A(net_6310) );
NAND2_X2 inst_10362 ( .ZN(net_10840), .A1(net_7427), .A2(net_4574) );
XNOR2_X2 inst_159 ( .ZN(net_17943), .A(net_17826), .B(net_980) );
NAND2_X4 inst_7042 ( .A2(net_20027), .A1(net_20026), .ZN(net_16510) );
INV_X4 inst_13220 ( .ZN(net_13628), .A(net_12783) );
INV_X2 inst_18680 ( .ZN(net_8805), .A(net_8804) );
NAND2_X2 inst_9572 ( .ZN(net_10957), .A1(net_10956), .A2(net_9200) );
INV_X4 inst_15281 ( .ZN(net_4196), .A(net_1849) );
AOI21_X4 inst_20104 ( .ZN(net_19200), .B1(net_16644), .A(net_16303), .B2(net_16196) );
NAND3_X2 inst_5759 ( .ZN(net_15994), .A3(net_15456), .A1(net_14710), .A2(net_10040) );
INV_X4 inst_13657 ( .A(net_8145), .ZN(net_8144) );
NAND2_X2 inst_11005 ( .A1(net_8115), .ZN(net_4885), .A2(net_2704) );
NAND3_X2 inst_6318 ( .ZN(net_12565), .A1(net_12564), .A3(net_12563), .A2(net_8306) );
NAND2_X4 inst_7379 ( .ZN(net_8949), .A1(net_4304), .A2(net_193) );
INV_X4 inst_15491 ( .ZN(net_12784), .A(net_2903) );
NAND2_X2 inst_8339 ( .ZN(net_17495), .A1(net_17494), .A2(net_17493) );
XOR2_X2 inst_19 ( .B(net_21135), .A(net_16885), .Z(net_16881) );
AOI211_X2 inst_21024 ( .ZN(net_14882), .A(net_14881), .B(net_12698), .C2(net_9382), .C1(net_4444) );
INV_X4 inst_13623 ( .A(net_8832), .ZN(net_8340) );
NAND2_X2 inst_11509 ( .ZN(net_9634), .A1(net_2326), .A2(net_1401) );
NAND2_X2 inst_10378 ( .A1(net_18025), .ZN(net_7388), .A2(net_669) );
INV_X4 inst_13599 ( .A(net_13655), .ZN(net_8738) );
NOR2_X2 inst_4268 ( .ZN(net_7584), .A1(net_3333), .A2(net_809) );
INV_X2 inst_18487 ( .A(net_12649), .ZN(net_12365) );
INV_X4 inst_14170 ( .A(net_13479), .ZN(net_5999) );
NOR2_X2 inst_3830 ( .A2(net_10251), .A1(net_10119), .ZN(net_9737) );
INV_X4 inst_16706 ( .A(net_15553), .ZN(net_15214) );
INV_X8 inst_12287 ( .ZN(net_2402), .A(net_1141) );
OAI21_X2 inst_1686 ( .ZN(net_15406), .B1(net_14600), .A(net_14344), .B2(net_13264) );
NAND2_X2 inst_10541 ( .A1(net_9937), .ZN(net_8103), .A2(net_6676) );
CLKBUF_X2 inst_22802 ( .A(net_22673), .Z(net_22674) );
INV_X4 inst_15732 ( .ZN(net_7862), .A(net_5387) );
INV_X4 inst_16724 ( .ZN(net_1771), .A(net_1054) );
OAI21_X2 inst_1789 ( .ZN(net_20163), .B2(net_11762), .B1(net_9912), .A(net_588) );
CLKBUF_X2 inst_22886 ( .A(net_21395), .Z(net_22758) );
INV_X4 inst_14664 ( .ZN(net_18863), .A(net_18025) );
NAND2_X4 inst_7192 ( .ZN(net_13173), .A2(net_8067), .A1(net_7880) );
INV_X4 inst_14832 ( .ZN(net_19816), .A(net_3873) );
INV_X4 inst_15803 ( .ZN(net_3389), .A(net_1887) );
INV_X4 inst_15951 ( .ZN(net_13076), .A(net_6733) );
INV_X4 inst_18251 ( .A(net_21101), .ZN(net_1511) );
NAND2_X2 inst_9437 ( .ZN(net_12677), .A1(net_11572), .A2(net_11571) );
NOR2_X2 inst_3441 ( .ZN(net_15054), .A2(net_13841), .A1(net_10349) );
NAND2_X4 inst_6955 ( .A2(net_20437), .ZN(net_18932), .A1(net_17363) );
CLKBUF_X2 inst_21925 ( .A(net_21444), .Z(net_21797) );
INV_X8 inst_12332 ( .A(net_990), .ZN(net_927) );
NAND2_X2 inst_9413 ( .ZN(net_11655), .A1(net_11654), .A2(net_9299) );
NAND2_X2 inst_8000 ( .ZN(net_18311), .A2(net_18310), .A1(net_17207) );
AND2_X2 inst_21350 ( .ZN(net_7519), .A1(net_1786), .A2(net_1771) );
NAND2_X2 inst_11535 ( .ZN(net_4950), .A2(net_2926), .A1(net_801) );
INV_X4 inst_15250 ( .A(net_3989), .ZN(net_2802) );
INV_X4 inst_17865 ( .ZN(net_309), .A(net_268) );
INV_X4 inst_16715 ( .ZN(net_11691), .A(net_10415) );
CLKBUF_X2 inst_21526 ( .A(net_21397), .Z(net_21398) );
INV_X4 inst_12516 ( .ZN(net_18599), .A(net_18595) );
INV_X4 inst_17791 ( .A(net_257), .ZN(net_135) );
NOR2_X2 inst_4860 ( .ZN(net_4174), .A1(net_3174), .A2(net_1695) );
INV_X4 inst_14923 ( .ZN(net_3561), .A(net_3560) );
INV_X8 inst_12226 ( .ZN(net_6233), .A(net_4473) );
NAND3_X2 inst_6770 ( .ZN(net_5293), .A2(net_5292), .A1(net_4987), .A3(net_3815) );
INV_X4 inst_16314 ( .ZN(net_1611), .A(net_1321) );
OAI221_X2 inst_1344 ( .ZN(net_13457), .C2(net_13456), .B1(net_11751), .C1(net_10864), .A(net_10589), .B2(net_5306) );
OAI21_X4 inst_1460 ( .B2(net_19390), .B1(net_19389), .ZN(net_15247), .A(net_1244) );
OAI21_X2 inst_2287 ( .ZN(net_6527), .A(net_6526), .B1(net_6525), .B2(net_6524) );
INV_X4 inst_17336 ( .ZN(net_2244), .A(net_319) );
NAND2_X2 inst_8968 ( .ZN(net_14523), .A2(net_13016), .A1(net_3828) );
NOR3_X4 inst_2630 ( .ZN(net_14611), .A1(net_13318), .A2(net_13018), .A3(net_12180) );
INV_X4 inst_15422 ( .A(net_9301), .ZN(net_8460) );
INV_X4 inst_17329 ( .ZN(net_4228), .A(net_2585) );
INV_X4 inst_17611 ( .A(net_21219), .ZN(net_949) );
OAI21_X4 inst_1443 ( .B2(net_20387), .B1(net_20386), .A(net_16394), .ZN(net_15762) );
SDFF_X2 inst_1028 ( .QN(net_21093), .D(net_452), .SE(net_263), .CK(net_22559), .SI(x1497) );
NAND3_X2 inst_5891 ( .ZN(net_20684), .A1(net_14485), .A3(net_14158), .A2(net_10663) );
NAND2_X2 inst_10107 ( .ZN(net_8433), .A2(net_5922), .A1(net_5206) );
NOR2_X2 inst_3935 ( .A1(net_11311), .ZN(net_10148), .A2(net_8702) );
NAND2_X2 inst_9645 ( .ZN(net_20835), .A1(net_10381), .A2(net_7760) );
OAI22_X2 inst_1271 ( .B1(net_21167), .A1(net_16879), .ZN(net_16875), .B2(net_16874), .A2(net_16521) );
NAND2_X2 inst_12110 ( .A2(net_2274), .ZN(net_706), .A1(net_308) );
OAI21_X2 inst_2321 ( .ZN(net_5666), .A(net_5665), .B1(net_5664), .B2(net_5256) );
INV_X4 inst_17503 ( .ZN(net_19718), .A(net_418) );
INV_X4 inst_13927 ( .ZN(net_10530), .A(net_6870) );
CLKBUF_X2 inst_22538 ( .A(net_22153), .Z(net_22410) );
NAND2_X2 inst_9928 ( .ZN(net_9187), .A2(net_9162), .A1(net_5635) );
NOR2_X2 inst_4425 ( .ZN(net_6110), .A2(net_4961), .A1(net_3852) );
CLKBUF_X2 inst_21423 ( .A(net_21294), .Z(net_21295) );
NAND2_X2 inst_9727 ( .ZN(net_13112), .A1(net_12070), .A2(net_11322) );
NOR2_X2 inst_4461 ( .ZN(net_20343), .A2(net_4530), .A1(net_2874) );
NAND3_X2 inst_6626 ( .ZN(net_9047), .A2(net_9046), .A3(net_9045), .A1(net_4787) );
INV_X4 inst_14332 ( .ZN(net_11679), .A(net_5410) );
NAND2_X4 inst_7407 ( .A1(net_19522), .ZN(net_6926), .A2(net_61) );
INV_X8 inst_12343 ( .ZN(net_1785), .A(net_1735) );
NAND2_X2 inst_10807 ( .A1(net_11016), .ZN(net_5531), .A2(net_2775) );
INV_X4 inst_17221 ( .ZN(net_3254), .A(net_154) );
OAI21_X2 inst_2236 ( .B1(net_11311), .ZN(net_7756), .B2(net_7755), .A(net_5280) );
NOR2_X2 inst_3368 ( .A2(net_17370), .ZN(net_16829), .A1(net_95) );
NAND2_X4 inst_7307 ( .ZN(net_6749), .A2(net_3909), .A1(net_143) );
CLKBUF_X2 inst_22388 ( .A(net_22259), .Z(net_22260) );
OAI21_X2 inst_1553 ( .ZN(net_17701), .B2(net_17607), .A(net_17449), .B1(net_17448) );
INV_X4 inst_13038 ( .ZN(net_16912), .A(net_16576) );
INV_X4 inst_13937 ( .ZN(net_8147), .A(net_6827) );
INV_X4 inst_16027 ( .ZN(net_11476), .A(net_10504) );
INV_X4 inst_15322 ( .ZN(net_12262), .A(net_2622) );
NAND2_X2 inst_10458 ( .A1(net_7723), .ZN(net_7022), .A2(net_7021) );
OAI21_X2 inst_1635 ( .ZN(net_19725), .A(net_15665), .B1(net_14460), .B2(net_12580) );
NOR2_X2 inst_4130 ( .A1(net_11681), .A2(net_10644), .ZN(net_6961) );
NAND2_X2 inst_12121 ( .ZN(net_2187), .A2(net_1697), .A1(net_193) );
INV_X4 inst_13102 ( .ZN(net_15825), .A(net_15647) );
INV_X4 inst_17515 ( .A(net_1529), .ZN(net_899) );
OAI21_X4 inst_1500 ( .ZN(net_13888), .B1(net_10089), .B2(net_10072), .A(net_9994) );
INV_X4 inst_14737 ( .A(net_5315), .ZN(net_4107) );
NAND2_X2 inst_11731 ( .A2(net_2950), .ZN(net_2215), .A1(net_2214) );
CLKBUF_X2 inst_22739 ( .A(net_22610), .Z(net_22611) );
NOR2_X4 inst_2805 ( .ZN(net_18075), .A2(net_18066), .A1(net_16044) );
NAND3_X2 inst_6438 ( .ZN(net_20602), .A3(net_9703), .A2(net_6827), .A1(net_5708) );
NOR2_X4 inst_2932 ( .ZN(net_10409), .A2(net_7472), .A1(net_7268) );
INV_X4 inst_17891 ( .ZN(net_166), .A(net_67) );
INV_X4 inst_18329 ( .A(net_20557), .ZN(net_20556) );
NAND2_X4 inst_6917 ( .A2(net_19730), .A1(net_19729), .ZN(net_17818) );
INV_X4 inst_17581 ( .A(net_14308), .ZN(net_14203) );
NAND2_X2 inst_9483 ( .ZN(net_14320), .A1(net_11751), .A2(net_9390) );
INV_X4 inst_15839 ( .ZN(net_1852), .A(net_1851) );
NOR2_X4 inst_3048 ( .ZN(net_8013), .A1(net_5034), .A2(net_952) );
NAND2_X2 inst_10911 ( .A2(net_9309), .ZN(net_5848), .A1(net_3250) );
NOR2_X2 inst_4854 ( .ZN(net_3759), .A2(net_1727), .A1(net_85) );
AOI21_X2 inst_20366 ( .ZN(net_15637), .B1(net_15636), .B2(net_14431), .A(net_11850) );
INV_X2 inst_19276 ( .ZN(net_2984), .A(net_2983) );
INV_X4 inst_13862 ( .ZN(net_12741), .A(net_4823) );
NOR2_X2 inst_3346 ( .ZN(net_18076), .A2(net_18065), .A1(net_16047) );
NOR2_X4 inst_2992 ( .ZN(net_10968), .A2(net_6077), .A1(net_142) );
OR2_X4 inst_1080 ( .ZN(net_9317), .A1(net_7903), .A2(net_5896) );
NAND3_X2 inst_6405 ( .A2(net_12945), .ZN(net_11973), .A3(net_9468), .A1(net_7431) );
OAI211_X4 inst_2374 ( .ZN(net_20434), .B(net_16396), .A(net_15939), .C2(net_13724), .C1(net_1111) );
NAND2_X4 inst_7473 ( .ZN(net_5234), .A2(net_3350), .A1(net_2516) );
INV_X4 inst_15723 ( .A(net_2521), .ZN(net_1966) );
OR2_X4 inst_1103 ( .A2(net_2681), .ZN(net_2466), .A1(net_2299) );
NAND3_X2 inst_6535 ( .ZN(net_10583), .A2(net_10582), .A3(net_5466), .A1(net_3325) );
NAND2_X2 inst_8620 ( .A2(net_16912), .ZN(net_16608), .A1(net_16607) );
AOI21_X4 inst_20212 ( .ZN(net_19117), .B1(net_14493), .A(net_12527), .B2(net_11524) );
INV_X4 inst_17709 ( .ZN(net_612), .A(net_257) );
NAND2_X2 inst_10678 ( .ZN(net_8906), .A1(net_6041), .A2(net_3587) );
NAND2_X2 inst_9256 ( .A1(net_13608), .ZN(net_12645), .A2(net_12644) );
NAND2_X4 inst_7494 ( .A2(net_19229), .ZN(net_4027), .A1(net_2365) );
CLKBUF_X2 inst_22556 ( .A(net_22427), .Z(net_22428) );
XNOR2_X2 inst_549 ( .B(net_17015), .ZN(net_720), .A(net_719) );
NOR2_X2 inst_4329 ( .ZN(net_7425), .A1(net_5785), .A2(net_3561) );
INV_X4 inst_12566 ( .ZN(net_18221), .A(net_18220) );
NOR2_X2 inst_4708 ( .ZN(net_4120), .A2(net_3038), .A1(net_2828) );
AOI21_X4 inst_20186 ( .B1(net_15362), .ZN(net_15219), .B2(net_14108), .A(net_13978) );
INV_X2 inst_18886 ( .ZN(net_6158), .A(net_6157) );
NAND4_X4 inst_5202 ( .A4(net_19481), .A1(net_19480), .ZN(net_16440), .A3(net_16317), .A2(net_13998) );
INV_X4 inst_13617 ( .A(net_8371), .ZN(net_8370) );
CLKBUF_X2 inst_21397 ( .A(net_21247), .Z(net_21269) );
NAND3_X2 inst_6231 ( .ZN(net_13225), .A3(net_12120), .A1(net_7172), .A2(net_6099) );
INV_X2 inst_19084 ( .ZN(net_4579), .A(net_4578) );
INV_X4 inst_16592 ( .ZN(net_6999), .A(net_2585) );
INV_X4 inst_16539 ( .ZN(net_3865), .A(net_107) );
INV_X4 inst_13776 ( .ZN(net_11017), .A(net_7588) );
NAND3_X2 inst_6331 ( .ZN(net_12469), .A1(net_9184), .A3(net_7561), .A2(net_7374) );
INV_X4 inst_16962 ( .ZN(net_9090), .A(net_608) );
NAND2_X2 inst_9737 ( .ZN(net_10104), .A2(net_7670), .A1(net_1964) );
NOR3_X2 inst_2673 ( .ZN(net_14808), .A1(net_13583), .A3(net_12380), .A2(net_9136) );
INV_X4 inst_13592 ( .ZN(net_8807), .A(net_8806) );
OAI21_X2 inst_1618 ( .A(net_20896), .ZN(net_16074), .B2(net_15535), .B1(net_13585) );
NOR2_X2 inst_5062 ( .ZN(net_10162), .A2(net_4329), .A1(net_910) );
INV_X4 inst_14166 ( .ZN(net_9341), .A(net_6009) );
OAI21_X2 inst_2126 ( .A(net_14837), .ZN(net_10007), .B2(net_10006), .B1(net_8047) );
INV_X2 inst_19216 ( .ZN(net_3477), .A(net_3476) );
NAND2_X2 inst_10484 ( .ZN(net_10774), .A1(net_6947), .A2(net_6946) );
INV_X2 inst_18917 ( .ZN(net_5957), .A(net_5956) );
NAND2_X2 inst_7776 ( .ZN(net_18733), .A2(net_18732), .A1(net_17409) );
CLKBUF_X2 inst_22658 ( .A(net_21534), .Z(net_22530) );
AND4_X2 inst_21105 ( .A4(net_12091), .ZN(net_11842), .A3(net_11841), .A2(net_5376), .A1(net_3142) );
INV_X2 inst_19615 ( .A(net_20961), .ZN(net_43) );
NOR3_X2 inst_2765 ( .A3(net_20836), .ZN(net_20150), .A2(net_20077), .A1(net_5018) );
NOR2_X2 inst_3600 ( .ZN(net_20827), .A2(net_9596), .A1(net_6910) );
XNOR2_X2 inst_219 ( .A(net_18211), .ZN(net_17525), .B(net_3581) );
AOI21_X2 inst_20390 ( .ZN(net_20101), .A(net_15742), .B2(net_14525), .B1(net_11306) );
CLKBUF_X2 inst_21380 ( .A(net_21251), .Z(net_21252) );
NOR2_X2 inst_4881 ( .ZN(net_4112), .A1(net_3033), .A2(net_1761) );
INV_X2 inst_19258 ( .A(net_3481), .ZN(net_3193) );
INV_X4 inst_15320 ( .ZN(net_3372), .A(net_2632) );
NAND2_X2 inst_8980 ( .ZN(net_14505), .A1(net_14051), .A2(net_12963) );
NAND4_X2 inst_5501 ( .ZN(net_11825), .A3(net_11824), .A1(net_11247), .A4(net_6749), .A2(net_5770) );
CLKBUF_X2 inst_22932 ( .A(net_22803), .Z(net_22804) );
OAI21_X2 inst_2204 ( .ZN(net_8544), .A(net_8543), .B1(net_8542), .B2(net_8541) );
INV_X4 inst_16785 ( .ZN(net_15463), .A(net_15178) );
INV_X4 inst_16595 ( .ZN(net_1713), .A(net_1254) );
OAI21_X2 inst_1609 ( .A(net_16260), .ZN(net_16144), .B1(net_15749), .B2(net_15234) );
NOR2_X2 inst_4105 ( .ZN(net_14936), .A1(net_7246), .A2(net_6607) );
INV_X4 inst_16530 ( .ZN(net_11376), .A(net_11311) );
INV_X4 inst_16984 ( .A(net_8224), .ZN(net_5701) );
XNOR2_X2 inst_408 ( .A(net_16721), .ZN(net_16625), .B(net_5757) );
NOR2_X2 inst_4701 ( .A1(net_10676), .ZN(net_4139), .A2(net_3171) );
INV_X2 inst_19649 ( .A(net_19464), .ZN(net_19463) );
NAND3_X2 inst_5644 ( .ZN(net_17225), .A3(net_16705), .A2(net_16038), .A1(net_12197) );
INV_X8 inst_12419 ( .A(net_20908), .ZN(net_110) );
NAND2_X2 inst_11212 ( .ZN(net_5808), .A1(net_4194), .A2(net_2297) );
INV_X4 inst_16524 ( .ZN(net_8334), .A(net_1182) );
NAND3_X4 inst_5596 ( .ZN(net_14749), .A3(net_12332), .A2(net_10227), .A1(net_4314) );
CLKBUF_X2 inst_21620 ( .A(net_21445), .Z(net_21492) );
INV_X4 inst_17374 ( .ZN(net_4030), .A(net_3861) );
NAND2_X2 inst_11591 ( .A1(net_3890), .ZN(net_2692), .A2(net_1782) );
NAND2_X2 inst_10719 ( .ZN(net_5885), .A1(net_5884), .A2(net_3504) );
NOR2_X2 inst_3814 ( .ZN(net_9826), .A1(net_6288), .A2(net_5917) );
INV_X4 inst_12968 ( .A(net_16520), .ZN(net_16519) );
NAND2_X2 inst_8498 ( .ZN(net_17077), .A1(net_16613), .A2(net_16475) );
INV_X4 inst_15605 ( .ZN(net_12564), .A(net_2200) );
NAND2_X2 inst_7871 ( .ZN(net_18545), .A2(net_18501), .A1(net_18330) );
NOR2_X2 inst_3514 ( .ZN(net_13821), .A2(net_13820), .A1(net_10167) );
NAND2_X2 inst_10826 ( .ZN(net_13062), .A1(net_8205), .A2(net_5076) );
AOI21_X4 inst_20190 ( .ZN(net_15207), .B2(net_14110), .A(net_12257), .B1(net_197) );
OAI21_X2 inst_1510 ( .ZN(net_18842), .B1(net_18840), .A(net_18808), .B2(net_18807) );
CLKBUF_X2 inst_21392 ( .A(net_21263), .Z(net_21264) );
XNOR2_X2 inst_121 ( .B(net_20378), .A(net_20377), .ZN(net_18402) );
INV_X4 inst_16659 ( .A(net_1789), .ZN(net_1475) );
INV_X8 inst_12449 ( .A(net_20557), .ZN(net_20554) );
OR3_X2 inst_1065 ( .ZN(net_1536), .A1(net_1535), .A3(net_252), .A2(net_112) );
NAND2_X2 inst_12002 ( .ZN(net_1652), .A2(net_1328), .A1(net_225) );
NOR2_X2 inst_4119 ( .ZN(net_8419), .A1(net_6207), .A2(net_4408) );
CLKBUF_X2 inst_22367 ( .A(net_21581), .Z(net_22239) );
CLKBUF_X2 inst_22335 ( .A(net_22206), .Z(net_22207) );
NOR2_X2 inst_4332 ( .ZN(net_10004), .A2(net_8881), .A1(net_6513) );
AOI211_X2 inst_21060 ( .A(net_13246), .ZN(net_10471), .C1(net_10470), .B(net_8795), .C2(net_4722) );
AOI21_X2 inst_20629 ( .ZN(net_13419), .B1(net_13418), .A(net_11675), .B2(net_8936) );
INV_X4 inst_13766 ( .A(net_12612), .ZN(net_10966) );
INV_X4 inst_14348 ( .ZN(net_5325), .A(net_4240) );
NAND2_X2 inst_9495 ( .ZN(net_12596), .A1(net_11430), .A2(net_9439) );
NAND4_X2 inst_5353 ( .ZN(net_15415), .A1(net_14661), .A3(net_14535), .A4(net_13805), .A2(net_11506) );
INV_X4 inst_14189 ( .A(net_9878), .ZN(net_7458) );
NAND2_X2 inst_9981 ( .A1(net_11964), .A2(net_10597), .ZN(net_8862) );
INV_X4 inst_16981 ( .ZN(net_5616), .A(net_1562) );
NOR2_X2 inst_4671 ( .ZN(net_3935), .A2(net_3131), .A1(net_777) );
INV_X4 inst_16860 ( .ZN(net_8376), .A(net_3254) );
XNOR2_X2 inst_530 ( .A(net_21194), .ZN(net_2555), .B(net_2554) );
NAND2_X2 inst_9009 ( .ZN(net_19727), .A2(net_13541), .A1(net_2718) );
NAND2_X2 inst_8004 ( .A1(net_20761), .A2(net_18315), .ZN(net_18305) );
INV_X2 inst_18417 ( .ZN(net_15837), .A(net_15671) );
INV_X2 inst_18994 ( .ZN(net_5080), .A(net_5079) );
OAI21_X4 inst_1353 ( .ZN(net_18426), .A(net_18309), .B2(net_18308), .B1(net_17205) );
NAND2_X4 inst_7370 ( .ZN(net_11766), .A2(net_6131), .A1(net_4280) );
INV_X4 inst_15483 ( .ZN(net_20334), .A(net_2444) );
SDFF_X2 inst_769 ( .Q(net_20906), .SE(net_18837), .SI(net_18469), .D(net_9005), .CK(net_22690) );
INV_X4 inst_13334 ( .ZN(net_12720), .A(net_11132) );
INV_X8 inst_12429 ( .A(net_20878), .ZN(net_525) );
OR2_X2 inst_1200 ( .A2(net_11225), .ZN(net_8500), .A1(net_3988) );
INV_X4 inst_15593 ( .ZN(net_2900), .A(net_1598) );
NAND2_X2 inst_10888 ( .ZN(net_9039), .A1(net_4299), .A2(net_3011) );
NAND2_X2 inst_10120 ( .ZN(net_8381), .A2(net_5227), .A1(net_3453) );
DFF_X1 inst_19820 ( .D(net_17780), .CK(net_22807), .Q(x1192) );
INV_X4 inst_17001 ( .A(net_14945), .ZN(net_869) );
INV_X4 inst_15473 ( .ZN(net_2888), .A(net_2462) );
NAND2_X2 inst_10918 ( .ZN(net_13532), .A2(net_5370), .A1(net_2469) );
NAND2_X2 inst_8523 ( .ZN(net_16905), .A1(net_16821), .A2(net_16654) );
NOR2_X4 inst_3021 ( .ZN(net_6656), .A2(net_4387), .A1(net_529) );
NAND3_X2 inst_6349 ( .A2(net_12932), .ZN(net_12222), .A3(net_12221), .A1(net_7218) );
INV_X4 inst_16037 ( .A(net_2294), .ZN(net_2147) );
NAND2_X4 inst_7365 ( .ZN(net_7309), .A2(net_4401), .A1(net_4400) );
NAND3_X2 inst_6474 ( .ZN(net_11287), .A3(net_9493), .A2(net_7588), .A1(net_2148) );
AOI21_X2 inst_20955 ( .B1(net_8543), .ZN(net_5338), .A(net_4175), .B2(net_2254) );
INV_X8 inst_12232 ( .ZN(net_5934), .A(net_3559) );
NAND2_X2 inst_11664 ( .ZN(net_3742), .A1(net_1049), .A2(net_817) );
INV_X2 inst_19491 ( .A(net_10377), .ZN(net_1306) );
INV_X4 inst_15084 ( .A(net_6400), .ZN(net_3261) );
INV_X2 inst_18794 ( .A(net_8697), .ZN(net_7442) );
INV_X4 inst_12618 ( .A(net_20880), .ZN(net_18070) );
INV_X4 inst_13045 ( .A(net_17767), .ZN(net_16815) );
INV_X2 inst_18628 ( .ZN(net_9544), .A(net_9543) );
CLKBUF_X2 inst_22198 ( .A(net_21375), .Z(net_22070) );
NAND2_X2 inst_11922 ( .A2(net_1778), .ZN(net_1506), .A1(net_1505) );
INV_X4 inst_14790 ( .ZN(net_4592), .A(net_4011) );
CLKBUF_X2 inst_21537 ( .A(net_21408), .Z(net_21409) );
NOR2_X2 inst_3911 ( .ZN(net_8858), .A1(net_7624), .A2(net_6499) );
DFF_X1 inst_19878 ( .D(net_17127), .CK(net_22060), .Q(x368) );
OAI21_X2 inst_1515 ( .ZN(net_18497), .A(net_18440), .B1(net_18439), .B2(net_18438) );
NAND3_X2 inst_6777 ( .ZN(net_4507), .A3(net_2632), .A1(net_1928), .A2(net_749) );
NAND2_X2 inst_9743 ( .ZN(net_10097), .A1(net_10096), .A2(net_7675) );
NAND2_X4 inst_7546 ( .ZN(net_2514), .A1(net_1803), .A2(net_299) );
CLKBUF_X2 inst_22437 ( .A(net_22308), .Z(net_22309) );
INV_X4 inst_13088 ( .ZN(net_15990), .A(net_15878) );
OAI21_X2 inst_1782 ( .A(net_15452), .ZN(net_14662), .B2(net_11937), .B1(net_10212) );
INV_X4 inst_15274 ( .ZN(net_6953), .A(net_3749) );
AOI21_X4 inst_20255 ( .ZN(net_6499), .B1(net_3692), .B2(net_2521), .A(net_735) );
NOR2_X2 inst_4472 ( .ZN(net_4412), .A2(net_4411), .A1(net_3224) );
NAND2_X4 inst_7513 ( .ZN(net_4066), .A1(net_2139), .A2(net_1730) );
SDFF_X2 inst_1015 ( .QN(net_21009), .D(net_533), .SE(net_263), .CK(net_22723), .SI(x2914) );
INV_X4 inst_15776 ( .A(net_9345), .ZN(net_5482) );
NAND2_X4 inst_7003 ( .ZN(net_20067), .A1(net_16711), .A2(net_16558) );
AOI21_X2 inst_20887 ( .ZN(net_7802), .A(net_7801), .B2(net_4162), .B1(net_3469) );
AOI22_X2 inst_19993 ( .B1(net_15205), .ZN(net_14573), .A1(net_14572), .A2(net_12002), .B2(net_6523) );
INV_X4 inst_14390 ( .A(net_14226), .ZN(net_5135) );
NOR2_X2 inst_3899 ( .ZN(net_10669), .A1(net_8361), .A2(net_7365) );
CLKBUF_X2 inst_21912 ( .A(net_21438), .Z(net_21784) );
INV_X4 inst_15940 ( .ZN(net_2130), .A(net_1718) );
INV_X4 inst_14226 ( .ZN(net_7365), .A(net_5834) );
NOR2_X4 inst_3213 ( .ZN(net_5743), .A2(net_3009), .A1(net_2514) );
CLKBUF_X2 inst_21717 ( .A(net_21348), .Z(net_21589) );
AND2_X4 inst_21243 ( .A2(net_3462), .ZN(net_2811), .A1(net_1582) );
INV_X4 inst_17254 ( .ZN(net_1331), .A(net_237) );
INV_X4 inst_15771 ( .ZN(net_4092), .A(net_1820) );
OAI21_X2 inst_1661 ( .B2(net_19793), .B1(net_19792), .ZN(net_19214), .A(net_14179) );
CLKBUF_X2 inst_22246 ( .A(net_21589), .Z(net_22118) );
INV_X4 inst_13583 ( .ZN(net_12875), .A(net_8978) );
XNOR2_X2 inst_283 ( .ZN(net_17165), .A(net_16822), .B(net_16759) );
INV_X4 inst_15193 ( .A(net_4232), .ZN(net_3415) );
OAI211_X2 inst_2519 ( .ZN(net_11887), .B(net_11886), .A(net_6815), .C1(net_5283), .C2(net_2908) );
NOR2_X2 inst_3406 ( .A1(net_19608), .A2(net_15969), .ZN(net_15808) );
OAI21_X2 inst_1597 ( .A(net_20952), .ZN(net_19502), .B2(net_15795), .B1(net_12926) );
NAND2_X4 inst_7574 ( .A1(net_19670), .ZN(net_3065), .A2(net_889) );
CLKBUF_X2 inst_22691 ( .A(net_22562), .Z(net_22563) );
INV_X4 inst_18000 ( .A(net_21096), .ZN(net_389) );
INV_X2 inst_18951 ( .ZN(net_5609), .A(net_4342) );
NAND2_X4 inst_7705 ( .ZN(net_418), .A2(net_137), .A1(net_35) );
XNOR2_X2 inst_431 ( .ZN(net_16480), .A(net_16479), .B(net_16096) );
NAND3_X2 inst_6063 ( .A1(net_20754), .ZN(net_20677), .A3(net_7556), .A2(net_3784) );
NAND2_X2 inst_11331 ( .ZN(net_4698), .A2(net_3730), .A1(net_112) );
CLKBUF_X2 inst_22116 ( .A(net_21987), .Z(net_21988) );
NAND2_X4 inst_6906 ( .ZN(net_17933), .A2(net_17714), .A1(net_17621) );
NAND2_X4 inst_7429 ( .ZN(net_6034), .A1(net_2168), .A2(net_1747) );
AND2_X4 inst_21154 ( .ZN(net_15749), .A2(net_15162), .A1(net_1850) );
INV_X4 inst_15657 ( .ZN(net_3856), .A(net_2091) );
OAI21_X4 inst_1364 ( .ZN(net_17853), .A(net_17604), .B1(net_17603), .B2(net_17602) );
CLKBUF_X2 inst_21712 ( .A(net_21407), .Z(net_21584) );
NAND2_X2 inst_11514 ( .ZN(net_3794), .A2(net_2998), .A1(net_1529) );
INV_X4 inst_18105 ( .A(net_21230), .ZN(net_77) );
INV_X4 inst_14460 ( .ZN(net_8207), .A(net_6829) );
NAND2_X4 inst_6847 ( .ZN(net_18654), .A2(net_18611), .A1(net_18606) );
INV_X4 inst_16417 ( .ZN(net_1255), .A(net_1254) );
CLKBUF_X2 inst_22252 ( .A(net_22055), .Z(net_22124) );
INV_X4 inst_14563 ( .ZN(net_8402), .A(net_4562) );
INV_X2 inst_19730 ( .A(net_20805), .ZN(net_20803) );
INV_X4 inst_14801 ( .ZN(net_7672), .A(net_3983) );
NAND2_X2 inst_11278 ( .ZN(net_6728), .A1(net_3867), .A2(net_3866) );
INV_X2 inst_18366 ( .ZN(net_17867), .A(net_17866) );
NAND2_X2 inst_9560 ( .ZN(net_13610), .A2(net_11535), .A1(net_10031) );
CLKBUF_X2 inst_22032 ( .A(net_21903), .Z(net_21904) );
OAI211_X2 inst_2544 ( .ZN(net_10825), .A(net_9569), .B(net_9090), .C2(net_4631), .C1(net_2633) );
INV_X4 inst_15329 ( .ZN(net_4681), .A(net_2615) );
INV_X2 inst_19118 ( .A(net_14551), .ZN(net_4437) );
INV_X4 inst_16854 ( .ZN(net_4526), .A(net_4158) );
INV_X4 inst_14364 ( .A(net_6914), .ZN(net_6313) );
AOI21_X2 inst_20479 ( .ZN(net_14909), .A(net_14908), .B2(net_13543), .B1(net_4358) );
XNOR2_X1 inst_685 ( .B(net_21143), .ZN(net_17282), .A(net_17162) );
CLKBUF_X2 inst_22302 ( .A(net_22173), .Z(net_22174) );
INV_X4 inst_13281 ( .ZN(net_12438), .A(net_11166) );
CLKBUF_X2 inst_21871 ( .A(net_21742), .Z(net_21743) );
NAND2_X2 inst_9586 ( .A2(net_11764), .ZN(net_10907), .A1(net_9106) );
INV_X4 inst_15478 ( .ZN(net_3609), .A(net_2486) );
INV_X4 inst_15236 ( .ZN(net_2835), .A(net_2834) );
INV_X4 inst_13829 ( .ZN(net_9171), .A(net_8592) );
AND2_X4 inst_21222 ( .ZN(net_8704), .A2(net_5534), .A1(net_5439) );
INV_X4 inst_17485 ( .A(net_2253), .ZN(net_2012) );
NAND2_X2 inst_9150 ( .ZN(net_13400), .A2(net_13399), .A1(net_9080) );
NAND3_X2 inst_6338 ( .ZN(net_12281), .A3(net_12280), .A2(net_12246), .A1(net_6219) );
CLKBUF_X2 inst_21976 ( .A(net_21847), .Z(net_21848) );
NAND2_X4 inst_7693 ( .ZN(net_769), .A2(net_301), .A1(net_282) );
NAND3_X2 inst_6561 ( .ZN(net_10486), .A1(net_8133), .A3(net_7920), .A2(net_7888) );
INV_X4 inst_12700 ( .A(net_17876), .ZN(net_17875) );
INV_X4 inst_12678 ( .ZN(net_17733), .A(net_17732) );
NAND2_X4 inst_6886 ( .ZN(net_18210), .A2(net_18104), .A1(net_18091) );
INV_X2 inst_19562 ( .A(net_14153), .ZN(net_829) );
XNOR2_X2 inst_427 ( .B(net_21139), .ZN(net_16484), .A(net_16482) );
CLKBUF_X2 inst_21886 ( .A(net_21757), .Z(net_21758) );
INV_X2 inst_18592 ( .ZN(net_10149), .A(net_10148) );
AND2_X4 inst_21264 ( .ZN(net_2495), .A2(net_1733), .A1(net_874) );
INV_X4 inst_13113 ( .ZN(net_20628), .A(net_15380) );
NAND2_X2 inst_11952 ( .ZN(net_3013), .A1(net_1433), .A2(net_1136) );
OAI21_X2 inst_2144 ( .ZN(net_9938), .B1(net_9937), .A(net_5544), .B2(net_5161) );
INV_X4 inst_15327 ( .ZN(net_4807), .A(net_2100) );
NAND3_X2 inst_5721 ( .ZN(net_16134), .A1(net_15901), .A3(net_13693), .A2(net_11626) );
NAND3_X2 inst_6121 ( .ZN(net_13853), .A2(net_13852), .A3(net_13851), .A1(net_9533) );
XNOR2_X2 inst_138 ( .B(net_21189), .A(net_20792), .ZN(net_18191) );
NAND3_X2 inst_6793 ( .A1(net_6318), .ZN(net_3885), .A2(net_2996), .A3(net_2497) );
AOI21_X4 inst_20164 ( .ZN(net_19782), .B1(net_14959), .A(net_14572), .B2(net_12213) );
NOR2_X4 inst_2810 ( .ZN(net_17632), .A1(net_17369), .A2(net_17238) );
INV_X4 inst_16969 ( .A(net_6604), .ZN(net_5435) );
SDFF_X2 inst_899 ( .Q(net_21166), .D(net_16772), .SE(net_263), .CK(net_21381), .SI(x5053) );
INV_X8 inst_12304 ( .ZN(net_3276), .A(net_868) );
INV_X4 inst_13346 ( .ZN(net_11069), .A(net_11068) );
INV_X4 inst_13256 ( .ZN(net_12718), .A(net_11660) );
NAND2_X2 inst_9889 ( .ZN(net_19460), .A2(net_9416), .A1(net_8462) );
CLKBUF_X2 inst_22776 ( .A(net_22647), .Z(net_22648) );
AOI21_X2 inst_20916 ( .A(net_10417), .ZN(net_7314), .B2(net_7313), .B1(net_2583) );
OAI21_X2 inst_2149 ( .A(net_10325), .ZN(net_9507), .B2(net_9506), .B1(net_3620) );
NAND2_X2 inst_8356 ( .A2(net_17578), .ZN(net_17461), .A1(net_17460) );
NAND2_X4 inst_6980 ( .ZN(net_17474), .A1(net_16906), .A2(net_16717) );
NOR2_X2 inst_5001 ( .A2(net_3035), .ZN(net_1360), .A1(net_824) );
NAND2_X2 inst_11875 ( .ZN(net_6426), .A2(net_1583), .A1(net_791) );
INV_X4 inst_17003 ( .A(net_12928), .ZN(net_1068) );
INV_X4 inst_14470 ( .A(net_5780), .ZN(net_4906) );
NAND2_X4 inst_7386 ( .ZN(net_10261), .A2(net_6752), .A1(net_4737) );
NAND2_X2 inst_9950 ( .A2(net_11594), .ZN(net_8940), .A1(net_8939) );
AOI21_X2 inst_20401 ( .ZN(net_15390), .B2(net_13972), .A(net_11093), .B1(net_10137) );
NAND2_X2 inst_9319 ( .ZN(net_12340), .A1(net_12339), .A2(net_8977) );
NAND2_X2 inst_8172 ( .ZN(net_17953), .A1(net_17952), .A2(net_17908) );
INV_X4 inst_13899 ( .ZN(net_7164), .A(net_7163) );
AOI211_X2 inst_21046 ( .ZN(net_12871), .B(net_12870), .C1(net_7903), .C2(net_7787), .A(net_7635) );
AOI211_X2 inst_21002 ( .ZN(net_15903), .C1(net_15858), .C2(net_15154), .B(net_14758), .A(net_11372) );
NAND2_X2 inst_8876 ( .ZN(net_20255), .A1(net_15248), .A2(net_14192) );
NOR2_X2 inst_4078 ( .A1(net_8246), .A2(net_7695), .ZN(net_7438) );
DFF_X1 inst_19860 ( .D(net_17256), .CK(net_22802), .Q(x1021) );
NOR2_X2 inst_4067 ( .ZN(net_7726), .A1(net_7725), .A2(net_4514) );
CLKBUF_X2 inst_22906 ( .A(net_22777), .Z(net_22778) );
INV_X2 inst_18846 ( .A(net_8571), .ZN(net_6657) );
NAND2_X2 inst_9109 ( .ZN(net_13601), .A2(net_13600), .A1(net_5068) );
NAND2_X2 inst_8894 ( .ZN(net_15111), .A1(net_15110), .A2(net_13957) );
NAND2_X2 inst_10175 ( .ZN(net_8203), .A1(net_8202), .A2(net_8201) );
INV_X4 inst_14972 ( .A(net_4503), .ZN(net_3423) );
INV_X4 inst_14180 ( .ZN(net_7834), .A(net_7832) );
NAND2_X2 inst_8885 ( .ZN(net_15148), .A2(net_14100), .A1(net_7300) );
NOR2_X2 inst_3883 ( .A1(net_11218), .ZN(net_9311), .A2(net_7846) );
NAND2_X2 inst_10020 ( .A1(net_10575), .ZN(net_8766), .A2(net_8027) );
INV_X2 inst_19632 ( .A(net_20889), .ZN(net_989) );
NAND2_X2 inst_11811 ( .ZN(net_1849), .A1(net_1848), .A2(net_1847) );
INV_X4 inst_13451 ( .ZN(net_12941), .A(net_9732) );
CLKBUF_X2 inst_21442 ( .A(net_21304), .Z(net_21314) );
NAND2_X2 inst_9096 ( .ZN(net_13783), .A1(net_13538), .A2(net_12469) );
NAND3_X2 inst_5818 ( .ZN(net_15596), .A2(net_15595), .A3(net_14268), .A1(net_13754) );
INV_X2 inst_19644 ( .ZN(net_19440), .A(net_2479) );
AOI21_X4 inst_20141 ( .ZN(net_19841), .B1(net_19758), .B2(net_15917), .A(net_13145) );
NAND4_X2 inst_5510 ( .A4(net_20403), .A1(net_20402), .ZN(net_11059), .A2(net_6693), .A3(net_5495) );
NAND2_X4 inst_7041 ( .ZN(net_16435), .A2(net_16406), .A1(net_16360) );
NAND2_X2 inst_8415 ( .ZN(net_17228), .A2(net_17227), .A1(net_13950) );
CLKBUF_X2 inst_22630 ( .A(net_21694), .Z(net_22502) );
INV_X4 inst_12632 ( .ZN(net_17970), .A(net_17921) );
NAND2_X2 inst_10308 ( .ZN(net_12056), .A1(net_7858), .A2(net_5981) );
OAI211_X2 inst_2577 ( .ZN(net_8479), .A(net_8478), .B(net_8377), .C1(net_3262), .C2(net_1325) );
INV_X4 inst_15319 ( .ZN(net_4930), .A(net_3850) );
NAND2_X4 inst_7565 ( .ZN(net_2068), .A2(net_1669), .A1(net_61) );
INV_X4 inst_16571 ( .ZN(net_10937), .A(net_9754) );
INV_X4 inst_17886 ( .A(net_386), .ZN(net_73) );
INV_X4 inst_13267 ( .ZN(net_12597), .A(net_12596) );
NAND3_X2 inst_6431 ( .ZN(net_11904), .A3(net_10351), .A1(net_7049), .A2(net_5659) );
INV_X4 inst_16759 ( .ZN(net_1761), .A(net_276) );
NAND2_X4 inst_7131 ( .ZN(net_20132), .A1(net_11941), .A2(net_4756) );
NOR2_X2 inst_3804 ( .ZN(net_9846), .A2(net_9845), .A1(net_5224) );
INV_X2 inst_19541 ( .ZN(net_1595), .A(net_1175) );
AOI21_X2 inst_20420 ( .ZN(net_15223), .B1(net_14981), .A(net_14437), .B2(net_14116) );
OAI21_X2 inst_2266 ( .ZN(net_20319), .B2(net_4341), .B1(net_3863), .A(net_86) );
INV_X4 inst_17741 ( .A(net_177), .ZN(net_176) );
INV_X4 inst_14331 ( .A(net_11718), .ZN(net_5416) );
NAND2_X4 inst_7148 ( .ZN(net_11068), .A2(net_9779), .A1(net_8709) );
INV_X4 inst_13206 ( .ZN(net_13822), .A(net_13131) );
INV_X4 inst_16250 ( .ZN(net_7865), .A(net_1358) );
INV_X4 inst_13440 ( .ZN(net_9809), .A(net_9808) );
AND2_X4 inst_21207 ( .ZN(net_7285), .A1(net_7284), .A2(net_5293) );
INV_X4 inst_15962 ( .ZN(net_2476), .A(net_817) );
NAND2_X2 inst_8744 ( .ZN(net_15988), .A2(net_15652), .A1(net_333) );
NAND2_X2 inst_12023 ( .A1(net_20946), .ZN(net_9289), .A2(net_154) );
INV_X4 inst_16814 ( .ZN(net_20065), .A(net_803) );
INV_X4 inst_13437 ( .ZN(net_11134), .A(net_8373) );
OAI211_X2 inst_2514 ( .ZN(net_12230), .B(net_12229), .A(net_11861), .C2(net_7545), .C1(net_5735) );
INV_X2 inst_19301 ( .ZN(net_2775), .A(net_2774) );
NAND2_X2 inst_7869 ( .ZN(net_18547), .A1(net_18474), .A2(net_17740) );
OR2_X4 inst_1128 ( .ZN(net_1980), .A2(net_168), .A1(net_52) );
NAND2_X2 inst_8009 ( .ZN(net_18298), .A2(net_18295), .A1(net_17745) );
NOR2_X4 inst_3222 ( .ZN(net_5351), .A1(net_3096), .A2(net_1848) );
NOR2_X2 inst_3759 ( .ZN(net_10357), .A1(net_9804), .A2(net_9414) );
CLKBUF_X2 inst_22429 ( .A(net_22300), .Z(net_22301) );
NAND2_X2 inst_10928 ( .ZN(net_6342), .A1(net_5220), .A2(net_3983) );
NAND2_X4 inst_7422 ( .ZN(net_4608), .A1(net_3513), .A2(net_2001) );
INV_X2 inst_19042 ( .ZN(net_4766), .A(net_4765) );
CLKBUF_X2 inst_21808 ( .A(net_21679), .Z(net_21680) );
INV_X2 inst_19344 ( .ZN(net_2438), .A(net_1546) );
CLKBUF_X2 inst_22221 ( .A(net_22092), .Z(net_22093) );
NOR2_X2 inst_4070 ( .A1(net_13848), .ZN(net_10648), .A2(net_4648) );
OAI21_X2 inst_1924 ( .ZN(net_13021), .B2(net_11487), .B1(net_5213), .A(net_1663) );
CLKBUF_X2 inst_21449 ( .A(net_21320), .Z(net_21321) );
NAND2_X2 inst_10502 ( .A1(net_11442), .ZN(net_8885), .A2(net_6919) );
INV_X2 inst_18452 ( .ZN(net_14197), .A(net_13571) );
NOR2_X2 inst_4748 ( .ZN(net_9897), .A1(net_3027), .A2(net_1565) );
AOI21_X2 inst_20538 ( .ZN(net_19245), .B1(net_13812), .A(net_10252), .B2(net_10223) );
NOR2_X2 inst_4160 ( .ZN(net_8824), .A2(net_5505), .A1(net_731) );
NAND3_X2 inst_5685 ( .A1(net_20448), .ZN(net_16301), .A3(net_15595), .A2(net_15546) );
SDFF_X2 inst_961 ( .QN(net_21033), .SE(net_2426), .D(net_463), .CK(net_22731), .SI(x2428) );
NOR2_X4 inst_3255 ( .A2(net_20478), .ZN(net_3263), .A1(net_1424) );
INV_X4 inst_13119 ( .ZN(net_15497), .A(net_15221) );
NAND2_X2 inst_11082 ( .A1(net_5818), .ZN(net_4446), .A2(net_3257) );
INV_X4 inst_12800 ( .ZN(net_17382), .A(net_17250) );
NAND2_X2 inst_8077 ( .A1(net_21187), .ZN(net_18154), .A2(net_18153) );
CLKBUF_X2 inst_22442 ( .A(net_21729), .Z(net_22314) );
NAND2_X2 inst_8332 ( .ZN(net_19189), .A2(net_17515), .A1(net_15957) );
NOR2_X2 inst_5103 ( .ZN(net_5259), .A1(net_765), .A2(net_493) );
CLKBUF_X2 inst_21849 ( .A(net_21290), .Z(net_21721) );
NAND2_X2 inst_11364 ( .A1(net_3715), .ZN(net_3599), .A2(net_3525) );
INV_X4 inst_16734 ( .ZN(net_1756), .A(net_1049) );
NAND2_X2 inst_8489 ( .A1(net_21156), .ZN(net_16958), .A2(net_16635) );
OAI21_X2 inst_2316 ( .ZN(net_5695), .A(net_5694), .B2(net_5485), .B1(net_1483) );
NOR3_X2 inst_2737 ( .ZN(net_12778), .A3(net_12777), .A2(net_10862), .A1(net_6741) );
NAND3_X2 inst_6654 ( .ZN(net_8509), .A2(net_8508), .A3(net_8507), .A1(net_4906) );
INV_X4 inst_14266 ( .ZN(net_5722), .A(net_4892) );
XNOR2_X2 inst_499 ( .A(net_17366), .ZN(net_9001), .B(net_1843) );
NAND3_X2 inst_6175 ( .ZN(net_13548), .A3(net_12505), .A1(net_12273), .A2(net_8333) );
NAND2_X2 inst_9468 ( .A1(net_13781), .ZN(net_13691), .A2(net_11481) );
OAI211_X2 inst_2400 ( .ZN(net_15956), .C1(net_15955), .B(net_15256), .A(net_11986), .C2(net_11325) );
AND2_X4 inst_21187 ( .ZN(net_11000), .A1(net_10999), .A2(net_10998) );
INV_X2 inst_18535 ( .A(net_12861), .ZN(net_11072) );
OAI21_X4 inst_1451 ( .B2(net_20010), .B1(net_20009), .ZN(net_15447), .A(net_14694) );
CLKBUF_X2 inst_21647 ( .A(net_21518), .Z(net_21519) );
NOR2_X2 inst_4082 ( .ZN(net_20237), .A1(net_7317), .A2(net_6615) );
NOR2_X2 inst_4781 ( .ZN(net_20225), .A2(net_2883), .A1(net_1224) );
INV_X4 inst_14207 ( .ZN(net_9574), .A(net_4866) );
INV_X4 inst_17779 ( .ZN(net_1961), .A(net_271) );
OAI21_X2 inst_2009 ( .ZN(net_11390), .A(net_11389), .B2(net_11388), .B1(net_2776) );
XNOR2_X2 inst_501 ( .ZN(net_8999), .A(net_6459), .B(net_2041) );
CLKBUF_X2 inst_22508 ( .A(net_22379), .Z(net_22380) );
OAI21_X2 inst_2093 ( .ZN(net_10154), .A(net_5716), .B2(net_5685), .B1(net_1069) );
OR2_X4 inst_1081 ( .A1(net_11050), .ZN(net_9314), .A2(net_5895) );
NOR2_X4 inst_3195 ( .ZN(net_3360), .A2(net_2399), .A1(net_955) );
NAND2_X2 inst_8873 ( .ZN(net_15259), .A2(net_14670), .A1(net_10066) );
NAND2_X2 inst_10731 ( .ZN(net_5807), .A2(net_4390), .A1(net_433) );
INV_X4 inst_17984 ( .A(net_21052), .ZN(net_736) );
INV_X4 inst_15888 ( .ZN(net_6861), .A(net_1298) );
INV_X4 inst_15828 ( .A(net_15677), .ZN(net_2547) );
NOR2_X4 inst_2905 ( .ZN(net_19106), .A1(net_7643), .A2(net_4225) );
INV_X2 inst_19222 ( .A(net_9929), .ZN(net_3444) );
NOR2_X4 inst_2819 ( .ZN(net_16506), .A1(net_16245), .A2(net_16220) );
CLKBUF_X2 inst_22040 ( .A(net_21911), .Z(net_21912) );
INV_X8 inst_12263 ( .ZN(net_2791), .A(net_1635) );
AOI21_X4 inst_20238 ( .ZN(net_11203), .B2(net_9509), .A(net_4426), .B1(net_2363) );
NAND3_X2 inst_6293 ( .ZN(net_12821), .A3(net_10933), .A2(net_10883), .A1(net_8116) );
INV_X4 inst_15016 ( .A(net_14315), .ZN(net_4447) );
DFF_X2 inst_19774 ( .QN(net_21219), .D(net_17264), .CK(net_22338) );
INV_X4 inst_17416 ( .ZN(net_5517), .A(net_5239) );
CLKBUF_X2 inst_21567 ( .A(net_21438), .Z(net_21439) );
NAND2_X2 inst_9963 ( .ZN(net_19721), .A2(net_8209), .A1(net_4733) );
AOI21_X2 inst_20270 ( .B1(net_18908), .ZN(net_16396), .B2(net_16395), .A(net_16253) );
OR2_X4 inst_1114 ( .ZN(net_4799), .A2(net_874), .A1(net_120) );
NAND2_X2 inst_7982 ( .ZN(net_18336), .A2(net_18335), .A1(net_17995) );
CLKBUF_X2 inst_22706 ( .A(net_22577), .Z(net_22578) );
NAND2_X2 inst_9327 ( .ZN(net_13558), .A1(net_12306), .A2(net_7475) );
NOR2_X2 inst_4163 ( .ZN(net_14996), .A1(net_12070), .A2(net_6518) );
INV_X4 inst_15391 ( .ZN(net_14166), .A(net_6513) );
NAND2_X2 inst_9020 ( .ZN(net_20674), .A1(net_14171), .A2(net_12235) );
AOI21_X1 inst_20987 ( .ZN(net_6438), .A(net_6437), .B1(net_2599), .B2(net_2192) );
INV_X4 inst_17244 ( .ZN(net_1044), .A(net_657) );
INV_X4 inst_17021 ( .ZN(net_8097), .A(net_986) );
OAI21_X2 inst_1982 ( .ZN(net_12111), .B2(net_8009), .A(net_6586), .B1(net_3787) );
AOI21_X2 inst_20656 ( .B1(net_14086), .ZN(net_13036), .A(net_12662), .B2(net_9308) );
INV_X4 inst_16246 ( .ZN(net_1361), .A(net_81) );
INV_X4 inst_15909 ( .ZN(net_1762), .A(net_1761) );
NAND2_X2 inst_11805 ( .A2(net_2235), .ZN(net_1904), .A1(net_1903) );
OAI21_X2 inst_1849 ( .ZN(net_14010), .A(net_14009), .B2(net_11301), .B1(net_11146) );
CLKBUF_X2 inst_22683 ( .A(net_22447), .Z(net_22555) );
INV_X2 inst_18378 ( .ZN(net_16949), .A(net_16948) );
NAND3_X4 inst_5540 ( .A3(net_19297), .A1(net_19296), .ZN(net_17312), .A2(net_13790) );
CLKBUF_X2 inst_22265 ( .A(net_22136), .Z(net_22137) );
NAND2_X2 inst_11123 ( .A1(net_20859), .ZN(net_10246), .A2(net_4289) );
OAI21_X2 inst_1976 ( .A(net_20889), .ZN(net_19304), .B1(net_11151), .B2(net_8253) );
NOR2_X2 inst_4932 ( .ZN(net_10379), .A1(net_7153), .A2(net_76) );
NOR3_X2 inst_2744 ( .ZN(net_12580), .A1(net_11365), .A3(net_11054), .A2(net_8541) );
NOR2_X2 inst_3681 ( .ZN(net_11424), .A2(net_10954), .A1(net_6600) );
NAND2_X4 inst_6909 ( .A2(net_19687), .A1(net_19686), .ZN(net_17858) );
AOI21_X2 inst_20982 ( .B2(net_20581), .B1(net_7878), .ZN(net_2947), .A(net_1079) );
INV_X4 inst_13238 ( .ZN(net_14813), .A(net_13439) );
NAND4_X2 inst_5277 ( .ZN(net_19102), .A2(net_19029), .A1(net_19028), .A4(net_14613), .A3(net_6802) );
OAI211_X2 inst_2384 ( .C2(net_20888), .C1(net_18954), .ZN(net_16708), .B(net_16172), .A(net_10368) );
NOR2_X2 inst_4614 ( .ZN(net_6349), .A2(net_2043), .A1(net_809) );
INV_X1 inst_19753 ( .A(net_10922), .ZN(net_9160) );
NAND2_X2 inst_9606 ( .ZN(net_10731), .A1(net_10730), .A2(net_8806) );
OR2_X2 inst_1212 ( .ZN(net_7082), .A2(net_3294), .A1(net_1660) );
XNOR2_X2 inst_670 ( .B(net_21188), .A(net_21124), .ZN(net_158) );
INV_X4 inst_17561 ( .ZN(net_5244), .A(net_365) );
CLKBUF_X2 inst_22764 ( .A(net_22635), .Z(net_22636) );
NOR2_X2 inst_4180 ( .A1(net_8874), .ZN(net_8104), .A2(net_4046) );
NAND3_X2 inst_5789 ( .ZN(net_15772), .A3(net_15130), .A2(net_13991), .A1(net_12703) );
NAND2_X2 inst_11105 ( .ZN(net_10620), .A2(net_6854), .A1(net_4330) );
NAND2_X2 inst_9612 ( .A1(net_10930), .ZN(net_10713), .A2(net_8487) );
NOR2_X2 inst_3901 ( .A1(net_10920), .A2(net_10834), .ZN(net_9092) );
INV_X2 inst_18425 ( .ZN(net_19977), .A(net_14690) );
INV_X2 inst_19071 ( .ZN(net_4628), .A(net_3333) );
INV_X4 inst_16901 ( .A(net_4183), .ZN(net_3760) );
INV_X4 inst_17979 ( .A(net_20920), .ZN(net_16259) );
NAND3_X2 inst_6679 ( .ZN(net_7742), .A2(net_6237), .A3(net_5142), .A1(net_2656) );
INV_X2 inst_19294 ( .ZN(net_5644), .A(net_3963) );
INV_X4 inst_15200 ( .A(net_3903), .ZN(net_3499) );
INV_X4 inst_14093 ( .ZN(net_12287), .A(net_6197) );
AOI222_X2 inst_20062 ( .ZN(net_14757), .C1(net_13700), .B1(net_11446), .C2(net_10853), .A2(net_10622), .B2(net_6470), .A1(net_2368) );
NAND3_X2 inst_5898 ( .ZN(net_15176), .A1(net_14565), .A2(net_10306), .A3(net_8942) );
CLKBUF_X2 inst_21416 ( .A(net_21287), .Z(net_21288) );
NAND2_X2 inst_8647 ( .A1(net_16718), .ZN(net_16566), .A2(net_16408) );
NAND2_X2 inst_10845 ( .ZN(net_5470), .A2(net_5469), .A1(net_3022) );
NAND2_X2 inst_9814 ( .A1(net_12958), .ZN(net_9664), .A2(net_9663) );
INV_X4 inst_14502 ( .ZN(net_5996), .A(net_4835) );
SDFF_X2 inst_807 ( .Q(net_20913), .SE(net_18862), .SI(net_17942), .D(net_740), .CK(net_21259) );
SDFF_X2 inst_705 ( .Q(net_20862), .SI(net_18834), .SE(net_18804), .D(net_645), .CK(net_22032) );
INV_X2 inst_18433 ( .ZN(net_19570), .A(net_14123) );
SDFF_X2 inst_911 ( .Q(net_21224), .SI(net_16682), .SE(net_125), .CK(net_21523), .D(x7235) );
AOI21_X2 inst_20863 ( .A(net_14463), .ZN(net_8750), .B2(net_4739), .B1(net_2838) );
NAND2_X2 inst_10921 ( .ZN(net_12447), .A1(net_7473), .A2(net_5291) );
AOI211_X2 inst_21012 ( .ZN(net_15685), .C1(net_15684), .C2(net_14930), .B(net_13407), .A(net_10100) );
INV_X4 inst_15746 ( .ZN(net_11441), .A(net_10875) );
SDFF_X2 inst_1003 ( .QN(net_21059), .D(net_626), .SE(net_263), .CK(net_21717), .SI(x2077) );
INV_X4 inst_14893 ( .ZN(net_6311), .A(net_5215) );
INV_X4 inst_13804 ( .ZN(net_12516), .A(net_7549) );
AOI21_X2 inst_20526 ( .ZN(net_14555), .B1(net_14554), .B2(net_11928), .A(net_5128) );
AOI21_X2 inst_20830 ( .ZN(net_9859), .B1(net_9450), .B2(net_7921), .A(net_2000) );
CLKBUF_X2 inst_22420 ( .A(net_21733), .Z(net_22292) );
INV_X4 inst_14889 ( .ZN(net_6336), .A(net_3661) );
NAND2_X2 inst_10284 ( .ZN(net_11727), .A1(net_9966), .A2(net_6178) );
NOR2_X2 inst_3469 ( .ZN(net_14510), .A1(net_14509), .A2(net_12848) );
NAND3_X2 inst_6026 ( .ZN(net_14372), .A1(net_12982), .A2(net_11037), .A3(net_10055) );
NAND4_X2 inst_5456 ( .A4(net_19748), .A1(net_19747), .ZN(net_13450), .A2(net_12031), .A3(net_9840) );
CLKBUF_X2 inst_21796 ( .A(net_21667), .Z(net_21668) );
OAI21_X2 inst_2080 ( .ZN(net_10518), .B1(net_8748), .A(net_7913), .B2(net_5326) );
OAI21_X2 inst_1625 ( .ZN(net_16044), .B1(net_15747), .B2(net_15475), .A(net_15394) );
NAND2_X2 inst_7710 ( .ZN(net_18855), .A2(net_18851), .A1(net_17039) );
CLKBUF_X2 inst_22158 ( .A(net_22029), .Z(net_22030) );
XNOR2_X2 inst_593 ( .ZN(net_559), .A(net_558), .B(net_557) );
NAND3_X2 inst_5707 ( .ZN(net_16201), .A1(net_16007), .A3(net_14838), .A2(net_10293) );
INV_X2 inst_18920 ( .ZN(net_5931), .A(net_5930) );
INV_X4 inst_15664 ( .A(net_3084), .ZN(net_2852) );
OAI21_X2 inst_2223 ( .ZN(net_8506), .A(net_8505), .B2(net_8504), .B1(net_1688) );
NOR2_X2 inst_4522 ( .ZN(net_19873), .A1(net_11681), .A2(net_11257) );
NAND3_X2 inst_6137 ( .ZN(net_19306), .A1(net_13012), .A2(net_6643), .A3(net_4445) );
INV_X8 inst_12426 ( .A(net_20926), .ZN(net_322) );
NAND2_X2 inst_10099 ( .ZN(net_19132), .A2(net_10506), .A1(net_8611) );
NAND3_X2 inst_5738 ( .ZN(net_19993), .A2(net_15498), .A3(net_15168), .A1(net_8319) );
NAND2_X2 inst_7845 ( .A1(net_20062), .ZN(net_18611), .A2(net_16425) );
NAND2_X2 inst_9065 ( .ZN(net_13988), .A2(net_11960), .A1(net_60) );
NAND2_X2 inst_10045 ( .ZN(net_13238), .A1(net_8709), .A2(net_8708) );
XNOR2_X2 inst_479 ( .A(net_16659), .ZN(net_11871), .B(net_1859) );
INV_X2 inst_19383 ( .ZN(net_3730), .A(net_3182) );
NAND2_X2 inst_10448 ( .ZN(net_7100), .A1(net_7099), .A2(net_4937) );
CLKBUF_X2 inst_22376 ( .A(net_22247), .Z(net_22248) );
INV_X4 inst_17271 ( .A(net_14483), .ZN(net_14033) );
OAI21_X2 inst_2344 ( .A(net_12564), .ZN(net_4379), .B2(net_4378), .B1(net_2307) );
NOR2_X4 inst_3326 ( .ZN(net_813), .A1(net_288), .A2(net_49) );
NAND2_X4 inst_7288 ( .ZN(net_19333), .A1(net_3424), .A2(net_3297) );
NAND2_X4 inst_7683 ( .ZN(net_1311), .A1(net_1270), .A2(net_930) );
INV_X4 inst_12892 ( .A(net_17019), .ZN(net_17011) );
NOR2_X2 inst_4387 ( .ZN(net_12890), .A1(net_7903), .A2(net_3168) );
NAND2_X2 inst_9420 ( .ZN(net_11634), .A2(net_11632), .A1(net_6978) );
INV_X1 inst_19749 ( .ZN(net_12389), .A(net_12388) );
INV_X4 inst_15068 ( .ZN(net_4368), .A(net_3286) );
NAND2_X4 inst_7113 ( .ZN(net_12705), .A1(net_11135), .A2(net_6091) );
AOI21_X2 inst_20264 ( .ZN(net_18068), .B2(net_18067), .B1(net_16014), .A(net_14855) );
NAND3_X2 inst_5780 ( .ZN(net_15823), .A1(net_15319), .A2(net_10790), .A3(net_10747) );
INV_X4 inst_16485 ( .A(net_10074), .ZN(net_1202) );
INV_X2 inst_19639 ( .A(net_19430), .ZN(net_19429) );
NAND2_X2 inst_10523 ( .ZN(net_6850), .A2(net_6849), .A1(net_6848) );
INV_X4 inst_17320 ( .A(net_935), .ZN(net_781) );
NOR2_X2 inst_4497 ( .ZN(net_19083), .A2(net_11962), .A1(net_11087) );
NOR3_X2 inst_2651 ( .A3(net_19382), .A1(net_19381), .ZN(net_15479), .A2(net_12660) );
NOR2_X2 inst_4756 ( .ZN(net_5071), .A2(net_1573), .A1(net_1228) );
NOR2_X2 inst_4201 ( .ZN(net_6685), .A2(net_6684), .A1(net_6443) );
NAND3_X2 inst_5658 ( .ZN(net_16429), .A3(net_16285), .A1(net_13414), .A2(net_12753) );
XOR2_X2 inst_48 ( .A(net_18141), .Z(net_444), .B(net_443) );
AOI21_X2 inst_20742 ( .A(net_20889), .B1(net_19196), .ZN(net_11417), .B2(net_9291) );
AOI21_X2 inst_20877 ( .ZN(net_8456), .B1(net_8455), .B2(net_6700), .A(net_3220) );
INV_X4 inst_16008 ( .ZN(net_5799), .A(net_1091) );
INV_X2 inst_19468 ( .A(net_6415), .ZN(net_1450) );
OAI21_X2 inst_2246 ( .A(net_10714), .ZN(net_7328), .B2(net_6920), .B1(net_2203) );
NAND2_X4 inst_7507 ( .ZN(net_7700), .A1(net_3026), .A2(net_1082) );
CLKBUF_X2 inst_22150 ( .A(net_22021), .Z(net_22022) );
XNOR2_X2 inst_443 ( .B(net_21112), .ZN(net_15589), .A(net_15588) );
INV_X4 inst_17114 ( .ZN(net_7394), .A(net_6314) );
INV_X2 inst_19633 ( .A(net_19418), .ZN(net_19417) );
NAND2_X2 inst_11022 ( .ZN(net_11276), .A1(net_8616), .A2(net_4708) );
NAND2_X2 inst_8766 ( .A1(net_15880), .ZN(net_15878), .A2(net_15422) );
NOR2_X2 inst_4259 ( .A1(net_6840), .ZN(net_6263), .A2(net_3179) );
CLKBUF_X2 inst_21744 ( .A(net_21615), .Z(net_21616) );
AOI21_X2 inst_20967 ( .ZN(net_5273), .B2(net_5272), .B1(net_4581), .A(net_4429) );
NAND2_X1 inst_12152 ( .ZN(net_10222), .A2(net_9723), .A1(net_6030) );
NAND2_X2 inst_9060 ( .ZN(net_13993), .A1(net_13091), .A2(net_11996) );
OAI21_X2 inst_1700 ( .ZN(net_15316), .A(net_14643), .B2(net_13611), .B1(net_7719) );
INV_X2 inst_19424 ( .A(net_15731), .ZN(net_1822) );
INV_X4 inst_15814 ( .ZN(net_2723), .A(net_1555) );
OAI211_X2 inst_2571 ( .C1(net_20531), .ZN(net_9016), .B(net_8976), .A(net_6307), .C2(net_1672) );
INV_X4 inst_12481 ( .ZN(net_18741), .A(net_18713) );
SDFF_X2 inst_730 ( .Q(net_20910), .SE(net_18858), .SI(net_18565), .D(net_3435), .CK(net_21916) );
NAND2_X2 inst_11430 ( .ZN(net_7985), .A2(net_3344), .A1(net_809) );
CLKBUF_X2 inst_22406 ( .A(net_22277), .Z(net_22278) );
NAND2_X2 inst_10116 ( .ZN(net_8400), .A1(net_8399), .A2(net_8398) );
NAND3_X2 inst_6754 ( .ZN(net_5711), .A3(net_5465), .A2(net_2996), .A1(net_112) );
XNOR2_X2 inst_321 ( .A(net_20212), .ZN(net_17163), .B(net_17036) );
INV_X16 inst_19745 ( .A(net_20568), .ZN(net_20567) );
INV_X2 inst_18831 ( .ZN(net_6775), .A(net_6774) );
NAND2_X2 inst_10977 ( .ZN(net_10010), .A2(net_4967), .A1(net_2420) );
CLKBUF_X2 inst_21754 ( .A(net_21329), .Z(net_21626) );
INV_X4 inst_18085 ( .A(net_20854), .ZN(net_128) );
AND2_X4 inst_21204 ( .ZN(net_7946), .A2(net_5643), .A1(net_5003) );
NOR2_X4 inst_3131 ( .ZN(net_7031), .A1(net_3847), .A2(net_3107) );
INV_X4 inst_12684 ( .ZN(net_17721), .A(net_17720) );
INV_X4 inst_14788 ( .ZN(net_8442), .A(net_4012) );
INV_X4 inst_13308 ( .ZN(net_11716), .A(net_10430) );
AOI21_X2 inst_20411 ( .B1(net_19565), .ZN(net_19280), .B2(net_11439), .A(net_9232) );
DFF_X1 inst_19881 ( .D(net_17135), .CK(net_21323), .Q(x233) );
NAND2_X2 inst_8264 ( .A1(net_21130), .ZN(net_19665), .A2(net_17455) );
INV_X4 inst_16049 ( .ZN(net_2189), .A(net_1090) );
CLKBUF_X2 inst_22849 ( .A(net_22720), .Z(net_22721) );
INV_X4 inst_16834 ( .ZN(net_1429), .A(net_985) );
OR2_X2 inst_1152 ( .ZN(net_9760), .A2(net_9759), .A1(net_8629) );
NAND2_X4 inst_6878 ( .ZN(net_18190), .A2(net_18119), .A1(net_16778) );
INV_X4 inst_15255 ( .ZN(net_5706), .A(net_4439) );
INV_X2 inst_19722 ( .A(net_20786), .ZN(net_20785) );
NAND3_X2 inst_6517 ( .A3(net_12011), .ZN(net_10651), .A1(net_6275), .A2(net_6170) );
INV_X2 inst_18582 ( .ZN(net_10304), .A(net_10303) );
NAND3_X1 inst_6823 ( .A2(net_13762), .ZN(net_9062), .A3(net_9061), .A1(net_5808) );
DFF_X1 inst_19896 ( .D(net_16940), .CK(net_22352), .Q(x912) );
NAND2_X2 inst_8670 ( .ZN(net_16468), .A2(net_16467), .A1(net_16422) );
XNOR2_X2 inst_182 ( .ZN(net_17766), .A(net_17334), .B(net_16701) );
CLKBUF_X2 inst_22282 ( .A(net_22153), .Z(net_22154) );
SDFF_X2 inst_931 ( .QN(net_20981), .D(net_2515), .SE(net_263), .CK(net_21859), .SI(x3311) );
NAND2_X2 inst_9205 ( .ZN(net_13063), .A1(net_13062), .A2(net_11256) );
NOR2_X4 inst_3174 ( .ZN(net_3145), .A1(net_1848), .A2(net_1549) );
OAI21_X2 inst_1674 ( .ZN(net_15547), .A(net_15248), .B2(net_14623), .B1(net_8610) );
NOR2_X2 inst_3824 ( .ZN(net_9775), .A2(net_9774), .A1(net_3996) );
NAND2_X4 inst_6895 ( .A2(net_20880), .ZN(net_18047), .A1(net_16008) );
INV_X4 inst_12807 ( .ZN(net_17321), .A(net_17212) );
NAND2_X2 inst_8438 ( .ZN(net_17272), .A1(net_16825), .A2(net_16671) );
INV_X4 inst_15983 ( .ZN(net_1899), .A(net_1400) );
NAND2_X2 inst_8315 ( .ZN(net_17575), .A2(net_17352), .A1(net_17229) );
AOI21_X2 inst_20762 ( .B1(net_11927), .ZN(net_10892), .A(net_10891), .B2(net_2931) );
INV_X4 inst_16226 ( .ZN(net_1870), .A(net_1380) );
NOR2_X2 inst_4089 ( .A1(net_15270), .A2(net_10465), .ZN(net_8783) );
INV_X4 inst_15929 ( .ZN(net_10920), .A(net_8328) );
INV_X4 inst_14320 ( .ZN(net_9878), .A(net_6572) );
OAI21_X4 inst_1415 ( .A(net_20904), .B2(net_18959), .B1(net_18958), .ZN(net_16150) );
AOI21_X2 inst_20741 ( .B1(net_19527), .ZN(net_11420), .B2(net_6474), .A(net_79) );
NAND2_X2 inst_12089 ( .ZN(net_830), .A2(net_312), .A1(net_71) );
INV_X4 inst_13631 ( .ZN(net_8275), .A(net_8274) );
NOR2_X4 inst_3301 ( .ZN(net_1781), .A1(net_1192), .A2(net_282) );
NAND3_X2 inst_5997 ( .ZN(net_14436), .A1(net_12761), .A3(net_11222), .A2(net_5447) );
NAND3_X2 inst_6469 ( .A2(net_11629), .ZN(net_11339), .A1(net_11338), .A3(net_11224) );
CLKBUF_X2 inst_21955 ( .A(net_21826), .Z(net_21827) );
AOI21_X2 inst_20695 ( .ZN(net_12180), .A(net_12179), .B1(net_8271), .B2(net_7946) );
INV_X2 inst_19483 ( .A(net_8961), .ZN(net_1378) );
INV_X4 inst_12571 ( .A(net_18256), .ZN(net_18199) );
INV_X2 inst_19164 ( .ZN(net_3921), .A(net_3920) );
INV_X2 inst_19317 ( .ZN(net_2625), .A(net_2624) );
INV_X4 inst_13433 ( .ZN(net_12160), .A(net_9869) );
NAND3_X4 inst_5578 ( .ZN(net_19921), .A1(net_15346), .A3(net_14611), .A2(net_9482) );
INV_X4 inst_13396 ( .ZN(net_10662), .A(net_10661) );
NAND2_X2 inst_8655 ( .A2(net_16701), .ZN(net_16542), .A1(net_3347) );
NAND2_X2 inst_11459 ( .ZN(net_3550), .A2(net_3216), .A1(net_1515) );
NOR2_X2 inst_4599 ( .ZN(net_6568), .A1(net_6135), .A2(net_3767) );
CLKBUF_X2 inst_22466 ( .A(net_22337), .Z(net_22338) );
NAND2_X2 inst_8147 ( .ZN(net_18018), .A2(net_17983), .A1(net_17860) );
NAND3_X2 inst_5906 ( .ZN(net_15066), .A3(net_13116), .A1(net_9853), .A2(net_9527) );
AOI21_X4 inst_20133 ( .B1(net_19160), .ZN(net_16079), .B2(net_15827), .A(net_14015) );
NOR2_X2 inst_4677 ( .ZN(net_3237), .A2(net_2530), .A1(net_222) );
AOI21_X2 inst_20281 ( .B2(net_19156), .B1(net_19155), .A(net_16347), .ZN(net_16277) );
CLKBUF_X2 inst_21962 ( .A(net_21524), .Z(net_21834) );
INV_X4 inst_14796 ( .ZN(net_3998), .A(net_3997) );
NAND4_X2 inst_5516 ( .ZN(net_9957), .A1(net_9956), .A2(net_9955), .A4(net_9954), .A3(net_3958) );
OAI21_X2 inst_1698 ( .B2(net_20450), .B1(net_20449), .ZN(net_19853), .A(net_1550) );
NAND2_X2 inst_11698 ( .ZN(net_3016), .A2(net_1748), .A1(net_170) );
SDFF_X2 inst_944 ( .QN(net_20988), .D(net_2473), .SE(net_253), .CK(net_22676), .SI(x3199) );
NAND4_X4 inst_5248 ( .ZN(net_19800), .A4(net_13472), .A1(net_9857), .A2(net_9147), .A3(net_7612) );
INV_X4 inst_15488 ( .A(net_7580), .ZN(net_2574) );
NAND2_X2 inst_7992 ( .ZN(net_18375), .A2(net_18267), .A1(net_18228) );
INV_X4 inst_16924 ( .ZN(net_2934), .A(net_2456) );
XNOR2_X2 inst_459 ( .B(net_15959), .ZN(net_13949), .A(net_9238) );
NAND2_X2 inst_8259 ( .ZN(net_17691), .A2(net_17690), .A1(net_17668) );
CLKBUF_X2 inst_22344 ( .A(net_21490), .Z(net_22216) );
NAND2_X2 inst_11737 ( .ZN(net_2182), .A1(net_2181), .A2(net_2180) );
NAND2_X2 inst_8532 ( .A1(net_20515), .ZN(net_16863), .A2(net_16786) );
DFF_X1 inst_19794 ( .D(net_18262), .CK(net_22829), .Q(x1068) );
NAND2_X2 inst_10084 ( .A2(net_10261), .ZN(net_8633), .A1(net_5903) );
NAND2_X4 inst_7461 ( .ZN(net_4951), .A2(net_2747), .A1(net_2636) );
INV_X4 inst_12861 ( .ZN(net_17039), .A(net_17038) );
INV_X4 inst_17396 ( .ZN(net_5241), .A(net_522) );
CLKBUF_X2 inst_22952 ( .A(net_21755), .Z(net_22824) );
AND2_X4 inst_21169 ( .ZN(net_19152), .A1(net_14782), .A2(net_10404) );
INV_X4 inst_13723 ( .ZN(net_7805), .A(net_7804) );
NOR2_X2 inst_3393 ( .ZN(net_19146), .A2(net_15732), .A1(net_15610) );
CLKBUF_X2 inst_21919 ( .A(net_21623), .Z(net_21791) );
NAND2_X2 inst_8613 ( .ZN(net_16616), .A2(net_16615), .A1(net_9712) );
CLKBUF_X2 inst_22117 ( .A(net_21732), .Z(net_21989) );
INV_X2 inst_18470 ( .ZN(net_12698), .A(net_12697) );
NAND2_X2 inst_8148 ( .ZN(net_18017), .A1(net_17972), .A2(net_17940) );
INV_X2 inst_18403 ( .A(net_16804), .ZN(net_16421) );
NOR2_X2 inst_4976 ( .A2(net_2773), .ZN(net_1551), .A1(net_222) );
AOI21_X4 inst_20132 ( .B1(net_19373), .ZN(net_19272), .B2(net_15550), .A(net_14077) );
NAND2_X2 inst_9657 ( .ZN(net_10336), .A2(net_7752), .A1(net_1267) );
NOR2_X2 inst_3409 ( .A2(net_20114), .A1(net_20113), .ZN(net_15734) );
CLKBUF_X2 inst_21695 ( .A(net_21480), .Z(net_21567) );
INV_X4 inst_13252 ( .ZN(net_12761), .A(net_11749) );
NOR2_X2 inst_3591 ( .A1(net_13348), .ZN(net_12608), .A2(net_12607) );
NAND3_X2 inst_5970 ( .A3(net_19416), .A1(net_19415), .ZN(net_14774), .A2(net_10123) );
INV_X4 inst_16888 ( .ZN(net_14788), .A(net_449) );
INV_X4 inst_16242 ( .ZN(net_1864), .A(net_1810) );
XNOR2_X2 inst_450 ( .ZN(net_14826), .A(net_14825), .B(net_2313) );
NAND2_X2 inst_9723 ( .A2(net_11874), .ZN(net_10145), .A1(net_10144) );
INV_X2 inst_18785 ( .ZN(net_7501), .A(net_7500) );
XNOR2_X2 inst_520 ( .A(net_18141), .ZN(net_4492), .B(net_4491) );
NAND3_X2 inst_5717 ( .ZN(net_20122), .A3(net_20000), .A1(net_19999), .A2(net_13708) );
NOR2_X2 inst_3658 ( .ZN(net_11628), .A2(net_11627), .A1(net_9121) );
CLKBUF_X2 inst_22411 ( .A(net_22282), .Z(net_22283) );
NAND2_X2 inst_10019 ( .ZN(net_8770), .A1(net_8769), .A2(net_8768) );
INV_X2 inst_18701 ( .ZN(net_8300), .A(net_8299) );
INV_X4 inst_17142 ( .ZN(net_1102), .A(net_170) );
NAND2_X2 inst_11667 ( .A2(net_6097), .A1(net_2686), .ZN(net_2383) );
NOR2_X2 inst_4554 ( .ZN(net_4956), .A2(net_3850), .A1(net_2630) );
INV_X4 inst_14850 ( .ZN(net_4892), .A(net_3828) );
NAND3_X2 inst_5977 ( .ZN(net_14624), .A3(net_12150), .A1(net_8385), .A2(net_6666) );
OAI21_X2 inst_2026 ( .ZN(net_11320), .A(net_10676), .B1(net_8867), .B2(net_7477) );
NOR2_X2 inst_3623 ( .ZN(net_13586), .A2(net_12378), .A1(net_10765) );
OAI21_X2 inst_1556 ( .B2(net_19458), .ZN(net_17708), .A(net_17181), .B1(net_16685) );
NAND2_X2 inst_9228 ( .ZN(net_19345), .A2(net_10159), .A1(net_6973) );
INV_X4 inst_14820 ( .ZN(net_5024), .A(net_3918) );
NAND3_X2 inst_6796 ( .A2(net_4990), .ZN(net_3453), .A1(net_3452), .A3(net_3451) );
INV_X4 inst_15636 ( .A(net_3061), .ZN(net_2878) );
NAND2_X2 inst_11243 ( .A1(net_4288), .ZN(net_3928), .A2(net_2905) );
INV_X4 inst_17450 ( .A(net_2221), .ZN(net_465) );
NAND2_X2 inst_12075 ( .ZN(net_1561), .A1(net_227), .A2(net_144) );
INV_X4 inst_14410 ( .ZN(net_8006), .A(net_3382) );
SDFF_X2 inst_862 ( .Q(net_21236), .D(net_17169), .SE(net_263), .CK(net_22440), .SI(x6797) );
NOR2_X2 inst_4358 ( .ZN(net_5569), .A2(net_4855), .A1(net_1335) );
NOR2_X2 inst_4390 ( .ZN(net_6303), .A1(net_5201), .A2(net_2865) );
INV_X4 inst_16387 ( .ZN(net_6598), .A(net_3750) );
INV_X4 inst_14618 ( .ZN(net_8050), .A(net_4410) );
INV_X4 inst_17383 ( .A(net_14308), .ZN(net_538) );
NAND2_X2 inst_10620 ( .A2(net_20782), .ZN(net_11956), .A1(net_6863) );
OAI21_X2 inst_1764 ( .A(net_14974), .ZN(net_14704), .B2(net_12159), .B1(net_6555) );
CLKBUF_X2 inst_22513 ( .A(net_21835), .Z(net_22385) );
INV_X4 inst_14024 ( .ZN(net_9705), .A(net_6290) );
NAND4_X2 inst_5271 ( .A4(net_20180), .A1(net_20179), .ZN(net_16119), .A2(net_14644), .A3(net_13794) );
INV_X4 inst_14799 ( .A(net_11279), .ZN(net_3987) );
NAND4_X2 inst_5323 ( .ZN(net_15727), .A4(net_14968), .A2(net_14145), .A1(net_14071), .A3(net_13815) );
INV_X4 inst_15366 ( .ZN(net_6548), .A(net_4491) );
INV_X2 inst_19409 ( .ZN(net_1978), .A(net_1977) );
NAND2_X4 inst_7472 ( .ZN(net_7096), .A1(net_1312), .A2(net_374) );
OR2_X2 inst_1159 ( .ZN(net_11393), .A2(net_7488), .A1(net_5153) );
NAND2_X2 inst_8740 ( .ZN(net_20052), .A1(net_15710), .A2(net_15424) );
NAND2_X2 inst_9550 ( .ZN(net_11030), .A2(net_11029), .A1(net_10623) );
NAND2_X2 inst_8659 ( .ZN(net_19143), .A2(net_16526), .A1(net_675) );
INV_X4 inst_16612 ( .ZN(net_6611), .A(net_809) );
NAND2_X2 inst_9835 ( .ZN(net_9580), .A1(net_9579), .A2(net_9578) );
SDFF_X2 inst_938 ( .QN(net_21054), .D(net_509), .SE(net_263), .CK(net_22534), .SI(x2139) );
INV_X4 inst_16420 ( .ZN(net_15046), .A(net_588) );
INV_X4 inst_14521 ( .ZN(net_5943), .A(net_4779) );
AOI21_X2 inst_20792 ( .ZN(net_18939), .B2(net_10506), .A(net_8417), .B1(net_8416) );
AOI21_X2 inst_20326 ( .ZN(net_20593), .B2(net_15325), .A(net_14305), .B1(net_1062) );
NAND2_X2 inst_11189 ( .ZN(net_7043), .A1(net_4508), .A2(net_4098) );
INV_X4 inst_12552 ( .ZN(net_18325), .A(net_18260) );
INV_X4 inst_12742 ( .ZN(net_17436), .A(net_17435) );
INV_X4 inst_16752 ( .ZN(net_1507), .A(net_806) );
AOI21_X2 inst_20522 ( .ZN(net_14561), .B2(net_11972), .A(net_8597), .B1(net_828) );
NAND3_X2 inst_6646 ( .ZN(net_8725), .A1(net_8724), .A3(net_5112), .A2(net_874) );
CLKBUF_X2 inst_21723 ( .A(net_21594), .Z(net_21595) );
DFF_X1 inst_19921 ( .Q(net_21111), .D(net_14379), .CK(net_21692) );
NAND2_X2 inst_9698 ( .ZN(net_19501), .A1(net_10922), .A2(net_10221) );
NOR2_X2 inst_3638 ( .ZN(net_12108), .A2(net_10039), .A1(net_8674) );
NAND2_X2 inst_8923 ( .ZN(net_14953), .A2(net_13729), .A1(net_3662) );
NOR2_X2 inst_4365 ( .ZN(net_5493), .A2(net_5492), .A1(net_3922) );
NAND2_X2 inst_9399 ( .ZN(net_11698), .A2(net_11697), .A1(net_9766) );
INV_X2 inst_18899 ( .ZN(net_10211), .A(net_6094) );
INV_X4 inst_16881 ( .A(net_7439), .ZN(net_5694) );
INV_X4 inst_18151 ( .A(net_21079), .ZN(net_406) );
NAND2_X2 inst_8957 ( .A1(net_14994), .ZN(net_14716), .A2(net_13210) );
AOI22_X2 inst_20021 ( .ZN(net_11149), .A1(net_11148), .B1(net_9247), .A2(net_8155), .B2(net_2961) );
NAND2_X2 inst_11320 ( .ZN(net_10520), .A1(net_6655), .A2(net_3759) );
INV_X4 inst_14253 ( .ZN(net_5757), .A(net_5756) );
INV_X2 inst_19124 ( .ZN(net_4390), .A(net_4389) );
NAND2_X4 inst_7426 ( .ZN(net_5074), .A1(net_4192), .A2(net_3505) );
OAI21_X2 inst_2102 ( .ZN(net_10064), .A(net_10063), .B1(net_8408), .B2(net_6168) );
INV_X4 inst_14070 ( .ZN(net_11273), .A(net_5515) );
INV_X2 inst_19298 ( .ZN(net_5057), .A(net_4081) );
NAND2_X2 inst_9762 ( .ZN(net_9839), .A2(net_9838), .A1(net_8495) );
NOR2_X2 inst_4908 ( .ZN(net_3595), .A1(net_2007), .A2(net_1949) );
NAND2_X4 inst_7160 ( .ZN(net_11603), .A1(net_9536), .A2(net_6358) );
NAND2_X4 inst_7619 ( .ZN(net_1665), .A2(net_1331), .A1(net_343) );
CLKBUF_X2 inst_22902 ( .A(net_22773), .Z(net_22774) );
NAND2_X2 inst_10343 ( .ZN(net_7526), .A2(net_5972), .A1(net_5840) );
INV_X4 inst_16806 ( .A(net_20875), .ZN(net_5591) );
NAND3_X2 inst_6168 ( .ZN(net_13618), .A2(net_13617), .A3(net_13616), .A1(net_12395) );
NAND2_X2 inst_8445 ( .ZN(net_17111), .A2(net_16929), .A1(net_16445) );
INV_X2 inst_19576 ( .ZN(net_919), .A(net_326) );
INV_X2 inst_18892 ( .ZN(net_9425), .A(net_6105) );
NAND2_X2 inst_11182 ( .ZN(net_8395), .A1(net_4179), .A2(net_2176) );
SDFF_X2 inst_784 ( .Q(net_20849), .SE(net_18581), .SI(net_18040), .D(net_728), .CK(net_22626) );
NOR2_X4 inst_3237 ( .ZN(net_5284), .A1(net_1475), .A2(net_1376) );
OAI22_X2 inst_1264 ( .B1(net_21142), .ZN(net_17142), .A1(net_17015), .A2(net_16785), .B2(net_16784) );
INV_X2 inst_19185 ( .A(net_4804), .ZN(net_3733) );
XNOR2_X1 inst_690 ( .A(net_17767), .ZN(net_16529), .B(net_11876) );
INV_X2 inst_19658 ( .ZN(net_20435), .A(net_20434) );
INV_X2 inst_18469 ( .ZN(net_12704), .A(net_11643) );
NAND2_X2 inst_11895 ( .A2(net_3696), .A1(net_2996), .ZN(net_2395) );
OAI21_X2 inst_2025 ( .ZN(net_11321), .B1(net_8249), .B2(net_7463), .A(net_731) );
CLKBUF_X2 inst_21445 ( .A(net_21316), .Z(net_21317) );
AOI21_X2 inst_20856 ( .ZN(net_20374), .A(net_11182), .B2(net_10644), .B1(net_4475) );
NAND2_X2 inst_7819 ( .ZN(net_18667), .A1(net_18625), .A2(net_18613) );
CLKBUF_X2 inst_21726 ( .A(net_21597), .Z(net_21598) );
NAND2_X2 inst_10607 ( .ZN(net_7869), .A1(net_4288), .A2(net_3869) );
NOR2_X2 inst_4717 ( .A2(net_6489), .ZN(net_5602), .A1(net_3133) );
INV_X4 inst_12722 ( .ZN(net_17718), .A(net_17611) );
CLKBUF_X2 inst_21772 ( .A(net_21253), .Z(net_21644) );
AOI21_X2 inst_20785 ( .B1(net_12440), .ZN(net_10552), .B2(net_6422), .A(net_6246) );
INV_X4 inst_18179 ( .A(net_21094), .ZN(net_746) );
NAND2_X2 inst_10969 ( .A1(net_5139), .ZN(net_5007), .A2(net_5006) );
NAND2_X2 inst_9666 ( .ZN(net_19749), .A1(net_10467), .A2(net_10314) );
AOI21_X2 inst_20331 ( .B1(net_19652), .ZN(net_15821), .B2(net_15186), .A(net_12879) );
XNOR2_X2 inst_75 ( .ZN(net_18712), .B(net_18664), .A(net_18017) );
CLKBUF_X2 inst_22580 ( .A(net_22451), .Z(net_22452) );
AOI21_X2 inst_20475 ( .A(net_20889), .ZN(net_19563), .B1(net_13810), .B2(net_12667) );
NAND2_X2 inst_7714 ( .ZN(net_18849), .A2(net_18832), .A1(net_18817) );
CLKBUF_X2 inst_22171 ( .A(net_22042), .Z(net_22043) );
INV_X4 inst_15656 ( .ZN(net_3945), .A(net_2098) );
NAND3_X2 inst_6386 ( .A2(net_14867), .ZN(net_12016), .A3(net_11792), .A1(net_11025) );
AOI22_X2 inst_20023 ( .B1(net_12320), .ZN(net_10513), .A1(net_10512), .A2(net_6522), .B2(net_5955) );
INV_X4 inst_16182 ( .A(net_2300), .ZN(net_1426) );
NAND2_X2 inst_7986 ( .ZN(net_18331), .A2(net_18330), .A1(net_17994) );
INV_X2 inst_19046 ( .ZN(net_4753), .A(net_4752) );
NAND2_X2 inst_9286 ( .A1(net_14972), .ZN(net_12539), .A2(net_12538) );
AND2_X4 inst_21181 ( .A1(net_11894), .ZN(net_11585), .A2(net_11584) );
NAND2_X4 inst_7600 ( .A2(net_2497), .ZN(net_1448), .A1(net_252) );
NAND2_X2 inst_7891 ( .ZN(net_18505), .A1(net_18443), .A2(net_18392) );
INV_X2 inst_18984 ( .ZN(net_5124), .A(net_5123) );
CLKBUF_X2 inst_22492 ( .A(net_22363), .Z(net_22364) );
NAND2_X2 inst_12082 ( .ZN(net_767), .A2(net_766), .A1(net_176) );
INV_X2 inst_19171 ( .A(net_5468), .ZN(net_3827) );
INV_X4 inst_13938 ( .ZN(net_8145), .A(net_7227) );
NAND2_X2 inst_10890 ( .A2(net_14334), .ZN(net_5404), .A1(net_5403) );
NAND2_X2 inst_10339 ( .ZN(net_11040), .A1(net_7538), .A2(net_4607) );
SDFF_X2 inst_1024 ( .QN(net_21079), .SE(net_2426), .D(net_406), .CK(net_22561), .SI(x1731) );
NAND3_X2 inst_5827 ( .A1(net_19843), .ZN(net_19346), .A3(net_10488), .A2(net_4178) );
NAND2_X1 inst_12144 ( .A2(net_17019), .ZN(net_16872), .A1(net_643) );
OAI21_X2 inst_2232 ( .ZN(net_8183), .A(net_3640), .B2(net_3605), .B1(net_2209) );
NOR2_X2 inst_4546 ( .A1(net_20555), .ZN(net_6940), .A2(net_2882) );
INV_X4 inst_13218 ( .ZN(net_20816), .A(net_12792) );
NAND2_X2 inst_12061 ( .ZN(net_876), .A1(net_875), .A2(net_722) );
INV_X4 inst_16716 ( .ZN(net_5204), .A(net_874) );
OAI21_X2 inst_1689 ( .ZN(net_15379), .A(net_14697), .B1(net_14141), .B2(net_12849) );
NAND2_X2 inst_8279 ( .ZN(net_17720), .A2(net_17489), .A1(net_17373) );
NOR2_X4 inst_2846 ( .ZN(net_14130), .A2(net_12267), .A1(net_6512) );
NOR2_X2 inst_3584 ( .ZN(net_14802), .A1(net_12658), .A2(net_12657) );
NAND2_X2 inst_11408 ( .A2(net_3614), .ZN(net_3432), .A1(net_2919) );
NAND2_X2 inst_9472 ( .A2(net_11582), .ZN(net_11473), .A1(net_11472) );
OAI21_X4 inst_1448 ( .B2(net_19091), .B1(net_19090), .ZN(net_18961), .A(net_15664) );
NAND2_X2 inst_8395 ( .ZN(net_20085), .A2(net_16972), .A1(net_16816) );
OAI21_X2 inst_1816 ( .ZN(net_14168), .B2(net_10731), .A(net_10389), .B1(net_6016) );
NAND2_X2 inst_11892 ( .ZN(net_4222), .A1(net_1593), .A2(net_1518) );
NAND2_X2 inst_11723 ( .A1(net_3713), .ZN(net_2236), .A2(net_2235) );
INV_X4 inst_14829 ( .ZN(net_10238), .A(net_3895) );
NOR2_X2 inst_5012 ( .A1(net_20851), .ZN(net_1265), .A2(net_1264) );
INV_X2 inst_19343 ( .A(net_6487), .ZN(net_2447) );
NOR2_X2 inst_3381 ( .ZN(net_20026), .A2(net_16254), .A1(net_15845) );
INV_X4 inst_17636 ( .ZN(net_13030), .A(net_277) );
INV_X4 inst_14123 ( .ZN(net_7534), .A(net_6125) );
OR2_X4 inst_1091 ( .ZN(net_9087), .A1(net_8273), .A2(net_5367) );
NAND2_X2 inst_9915 ( .ZN(net_13607), .A2(net_9430), .A1(net_9310) );
NOR2_X2 inst_4837 ( .ZN(net_2373), .A2(net_1137), .A1(net_117) );
NOR2_X2 inst_5059 ( .ZN(net_1003), .A2(net_856), .A1(net_153) );
NAND2_X2 inst_8206 ( .ZN(net_17871), .A2(net_17713), .A1(net_17620) );
NAND2_X2 inst_10450 ( .ZN(net_7061), .A1(net_7054), .A2(net_4381) );
INV_X4 inst_16308 ( .ZN(net_2345), .A(net_1221) );
INV_X4 inst_13800 ( .A(net_10598), .ZN(net_7557) );
INV_X2 inst_18525 ( .A(net_13220), .ZN(net_11130) );
NOR2_X2 inst_4154 ( .ZN(net_6897), .A1(net_6896), .A2(net_6895) );
NAND2_X2 inst_10374 ( .ZN(net_12513), .A2(net_7392), .A1(net_70) );
NAND4_X2 inst_5398 ( .ZN(net_19078), .A3(net_14798), .A4(net_12931), .A1(net_11410), .A2(net_10684) );
AOI21_X2 inst_20680 ( .ZN(net_19114), .B1(net_12382), .B2(net_7359), .A(net_6359) );
NOR2_X2 inst_4816 ( .ZN(net_4266), .A2(net_2569), .A1(net_2568) );
CLKBUF_X2 inst_22883 ( .A(net_21246), .Z(net_22755) );
NOR2_X4 inst_3179 ( .ZN(net_5611), .A1(net_3136), .A2(net_2012) );
AOI21_X2 inst_20288 ( .B1(net_19219), .B2(net_16347), .ZN(net_16215), .A(net_15261) );
NOR2_X4 inst_3059 ( .ZN(net_6109), .A2(net_4833), .A1(net_1357) );
INV_X4 inst_15297 ( .ZN(net_2704), .A(net_1909) );
NAND2_X2 inst_11357 ( .ZN(net_20679), .A2(net_3658), .A1(net_3617) );
CLKBUF_X2 inst_21407 ( .A(net_21278), .Z(net_21279) );
AOI21_X2 inst_20570 ( .ZN(net_14147), .B1(net_12864), .B2(net_10771), .A(net_5404) );
INV_X4 inst_15660 ( .A(net_2481), .ZN(net_2087) );
AND3_X4 inst_21119 ( .ZN(net_13160), .A3(net_13159), .A2(net_12807), .A1(net_9503) );
NAND2_X2 inst_9390 ( .ZN(net_11715), .A2(net_9577), .A1(net_7028) );
OAI211_X2 inst_2587 ( .ZN(net_6388), .B(net_6387), .A(net_4606), .C1(net_4511), .C2(net_1840) );
NAND3_X2 inst_6680 ( .ZN(net_7737), .A3(net_5564), .A1(net_4547), .A2(net_3571) );
NAND2_X2 inst_8868 ( .ZN(net_19569), .A1(net_14974), .A2(net_14246) );
AOI21_X2 inst_20586 ( .ZN(net_14023), .A(net_14022), .B2(net_11298), .B1(net_9856) );
INV_X2 inst_19664 ( .A(net_20472), .ZN(net_20471) );
INV_X4 inst_13072 ( .ZN(net_16339), .A(net_16185) );
AOI21_X2 inst_20268 ( .A(net_18067), .ZN(net_18056), .B2(net_15855), .B1(net_10953) );
NAND2_X2 inst_8883 ( .ZN(net_15153), .A1(net_14352), .A2(net_14152) );
NOR2_X4 inst_3031 ( .ZN(net_6310), .A2(net_5204), .A1(net_3979) );
INV_X4 inst_18218 ( .A(net_21205), .ZN(net_15294) );
OAI22_X2 inst_1257 ( .B1(net_21120), .A2(net_20713), .B2(net_20712), .ZN(net_17523), .A1(net_17522) );
SDFF_X2 inst_875 ( .Q(net_21180), .SI(net_17042), .SE(net_125), .CK(net_22230), .D(x6600) );
NOR2_X4 inst_3298 ( .ZN(net_2178), .A2(net_540), .A1(net_221) );
NOR2_X2 inst_3482 ( .ZN(net_14310), .A2(net_13522), .A1(net_11407) );
NOR2_X2 inst_5075 ( .ZN(net_908), .A2(net_766), .A1(net_63) );
INV_X2 inst_19330 ( .A(net_3609), .ZN(net_2544) );
INV_X4 inst_17680 ( .A(net_307), .ZN(net_235) );
OAI21_X2 inst_2069 ( .A(net_12298), .ZN(net_10658), .B2(net_8657), .B1(net_6343) );
AOI21_X2 inst_20704 ( .A(net_14203), .ZN(net_12127), .B2(net_8396), .B1(net_5331) );
CLKBUF_X2 inst_21842 ( .A(net_21713), .Z(net_21714) );
AOI22_X2 inst_20057 ( .A1(net_4751), .A2(net_3045), .ZN(net_2949), .B2(net_2948), .B1(net_1415) );
INV_X4 inst_15032 ( .ZN(net_4768), .A(net_3361) );
NOR2_X2 inst_4098 ( .A1(net_11691), .ZN(net_7228), .A2(net_7227) );
NAND2_X2 inst_11220 ( .A2(net_8537), .A1(net_5472), .ZN(net_4994) );
NAND3_X2 inst_5703 ( .A3(net_19742), .A1(net_19741), .ZN(net_16217), .A2(net_13795) );
NOR2_X4 inst_2978 ( .A1(net_20315), .ZN(net_7573), .A2(net_3800) );
AND2_X2 inst_21298 ( .ZN(net_20594), .A2(net_10117), .A1(net_9967) );
INV_X2 inst_19622 ( .A(net_20971), .ZN(net_94) );
INV_X4 inst_14817 ( .ZN(net_5538), .A(net_3930) );
INV_X4 inst_14239 ( .ZN(net_5805), .A(net_5804) );
NAND2_X2 inst_11033 ( .ZN(net_9676), .A1(net_4751), .A2(net_2833) );
NAND2_X2 inst_11393 ( .ZN(net_7750), .A2(net_3409), .A1(net_547) );
NAND2_X2 inst_10269 ( .ZN(net_19055), .A1(net_13353), .A2(net_5103) );
INV_X4 inst_14352 ( .ZN(net_5283), .A(net_5282) );
OAI21_X2 inst_2019 ( .ZN(net_11344), .A(net_11311), .B1(net_11218), .B2(net_6944) );
INV_X4 inst_13679 ( .ZN(net_10101), .A(net_8712) );
NAND2_X2 inst_8323 ( .ZN(net_17556), .A1(net_17304), .A2(net_17292) );
NAND4_X4 inst_5186 ( .A4(net_18970), .A1(net_18969), .ZN(net_17052), .A3(net_16345), .A2(net_14042) );
CLKBUF_X2 inst_22230 ( .A(net_22101), .Z(net_22102) );
INV_X4 inst_15061 ( .ZN(net_4520), .A(net_3300) );
XNOR2_X2 inst_69 ( .B(net_19557), .ZN(net_18802), .A(net_18752) );
INV_X2 inst_18854 ( .ZN(net_6368), .A(net_6367) );
INV_X4 inst_18077 ( .A(net_20970), .ZN(net_602) );
INV_X4 inst_15542 ( .ZN(net_6402), .A(net_1673) );
INV_X4 inst_14448 ( .ZN(net_6123), .A(net_4973) );
NOR3_X2 inst_2669 ( .A3(net_19801), .A1(net_19800), .ZN(net_14830), .A2(net_9347) );
INV_X4 inst_15396 ( .A(net_3949), .ZN(net_2542) );
INV_X4 inst_17278 ( .A(net_11395), .ZN(net_10686) );
INV_X4 inst_12844 ( .A(net_17633), .ZN(net_17204) );
INV_X4 inst_17319 ( .ZN(net_15454), .A(net_10122) );
SDFF_X2 inst_844 ( .Q(net_21176), .SI(net_17316), .SE(net_125), .CK(net_21660), .D(x4668) );
OAI211_X2 inst_2489 ( .C1(net_14185), .ZN(net_13197), .A(net_13196), .B(net_13149), .C2(net_4984) );
INV_X4 inst_14712 ( .ZN(net_5179), .A(net_3152) );
NAND2_X4 inst_6968 ( .ZN(net_17413), .A1(net_17005), .A2(net_16863) );
CLKBUF_X2 inst_22237 ( .A(net_22108), .Z(net_22109) );
NOR2_X2 inst_3619 ( .ZN(net_12354), .A1(net_12353), .A2(net_8972) );
NAND3_X2 inst_6709 ( .ZN(net_7110), .A3(net_7109), .A1(net_3916), .A2(net_3029) );
NAND3_X2 inst_5805 ( .ZN(net_15658), .A2(net_14941), .A3(net_14524), .A1(net_11636) );
NAND2_X4 inst_6939 ( .A2(net_19352), .A1(net_19351), .ZN(net_17851) );
NOR2_X2 inst_4641 ( .A1(net_3452), .ZN(net_3401), .A2(net_3238) );
NAND2_X4 inst_7056 ( .A2(net_20864), .A1(net_20095), .ZN(net_16360) );
NAND2_X2 inst_11038 ( .ZN(net_12523), .A1(net_5204), .A2(net_3948) );
XNOR2_X2 inst_460 ( .ZN(net_13292), .B(net_13291), .A(net_9195) );
NAND2_X2 inst_10877 ( .ZN(net_5983), .A2(net_5422), .A1(net_3947) );
OAI21_X4 inst_1455 ( .ZN(net_20645), .B2(net_20081), .B1(net_20080), .A(net_1046) );
NAND2_X4 inst_7135 ( .ZN(net_14303), .A1(net_10189), .A2(net_8202) );
OAI211_X2 inst_2497 ( .ZN(net_12867), .B(net_12866), .A(net_11124), .C1(net_9498), .C2(net_4651) );
NOR2_X2 inst_3660 ( .ZN(net_11601), .A2(net_11548), .A1(net_8824) );
INV_X4 inst_16975 ( .ZN(net_2686), .A(net_514) );
INV_X4 inst_15678 ( .ZN(net_11204), .A(net_2044) );
INV_X4 inst_16274 ( .ZN(net_8048), .A(net_732) );
NOR2_X2 inst_4230 ( .ZN(net_8733), .A1(net_6589), .A2(net_6588) );
INV_X4 inst_15316 ( .ZN(net_4814), .A(net_2640) );
INV_X4 inst_16771 ( .ZN(net_6840), .A(net_5277) );
NAND3_X4 inst_5571 ( .ZN(net_20352), .A3(net_15302), .A2(net_14722), .A1(net_14647) );
INV_X4 inst_13455 ( .A(net_11865), .ZN(net_9726) );
SDFF_X2 inst_950 ( .QN(net_20991), .D(net_2458), .SE(net_263), .CK(net_21851), .SI(x3153) );
NOR2_X2 inst_3955 ( .A1(net_9532), .ZN(net_8599), .A2(net_6483) );
OR2_X2 inst_1218 ( .ZN(net_2752), .A1(net_2751), .A2(net_2750) );
NAND2_X2 inst_8458 ( .A1(net_21133), .ZN(net_19041), .A2(net_17441) );
NAND3_X2 inst_6414 ( .A3(net_13941), .ZN(net_11950), .A2(net_6794), .A1(net_6380) );
INV_X4 inst_15842 ( .ZN(net_15688), .A(net_828) );
NAND2_X2 inst_9541 ( .A1(net_11925), .ZN(net_11056), .A2(net_11055) );
INV_X2 inst_19464 ( .ZN(net_3160), .A(net_1465) );
XNOR2_X2 inst_101 ( .ZN(net_18534), .A(net_18425), .B(net_17536) );
INV_X2 inst_19526 ( .ZN(net_1940), .A(net_1055) );
CLKBUF_X2 inst_21461 ( .A(net_21332), .Z(net_21333) );
INV_X2 inst_19697 ( .ZN(net_20552), .A(net_20548) );
INV_X4 inst_17696 ( .ZN(net_3350), .A(net_218) );
INV_X4 inst_14033 ( .A(net_6276), .ZN(net_6275) );
NOR2_X2 inst_3555 ( .ZN(net_13034), .A2(net_10419), .A1(net_10181) );
CLKBUF_X2 inst_22249 ( .A(net_22120), .Z(net_22121) );
NAND2_X2 inst_10234 ( .ZN(net_9583), .A2(net_8044), .A1(net_7121) );
INV_X4 inst_14377 ( .ZN(net_8120), .A(net_5174) );
CLKBUF_X2 inst_22212 ( .A(net_22083), .Z(net_22084) );
AND2_X2 inst_21291 ( .ZN(net_20168), .A1(net_12126), .A2(net_12125) );
CLKBUF_X2 inst_21630 ( .A(net_21501), .Z(net_21502) );
NAND2_X2 inst_11388 ( .ZN(net_6826), .A1(net_3516), .A2(net_1201) );
NOR2_X2 inst_4722 ( .ZN(net_4122), .A2(net_3113), .A1(net_966) );
XNOR2_X2 inst_510 ( .B(net_21207), .ZN(net_7353), .A(net_4447) );
AOI21_X4 inst_20123 ( .B2(net_19414), .B1(net_19413), .ZN(net_16212), .A(net_15667) );
INV_X8 inst_12194 ( .ZN(net_16718), .A(net_16382) );
NAND3_X2 inst_6505 ( .ZN(net_10806), .A3(net_7070), .A2(net_6971), .A1(net_5609) );
CLKBUF_X2 inst_21920 ( .A(net_21791), .Z(net_21792) );
OAI21_X2 inst_1677 ( .ZN(net_15494), .B2(net_14579), .A(net_14341), .B1(net_13089) );
SDFF_X2 inst_830 ( .Q(net_21226), .SI(net_17538), .SE(net_125), .CK(net_21407), .D(x7158) );
NAND2_X2 inst_8433 ( .ZN(net_17450), .A1(net_16855), .A2(net_16686) );
INV_X4 inst_15646 ( .ZN(net_5852), .A(net_2113) );
NOR2_X4 inst_2878 ( .ZN(net_11566), .A1(net_9587), .A2(net_5479) );
OAI211_X2 inst_2494 ( .ZN(net_13153), .B(net_13152), .A(net_11748), .C1(net_8791), .C2(net_5980) );
SDFF_X2 inst_776 ( .Q(net_20896), .SE(net_18864), .SI(net_18431), .D(net_427), .CK(net_21428) );
INV_X2 inst_18480 ( .ZN(net_12587), .A(net_11405) );
OAI211_X2 inst_2526 ( .ZN(net_11785), .A(net_11784), .C1(net_11783), .C2(net_9658), .B(net_7275) );
NOR2_X2 inst_5047 ( .ZN(net_2303), .A1(net_1065), .A2(net_1031) );
CLKBUF_X2 inst_21777 ( .A(net_21648), .Z(net_21649) );
NAND2_X2 inst_10787 ( .ZN(net_5589), .A1(net_5588), .A2(net_5587) );
NAND4_X2 inst_5313 ( .A4(net_20164), .A1(net_20163), .ZN(net_19578), .A3(net_14902), .A2(net_13796) );
OAI21_X2 inst_1972 ( .A(net_20889), .ZN(net_12201), .B2(net_7802), .B1(net_5871) );
XNOR2_X2 inst_558 ( .B(net_9193), .ZN(net_689), .A(net_688) );
CLKBUF_X2 inst_22961 ( .A(net_22832), .Z(net_22833) );
NAND3_X2 inst_6167 ( .ZN(net_13627), .A3(net_12665), .A2(net_10406), .A1(net_8208) );
INV_X4 inst_12704 ( .ZN(net_17595), .A(net_17594) );
CLKBUF_X2 inst_21612 ( .A(net_21483), .Z(net_21484) );
NAND2_X2 inst_10591 ( .A1(net_10191), .ZN(net_6645), .A2(net_6644) );
XNOR2_X2 inst_389 ( .ZN(net_16772), .A(net_16766), .B(net_13291) );
NAND4_X4 inst_5179 ( .A4(net_19187), .A1(net_19186), .ZN(net_16656), .A3(net_16316), .A2(net_14043) );
INV_X4 inst_14301 ( .A(net_5768), .ZN(net_5535) );
INV_X4 inst_13460 ( .ZN(net_11501), .A(net_10235) );
NOR3_X2 inst_2712 ( .ZN(net_13614), .A3(net_12794), .A1(net_11529), .A2(net_5987) );
INV_X4 inst_16257 ( .ZN(net_14759), .A(net_13514) );
NAND2_X2 inst_10252 ( .A1(net_12504), .ZN(net_9545), .A2(net_5406) );
NAND3_X2 inst_6152 ( .ZN(net_13675), .A1(net_12270), .A3(net_11082), .A2(net_7551) );
CLKBUF_X2 inst_22578 ( .A(net_22449), .Z(net_22450) );
NAND2_X2 inst_8650 ( .A2(net_16912), .ZN(net_16561), .A1(net_16560) );
OAI21_X4 inst_1382 ( .A(net_20904), .B2(net_19178), .B1(net_19177), .ZN(net_16354) );
CLKBUF_X2 inst_22219 ( .A(net_22090), .Z(net_22091) );
NAND2_X2 inst_8841 ( .ZN(net_15445), .A1(net_15158), .A2(net_15014) );
NOR3_X2 inst_2795 ( .A2(net_3867), .ZN(net_3236), .A1(net_3235), .A3(net_1376) );
CLKBUF_X2 inst_21618 ( .A(net_21325), .Z(net_21490) );
NAND4_X2 inst_5266 ( .A4(net_19761), .A1(net_19760), .ZN(net_19302), .A2(net_13857), .A3(net_13792) );
NOR2_X2 inst_4766 ( .A1(net_9937), .ZN(net_7159), .A2(net_2510) );
INV_X2 inst_19240 ( .ZN(net_3303), .A(net_3302) );
NOR2_X2 inst_4445 ( .ZN(net_5956), .A2(net_4793), .A1(net_526) );
NAND3_X2 inst_5895 ( .A2(net_20330), .A1(net_20329), .A3(net_20178), .ZN(net_15181) );
INV_X4 inst_16545 ( .A(net_11442), .ZN(net_9727) );
INV_X4 inst_17726 ( .A(net_14029), .ZN(net_10122) );
INV_X4 inst_15898 ( .ZN(net_16214), .A(net_15880) );
NAND2_X2 inst_11785 ( .ZN(net_2002), .A1(net_2001), .A2(net_1206) );
NAND2_X2 inst_9977 ( .ZN(net_8871), .A1(net_8870), .A2(net_6514) );
INV_X4 inst_12866 ( .ZN(net_17287), .A(net_17014) );
INV_X4 inst_12766 ( .ZN(net_17673), .A(net_17225) );
NAND2_X2 inst_8365 ( .ZN(net_19641), .A2(net_17374), .A1(net_17107) );
INV_X4 inst_14195 ( .ZN(net_10454), .A(net_5975) );
INV_X2 inst_19108 ( .ZN(net_4485), .A(net_2058) );
CLKBUF_X2 inst_22742 ( .A(net_22613), .Z(net_22614) );
AOI21_X2 inst_20462 ( .ZN(net_15008), .B1(net_14962), .B2(net_13003), .A(net_7299) );
NAND2_X4 inst_7105 ( .ZN(net_12189), .A1(net_11297), .A2(net_9907) );
NAND2_X2 inst_10843 ( .ZN(net_6758), .A1(net_4890), .A2(net_4353) );
INV_X4 inst_18064 ( .A(net_20966), .ZN(net_87) );
INV_X4 inst_16789 ( .ZN(net_1755), .A(net_1013) );
NAND2_X2 inst_11613 ( .ZN(net_5035), .A1(net_2600), .A2(net_1094) );
NAND2_X4 inst_7687 ( .A1(net_19376), .ZN(net_753), .A2(net_275) );
AOI21_X2 inst_20860 ( .ZN(net_8898), .A(net_7394), .B2(net_6260), .B1(net_3619) );
NAND2_X2 inst_11133 ( .ZN(net_8947), .A2(net_4303), .A1(net_4205) );
INV_X4 inst_16067 ( .ZN(net_1889), .A(net_761) );
NAND2_X2 inst_11724 ( .A1(net_5169), .A2(net_2255), .ZN(net_2234) );
AOI21_X2 inst_20904 ( .B1(net_20806), .ZN(net_7696), .B2(net_3970), .A(net_2092) );
INV_X2 inst_19015 ( .A(net_6926), .ZN(net_4997) );
INV_X4 inst_17837 ( .ZN(net_890), .A(net_156) );
INV_X4 inst_13321 ( .ZN(net_13824), .A(net_11503) );
NAND2_X2 inst_9446 ( .ZN(net_11533), .A1(net_11532), .A2(net_5442) );
INV_X2 inst_18685 ( .ZN(net_8673), .A(net_8672) );
CLKBUF_X2 inst_22862 ( .A(net_22733), .Z(net_22734) );
INV_X4 inst_13467 ( .A(net_9672), .ZN(net_9671) );
NOR2_X2 inst_4212 ( .ZN(net_8625), .A2(net_7018), .A1(net_6736) );
AOI21_X2 inst_20633 ( .ZN(net_13372), .B2(net_8643), .B1(net_7011), .A(net_3803) );
AOI21_X2 inst_20795 ( .B2(net_20772), .A(net_11550), .ZN(net_10420), .B1(net_4649) );
INV_X4 inst_15257 ( .A(net_3753), .ZN(net_2785) );
INV_X4 inst_15716 ( .ZN(net_13554), .A(net_7004) );
NAND2_X2 inst_11231 ( .ZN(net_6794), .A2(net_3866), .A1(net_1724) );
INV_X4 inst_12912 ( .ZN(net_17216), .A(net_16684) );
NAND2_X2 inst_11759 ( .ZN(net_2851), .A2(net_2093), .A1(net_168) );
NAND2_X2 inst_9594 ( .ZN(net_10849), .A2(net_7732), .A1(net_269) );
INV_X4 inst_16238 ( .ZN(net_4150), .A(net_1157) );
OAI21_X2 inst_2309 ( .ZN(net_5751), .B2(net_5571), .B1(net_2194), .A(net_1173) );
DFF_X1 inst_19916 ( .D(net_16534), .CK(net_22070), .Q(x402) );
INV_X4 inst_15011 ( .ZN(net_11779), .A(net_10690) );
NAND2_X4 inst_7644 ( .ZN(net_1393), .A2(net_954), .A1(net_821) );
CLKBUF_X2 inst_21933 ( .A(net_21308), .Z(net_21805) );
INV_X4 inst_16285 ( .ZN(net_2114), .A(net_767) );
NAND2_X4 inst_7196 ( .ZN(net_14904), .A2(net_8304), .A1(net_8245) );
INV_X4 inst_18225 ( .A(net_21027), .ZN(net_648) );
NAND2_X2 inst_11283 ( .ZN(net_8438), .A1(net_5476), .A2(net_3856) );
NOR3_X4 inst_2603 ( .ZN(net_19898), .A3(net_16061), .A1(net_15760), .A2(net_6396) );
INV_X4 inst_15792 ( .ZN(net_2938), .A(net_1408) );
NAND2_X2 inst_11335 ( .ZN(net_3716), .A1(net_3715), .A2(net_1975) );
NOR2_X2 inst_4603 ( .ZN(net_6553), .A2(net_4269), .A1(net_1931) );
NAND2_X2 inst_9339 ( .ZN(net_12219), .A2(net_9280), .A1(net_278) );
OAI21_X2 inst_2153 ( .ZN(net_9302), .B1(net_9301), .A(net_5297), .B2(net_4593) );
CLKBUF_X2 inst_22910 ( .A(net_22781), .Z(net_22782) );
INV_X2 inst_18808 ( .ZN(net_7371), .A(net_7370) );
NAND2_X2 inst_11271 ( .ZN(net_3889), .A2(net_2429), .A1(net_193) );
NAND2_X2 inst_11904 ( .A2(net_1689), .ZN(net_1565), .A1(net_900) );
NAND2_X2 inst_11798 ( .ZN(net_1929), .A2(net_1216), .A1(net_1088) );
AND2_X4 inst_21268 ( .ZN(net_7077), .A1(net_790), .A2(net_165) );
INV_X2 inst_18759 ( .A(net_10348), .ZN(net_7635) );
INV_X4 inst_16996 ( .ZN(net_11461), .A(net_2344) );
NAND4_X2 inst_5494 ( .ZN(net_12234), .A2(net_12233), .A4(net_8534), .A3(net_6710), .A1(net_4861) );
AOI21_X2 inst_20776 ( .ZN(net_10615), .B2(net_6462), .A(net_5593), .B1(net_3886) );
NAND2_X2 inst_10586 ( .A1(net_8252), .ZN(net_6661), .A2(net_4779) );
AOI21_X2 inst_20825 ( .ZN(net_9872), .B1(net_9785), .A(net_5817), .B2(net_4486) );
NAND2_X4 inst_7674 ( .A1(net_1192), .ZN(net_1172), .A2(net_836) );
NAND4_X2 inst_5441 ( .ZN(net_13891), .A3(net_12835), .A4(net_11346), .A1(net_11158), .A2(net_9809) );
NAND2_X2 inst_9906 ( .ZN(net_9340), .A1(net_9339), .A2(net_9338) );
NAND2_X4 inst_6874 ( .A2(net_19002), .A1(net_19001), .ZN(net_18315) );
NOR2_X2 inst_3485 ( .ZN(net_14294), .A1(net_14293), .A2(net_12630) );
NAND3_X2 inst_5854 ( .ZN(net_15409), .A3(net_14477), .A2(net_11740), .A1(net_11500) );
NAND2_X2 inst_8587 ( .A1(net_19443), .ZN(net_16713), .A2(net_16439) );
NAND2_X2 inst_8680 ( .A1(net_20215), .A2(net_16774), .ZN(net_16453) );
CLKBUF_X2 inst_22763 ( .A(net_22101), .Z(net_22635) );
HA_X1 inst_19766 ( .S(net_13206), .CO(net_1351), .A(net_55), .B(net_42) );
NAND3_X2 inst_6678 ( .ZN(net_7746), .A2(net_7745), .A1(net_5896), .A3(net_4857) );
INV_X4 inst_17646 ( .A(net_3745), .ZN(net_662) );
INV_X4 inst_16451 ( .ZN(net_15858), .A(net_14593) );
CLKBUF_X2 inst_21942 ( .A(net_21813), .Z(net_21814) );
NAND2_X2 inst_9616 ( .ZN(net_10697), .A2(net_9979), .A1(net_5203) );
INV_X4 inst_12798 ( .ZN(net_17527), .A(net_17278) );
INV_X4 inst_16367 ( .A(net_1363), .ZN(net_1283) );
NAND2_X4 inst_7011 ( .A2(net_19130), .A1(net_19129), .ZN(net_17139) );
CLKBUF_X2 inst_22936 ( .A(net_21873), .Z(net_22808) );
NAND2_X4 inst_7201 ( .A1(net_20412), .ZN(net_9721), .A2(net_874) );
NAND2_X2 inst_11049 ( .A2(net_12262), .ZN(net_7791), .A1(net_4711) );
NAND2_X2 inst_9649 ( .ZN(net_10366), .A1(net_10365), .A2(net_10364) );
INV_X2 inst_19204 ( .A(net_4736), .ZN(net_3547) );
NAND2_X2 inst_9320 ( .ZN(net_12332), .A2(net_9069), .A1(net_5509) );
XNOR2_X2 inst_620 ( .B(net_16759), .ZN(net_478), .A(net_477) );
NAND3_X2 inst_6496 ( .ZN(net_10856), .A1(net_7748), .A2(net_6898), .A3(net_5825) );
NOR2_X4 inst_3118 ( .A1(net_20474), .ZN(net_6846), .A2(net_2879) );
AOI21_X2 inst_20659 ( .ZN(net_12990), .B2(net_12989), .B1(net_12283), .A(net_9636) );
NAND3_X2 inst_6401 ( .ZN(net_11982), .A1(net_7601), .A3(net_6820), .A2(net_5921) );
INV_X2 inst_18944 ( .A(net_6732), .ZN(net_5684) );
CLKBUF_X2 inst_22479 ( .A(net_22350), .Z(net_22351) );
NAND2_X4 inst_6869 ( .ZN(net_18328), .A2(net_18190), .A1(net_18165) );
INV_X4 inst_14597 ( .A(net_6725), .ZN(net_6241) );
INV_X4 inst_14514 ( .A(net_11729), .ZN(net_5979) );
CLKBUF_X2 inst_21818 ( .A(net_21689), .Z(net_21690) );
OAI21_X4 inst_1409 ( .A(net_20864), .B2(net_19972), .B1(net_19971), .ZN(net_18877) );
NAND2_X2 inst_10757 ( .ZN(net_8087), .A2(net_2724), .A1(net_1058) );
NAND2_X2 inst_11570 ( .ZN(net_2767), .A2(net_2642), .A1(net_1391) );
INV_X4 inst_13752 ( .A(net_9673), .ZN(net_7620) );
INV_X4 inst_15613 ( .ZN(net_8457), .A(net_4820) );
INV_X2 inst_19325 ( .ZN(net_2588), .A(net_2587) );
INV_X4 inst_13509 ( .ZN(net_12870), .A(net_9409) );
NOR2_X4 inst_2996 ( .ZN(net_9512), .A1(net_5909), .A2(net_1103) );
NOR2_X2 inst_5037 ( .ZN(net_1716), .A1(net_227), .A2(net_192) );
NAND2_X2 inst_10601 ( .A1(net_11292), .ZN(net_6621), .A2(net_5375) );
CLKBUF_X2 inst_22384 ( .A(net_22255), .Z(net_22256) );
INV_X4 inst_16261 ( .ZN(net_7890), .A(net_5570) );
INV_X2 inst_19539 ( .ZN(net_960), .A(net_959) );
INV_X4 inst_16762 ( .ZN(net_9098), .A(net_732) );
NAND2_X2 inst_11946 ( .ZN(net_1436), .A1(net_1435), .A2(net_1434) );
AOI21_X4 inst_20222 ( .B2(net_20732), .B1(net_20731), .ZN(net_14082), .A(net_14022) );
NAND2_X2 inst_9517 ( .ZN(net_11144), .A2(net_7423), .A1(net_6320) );
CLKBUF_X2 inst_22480 ( .A(net_22125), .Z(net_22352) );
INV_X2 inst_19629 ( .A(net_21231), .ZN(net_31) );
AOI21_X2 inst_20801 ( .ZN(net_10362), .B2(net_10361), .B1(net_5843), .A(net_5330) );
INV_X4 inst_14002 ( .ZN(net_10754), .A(net_6365) );
NAND2_X2 inst_8763 ( .A1(net_16260), .ZN(net_15883), .A2(net_15644) );
XOR2_X2 inst_4 ( .B(net_21191), .A(net_20217), .Z(net_18156) );
NOR2_X2 inst_3795 ( .ZN(net_10028), .A1(net_6909), .A2(net_6763) );
INV_X4 inst_18323 ( .A(net_20923), .ZN(net_20538) );
NOR2_X4 inst_3272 ( .ZN(net_4289), .A1(net_1842), .A2(net_1544) );
NAND2_X2 inst_9846 ( .ZN(net_9539), .A2(net_7510), .A1(net_5019) );
NAND2_X2 inst_9455 ( .A1(net_14365), .ZN(net_11507), .A2(net_9613) );
NAND2_X2 inst_10494 ( .A1(net_9972), .ZN(net_8299), .A2(net_4433) );
CLKBUF_X2 inst_22318 ( .A(net_22189), .Z(net_22190) );
INV_X4 inst_14232 ( .ZN(net_7364), .A(net_4878) );
OAI21_X2 inst_1866 ( .ZN(net_13755), .B2(net_13707), .A(net_12496), .B1(net_6809) );
INV_X4 inst_15230 ( .ZN(net_4920), .A(net_2851) );
NAND2_X2 inst_8795 ( .ZN(net_15712), .A2(net_15193), .A1(net_14933) );
AOI21_X4 inst_20108 ( .ZN(net_19059), .B1(net_16210), .B2(net_16168), .A(net_16143) );
OAI21_X2 inst_1878 ( .ZN(net_13667), .B2(net_13644), .B1(net_11645), .A(net_4352) );
INV_X2 inst_19569 ( .ZN(net_1925), .A(net_1195) );
NOR2_X2 inst_5136 ( .A2(net_2585), .ZN(net_341), .A1(net_156) );
INV_X4 inst_18240 ( .A(net_20888), .ZN(net_16347) );
NAND3_X2 inst_6016 ( .ZN(net_14392), .A2(net_14391), .A3(net_14342), .A1(net_13539) );
INV_X4 inst_16459 ( .A(net_5153), .ZN(net_4039) );
NAND2_X2 inst_10290 ( .A1(net_8741), .ZN(net_7928), .A2(net_6367) );
SDFF_X2 inst_765 ( .Q(net_20963), .SE(net_18847), .SI(net_18513), .D(net_579), .CK(net_22256) );
NAND2_X2 inst_10790 ( .A1(net_8190), .ZN(net_6287), .A2(net_5582) );
NAND2_X2 inst_9870 ( .ZN(net_9477), .A2(net_9476), .A1(net_5454) );
INV_X4 inst_17434 ( .ZN(net_8115), .A(net_761) );
NAND2_X2 inst_10664 ( .ZN(net_12248), .A2(net_7124), .A1(net_1103) );
INV_X4 inst_14247 ( .A(net_6459), .ZN(net_5761) );
NOR2_X2 inst_3422 ( .ZN(net_18923), .A2(net_15131), .A1(net_14040) );
INV_X4 inst_13266 ( .ZN(net_12610), .A(net_11467) );
NOR2_X2 inst_3832 ( .ZN(net_19407), .A1(net_9727), .A2(net_9053) );
NAND3_X2 inst_6618 ( .A2(net_14669), .ZN(net_9063), .A3(net_8965), .A1(net_8233) );
AND2_X4 inst_21256 ( .ZN(net_10756), .A1(net_6849), .A2(net_761) );
NOR2_X2 inst_4039 ( .ZN(net_9443), .A2(net_6056), .A1(net_809) );
NOR2_X4 inst_2967 ( .ZN(net_9356), .A1(net_4578), .A2(net_3904) );
INV_X4 inst_16681 ( .ZN(net_1949), .A(net_1752) );
INV_X4 inst_13279 ( .ZN(net_12439), .A(net_11170) );
CLKBUF_X2 inst_22353 ( .A(net_22150), .Z(net_22225) );
NAND3_X2 inst_5674 ( .ZN(net_20694), .A3(net_19838), .A1(net_19837), .A2(net_12751) );
NAND2_X2 inst_9029 ( .ZN(net_14074), .A1(net_13348), .A2(net_11899) );
INV_X4 inst_14873 ( .A(net_4666), .ZN(net_3691) );
SDFF_X2 inst_699 ( .Q(net_20857), .SE(net_18863), .SI(net_18846), .D(net_620), .CK(net_22040) );
NAND2_X2 inst_8377 ( .ZN(net_17352), .A2(net_17350), .A1(net_15959) );
AOI21_X2 inst_20456 ( .ZN(net_15047), .B1(net_15046), .B2(net_12971), .A(net_10994) );
NAND2_X2 inst_9921 ( .A1(net_10610), .ZN(net_9271), .A2(net_4873) );
INV_X4 inst_18025 ( .A(net_21050), .ZN(net_413) );
NAND2_X2 inst_9514 ( .ZN(net_11147), .A2(net_10840), .A1(net_2360) );
AOI21_X2 inst_20892 ( .ZN(net_7785), .B2(net_6366), .A(net_6347), .B1(net_1670) );
AOI21_X4 inst_20176 ( .B1(net_19802), .ZN(net_15500), .B2(net_15499), .A(net_12415) );
INV_X4 inst_13823 ( .ZN(net_11006), .A(net_9631) );
INV_X2 inst_18644 ( .ZN(net_9336), .A(net_9335) );
INV_X4 inst_14880 ( .ZN(net_6362), .A(net_2725) );
CLKBUF_X2 inst_22398 ( .A(net_21495), .Z(net_22270) );
INV_X2 inst_19592 ( .A(net_20897), .ZN(net_269) );
INV_X4 inst_13144 ( .ZN(net_15067), .A(net_14641) );
OAI211_X2 inst_2426 ( .ZN(net_15180), .C1(net_14751), .B(net_13813), .A(net_13177), .C2(net_13017) );
CLKBUF_X2 inst_21665 ( .A(net_21536), .Z(net_21537) );
INV_X4 inst_14211 ( .ZN(net_9509), .A(net_5901) );
NAND3_X2 inst_6377 ( .ZN(net_12039), .A1(net_12038), .A3(net_9817), .A2(net_6418) );
INV_X4 inst_14528 ( .ZN(net_7448), .A(net_6076) );
INV_X4 inst_18304 ( .A(net_20495), .ZN(net_20488) );
INV_X4 inst_18260 ( .A(net_19423), .ZN(net_19422) );
INV_X4 inst_17547 ( .A(net_14678), .ZN(net_14151) );
OAI21_X4 inst_1485 ( .ZN(net_19905), .A(net_12363), .B1(net_11019), .B2(net_7996) );
INV_X4 inst_17283 ( .ZN(net_4093), .A(net_1376) );
INV_X8 inst_12259 ( .ZN(net_4229), .A(net_1702) );
AOI21_X4 inst_20195 ( .ZN(net_19642), .B1(net_15119), .B2(net_13217), .A(net_13051) );
SDFF_X2 inst_750 ( .Q(net_20903), .SE(net_18859), .SI(net_18535), .D(net_725), .CK(net_21491) );
XNOR2_X2 inst_317 ( .B(net_21165), .A(net_17445), .ZN(net_17065) );
NAND2_X2 inst_10561 ( .ZN(net_8712), .A2(net_6853), .A1(net_4179) );
NAND2_X2 inst_8947 ( .ZN(net_19282), .A2(net_13241), .A1(net_750) );
XNOR2_X2 inst_278 ( .ZN(net_17173), .A(net_17168), .B(net_15798) );
NOR2_X2 inst_4429 ( .ZN(net_6059), .A2(net_4917), .A1(net_4916) );
AOI21_X2 inst_20277 ( .B1(net_20952), .ZN(net_16322), .B2(net_16062), .A(net_12132) );
XNOR2_X2 inst_467 ( .B(net_21199), .ZN(net_12873), .A(net_12872) );
AOI21_X2 inst_20293 ( .B1(net_20191), .B2(net_16368), .ZN(net_16160), .A(net_14853) );
INV_X4 inst_16117 ( .A(net_4025), .ZN(net_3459) );
NOR2_X2 inst_3677 ( .ZN(net_11434), .A2(net_9515), .A1(net_9400) );
NOR2_X2 inst_3456 ( .ZN(net_20173), .A2(net_13587), .A1(net_12651) );
INV_X4 inst_17370 ( .ZN(net_4374), .A(net_3861) );
NOR2_X4 inst_2963 ( .ZN(net_7860), .A2(net_4841), .A1(net_2585) );
NAND2_X2 inst_7923 ( .ZN(net_18450), .A2(net_18336), .A1(net_18282) );
NAND2_X2 inst_10535 ( .ZN(net_6811), .A2(net_6810), .A1(net_3847) );
OAI221_X2 inst_1329 ( .ZN(net_15845), .C2(net_14935), .B2(net_14361), .B1(net_14070), .A(net_12346), .C1(net_12208) );
OR2_X2 inst_1204 ( .ZN(net_3544), .A1(net_3543), .A2(net_2285) );
NAND2_X2 inst_8687 ( .ZN(net_16418), .A1(net_16348), .A2(net_16151) );
NOR2_X2 inst_4066 ( .ZN(net_7778), .A2(net_7777), .A1(net_1368) );
INV_X4 inst_17974 ( .A(net_20942), .ZN(net_246) );
NAND2_X4 inst_7669 ( .ZN(net_1096), .A2(net_879), .A1(net_234) );
INV_X4 inst_13568 ( .ZN(net_12788), .A(net_9134) );
INV_X4 inst_13158 ( .ZN(net_14869), .A(net_14324) );
NAND2_X2 inst_10162 ( .ZN(net_8255), .A2(net_8254), .A1(net_918) );
INV_X4 inst_17687 ( .ZN(net_10683), .A(net_1815) );
NAND2_X2 inst_11015 ( .ZN(net_12444), .A1(net_3814), .A2(net_2708) );
NAND2_X2 inst_11718 ( .A2(net_2846), .ZN(net_2262), .A1(net_1596) );
NOR3_X4 inst_2618 ( .ZN(net_19856), .A1(net_15082), .A3(net_14575), .A2(net_10542) );
INV_X4 inst_15065 ( .ZN(net_15561), .A(net_3296) );
NAND2_X2 inst_10952 ( .ZN(net_7781), .A2(net_5032), .A1(net_4795) );
NOR2_X2 inst_4950 ( .A1(net_20529), .ZN(net_2346), .A2(net_1664) );
INV_X4 inst_14726 ( .ZN(net_6874), .A(net_4012) );
NAND2_X2 inst_8853 ( .ZN(net_15381), .A1(net_14514), .A2(net_14162) );
NAND2_X2 inst_11443 ( .ZN(net_8492), .A1(net_5516), .A2(net_2973) );
NAND2_X2 inst_9241 ( .ZN(net_12691), .A2(net_12388), .A1(net_12374) );
INV_X2 inst_19053 ( .ZN(net_4733), .A(net_4732) );
CLKBUF_X2 inst_22431 ( .A(net_22302), .Z(net_22303) );
INV_X4 inst_17943 ( .A(net_21174), .ZN(net_16470) );
CLKBUF_X2 inst_22453 ( .A(net_21530), .Z(net_22325) );
INV_X4 inst_16916 ( .ZN(net_3750), .A(net_417) );
INV_X4 inst_14428 ( .A(net_11258), .ZN(net_5033) );
OAI21_X2 inst_1729 ( .A(net_15677), .ZN(net_15085), .B2(net_12897), .B1(net_8907) );
NAND2_X2 inst_8346 ( .A2(net_17651), .ZN(net_17481), .A1(net_17480) );
INV_X4 inst_13175 ( .ZN(net_14377), .A(net_13912) );
NAND3_X2 inst_6126 ( .ZN(net_13745), .A3(net_13744), .A1(net_10613), .A2(net_8342) );
NAND2_X4 inst_6996 ( .ZN(net_17554), .A1(net_16735), .A2(net_16581) );
CLKBUF_X2 inst_22939 ( .A(net_22810), .Z(net_22811) );
INV_X4 inst_13576 ( .ZN(net_9121), .A(net_6978) );
INV_X4 inst_15202 ( .ZN(net_9819), .A(net_2450) );
NOR2_X2 inst_4648 ( .ZN(net_5095), .A1(net_4401), .A2(net_2006) );
NAND2_X2 inst_10469 ( .A1(net_9109), .ZN(net_8879), .A2(net_6997) );
NAND2_X2 inst_10297 ( .A2(net_8393), .ZN(net_7898), .A1(net_3336) );
NAND2_X2 inst_11460 ( .A1(net_3331), .ZN(net_3207), .A2(net_3206) );
NAND2_X4 inst_7595 ( .ZN(net_3173), .A2(net_2590), .A1(net_420) );
XNOR2_X2 inst_165 ( .ZN(net_17848), .A(net_17672), .B(net_943) );
NOR2_X2 inst_3733 ( .A1(net_11468), .ZN(net_10866), .A2(net_10865) );
NAND4_X2 inst_5376 ( .A2(net_18992), .A1(net_18991), .ZN(net_15220), .A4(net_14013), .A3(net_11683) );
OR2_X2 inst_1176 ( .A2(net_11279), .A1(net_10515), .ZN(net_5580) );
INV_X4 inst_17102 ( .ZN(net_11018), .A(net_8220) );
INV_X4 inst_12537 ( .ZN(net_18374), .A(net_18373) );
NAND2_X2 inst_8159 ( .ZN(net_17986), .A1(net_17928), .A2(net_17884) );
INV_X4 inst_18127 ( .A(net_21177), .ZN(net_466) );
AOI21_X2 inst_20412 ( .ZN(net_20193), .B2(net_13572), .A(net_13534), .B1(net_9797) );
INV_X4 inst_12696 ( .ZN(net_17637), .A(net_17636) );
NAND4_X2 inst_5450 ( .ZN(net_20337), .A2(net_9149), .A1(net_7060), .A4(net_5074), .A3(net_3307) );
AOI21_X2 inst_20961 ( .B1(net_9131), .ZN(net_5328), .B2(net_5327), .A(net_3155) );
INV_X4 inst_15706 ( .ZN(net_1995), .A(net_1994) );
NAND2_X2 inst_11340 ( .ZN(net_3679), .A1(net_3678), .A2(net_2535) );
NOR2_X2 inst_4172 ( .ZN(net_8155), .A2(net_3557), .A1(net_809) );
INV_X4 inst_13388 ( .A(net_10740), .ZN(net_10739) );
NOR3_X4 inst_2605 ( .ZN(net_16199), .A1(net_16000), .A3(net_14454), .A2(net_4946) );
INV_X4 inst_14423 ( .A(net_6908), .ZN(net_5049) );
INV_X4 inst_14147 ( .ZN(net_7202), .A(net_6049) );
AOI22_X2 inst_20007 ( .ZN(net_19849), .B1(net_13873), .B2(net_12890), .A2(net_12847), .A1(net_3379) );
INV_X4 inst_13759 ( .ZN(net_10080), .A(net_7612) );
NAND2_X4 inst_7252 ( .ZN(net_11589), .A2(net_6740), .A1(net_2585) );
AOI21_X2 inst_20736 ( .A(net_13350), .ZN(net_11573), .B2(net_7413), .B1(net_4763) );
INV_X4 inst_13717 ( .ZN(net_11744), .A(net_7826) );
NOR3_X2 inst_2703 ( .A3(net_15804), .ZN(net_13923), .A2(net_13922), .A1(net_12018) );
INV_X4 inst_17464 ( .A(net_6524), .ZN(net_447) );
INV_X4 inst_13857 ( .ZN(net_13486), .A(net_7462) );
NAND2_X2 inst_9784 ( .ZN(net_15018), .A1(net_9421), .A2(net_7552) );
XNOR2_X2 inst_143 ( .B(net_19422), .ZN(net_18157), .A(net_18124) );
INV_X4 inst_15958 ( .ZN(net_2860), .A(net_1703) );
INV_X4 inst_16698 ( .ZN(net_5551), .A(net_1085) );
NAND4_X2 inst_5286 ( .ZN(net_15944), .A4(net_15196), .A1(net_15028), .A2(net_14707), .A3(net_10045) );
NAND3_X2 inst_6260 ( .ZN(net_19774), .A2(net_12994), .A1(net_9702), .A3(net_9413) );
NOR2_X2 inst_4272 ( .ZN(net_11042), .A1(net_6899), .A2(net_6130) );
INV_X4 inst_16403 ( .ZN(net_14227), .A(net_5415) );
INV_X4 inst_16878 ( .A(net_1022), .ZN(net_957) );
OAI21_X2 inst_2337 ( .ZN(net_4682), .A(net_4681), .B1(net_3234), .B2(net_2229) );
NOR2_X4 inst_3250 ( .ZN(net_2742), .A2(net_1362), .A1(net_629) );
INV_X4 inst_15052 ( .ZN(net_4385), .A(net_1916) );
NAND2_X2 inst_9357 ( .A1(net_13095), .ZN(net_12153), .A2(net_8807) );
OAI21_X2 inst_1778 ( .B2(net_20673), .B1(net_20672), .ZN(net_14671), .A(net_14022) );
INV_X2 inst_18991 ( .ZN(net_5087), .A(net_5086) );
INV_X4 inst_16158 ( .ZN(net_2140), .A(net_2045) );
NAND2_X1 inst_12132 ( .A1(net_21201), .ZN(net_19864), .A2(net_18170) );
NAND2_X2 inst_8091 ( .A1(net_18214), .ZN(net_18131), .A2(net_18092) );
OAI21_X2 inst_1736 ( .ZN(net_15069), .A(net_14687), .B1(net_13501), .B2(net_10468) );
SDFF_X2 inst_1040 ( .QN(net_21006), .D(net_1865), .SE(net_263), .CK(net_21874), .SI(x2971) );
NOR2_X2 inst_4027 ( .ZN(net_8010), .A2(net_6679), .A1(net_5094) );
INV_X4 inst_16648 ( .ZN(net_15312), .A(net_14788) );
INV_X4 inst_15218 ( .ZN(net_4373), .A(net_2881) );
NAND2_X2 inst_9158 ( .ZN(net_13384), .A1(net_13383), .A2(net_10438) );
NAND3_X2 inst_6009 ( .ZN(net_20396), .A3(net_12554), .A2(net_11616), .A1(net_10358) );
NOR2_X2 inst_5042 ( .A1(net_1328), .ZN(net_1089), .A2(net_1043) );
INV_X4 inst_17032 ( .ZN(net_1163), .A(net_222) );
INV_X4 inst_16218 ( .ZN(net_7610), .A(net_6601) );
INV_X2 inst_19645 ( .A(net_19444), .ZN(net_19442) );
NOR2_X4 inst_3146 ( .ZN(net_3621), .A1(net_3459), .A2(net_1939) );
NAND2_X2 inst_10246 ( .ZN(net_10194), .A2(net_6252), .A1(net_948) );
NAND2_X4 inst_7303 ( .A1(net_19202), .ZN(net_6820), .A2(net_1358) );
NAND2_X2 inst_11651 ( .ZN(net_2450), .A2(net_2449), .A1(net_921) );
CLKBUF_X2 inst_22011 ( .A(net_21882), .Z(net_21883) );
OAI21_X2 inst_2056 ( .ZN(net_10741), .B1(net_5867), .B2(net_4909), .A(net_1815) );
OAI21_X2 inst_2116 ( .ZN(net_10032), .A(net_10031), .B1(net_10030), .B2(net_7008) );
AOI21_X2 inst_20569 ( .ZN(net_19938), .B1(net_14164), .B2(net_10717), .A(net_1864) );
NOR2_X4 inst_2825 ( .ZN(net_18975), .A2(net_15983), .A1(net_15808) );
NOR2_X2 inst_5071 ( .A2(net_2123), .ZN(net_1567), .A1(net_170) );
INV_X4 inst_17135 ( .ZN(net_6131), .A(net_912) );
NOR2_X2 inst_4031 ( .A2(net_20779), .ZN(net_7980), .A1(net_7979) );
AND2_X2 inst_21303 ( .A2(net_9981), .ZN(net_9831), .A1(net_6297) );
INV_X2 inst_19262 ( .ZN(net_3141), .A(net_3140) );
INV_X4 inst_16607 ( .A(net_10914), .ZN(net_7901) );
INV_X4 inst_15370 ( .ZN(net_5786), .A(net_2571) );
NAND2_X2 inst_8135 ( .ZN(net_18035), .A1(net_18021), .A2(net_18000) );
XNOR2_X2 inst_346 ( .B(net_21123), .ZN(net_16942), .A(net_16562) );
NAND2_X2 inst_8755 ( .A1(net_16210), .ZN(net_15912), .A2(net_15511) );
NAND2_X2 inst_10711 ( .ZN(net_5985), .A1(net_5984), .A2(net_4557) );
NAND2_X2 inst_12058 ( .ZN(net_19426), .A1(net_889), .A2(net_322) );
AND4_X2 inst_21095 ( .ZN(net_14616), .A4(net_14312), .A1(net_13320), .A3(net_11799), .A2(net_11343) );
NAND3_X2 inst_6195 ( .ZN(net_13314), .A3(net_9873), .A1(net_9389), .A2(net_3526) );
CLKBUF_X2 inst_21819 ( .A(net_21690), .Z(net_21691) );
NAND2_X2 inst_9777 ( .ZN(net_11120), .A2(net_9813), .A1(net_154) );
NAND2_X2 inst_11347 ( .ZN(net_8440), .A2(net_3263), .A1(net_3063) );
INV_X4 inst_12972 ( .A(net_16515), .ZN(net_16514) );
NOR2_X2 inst_3929 ( .A1(net_13187), .ZN(net_8743), .A2(net_8045) );
NAND2_X2 inst_8856 ( .ZN(net_15361), .A1(net_15360), .A2(net_14409) );
INV_X8 inst_12312 ( .A(net_3297), .ZN(net_1477) );
NAND2_X2 inst_10506 ( .ZN(net_11556), .A2(net_6908), .A1(net_6861) );
NOR2_X2 inst_3852 ( .ZN(net_9526), .A1(net_9525), .A2(net_7573) );
CLKBUF_X2 inst_21603 ( .A(net_21474), .Z(net_21475) );
INV_X2 inst_18549 ( .ZN(net_10934), .A(net_10933) );
INV_X4 inst_15131 ( .ZN(net_13196), .A(net_7080) );
INV_X4 inst_14168 ( .ZN(net_9445), .A(net_6007) );
SDFF_X2 inst_1051 ( .QN(net_20983), .D(net_1855), .SE(net_263), .CK(net_22643), .SI(x3279) );
OAI211_X2 inst_2566 ( .ZN(net_9287), .B(net_8594), .A(net_2678), .C1(net_2517), .C2(net_1960) );
CLKBUF_X2 inst_21995 ( .A(net_21866), .Z(net_21867) );
INV_X2 inst_19024 ( .ZN(net_4933), .A(net_4932) );
NAND3_X2 inst_6102 ( .A3(net_20055), .A1(net_20054), .ZN(net_13906), .A2(net_9707) );
CLKBUF_X2 inst_21507 ( .A(net_21378), .Z(net_21379) );
INV_X2 inst_18690 ( .ZN(net_8606), .A(net_7178) );
INV_X4 inst_12901 ( .ZN(net_17254), .A(net_16783) );
NOR2_X2 inst_3603 ( .ZN(net_12464), .A1(net_9624), .A2(net_6715) );
NAND2_X2 inst_11076 ( .A2(net_12939), .A1(net_9313), .ZN(net_4476) );
NOR2_X4 inst_3043 ( .ZN(net_5073), .A1(net_2391), .A2(net_950) );
CLKBUF_X2 inst_22685 ( .A(net_22556), .Z(net_22557) );
NAND2_X2 inst_8063 ( .ZN(net_18222), .A2(net_18132), .A1(net_18115) );
AOI21_X2 inst_20448 ( .ZN(net_15095), .A(net_13070), .B2(net_12978), .B1(net_8347) );
INV_X4 inst_13665 ( .ZN(net_11863), .A(net_8098) );
NAND3_X2 inst_5752 ( .ZN(net_16004), .A1(net_15689), .A3(net_15195), .A2(net_14389) );
INV_X4 inst_14969 ( .ZN(net_3429), .A(net_3428) );
NAND2_X2 inst_10548 ( .ZN(net_13774), .A1(net_11541), .A2(net_6752) );
CLKBUF_X2 inst_22123 ( .A(net_21994), .Z(net_21995) );
INV_X4 inst_13781 ( .ZN(net_11104), .A(net_10582) );
NAND2_X2 inst_11360 ( .ZN(net_3613), .A2(net_3258), .A1(net_2576) );
XNOR2_X2 inst_573 ( .A(net_9235), .B(net_738), .ZN(net_623) );
NAND2_X2 inst_7736 ( .ZN(net_18812), .A2(net_18784), .A1(net_17737) );
INV_X4 inst_17735 ( .A(net_21238), .ZN(net_5415) );
INV_X4 inst_17123 ( .ZN(net_1921), .A(net_779) );
INV_X4 inst_17757 ( .A(net_890), .ZN(net_522) );
NAND2_X2 inst_9041 ( .ZN(net_14057), .A1(net_12881), .A2(net_12022) );
NAND2_X2 inst_8088 ( .ZN(net_20323), .A2(net_18107), .A1(net_17104) );
NAND4_X2 inst_5364 ( .A2(net_20049), .A1(net_20048), .ZN(net_15273), .A4(net_9046), .A3(net_3732) );
INV_X2 inst_18669 ( .ZN(net_9168), .A(net_9167) );
NOR2_X2 inst_4245 ( .A1(net_9421), .ZN(net_6510), .A2(net_6509) );
AND2_X4 inst_21172 ( .A1(net_12705), .ZN(net_12700), .A2(net_6796) );
INV_X4 inst_18169 ( .ZN(net_1097), .A(net_27) );
INV_X4 inst_17868 ( .ZN(net_169), .A(net_110) );
INV_X8 inst_12391 ( .A(net_20870), .ZN(net_258) );
NAND2_X2 inst_8978 ( .ZN(net_14508), .A1(net_14166), .A2(net_12841) );
CLKBUF_X2 inst_21372 ( .A(x7698), .Z(net_21244) );
CLKBUF_X2 inst_22750 ( .A(net_22621), .Z(net_22622) );
NOR2_X2 inst_3544 ( .ZN(net_13134), .A2(net_11268), .A1(net_1471) );
NAND2_X2 inst_10973 ( .A1(net_8877), .A2(net_7348), .ZN(net_4971) );
INV_X2 inst_18871 ( .ZN(net_10546), .A(net_6245) );
CLKBUF_X2 inst_22201 ( .A(net_22072), .Z(net_22073) );
CLKBUF_X2 inst_21464 ( .A(net_21335), .Z(net_21336) );
INV_X4 inst_17558 ( .ZN(net_9984), .A(net_401) );
NAND2_X2 inst_7970 ( .ZN(net_18361), .A2(net_18360), .A1(net_17297) );
INV_X4 inst_13607 ( .ZN(net_8464), .A(net_7108) );
INV_X2 inst_19678 ( .A(net_20512), .ZN(net_20511) );
INV_X4 inst_17404 ( .ZN(net_14153), .A(net_10216) );
CLKBUF_X2 inst_21451 ( .A(net_21322), .Z(net_21323) );
NAND2_X2 inst_9362 ( .ZN(net_12141), .A1(net_12140), .A2(net_9933) );
INV_X4 inst_18351 ( .A(net_20799), .ZN(net_20797) );
NAND3_X2 inst_6367 ( .ZN(net_12077), .A3(net_12076), .A1(net_7333), .A2(net_3785) );
INV_X2 inst_19265 ( .ZN(net_3106), .A(net_3105) );
CLKBUF_X2 inst_22276 ( .A(net_22147), .Z(net_22148) );
CLKBUF_X2 inst_22208 ( .A(net_22079), .Z(net_22080) );
INV_X2 inst_18656 ( .A(net_11017), .ZN(net_9213) );
INV_X4 inst_15876 ( .ZN(net_1792), .A(net_1791) );
NAND3_X4 inst_5553 ( .A3(net_20373), .A1(net_20372), .ZN(net_19165), .A2(net_5805) );
NAND2_X2 inst_11518 ( .ZN(net_3785), .A2(net_2147), .A1(net_547) );
NAND3_X2 inst_6111 ( .ZN(net_13889), .A3(net_13888), .A2(net_13442), .A1(net_8292) );
NOR2_X2 inst_3522 ( .ZN(net_18962), .A1(net_11579), .A2(net_8757) );
INV_X4 inst_15795 ( .ZN(net_4247), .A(net_2836) );
NAND3_X2 inst_6306 ( .ZN(net_12783), .A2(net_12782), .A3(net_12254), .A1(net_8725) );
INV_X4 inst_14119 ( .ZN(net_7544), .A(net_6140) );
INV_X2 inst_18475 ( .ZN(net_12634), .A(net_12633) );
OAI21_X2 inst_1758 ( .ZN(net_14786), .B2(net_13270), .B1(net_6833), .A(net_1471) );
OR2_X2 inst_1142 ( .A1(net_11468), .ZN(net_11119), .A2(net_11118) );
NAND3_X2 inst_6280 ( .ZN(net_12901), .A2(net_12900), .A3(net_12899), .A1(net_9895) );
CLKBUF_X2 inst_21545 ( .A(net_21253), .Z(net_21417) );
NOR2_X2 inst_3816 ( .ZN(net_9803), .A2(net_9688), .A1(net_8958) );
AOI21_X2 inst_20348 ( .ZN(net_15751), .B2(net_15043), .B1(net_4285), .A(net_864) );
NAND2_X2 inst_11138 ( .ZN(net_8261), .A1(net_4252), .A2(net_3087) );
INV_X4 inst_14914 ( .ZN(net_6119), .A(net_4870) );
INV_X4 inst_15979 ( .ZN(net_2213), .A(net_1680) );
INV_X2 inst_19335 ( .ZN(net_3516), .A(net_2483) );
INV_X4 inst_14772 ( .ZN(net_6643), .A(net_5451) );
NAND4_X2 inst_5418 ( .A4(net_20277), .A2(net_19463), .ZN(net_19343), .A3(net_11713), .A1(net_11712) );
INV_X2 inst_19152 ( .A(net_4051), .ZN(net_4050) );
OAI21_X4 inst_1381 ( .A(net_20848), .ZN(net_19162), .B2(net_18981), .B1(net_18980) );
AOI21_X2 inst_20431 ( .ZN(net_15182), .B2(net_13964), .B1(net_12102), .A(net_1052) );
INV_X4 inst_15527 ( .ZN(net_13940), .A(net_12006) );
XNOR2_X2 inst_643 ( .B(net_17036), .ZN(net_16267), .A(net_430) );
AOI21_X4 inst_20109 ( .B1(net_19380), .ZN(net_18938), .B2(net_16041), .A(net_15964) );
INV_X4 inst_12471 ( .ZN(net_18765), .A(net_18764) );
INV_X2 inst_19701 ( .A(net_20564), .ZN(net_20563) );
INV_X4 inst_13726 ( .ZN(net_10179), .A(net_7798) );
NAND2_X2 inst_9430 ( .ZN(net_11608), .A1(net_11607), .A2(net_11606) );
NAND2_X2 inst_10745 ( .ZN(net_12243), .A1(net_8874), .A2(net_5713) );
NAND2_X2 inst_7763 ( .ZN(net_18750), .A2(net_18722), .A1(net_18698) );
NAND2_X2 inst_12117 ( .ZN(net_217), .A1(net_203), .A2(net_202) );
AOI22_X2 inst_19983 ( .ZN(net_15371), .A1(net_15370), .B1(net_15369), .A2(net_13884), .B2(net_9960) );
INV_X8 inst_12220 ( .ZN(net_8250), .A(net_5179) );
NOR2_X2 inst_4961 ( .A2(net_2978), .ZN(net_1616), .A1(net_112) );
AOI21_X2 inst_20548 ( .ZN(net_14371), .B2(net_12000), .B1(net_8968), .A(net_253) );
NAND2_X2 inst_8588 ( .A1(net_20659), .A2(net_19444), .ZN(net_16712) );
CLKBUF_X2 inst_22309 ( .A(net_22180), .Z(net_22181) );
NAND3_X2 inst_6466 ( .ZN(net_11360), .A3(net_11359), .A1(net_9118), .A2(net_9041) );
MUX2_X2 inst_12165 ( .Z(net_19804), .B(net_11908), .S(net_11907), .A(net_11839) );
NAND2_X2 inst_8581 ( .A2(net_16729), .ZN(net_16722), .A1(net_16721) );
NAND4_X2 inst_5447 ( .A3(net_20642), .ZN(net_13611), .A1(net_13610), .A2(net_13431), .A4(net_9561) );
NAND3_X2 inst_6371 ( .ZN(net_12062), .A1(net_12061), .A2(net_11764), .A3(net_10525) );
INV_X4 inst_17538 ( .ZN(net_1158), .A(net_302) );
NOR2_X2 inst_4146 ( .A1(net_9325), .ZN(net_6910), .A2(net_5069) );
INV_X4 inst_12526 ( .ZN(net_18436), .A(net_18435) );
INV_X4 inst_17220 ( .A(net_1662), .ZN(net_691) );
INV_X4 inst_12959 ( .ZN(net_16922), .A(net_16742) );
CLKBUF_X2 inst_21555 ( .A(net_21362), .Z(net_21427) );
OAI21_X2 inst_1997 ( .ZN(net_11867), .B1(net_11866), .B2(net_11865), .A(net_8362) );
NAND2_X4 inst_6971 ( .ZN(net_17421), .A1(net_16968), .A2(net_16809) );
INV_X4 inst_12669 ( .ZN(net_17785), .A(net_17784) );
OAI21_X2 inst_2297 ( .ZN(net_6435), .A(net_6434), .B1(net_6433), .B2(net_6432) );
NOR2_X2 inst_3736 ( .ZN(net_10721), .A1(net_10720), .A2(net_8540) );
NOR2_X2 inst_3341 ( .ZN(net_19626), .A1(net_18539), .A2(net_16703) );
NAND2_X2 inst_8500 ( .ZN(net_17075), .A1(net_16609), .A2(net_16473) );
AOI22_X2 inst_20044 ( .B1(net_6669), .ZN(net_6380), .B2(net_6379), .A2(net_2721), .A1(net_1790) );
INV_X4 inst_13411 ( .ZN(net_10331), .A(net_10330) );
NAND3_X2 inst_6374 ( .A1(net_16009), .A3(net_13747), .ZN(net_12046), .A2(net_11629) );
INV_X4 inst_15296 ( .A(net_3879), .ZN(net_2708) );
INV_X4 inst_14913 ( .A(net_4870), .ZN(net_3572) );
OAI211_X2 inst_2508 ( .ZN(net_12506), .A(net_12505), .C1(net_12504), .C2(net_6538), .B(net_4693) );
NAND2_X2 inst_10207 ( .ZN(net_10264), .A1(net_9917), .A2(net_3421) );
INV_X4 inst_14642 ( .A(net_5706), .ZN(net_4376) );
SDFF_X2 inst_773 ( .Q(net_20971), .SE(net_18864), .SI(net_18475), .D(net_11885), .CK(net_22739) );
NAND2_X2 inst_10776 ( .A1(net_20546), .A2(net_7146), .ZN(net_7014) );
INV_X4 inst_15642 ( .ZN(net_9024), .A(net_2120) );
INV_X4 inst_13091 ( .ZN(net_15968), .A(net_15846) );
NAND2_X2 inst_10074 ( .A1(net_9909), .ZN(net_8652), .A2(net_8651) );
NOR2_X2 inst_3620 ( .ZN(net_12338), .A1(net_12337), .A2(net_9338) );
INV_X4 inst_14134 ( .A(net_7957), .ZN(net_6103) );
INV_X4 inst_14763 ( .ZN(net_10361), .A(net_4057) );
NAND2_X2 inst_9798 ( .ZN(net_11683), .A2(net_9774), .A1(net_8020) );
XNOR2_X2 inst_260 ( .A(net_20789), .ZN(net_17263), .B(net_17262) );
NAND2_X2 inst_11277 ( .ZN(net_12431), .A2(net_3872), .A1(net_405) );
NAND2_X2 inst_9371 ( .A1(net_18025), .ZN(net_12083), .A2(net_8999) );
NAND2_X2 inst_11597 ( .A1(net_8278), .ZN(net_2670), .A2(net_2669) );
NOR2_X2 inst_4973 ( .ZN(net_3088), .A1(net_1376), .A2(net_1055) );
NOR2_X2 inst_4139 ( .ZN(net_19895), .A2(net_6875), .A1(net_5067) );
INV_X2 inst_19284 ( .A(net_4125), .ZN(net_2907) );
NAND3_X2 inst_6762 ( .A1(net_8865), .ZN(net_5395), .A2(net_3804), .A3(net_2028) );
CLKBUF_X2 inst_22100 ( .A(net_21971), .Z(net_21972) );
NOR2_X2 inst_4611 ( .ZN(net_6574), .A1(net_4874), .A2(net_1544) );
INV_X4 inst_13839 ( .ZN(net_11055), .A(net_7484) );
NAND2_X2 inst_10725 ( .A1(net_6097), .ZN(net_5868), .A2(net_3511) );
NOR2_X2 inst_4567 ( .A1(net_7597), .ZN(net_4570), .A2(net_3882) );
NOR2_X2 inst_3889 ( .ZN(net_9243), .A2(net_5965), .A1(net_4220) );
INV_X4 inst_17093 ( .ZN(net_11460), .A(net_6668) );
CLKBUF_X2 inst_21679 ( .A(net_21511), .Z(net_21551) );
AND2_X4 inst_21164 ( .ZN(net_20203), .A1(net_15356), .A2(net_13578) );
INV_X4 inst_16746 ( .ZN(net_10252), .A(net_816) );
NAND2_X2 inst_9880 ( .A1(net_10233), .ZN(net_9447), .A2(net_8632) );
NAND2_X2 inst_8739 ( .ZN(net_19933), .A2(net_15748), .A1(net_14899) );
XNOR2_X2 inst_516 ( .ZN(net_5787), .B(net_5786), .A(net_1900) );
AOI21_X2 inst_20376 ( .ZN(net_15590), .B2(net_14258), .A(net_11416), .B1(net_872) );
INV_X4 inst_18196 ( .A(net_20976), .ZN(net_560) );
INV_X8 inst_12243 ( .ZN(net_4833), .A(net_4242) );
OAI21_X2 inst_2258 ( .ZN(net_7236), .B2(net_6634), .A(net_5482), .B1(net_3926) );
AOI21_X2 inst_20512 ( .ZN(net_14613), .B1(net_14612), .B2(net_12014), .A(net_11571) );
INV_X4 inst_13986 ( .ZN(net_7810), .A(net_5352) );
XNOR2_X2 inst_190 ( .B(net_21121), .ZN(net_17684), .A(net_17683) );
INV_X4 inst_16174 ( .ZN(net_16076), .A(net_15214) );
NAND2_X2 inst_9602 ( .A1(net_15450), .ZN(net_10752), .A2(net_8491) );
AOI21_X2 inst_20516 ( .ZN(net_14594), .B1(net_14593), .A(net_13250), .B2(net_6424) );
NOR2_X2 inst_4873 ( .ZN(net_2220), .A1(net_2219), .A2(net_2218) );
INV_X4 inst_13484 ( .ZN(net_11444), .A(net_10155) );
NAND2_X2 inst_9932 ( .ZN(net_9155), .A2(net_7110), .A1(net_3201) );
CLKBUF_X2 inst_22584 ( .A(net_22455), .Z(net_22456) );
NAND3_X2 inst_6424 ( .A3(net_12099), .ZN(net_11939), .A2(net_11379), .A1(net_7655) );
OAI21_X2 inst_2062 ( .ZN(net_10694), .B2(net_6887), .B1(net_6818), .A(net_333) );
AOI21_X4 inst_20217 ( .B1(net_18893), .ZN(net_14196), .B2(net_14195), .A(net_7942) );
INV_X4 inst_15442 ( .ZN(net_4502), .A(net_573) );
OAI21_X2 inst_2350 ( .ZN(net_3723), .B2(net_3654), .A(net_3206), .B1(net_2840) );
INV_X4 inst_15168 ( .ZN(net_5076), .A(net_4226) );
AOI21_X2 inst_20439 ( .ZN(net_15138), .B2(net_13327), .B1(net_10945), .A(net_8280) );
INV_X4 inst_17471 ( .A(net_6002), .ZN(net_5374) );
INV_X4 inst_15363 ( .A(net_4581), .ZN(net_4377) );
AOI21_X4 inst_20246 ( .ZN(net_9895), .B1(net_9894), .B2(net_6695), .A(net_6047) );
AND3_X4 inst_21127 ( .ZN(net_11722), .A2(net_11721), .A3(net_11720), .A1(net_9488) );
AOI21_X4 inst_20229 ( .ZN(net_19223), .B2(net_11059), .A(net_10678), .B1(net_10216) );
NAND2_X2 inst_11911 ( .A2(net_19027), .ZN(net_3057), .A1(net_2283) );
NOR2_X2 inst_3435 ( .ZN(net_15267), .A1(net_14198), .A2(net_13047) );
NAND2_X4 inst_6934 ( .A2(net_19044), .A1(net_19043), .ZN(net_17627) );
AOI21_X4 inst_20152 ( .B1(net_19912), .ZN(net_15793), .B2(net_15501), .A(net_12886) );
SDFF_X2 inst_829 ( .Q(net_21162), .SI(net_17540), .SE(net_125), .CK(net_21253), .D(x5244) );
INV_X4 inst_15697 ( .ZN(net_3409), .A(net_2017) );
XNOR2_X2 inst_197 ( .B(net_21169), .A(net_17673), .ZN(net_17672) );
NAND2_X4 inst_7277 ( .ZN(net_7441), .A2(net_6604), .A1(net_5945) );
NOR2_X2 inst_4702 ( .A1(net_20859), .ZN(net_4130), .A2(net_2217) );
INV_X4 inst_17628 ( .ZN(net_3309), .A(net_293) );
NAND2_X2 inst_10129 ( .ZN(net_8349), .A2(net_8348), .A1(net_7021) );
INV_X4 inst_14866 ( .ZN(net_4729), .A(net_3873) );
CLKBUF_X2 inst_21524 ( .A(net_21395), .Z(net_21396) );
INV_X4 inst_12830 ( .ZN(net_17140), .A(net_17139) );
INV_X4 inst_17933 ( .A(net_21134), .ZN(net_675) );
NAND2_X2 inst_11155 ( .ZN(net_5336), .A1(net_5008), .A2(net_3609) );
NAND2_X2 inst_8558 ( .A1(net_21203), .ZN(net_16751), .A2(net_16750) );
XNOR2_X2 inst_150 ( .ZN(net_18008), .A(net_17948), .B(net_17598) );
NAND3_X2 inst_6743 ( .ZN(net_6401), .A2(net_6400), .A3(net_6399), .A1(net_3699) );
NAND4_X2 inst_5358 ( .ZN(net_15322), .A2(net_13717), .A4(net_9951), .A1(net_9557), .A3(net_6727) );
NOR2_X2 inst_4540 ( .A1(net_7661), .ZN(net_5062), .A2(net_2126) );
SDFF_X2 inst_887 ( .Q(net_21127), .SI(net_16878), .SE(net_125), .CK(net_22224), .D(x4139) );
INV_X2 inst_18561 ( .ZN(net_10797), .A(net_10796) );
INV_X4 inst_16016 ( .ZN(net_2795), .A(net_1651) );
NAND4_X4 inst_5175 ( .A4(net_19064), .A1(net_19063), .ZN(net_16911), .A3(net_14954), .A2(net_10719) );
NAND2_X2 inst_8036 ( .ZN(net_18257), .A2(net_18256), .A1(net_17743) );
INV_X4 inst_17495 ( .ZN(net_14791), .A(net_10683) );
INV_X4 inst_15630 ( .ZN(net_9762), .A(net_8952) );
NAND2_X2 inst_8547 ( .A1(net_21188), .A2(net_16965), .ZN(net_16797) );
INV_X4 inst_13647 ( .ZN(net_13934), .A(net_8158) );
NOR2_X2 inst_4316 ( .A1(net_11550), .ZN(net_5888), .A2(net_5887) );
OAI21_X2 inst_2357 ( .A(net_7703), .B2(net_3393), .ZN(net_2958), .B1(net_2957) );
INV_X4 inst_13911 ( .ZN(net_8847), .A(net_6970) );
NAND3_X2 inst_6541 ( .ZN(net_10571), .A2(net_10442), .A1(net_7978), .A3(net_3806) );
INV_X4 inst_18180 ( .A(net_21004), .ZN(net_2041) );
INV_X8 inst_12248 ( .A(net_3791), .ZN(net_3512) );
OAI21_X2 inst_1961 ( .ZN(net_12490), .B2(net_10361), .A(net_9803), .B1(net_8667) );
INV_X4 inst_14343 ( .ZN(net_8122), .A(net_5357) );
NAND3_X2 inst_5799 ( .ZN(net_15717), .A3(net_15055), .A2(net_10863), .A1(net_3154) );
NAND3_X2 inst_5954 ( .ZN(net_14860), .A1(net_14089), .A3(net_13919), .A2(net_13617) );
DFF_X1 inst_19834 ( .D(net_18871), .CK(net_21990), .Q(x1005) );
SDFF_X2 inst_1010 ( .QN(net_20976), .D(net_560), .SE(net_253), .CK(net_22659), .SI(x3354) );
NAND2_X2 inst_7934 ( .ZN(net_18434), .A2(net_18320), .A1(net_18272) );
INV_X4 inst_14939 ( .ZN(net_11841), .A(net_3533) );
AOI21_X2 inst_20949 ( .ZN(net_5855), .B2(net_4580), .A(net_3638), .B1(net_1016) );
INV_X4 inst_14979 ( .ZN(net_8472), .A(net_3415) );
SDFF_X2 inst_867 ( .Q(net_21131), .D(net_17095), .SE(net_263), .CK(net_21398), .SI(x3951) );
INV_X4 inst_14179 ( .ZN(net_19984), .A(net_7832) );
INV_X4 inst_18132 ( .A(net_20906), .ZN(net_117) );
NOR2_X2 inst_3568 ( .ZN(net_12790), .A2(net_11333), .A1(net_8797) );
NAND3_X2 inst_6202 ( .ZN(net_13303), .A3(net_9865), .A1(net_7003), .A2(net_3245) );
AOI21_X2 inst_20809 ( .ZN(net_10184), .A(net_10183), .B2(net_5990), .B1(net_4191) );
INV_X4 inst_16400 ( .ZN(net_5173), .A(net_1262) );
AND2_X4 inst_21214 ( .ZN(net_20119), .A2(net_6348), .A1(net_242) );
INV_X2 inst_18544 ( .ZN(net_10982), .A(net_10981) );
NAND2_X2 inst_10760 ( .A1(net_6604), .ZN(net_6061), .A2(net_4814) );
NAND2_X2 inst_8963 ( .ZN(net_14685), .A1(net_14684), .A2(net_13314) );
INV_X4 inst_15449 ( .ZN(net_2736), .A(net_1443) );
INV_X8 inst_12364 ( .A(net_20875), .ZN(net_765) );
NAND2_X2 inst_9342 ( .ZN(net_12210), .A2(net_10403), .A1(net_1902) );
NOR2_X2 inst_4158 ( .ZN(net_6890), .A1(net_6889), .A2(net_6888) );
NAND2_X2 inst_11481 ( .ZN(net_5584), .A2(net_3092), .A1(net_703) );
OAI21_X2 inst_1643 ( .B2(net_19542), .B1(net_19541), .ZN(net_15946), .A(net_15027) );
NOR2_X2 inst_4660 ( .ZN(net_4058), .A2(net_2165), .A1(net_154) );
INV_X4 inst_14537 ( .ZN(net_5850), .A(net_4654) );
OAI21_X2 inst_2120 ( .A(net_10714), .ZN(net_10021), .B2(net_7960), .B1(net_5778) );
NOR3_X2 inst_2678 ( .ZN(net_14665), .A2(net_13702), .A1(net_13436), .A3(net_9993) );
NAND2_X2 inst_9196 ( .ZN(net_13094), .A1(net_13093), .A2(net_11242) );
INV_X4 inst_16898 ( .ZN(net_5537), .A(net_2273) );
INV_X4 inst_15079 ( .A(net_11861), .ZN(net_7725) );
NOR3_X4 inst_2613 ( .ZN(net_19716), .A3(net_15169), .A1(net_15073), .A2(net_14284) );
INV_X4 inst_15003 ( .A(net_3478), .ZN(net_3388) );
CLKBUF_X2 inst_22941 ( .A(net_22413), .Z(net_22813) );
NAND2_X2 inst_10577 ( .A1(net_11770), .ZN(net_6686), .A2(net_3971) );
NAND2_X4 inst_7143 ( .ZN(net_12833), .A1(net_9285), .A2(net_7394) );
INV_X8 inst_12239 ( .ZN(net_4396), .A(net_1952) );
NOR2_X2 inst_3866 ( .ZN(net_10893), .A2(net_9467), .A1(net_9378) );
CLKBUF_X2 inst_22673 ( .A(net_22102), .Z(net_22545) );
INV_X2 inst_19586 ( .ZN(net_939), .A(net_274) );
AOI21_X2 inst_20562 ( .ZN(net_14252), .B2(net_12420), .A(net_10683), .B1(net_5883) );
NAND2_X2 inst_10460 ( .ZN(net_7017), .A1(net_6732), .A2(net_2347) );
AOI21_X2 inst_20816 ( .B2(net_11224), .ZN(net_10047), .A(net_8556), .B1(net_7714) );
NAND2_X2 inst_8186 ( .ZN(net_17950), .A2(net_17816), .A1(net_17753) );
NAND2_X2 inst_7976 ( .ZN(net_18348), .A2(net_18243), .A1(net_17384) );
INV_X4 inst_17082 ( .A(net_5517), .ZN(net_3293) );
NOR2_X2 inst_4371 ( .A2(net_9322), .ZN(net_6734), .A1(net_4047) );
NAND4_X2 inst_5253 ( .ZN(net_18079), .A2(net_18059), .A1(net_18052), .A4(net_16067), .A3(net_15792) );
AOI21_X2 inst_20441 ( .B1(net_15186), .ZN(net_15124), .B2(net_13222), .A(net_12127) );
INV_X4 inst_17180 ( .ZN(net_4020), .A(net_3491) );
OAI21_X2 inst_1649 ( .A(net_16187), .ZN(net_15888), .B2(net_15321), .B1(net_14299) );
NAND2_X2 inst_7756 ( .ZN(net_18785), .A1(net_18743), .A2(net_18717) );
INV_X4 inst_12921 ( .ZN(net_17029), .A(net_16662) );
INV_X4 inst_13594 ( .ZN(net_8778), .A(net_8777) );
NAND3_X2 inst_5815 ( .ZN(net_15642), .A2(net_14423), .A3(net_13275), .A1(net_9424) );
NAND3_X2 inst_5873 ( .A3(net_19723), .A1(net_19722), .ZN(net_15306), .A2(net_11239) );
CLKBUF_X2 inst_22759 ( .A(net_21476), .Z(net_22631) );
INV_X2 inst_18557 ( .ZN(net_10881), .A(net_10880) );
NAND2_X2 inst_8697 ( .ZN(net_16344), .A1(net_16259), .A2(net_16186) );
XNOR2_X2 inst_669 ( .A(net_21170), .B(net_21138), .ZN(net_5236) );
NAND2_X2 inst_9214 ( .ZN(net_13039), .A2(net_11356), .A1(net_3725) );
AND2_X2 inst_21321 ( .A2(net_8467), .ZN(net_6791), .A1(net_6790) );
NAND2_X2 inst_10024 ( .A1(net_9658), .A2(net_9099), .ZN(net_8761) );
INV_X4 inst_16092 ( .ZN(net_3697), .A(net_1808) );
NAND2_X2 inst_8988 ( .ZN(net_14471), .A1(net_14395), .A2(net_12905) );
CLKBUF_X2 inst_21487 ( .A(net_21358), .Z(net_21359) );
INV_X4 inst_14633 ( .A(net_11893), .ZN(net_4386) );
INV_X4 inst_14530 ( .ZN(net_6021), .A(net_4729) );
AOI21_X2 inst_20980 ( .ZN(net_3209), .B2(net_3208), .A(net_2063), .B1(net_60) );
INV_X4 inst_17817 ( .ZN(net_171), .A(net_130) );
NAND2_X2 inst_10532 ( .ZN(net_6816), .A2(net_6815), .A1(net_4438) );
NAND2_X2 inst_8236 ( .A2(net_17754), .ZN(net_17751), .A1(net_17653) );
INV_X4 inst_18056 ( .A(net_21070), .ZN(net_644) );
INV_X4 inst_17798 ( .A(net_874), .ZN(net_194) );
AND2_X2 inst_21341 ( .ZN(net_8526), .A2(net_2891), .A1(net_2634) );
NOR2_X2 inst_4897 ( .A1(net_3984), .ZN(net_2019), .A2(net_1793) );
NAND2_X4 inst_7603 ( .ZN(net_3196), .A1(net_774), .A2(net_187) );
AOI21_X4 inst_20097 ( .B2(net_20936), .ZN(net_19058), .B1(net_16272), .A(net_13765) );
OAI21_X2 inst_1844 ( .ZN(net_19540), .B2(net_11299), .B1(net_11147), .A(net_1744) );
OAI21_X2 inst_1913 ( .A(net_20897), .ZN(net_19819), .B1(net_19407), .B2(net_12532) );
NAND4_X4 inst_5209 ( .ZN(net_16526), .A1(net_16239), .A4(net_16136), .A2(net_15762), .A3(net_10826) );
OAI21_X2 inst_1990 ( .ZN(net_12026), .A(net_12025), .B1(net_9579), .B2(net_7671) );
NAND3_X2 inst_5700 ( .ZN(net_16224), .A1(net_16026), .A3(net_15787), .A2(net_15638) );
XOR2_X2 inst_36 ( .A(net_17036), .Z(net_669), .B(net_668) );
INV_X4 inst_12770 ( .A(net_17747), .ZN(net_17336) );
INV_X4 inst_14658 ( .ZN(net_6958), .A(net_4360) );
INV_X4 inst_13686 ( .ZN(net_11970), .A(net_7966) );
NAND2_X2 inst_9039 ( .A1(net_14460), .ZN(net_14059), .A2(net_11840) );
INV_X2 inst_19242 ( .ZN(net_3288), .A(net_2439) );
AND2_X2 inst_21319 ( .ZN(net_7024), .A1(net_7023), .A2(net_6430) );
NAND2_X2 inst_9652 ( .ZN(net_10352), .A2(net_10351), .A1(net_6235) );
INV_X4 inst_15175 ( .A(net_4132), .ZN(net_3006) );
INV_X2 inst_18564 ( .ZN(net_20754), .A(net_12372) );
INV_X4 inst_13040 ( .ZN(net_16614), .A(net_16562) );
AOI21_X2 inst_20313 ( .ZN(net_15977), .B1(net_15976), .B2(net_15594), .A(net_6724) );
INV_X4 inst_18011 ( .A(net_20855), .ZN(net_598) );
INV_X4 inst_16663 ( .A(net_3990), .ZN(net_3381) );
NAND2_X2 inst_10721 ( .ZN(net_19173), .A1(net_10819), .A2(net_3488) );
NAND2_X2 inst_7998 ( .ZN(net_18316), .A2(net_18315), .A1(net_17867) );
INV_X2 inst_19075 ( .ZN(net_4605), .A(net_4604) );
INV_X2 inst_19609 ( .A(net_21215), .ZN(net_52) );
NAND2_X2 inst_7954 ( .ZN(net_18397), .A2(net_18357), .A1(net_17401) );
INV_X4 inst_13284 ( .ZN(net_14188), .A(net_12681) );
NOR2_X4 inst_3067 ( .A2(net_7096), .ZN(net_5982), .A1(net_4820) );
INV_X4 inst_13023 ( .A(net_16778), .ZN(net_16757) );
INV_X4 inst_14456 ( .ZN(net_8163), .A(net_4948) );
NAND2_X2 inst_9877 ( .ZN(net_9453), .A1(net_9349), .A2(net_7415) );
CLKBUF_X2 inst_21799 ( .A(net_21670), .Z(net_21671) );
INV_X4 inst_17579 ( .A(net_10676), .ZN(net_4995) );
NAND2_X2 inst_9142 ( .A1(net_13871), .ZN(net_13414), .A2(net_10500) );
INV_X4 inst_13737 ( .ZN(net_11406), .A(net_7647) );
AOI21_X2 inst_20596 ( .ZN(net_13900), .B2(net_11371), .A(net_5096), .B1(net_4113) );
INV_X4 inst_17572 ( .A(net_612), .ZN(net_348) );
AND2_X2 inst_21353 ( .ZN(net_2152), .A1(net_1280), .A2(net_1174) );
NAND2_X2 inst_10058 ( .A1(net_11907), .ZN(net_8686), .A2(net_6767) );
NAND4_X2 inst_5307 ( .A2(net_20723), .A1(net_20722), .ZN(net_20416), .A4(net_13048), .A3(net_7270) );
INV_X4 inst_13188 ( .ZN(net_14219), .A(net_13615) );
XNOR2_X2 inst_676 ( .ZN(net_18871), .B(net_16967), .A(net_9002) );
INV_X4 inst_17183 ( .A(net_879), .ZN(net_780) );
NAND2_X2 inst_9755 ( .A1(net_10947), .ZN(net_10019), .A2(net_6836) );
INV_X4 inst_16642 ( .ZN(net_11270), .A(net_5162) );
INV_X4 inst_15930 ( .ZN(net_9023), .A(net_7812) );
INV_X2 inst_18660 ( .ZN(net_9198), .A(net_6213) );
NOR2_X2 inst_4222 ( .ZN(net_11492), .A1(net_6626), .A2(net_6421) );
NAND3_X2 inst_6669 ( .A3(net_14465), .A2(net_14046), .A1(net_8397), .ZN(net_7775) );
NOR2_X2 inst_4859 ( .ZN(net_4170), .A1(net_2264), .A2(net_1188) );
INV_X4 inst_12588 ( .A(net_18192), .ZN(net_18119) );
NAND2_X2 inst_10193 ( .ZN(net_13265), .A2(net_7892), .A1(net_6161) );
OAI21_X2 inst_2255 ( .ZN(net_7266), .B2(net_4006), .B1(net_2261), .A(net_365) );
NOR2_X2 inst_4560 ( .ZN(net_5641), .A1(net_5438), .A2(net_3884) );
OR2_X4 inst_1076 ( .ZN(net_7936), .A2(net_7935), .A1(net_1147) );
NAND3_X2 inst_6360 ( .A3(net_12246), .ZN(net_12086), .A1(net_9100), .A2(net_4753) );
NAND3_X2 inst_6078 ( .ZN(net_13981), .A3(net_13980), .A2(net_9942), .A1(net_4980) );
INV_X4 inst_17660 ( .ZN(net_13362), .A(net_1815) );
INV_X4 inst_13292 ( .ZN(net_12387), .A(net_12386) );
NAND2_X2 inst_9264 ( .ZN(net_19178), .A2(net_12617), .A1(net_9179) );
OAI21_X2 inst_2000 ( .B1(net_13350), .ZN(net_11848), .B2(net_11847), .A(net_5603) );
NOR2_X2 inst_3748 ( .ZN(net_20413), .A2(net_7271), .A1(net_7241) );
AOI21_X4 inst_20153 ( .B1(net_19619), .ZN(net_15791), .A(net_10505), .B2(net_1046) );
NAND3_X2 inst_6732 ( .ZN(net_6481), .A2(net_6480), .A1(net_3454), .A3(net_1618) );
NAND2_X2 inst_10223 ( .ZN(net_8069), .A1(net_8068), .A2(net_8014) );
OR2_X2 inst_1195 ( .ZN(net_4036), .A2(net_3245), .A1(net_1898) );
NAND3_X2 inst_6222 ( .ZN(net_13240), .A3(net_10152), .A2(net_9477), .A1(net_5633) );
INV_X4 inst_16057 ( .ZN(net_2506), .A(net_1332) );
NAND2_X2 inst_9699 ( .A2(net_12099), .ZN(net_10215), .A1(net_9739) );
INV_X8 inst_12252 ( .ZN(net_3565), .A(net_2284) );
NAND2_X2 inst_11829 ( .ZN(net_7745), .A1(net_1776), .A2(net_200) );
NAND2_X4 inst_6839 ( .A2(net_21169), .ZN(net_18737), .A1(net_18669) );
OAI21_X2 inst_2248 ( .ZN(net_7326), .A(net_7325), .B2(net_6918), .B1(net_2201) );
INV_X4 inst_16740 ( .ZN(net_15550), .A(net_14159) );
OAI211_X2 inst_2453 ( .ZN(net_14432), .C2(net_13744), .C1(net_13095), .B(net_11335), .A(net_10371) );
OAI22_X2 inst_1312 ( .B1(net_20551), .A2(net_8504), .ZN(net_8471), .B2(net_6402), .A1(net_3230) );
CLKBUF_X2 inst_22505 ( .A(net_21856), .Z(net_22377) );
INV_X4 inst_17166 ( .ZN(net_741), .A(net_221) );
INV_X2 inst_18737 ( .ZN(net_7924), .A(net_7923) );
INV_X4 inst_16193 ( .ZN(net_15205), .A(net_8128) );
INV_X4 inst_15145 ( .ZN(net_3099), .A(net_3098) );
INV_X2 inst_18447 ( .ZN(net_19292), .A(net_12691) );
CLKBUF_X2 inst_22521 ( .A(net_22126), .Z(net_22393) );
NAND3_X2 inst_5785 ( .A2(net_20251), .ZN(net_15781), .A1(net_15249), .A3(net_10620) );
INV_X4 inst_18141 ( .A(net_21076), .ZN(net_665) );
NOR2_X2 inst_3419 ( .ZN(net_15576), .A2(net_14806), .A1(net_8734) );
INV_X4 inst_17423 ( .ZN(net_8820), .A(net_499) );
INV_X4 inst_13749 ( .ZN(net_9223), .A(net_7622) );
NAND2_X2 inst_8406 ( .ZN(net_18995), .A1(net_17244), .A2(net_17243) );
NOR2_X2 inst_4951 ( .ZN(net_7653), .A2(net_1304), .A1(net_338) );
INV_X4 inst_14954 ( .ZN(net_5970), .A(net_2754) );
INV_X4 inst_17637 ( .A(net_20876), .ZN(net_2629) );
SDFF_X2 inst_971 ( .QN(net_21022), .D(net_694), .SE(net_263), .CK(net_21968), .SI(x2650) );
OR2_X2 inst_1219 ( .ZN(net_2749), .A2(net_2687), .A1(net_2204) );
INV_X4 inst_18246 ( .A(net_21051), .ZN(net_350) );
NAND2_X2 inst_8018 ( .ZN(net_19947), .A2(net_18280), .A1(net_17327) );
NOR2_X2 inst_3459 ( .ZN(net_14736), .A2(net_13459), .A1(net_11447) );
INV_X4 inst_18345 ( .A(net_20778), .ZN(net_20777) );
INV_X4 inst_16362 ( .ZN(net_9968), .A(net_5694) );
CLKBUF_X2 inst_22549 ( .A(net_22420), .Z(net_22421) );
NOR2_X2 inst_4488 ( .ZN(net_5713), .A1(net_4288), .A2(net_3191) );
INV_X2 inst_18587 ( .ZN(net_10271), .A(net_10270) );
NAND2_X4 inst_7633 ( .A2(net_3704), .ZN(net_2107), .A1(net_856) );
INV_X4 inst_15357 ( .A(net_16287), .ZN(net_15936) );
INV_X4 inst_12716 ( .A(net_17775), .ZN(net_17756) );
NAND2_X2 inst_11732 ( .ZN(net_2689), .A2(net_2315), .A1(net_2199) );
NAND2_X2 inst_11741 ( .ZN(net_4269), .A1(net_2171), .A2(net_1805) );
INV_X4 inst_15992 ( .ZN(net_12708), .A(net_9313) );
INV_X4 inst_15123 ( .ZN(net_16125), .A(net_3164) );
INV_X2 inst_19502 ( .A(net_10335), .ZN(net_1257) );
NAND2_X2 inst_9454 ( .ZN(net_14316), .A2(net_11510), .A1(net_1361) );
NAND2_X4 inst_7222 ( .ZN(net_19527), .A2(net_7487), .A1(net_4396) );
INV_X2 inst_18380 ( .A(net_16919), .ZN(net_16824) );
INV_X4 inst_12628 ( .ZN(net_17925), .A(net_17924) );
INV_X4 inst_12991 ( .ZN(net_16965), .A(net_16491) );
INV_X4 inst_18038 ( .A(net_21180), .ZN(net_16607) );
NAND3_X2 inst_5842 ( .ZN(net_15471), .A3(net_14585), .A1(net_13408), .A2(net_12574) );
INV_X4 inst_16206 ( .ZN(net_2469), .A(net_1405) );
NAND2_X2 inst_10135 ( .ZN(net_8331), .A1(net_8330), .A2(net_6276) );
NOR2_X4 inst_3286 ( .ZN(net_2125), .A1(net_1248), .A2(net_1002) );
NOR2_X2 inst_4225 ( .ZN(net_7891), .A1(net_6624), .A2(net_955) );
NAND3_X4 inst_5625 ( .ZN(net_10943), .A2(net_9459), .A3(net_8720), .A1(net_5834) );
NAND2_X2 inst_11371 ( .ZN(net_3576), .A2(net_2606), .A1(net_2505) );
NAND2_X2 inst_11421 ( .ZN(net_11353), .A1(net_7007), .A2(net_2822) );
NAND2_X2 inst_9533 ( .ZN(net_12414), .A1(net_11087), .A2(net_11086) );
NOR2_X2 inst_4141 ( .A1(net_12006), .ZN(net_6928), .A2(net_6927) );
CLKBUF_X2 inst_22291 ( .A(net_21295), .Z(net_22163) );
AOI21_X2 inst_20308 ( .A(net_20889), .B2(net_18924), .B1(net_18923), .ZN(net_16065) );
INV_X4 inst_14293 ( .ZN(net_5568), .A(net_5567) );
NOR2_X2 inst_4591 ( .ZN(net_12952), .A1(net_3790), .A2(net_2585) );
INV_X4 inst_16470 ( .ZN(net_9728), .A(net_8616) );
NAND4_X2 inst_5318 ( .ZN(net_15770), .A2(net_15122), .A4(net_15000), .A1(net_12663), .A3(net_7296) );
INV_X4 inst_12493 ( .A(net_18670), .ZN(net_18653) );
NAND2_X2 inst_9865 ( .ZN(net_9489), .A1(net_8700), .A2(net_7555) );
INV_X4 inst_17119 ( .ZN(net_5008), .A(net_1776) );
NAND2_X2 inst_9162 ( .ZN(net_19891), .A1(net_13462), .A2(net_10436) );
NAND2_X2 inst_11290 ( .A1(net_7850), .A2(net_4092), .ZN(net_3833) );
XNOR2_X2 inst_188 ( .B(net_20411), .A(net_20410), .ZN(net_17807) );
NOR2_X2 inst_4528 ( .A2(net_19462), .ZN(net_4064), .A1(net_107) );
INV_X4 inst_13534 ( .ZN(net_12370), .A(net_9212) );
NAND3_X2 inst_6093 ( .ZN(net_13931), .A2(net_11000), .A3(net_8859), .A1(net_8059) );
INV_X4 inst_14586 ( .ZN(net_7984), .A(net_4486) );
AOI21_X2 inst_20423 ( .ZN(net_15218), .B1(net_15217), .B2(net_14115), .A(net_13974) );
INV_X2 inst_18732 ( .ZN(net_8016), .A(net_8015) );
NOR2_X4 inst_3011 ( .A2(net_19648), .ZN(net_6068), .A1(net_4991) );
INV_X2 inst_19555 ( .ZN(net_2181), .A(net_860) );
INV_X2 inst_18761 ( .ZN(net_7629), .A(net_7628) );
INV_X4 inst_16585 ( .ZN(net_6587), .A(net_6433) );
NOR2_X2 inst_4826 ( .ZN(net_2509), .A1(net_1848), .A2(net_1684) );
NAND3_X2 inst_6695 ( .ZN(net_7675), .A2(net_6100), .A3(net_4908), .A1(net_3576) );
OAI21_X2 inst_1537 ( .ZN(net_17922), .A(net_17748), .B2(net_17747), .B1(net_17746) );
OAI21_X2 inst_2041 ( .ZN(net_13842), .A(net_11296), .B1(net_11295), .B2(net_3775) );
NAND3_X2 inst_6323 ( .A3(net_14209), .ZN(net_12517), .A2(net_12516), .A1(net_9273) );
NAND4_X4 inst_5235 ( .A1(net_19633), .ZN(net_19006), .A4(net_15565), .A2(net_14204), .A3(net_10710) );
INV_X4 inst_15509 ( .ZN(net_3228), .A(net_2413) );
NOR2_X2 inst_4589 ( .ZN(net_12935), .A2(net_3542), .A1(net_2808) );
NAND3_X2 inst_6768 ( .ZN(net_5301), .A2(net_5300), .A3(net_5299), .A1(net_3767) );
INV_X2 inst_18443 ( .ZN(net_20739), .A(net_12817) );
NAND2_X2 inst_11550 ( .A1(net_20868), .ZN(net_18976), .A2(net_1387) );
NOR2_X4 inst_3325 ( .A2(net_19484), .ZN(net_820), .A1(net_163) );
INV_X4 inst_13393 ( .ZN(net_14711), .A(net_10711) );
NAND2_X2 inst_11145 ( .ZN(net_5380), .A1(net_3780), .A2(net_2487) );
NAND2_X2 inst_11085 ( .ZN(net_4404), .A1(net_4403), .A2(net_3756) );
NAND2_X2 inst_9083 ( .ZN(net_19031), .A1(net_13815), .A2(net_13814) );
INV_X4 inst_13991 ( .A(net_9006), .ZN(net_7774) );
NOR2_X2 inst_4168 ( .ZN(net_8166), .A2(net_4903), .A1(net_3842) );
XNOR2_X2 inst_195 ( .ZN(net_17676), .A(net_17675), .B(net_482) );
INV_X2 inst_18507 ( .A(net_13127), .ZN(net_11689) );
NAND2_X2 inst_11835 ( .A1(net_20923), .ZN(net_4214), .A2(net_1751) );
INV_X4 inst_12839 ( .A(net_17237), .ZN(net_17212) );
OAI21_X2 inst_1987 ( .ZN(net_12047), .B1(net_10046), .B2(net_7744), .A(net_6038) );
AOI21_X2 inst_20874 ( .ZN(net_8503), .A(net_8502), .B1(net_8501), .B2(net_8500) );
INV_X4 inst_13418 ( .ZN(net_10263), .A(net_8773) );
INV_X2 inst_19602 ( .A(net_238), .ZN(net_145) );
INV_X4 inst_14372 ( .ZN(net_6294), .A(net_5181) );
NAND3_X4 inst_5605 ( .ZN(net_19308), .A3(net_13772), .A2(net_10963), .A1(net_8608) );
NAND2_X4 inst_7070 ( .A2(net_20888), .A1(net_20395), .ZN(net_20250) );
NAND2_X4 inst_7106 ( .A1(net_20245), .ZN(net_13803), .A2(net_11645) );
AND2_X4 inst_21239 ( .A2(net_7667), .ZN(net_6052), .A1(net_1376) );
AOI211_X2 inst_21007 ( .ZN(net_15843), .C1(net_15842), .C2(net_15284), .B(net_10934), .A(net_8648) );
NOR2_X2 inst_4780 ( .ZN(net_19327), .A1(net_2887), .A2(net_2886) );
INV_X4 inst_12981 ( .A(net_17815), .ZN(net_17752) );
INV_X4 inst_15468 ( .ZN(net_9064), .A(net_2460) );
NOR2_X2 inst_4658 ( .ZN(net_3801), .A1(net_3297), .A2(net_2386) );
NAND3_X2 inst_5916 ( .ZN(net_20190), .A3(net_18949), .A1(net_18948), .A2(net_12486) );
NAND2_X4 inst_7154 ( .A1(net_20528), .ZN(net_12989), .A2(net_8590) );
OAI21_X2 inst_1589 ( .A(net_21212), .ZN(net_16258), .B2(net_15929), .B1(net_11375) );
NAND2_X2 inst_11994 ( .ZN(net_1208), .A1(net_366), .A2(net_74) );
NAND2_X2 inst_8926 ( .ZN(net_14940), .A2(net_13690), .A1(net_13093) );
INV_X4 inst_14114 ( .ZN(net_11290), .A(net_8044) );
NAND3_X4 inst_5607 ( .ZN(net_14122), .A3(net_10600), .A1(net_8872), .A2(net_8630) );
CLKBUF_X2 inst_21783 ( .A(net_21654), .Z(net_21655) );
INV_X4 inst_14095 ( .ZN(net_6192), .A(net_6191) );
INV_X4 inst_16499 ( .ZN(net_10134), .A(net_7121) );
INV_X4 inst_15263 ( .A(net_3264), .ZN(net_2768) );
INV_X4 inst_15160 ( .ZN(net_4910), .A(net_2115) );
XNOR2_X2 inst_335 ( .B(net_17404), .A(net_17000), .ZN(net_16988) );
INV_X4 inst_15244 ( .ZN(net_3563), .A(net_2810) );
INV_X4 inst_12827 ( .ZN(net_17155), .A(net_17154) );
INV_X4 inst_14406 ( .ZN(net_5099), .A(net_4422) );
NAND2_X4 inst_6862 ( .ZN(net_18411), .A2(net_18253), .A1(net_18206) );
NAND2_X2 inst_8420 ( .ZN(net_17303), .A1(net_16925), .A2(net_16749) );
NAND2_X2 inst_9336 ( .ZN(net_12279), .A2(net_8873), .A1(net_7363) );
CLKBUF_X2 inst_22712 ( .A(net_22583), .Z(net_22584) );
NAND2_X2 inst_11562 ( .ZN(net_3441), .A1(net_2470), .A2(net_797) );
INV_X4 inst_14045 ( .A(net_8333), .ZN(net_6258) );
INV_X4 inst_16155 ( .A(net_14227), .ZN(net_2368) );
INV_X4 inst_14276 ( .ZN(net_6257), .A(net_5657) );
XNOR2_X2 inst_438 ( .ZN(net_16094), .A(net_16093), .B(net_15587) );
AOI21_X2 inst_20870 ( .B2(net_9076), .ZN(net_8569), .A(net_8568), .B1(net_8567) );
INV_X4 inst_13311 ( .ZN(net_11666), .A(net_10374) );
CLKBUF_X2 inst_22620 ( .A(net_22491), .Z(net_22492) );
NAND2_X4 inst_7326 ( .ZN(net_6009), .A2(net_3512), .A1(net_3184) );
NAND3_X2 inst_6351 ( .ZN(net_12161), .A1(net_12160), .A3(net_11766), .A2(net_7264) );
INV_X2 inst_19516 ( .ZN(net_1130), .A(net_1129) );
NAND2_X2 inst_10769 ( .ZN(net_19750), .A1(net_8700), .A2(net_4126) );
INV_X4 inst_14336 ( .ZN(net_5987), .A(net_5390) );
NAND2_X2 inst_9692 ( .ZN(net_19908), .A1(net_10236), .A2(net_10235) );
XNOR2_X2 inst_324 ( .B(net_21199), .ZN(net_17028), .A(net_16667) );
NAND2_X2 inst_11640 ( .ZN(net_2501), .A2(net_1737), .A1(net_703) );
NOR2_X2 inst_3550 ( .ZN(net_13097), .A2(net_11180), .A1(net_1286) );
NAND3_X2 inst_6046 ( .ZN(net_20351), .A1(net_13488), .A2(net_11878), .A3(net_9334) );
AOI21_X2 inst_20746 ( .A(net_12916), .ZN(net_11401), .B2(net_10631), .B1(net_5795) );
NOR2_X2 inst_4083 ( .A1(net_12320), .A2(net_10595), .ZN(net_7307) );
INV_X4 inst_17240 ( .ZN(net_1136), .A(net_231) );
XOR2_X2 inst_43 ( .A(net_21170), .Z(net_542), .B(net_541) );
NAND3_X2 inst_5936 ( .ZN(net_14922), .A3(net_14921), .A2(net_13885), .A1(net_13626) );
OAI21_X2 inst_1707 ( .ZN(net_20644), .B2(net_14107), .B1(net_13536), .A(net_1832) );
INV_X4 inst_17955 ( .A(net_21133), .ZN(net_16921) );
NAND2_X4 inst_7213 ( .A2(net_20541), .ZN(net_12284), .A1(net_5764) );
NAND3_X2 inst_6715 ( .ZN(net_7092), .A2(net_7091), .A3(net_7090), .A1(net_3858) );
NAND2_X2 inst_8115 ( .ZN(net_18100), .A2(net_18099), .A1(net_17767) );
XNOR2_X2 inst_375 ( .A(net_17760), .ZN(net_16840), .B(net_16839) );
NAND2_X2 inst_11241 ( .ZN(net_6521), .A1(net_4212), .A2(net_3933) );
NAND2_X2 inst_9959 ( .ZN(net_19966), .A2(net_8915), .A1(net_6228) );
NAND2_X2 inst_8606 ( .A2(net_20075), .ZN(net_19105), .A1(net_17483) );
NOR2_X2 inst_3490 ( .ZN(net_19612), .A1(net_14200), .A2(net_10420) );
NAND2_X4 inst_7039 ( .ZN(net_16449), .A1(net_16423), .A2(net_16380) );
INV_X4 inst_15780 ( .ZN(net_19825), .A(net_3075) );
NAND2_X2 inst_10933 ( .ZN(net_6330), .A2(net_2915), .A1(net_2585) );
XNOR2_X2 inst_285 ( .B(net_21207), .ZN(net_17160), .A(net_16814) );
NAND2_X4 inst_7215 ( .ZN(net_9395), .A1(net_7865), .A2(net_3874) );
OAI21_X2 inst_1830 ( .ZN(net_14134), .B1(net_11238), .B2(net_10455), .A(net_512) );
INV_X2 inst_18515 ( .ZN(net_11569), .A(net_11568) );
NAND2_X2 inst_11780 ( .ZN(net_2023), .A2(net_253), .A1(x6494) );
NAND3_X4 inst_5563 ( .ZN(net_15999), .A1(net_15696), .A3(net_14756), .A2(net_10018) );
OAI21_X2 inst_1563 ( .ZN(net_17502), .B1(net_17091), .B2(net_16935), .A(net_16710) );
NAND3_X2 inst_6363 ( .ZN(net_12081), .A3(net_10106), .A1(net_9008), .A2(net_8239) );
INV_X4 inst_17044 ( .ZN(net_8724), .A(net_6631) );
AOI21_X2 inst_20712 ( .ZN(net_12054), .B1(net_12053), .A(net_11057), .B2(net_7746) );
NOR2_X4 inst_3242 ( .A2(net_5043), .ZN(net_3374), .A1(net_2328) );
NAND2_X4 inst_7398 ( .ZN(net_11995), .A2(net_4305), .A1(net_4089) );
NAND2_X2 inst_10638 ( .ZN(net_6422), .A2(net_6421), .A1(net_2691) );
AOI21_X2 inst_20351 ( .B1(net_19918), .ZN(net_15716), .B2(net_14738), .A(net_8570) );
NAND2_X2 inst_9895 ( .ZN(net_9402), .A1(net_9401), .A2(net_9400) );
SDFF_X2 inst_982 ( .QN(net_21048), .D(net_581), .SE(net_263), .CK(net_22518), .SI(x2219) );
NOR2_X4 inst_3138 ( .ZN(net_5066), .A1(net_3780), .A2(net_3329) );
INV_X4 inst_17451 ( .A(net_10345), .ZN(net_458) );
NAND2_X2 inst_10864 ( .ZN(net_12752), .A1(net_7432), .A2(net_5433) );
XNOR2_X2 inst_299 ( .B(net_21124), .A(net_19444), .ZN(net_17346) );
INV_X4 inst_13871 ( .A(net_11629), .ZN(net_7437) );
NAND2_X2 inst_10567 ( .ZN(net_7978), .A1(net_4940), .A2(net_874) );
NAND2_X4 inst_7656 ( .ZN(net_1248), .A1(net_875), .A2(net_234) );
OAI21_X2 inst_1798 ( .ZN(net_14501), .A(net_14500), .B2(net_11563), .B1(net_11522) );
NOR2_X4 inst_2927 ( .ZN(net_9411), .A2(net_7874), .A1(net_7873) );
CLKBUF_X2 inst_22528 ( .A(net_22399), .Z(net_22400) );
NAND2_X2 inst_10336 ( .ZN(net_10407), .A1(net_5845), .A2(net_5824) );
CLKBUF_X2 inst_22330 ( .A(net_22201), .Z(net_22202) );
CLKBUF_X2 inst_22744 ( .A(net_22615), .Z(net_22616) );
CLKBUF_X2 inst_21576 ( .A(net_21447), .Z(net_21448) );
NAND3_X2 inst_5853 ( .ZN(net_15419), .A3(net_14491), .A1(net_14356), .A2(net_7770) );
NAND2_X2 inst_10383 ( .ZN(net_7339), .A1(net_7338), .A2(net_7337) );
INV_X4 inst_17826 ( .ZN(net_992), .A(net_107) );
INV_X4 inst_17016 ( .ZN(net_7397), .A(net_554) );
NAND2_X2 inst_8727 ( .ZN(net_16067), .A2(net_15774), .A1(net_15677) );
NOR3_X2 inst_2760 ( .ZN(net_11193), .A3(net_11192), .A2(net_8419), .A1(net_6621) );
NAND3_X2 inst_6452 ( .ZN(net_11756), .A1(net_9691), .A2(net_9630), .A3(net_8912) );
INV_X2 inst_18838 ( .ZN(net_6735), .A(net_6734) );
INV_X4 inst_15213 ( .ZN(net_4409), .A(net_2889) );
NAND2_X4 inst_7098 ( .ZN(net_13593), .A2(net_13556), .A1(net_13440) );
INV_X4 inst_17596 ( .ZN(net_596), .A(net_329) );
NAND3_X2 inst_6288 ( .A2(net_19895), .ZN(net_12841), .A3(net_11425), .A1(net_6820) );
NAND2_X4 inst_7030 ( .A1(net_20517), .ZN(net_19959), .A2(net_17008) );
INV_X4 inst_15581 ( .ZN(net_3955), .A(net_3096) );
NOR2_X2 inst_5129 ( .ZN(net_250), .A2(net_230), .A1(net_227) );
INV_X4 inst_13524 ( .ZN(net_12807), .A(net_9333) );
INV_X4 inst_14841 ( .ZN(net_8473), .A(net_3854) );
NAND2_X2 inst_10656 ( .ZN(net_9847), .A1(net_6316), .A2(net_6315) );
NOR2_X2 inst_4995 ( .ZN(net_1373), .A2(net_1196), .A1(net_221) );
NOR2_X4 inst_3260 ( .ZN(net_2966), .A1(net_1507), .A2(net_85) );
NOR2_X4 inst_3158 ( .A1(net_20545), .ZN(net_5475), .A2(net_2546) );
NOR2_X2 inst_4190 ( .ZN(net_11324), .A2(net_8035), .A1(net_3289) );
INV_X4 inst_17878 ( .A(net_1469), .ZN(net_238) );
INV_X4 inst_13894 ( .ZN(net_9747), .A(net_7292) );
NAND2_X2 inst_11248 ( .ZN(net_8831), .A1(net_5595), .A2(net_3872) );
CLKBUF_X2 inst_22635 ( .A(net_21514), .Z(net_22507) );
CLKBUF_X2 inst_21482 ( .A(net_21353), .Z(net_21354) );
NAND4_X2 inst_5387 ( .ZN(net_19775), .A2(net_19710), .A1(net_19709), .A4(net_12684), .A3(net_8723) );
AOI21_X2 inst_20402 ( .B1(net_15708), .ZN(net_15377), .A(net_14273), .B2(net_13891) );
INV_X4 inst_14067 ( .A(net_6241), .ZN(net_6240) );
OAI21_X2 inst_2186 ( .ZN(net_19215), .B1(net_7519), .A(net_6570), .B2(net_4964) );
NOR2_X4 inst_3269 ( .ZN(net_3590), .A1(net_1934), .A2(net_1933) );
INV_X4 inst_15745 ( .A(net_15924), .ZN(net_1946) );
OAI21_X2 inst_1944 ( .ZN(net_12650), .A(net_11088), .B2(net_9103), .B1(net_2845) );
NAND2_X2 inst_9079 ( .A1(net_15810), .ZN(net_13830), .A2(net_11689) );
XNOR2_X2 inst_210 ( .ZN(net_17569), .B(net_17378), .A(net_17199) );
INV_X4 inst_13763 ( .A(net_9635), .ZN(net_7609) );
NAND2_X2 inst_11675 ( .ZN(net_2356), .A2(net_1590), .A1(net_198) );
NOR2_X4 inst_3101 ( .A2(net_7700), .ZN(net_5225), .A1(net_4268) );
INV_X4 inst_16142 ( .ZN(net_2827), .A(net_1796) );
NOR2_X2 inst_4942 ( .ZN(net_3071), .A2(net_2202), .A1(net_606) );
INV_X4 inst_14998 ( .A(net_13095), .ZN(net_13032) );
AOI21_X4 inst_20169 ( .B2(net_19833), .B1(net_19832), .A(net_15616), .ZN(net_15597) );
NAND4_X2 inst_5331 ( .ZN(net_20311), .A4(net_19093), .A1(net_19092), .A3(net_14407), .A2(net_13092) );
NAND2_X2 inst_8164 ( .ZN(net_17968), .A1(net_17967), .A2(net_17853) );
AOI21_X2 inst_20616 ( .ZN(net_13587), .A(net_12542), .B2(net_10665), .B1(net_4603) );
NAND2_X4 inst_7123 ( .ZN(net_12617), .A1(net_9203), .A2(net_1903) );
OAI22_X2 inst_1294 ( .ZN(net_12473), .A2(net_11021), .B1(net_10989), .B2(net_4659), .A1(net_1410) );
INV_X4 inst_16865 ( .A(net_4163), .ZN(net_2199) );
OAI21_X2 inst_1712 ( .ZN(net_15195), .A(net_14643), .B2(net_13680), .B1(net_13413) );
NAND4_X4 inst_5238 ( .A4(net_19675), .A1(net_19674), .ZN(net_19353), .A2(net_11229), .A3(net_10675) );
INV_X4 inst_14605 ( .ZN(net_16041), .A(net_4436) );
NOR2_X4 inst_3108 ( .ZN(net_9558), .A1(net_4074), .A2(net_2549) );
INV_X4 inst_12626 ( .ZN(net_20128), .A(net_17964) );
NOR2_X4 inst_2853 ( .ZN(net_20429), .A2(net_10262), .A1(net_7242) );
NAND2_X4 inst_7267 ( .A1(net_19299), .ZN(net_7588), .A2(net_3086) );
INV_X4 inst_15331 ( .A(net_5385), .ZN(net_4419) );
NAND2_X2 inst_10291 ( .A1(net_20560), .ZN(net_10106), .A2(net_5115) );
NAND3_X2 inst_6546 ( .ZN(net_10561), .A1(net_9500), .A3(net_6806), .A2(net_5905) );
MUX2_X2 inst_12166 ( .Z(net_20690), .S(net_12763), .A(net_11855), .B(net_11854) );
NAND2_X2 inst_7855 ( .A1(net_18582), .ZN(net_18578), .A2(net_18560) );
INV_X4 inst_15055 ( .ZN(net_3854), .A(net_3678) );
NAND2_X2 inst_8553 ( .ZN(net_16779), .A1(net_16778), .A2(net_16777) );
NAND2_X2 inst_11658 ( .ZN(net_2425), .A2(net_2424), .A1(net_1690) );
NAND2_X2 inst_10853 ( .ZN(net_13456), .A2(net_3881), .A1(net_3812) );
INV_X2 inst_18651 ( .A(net_10974), .ZN(net_10787) );
CLKBUF_X2 inst_22573 ( .A(net_21734), .Z(net_22445) );
NAND3_X2 inst_6291 ( .ZN(net_12832), .A1(net_11043), .A2(net_10192), .A3(net_8301) );
INV_X4 inst_14848 ( .ZN(net_5405), .A(net_4448) );
INV_X4 inst_12476 ( .ZN(net_18702), .A(net_18701) );
INV_X4 inst_14547 ( .ZN(net_4613), .A(net_4612) );
NAND3_X2 inst_5740 ( .A3(net_19289), .A1(net_19288), .ZN(net_19174), .A2(net_14800) );
NAND2_X2 inst_10602 ( .A1(net_9575), .ZN(net_6619), .A2(net_6618) );
NAND2_X2 inst_10993 ( .A2(net_20807), .ZN(net_9294), .A1(net_6274) );
NAND3_X2 inst_6227 ( .ZN(net_13233), .A3(net_10166), .A1(net_9844), .A2(net_9464) );
INV_X4 inst_13489 ( .ZN(net_9521), .A(net_9520) );
INV_X4 inst_14930 ( .ZN(net_6627), .A(net_4366) );
INV_X4 inst_15511 ( .ZN(net_3481), .A(net_2409) );
INV_X2 inst_18613 ( .ZN(net_12899), .A(net_9672) );
INV_X4 inst_14898 ( .A(net_13355), .ZN(net_3628) );
CLKBUF_X2 inst_21573 ( .A(net_21378), .Z(net_21445) );
NAND2_X2 inst_11620 ( .ZN(net_4849), .A2(net_2726), .A1(net_2123) );
NAND2_X2 inst_11605 ( .ZN(net_4563), .A1(net_2630), .A2(net_2504) );
AOI21_X2 inst_20940 ( .A(net_8455), .ZN(net_6427), .B2(net_6426), .B1(net_4563) );
SDFF_X2 inst_907 ( .Q(net_21218), .SI(net_16847), .SE(net_125), .CK(net_22208), .D(x7443) );
CLKBUF_X2 inst_22485 ( .A(net_21302), .Z(net_22357) );
SDFF_X2 inst_922 ( .Q(net_21211), .D(net_16480), .SE(net_263), .CK(net_22134), .SI(x5787) );
NAND2_X2 inst_11323 ( .ZN(net_8501), .A2(net_3753), .A1(net_90) );
INV_X4 inst_18095 ( .A(net_20943), .ZN(net_386) );
NAND2_X2 inst_8225 ( .ZN(net_17798), .A2(net_17797), .A1(net_17658) );
AOI21_X2 inst_20719 ( .ZN(net_11998), .B1(net_11997), .B2(net_7704), .A(net_7140) );
INV_X2 inst_18387 ( .A(net_17126), .ZN(net_16640) );
NAND2_X2 inst_8773 ( .ZN(net_15830), .A2(net_15596), .A1(net_1046) );
INV_X2 inst_19111 ( .A(net_5282), .ZN(net_4460) );
INV_X4 inst_15072 ( .A(net_9487), .ZN(net_3274) );
INV_X8 inst_12435 ( .ZN(net_20443), .A(net_20442) );
NAND2_X2 inst_10693 ( .ZN(net_10431), .A2(net_6076), .A1(net_90) );
NAND2_X2 inst_9475 ( .ZN(net_11462), .A2(net_10988), .A1(net_10598) );
INV_X4 inst_14418 ( .A(net_8553), .ZN(net_6011) );
NAND2_X2 inst_8516 ( .A1(net_17031), .ZN(net_16914), .A2(net_16562) );
INV_X4 inst_12621 ( .ZN(net_17996), .A(net_17995) );
INV_X4 inst_13231 ( .ZN(net_20832), .A(net_12491) );
NOR2_X2 inst_3907 ( .ZN(net_13114), .A1(net_11747), .A2(net_10774) );
NAND2_X2 inst_9619 ( .ZN(net_10691), .A1(net_10690), .A2(net_8477) );
DFF_X1 inst_19914 ( .D(net_16547), .CK(net_22785), .Q(x1299) );
INV_X4 inst_14752 ( .ZN(net_4072), .A(net_4071) );
INV_X8 inst_12383 ( .ZN(net_161), .A(net_116) );
NOR2_X2 inst_3692 ( .ZN(net_11323), .A1(net_11322), .A2(net_6824) );
INV_X4 inst_18033 ( .A(net_21028), .ZN(net_593) );
XNOR2_X2 inst_653 ( .B(net_16402), .ZN(net_362), .A(net_361) );
NAND2_X2 inst_8304 ( .ZN(net_17668), .A2(net_17397), .A1(net_17265) );
OAI21_X2 inst_1746 ( .ZN(net_20643), .B2(net_13535), .B1(net_13470), .A(net_1402) );
NAND2_X2 inst_11099 ( .ZN(net_5606), .A1(net_4340), .A2(net_4330) );
AOI22_X2 inst_20014 ( .ZN(net_11772), .A1(net_11771), .B1(net_11770), .A2(net_7896), .B2(net_4500) );
INV_X4 inst_18274 ( .ZN(net_19454), .A(net_16932) );
INV_X4 inst_13406 ( .A(net_12193), .ZN(net_10401) );
NAND2_X2 inst_8233 ( .ZN(net_19119), .A1(net_17756), .A2(net_466) );
CLKBUF_X2 inst_21760 ( .A(net_21331), .Z(net_21632) );
INV_X4 inst_15817 ( .A(net_11426), .ZN(net_6513) );
NOR2_X2 inst_3649 ( .ZN(net_11674), .A2(net_11673), .A1(net_8104) );
INV_X4 inst_17131 ( .ZN(net_6394), .A(net_3310) );
NOR2_X2 inst_4609 ( .A1(net_13538), .A2(net_11902), .ZN(net_3738) );
NAND3_X2 inst_6526 ( .ZN(net_10614), .A3(net_10613), .A1(net_10440), .A2(net_5101) );
NAND2_X2 inst_11843 ( .A1(net_20923), .ZN(net_1875), .A2(net_61) );
NOR3_X2 inst_2656 ( .ZN(net_15281), .A3(net_15280), .A1(net_14228), .A2(net_8321) );
INV_X4 inst_16165 ( .ZN(net_2891), .A(net_1039) );
NAND2_X2 inst_8301 ( .ZN(net_17692), .A1(net_17425), .A2(net_17291) );
OAI21_X2 inst_1604 ( .A(net_20944), .ZN(net_16152), .B2(net_15740), .B1(net_10173) );
CLKBUF_X2 inst_21902 ( .A(net_21773), .Z(net_21774) );
INV_X4 inst_18146 ( .A(net_21031), .ZN(net_724) );
NAND2_X2 inst_9426 ( .ZN(net_13811), .A1(net_12888), .A2(net_11048) );
AOI211_X2 inst_21067 ( .ZN(net_8484), .B(net_8483), .A(net_5641), .C1(net_5616), .C2(net_2271) );
INV_X2 inst_18818 ( .A(net_10525), .ZN(net_7013) );
INV_X4 inst_13854 ( .ZN(net_11767), .A(net_7464) );
INV_X4 inst_14441 ( .A(net_14974), .ZN(net_8031) );
INV_X2 inst_19608 ( .A(net_21243), .ZN(net_53) );
NAND2_X2 inst_8592 ( .ZN(net_16695), .A2(net_16694), .A1(net_2571) );
INV_X4 inst_16934 ( .ZN(net_1224), .A(net_927) );
XOR2_X2 inst_7 ( .A(net_21117), .B(net_17312), .Z(net_17296) );
INV_X2 inst_18642 ( .ZN(net_11481), .A(net_9375) );
NAND2_X2 inst_9672 ( .ZN(net_20730), .A1(net_12454), .A2(net_8049) );
AOI21_X4 inst_20251 ( .B2(net_20094), .A(net_8924), .ZN(net_7315), .B1(net_5627) );
INV_X4 inst_16465 ( .ZN(net_15289), .A(net_9518) );
AOI21_X2 inst_20929 ( .B1(net_10864), .ZN(net_7081), .B2(net_7080), .A(net_3623) );
NOR2_X2 inst_3450 ( .ZN(net_14914), .A1(net_14913), .A2(net_13759) );
NAND2_X2 inst_9707 ( .ZN(net_13810), .A1(net_10398), .A2(net_10197) );
INV_X4 inst_13742 ( .A(net_11927), .ZN(net_7636) );
NAND4_X2 inst_5408 ( .ZN(net_14641), .A3(net_13840), .A2(net_12182), .A1(net_9858), .A4(net_9751) );
INV_X4 inst_17074 ( .ZN(net_1786), .A(net_374) );
NAND2_X2 inst_12036 ( .A1(net_1614), .ZN(net_1050), .A2(net_493) );
OR2_X2 inst_1136 ( .A2(net_12957), .ZN(net_12697), .A1(net_60) );
AOI22_X2 inst_19963 ( .B1(net_16054), .ZN(net_16040), .A2(net_15523), .B2(net_13155), .A1(net_4189) );
CLKBUF_X2 inst_21501 ( .A(net_21372), .Z(net_21373) );
CLKBUF_X2 inst_21656 ( .A(net_21527), .Z(net_21528) );
NAND2_X2 inst_10402 ( .ZN(net_7276), .A2(net_7275), .A1(net_6714) );
AOI21_X2 inst_20835 ( .ZN(net_9319), .A(net_7489), .B2(net_6387), .B1(net_4521) );
INV_X4 inst_13360 ( .ZN(net_12348), .A(net_10943) );
NAND2_X2 inst_11262 ( .ZN(net_13203), .A1(net_7858), .A2(net_3905) );
INV_X2 inst_19069 ( .ZN(net_4631), .A(net_4630) );
INV_X4 inst_16141 ( .ZN(net_2502), .A(net_1791) );
NAND2_X2 inst_9621 ( .ZN(net_10685), .A2(net_8493), .A1(net_816) );
INV_X4 inst_14474 ( .ZN(net_8171), .A(net_4895) );
NOR2_X4 inst_3311 ( .ZN(net_2519), .A2(net_982), .A1(net_221) );
INV_X4 inst_13598 ( .ZN(net_14745), .A(net_7255) );
INV_X4 inst_13339 ( .ZN(net_11103), .A(net_11102) );
NOR2_X2 inst_5081 ( .ZN(net_10158), .A2(net_4915), .A1(net_862) );
NOR2_X2 inst_5117 ( .ZN(net_319), .A1(net_318), .A2(net_317) );
NOR2_X2 inst_4929 ( .ZN(net_1779), .A2(net_1370), .A1(net_61) );
NOR2_X2 inst_5114 ( .ZN(net_849), .A2(net_508), .A1(net_62) );
INV_X4 inst_13942 ( .ZN(net_6806), .A(net_6805) );
CLKBUF_X2 inst_21637 ( .A(net_21508), .Z(net_21509) );
INV_X4 inst_14885 ( .ZN(net_6323), .A(net_3669) );
CLKBUF_X2 inst_21984 ( .A(net_21855), .Z(net_21856) );
NAND2_X2 inst_10423 ( .A1(net_13651), .ZN(net_7224), .A2(net_5502) );
NAND2_X4 inst_7341 ( .A2(net_19314), .ZN(net_10144), .A1(net_4821) );
AOI21_X2 inst_20393 ( .ZN(net_15461), .B1(net_14461), .B2(net_13337), .A(net_1774) );
NAND3_X2 inst_6268 ( .ZN(net_12961), .A2(net_12960), .A3(net_5484), .A1(net_2895) );
INV_X4 inst_17753 ( .ZN(net_417), .A(net_90) );
NOR2_X2 inst_3713 ( .ZN(net_10994), .A1(net_10993), .A2(net_7899) );
NAND3_X2 inst_5681 ( .ZN(net_16330), .A3(net_16079), .A2(net_14221), .A1(net_14084) );
OAI211_X2 inst_2394 ( .ZN(net_16132), .A(net_15850), .C2(net_15428), .B(net_14894), .C1(net_1923) );
DFF_X1 inst_19874 ( .D(net_17027), .CK(net_21334), .Q(x246) );
NOR2_X2 inst_4574 ( .A1(net_5594), .ZN(net_5039), .A2(net_3286) );
AOI21_X2 inst_20878 ( .ZN(net_8454), .B2(net_7256), .B1(net_4032), .A(net_3240) );
NAND2_X2 inst_8562 ( .A1(net_21195), .ZN(net_16746), .A2(net_16576) );
NAND2_X2 inst_9404 ( .ZN(net_11684), .A2(net_11683), .A1(net_6183) );
NAND2_X2 inst_10681 ( .ZN(net_7545), .A1(net_7075), .A2(net_6052) );
NAND2_X2 inst_10612 ( .ZN(net_10446), .A1(net_6598), .A2(net_6597) );
NAND4_X2 inst_5294 ( .ZN(net_15929), .A2(net_15204), .A1(net_14005), .A4(net_8702), .A3(net_5533) );
INV_X4 inst_17962 ( .A(net_21002), .ZN(net_2437) );
NAND4_X4 inst_5251 ( .A3(net_12076), .ZN(net_11823), .A2(net_11822), .A4(net_11240), .A1(net_10762) );
NOR2_X2 inst_4422 ( .ZN(net_12396), .A1(net_9278), .A2(net_4974) );
INV_X4 inst_12578 ( .ZN(net_18251), .A(net_18204) );
INV_X8 inst_12219 ( .ZN(net_10467), .A(net_5993) );
CLKBUF_X2 inst_22402 ( .A(net_22273), .Z(net_22274) );
INV_X2 inst_19595 ( .A(net_314), .ZN(net_207) );
CLKBUF_X2 inst_22224 ( .A(net_22095), .Z(net_22096) );
INV_X4 inst_14056 ( .ZN(net_9647), .A(net_8023) );
NAND2_X2 inst_11905 ( .ZN(net_1564), .A2(net_1563), .A1(net_221) );
NAND2_X2 inst_8623 ( .ZN(net_16603), .A2(net_16602), .A1(net_16488) );
NOR2_X2 inst_5092 ( .A1(net_1339), .ZN(net_827), .A2(net_103) );
AOI21_X2 inst_20551 ( .B2(net_19574), .B1(net_19573), .A(net_15301), .ZN(net_14306) );
INV_X4 inst_15330 ( .A(net_3829), .ZN(net_2611) );
NAND4_X2 inst_5342 ( .ZN(net_15458), .A1(net_14745), .A2(net_14468), .A3(net_11577), .A4(net_8838) );
OAI21_X2 inst_1670 ( .ZN(net_15618), .B2(net_14277), .B1(net_11798), .A(net_1528) );
INV_X2 inst_19374 ( .ZN(net_2185), .A(net_2184) );
INV_X4 inst_12932 ( .ZN(net_16787), .A(net_16495) );
NAND2_X2 inst_11491 ( .A1(net_4762), .ZN(net_3997), .A2(net_3090) );
AOI21_X4 inst_20171 ( .B2(net_19114), .B1(net_19113), .ZN(net_19019), .A(net_15550) );
NAND2_X2 inst_10352 ( .ZN(net_12446), .A1(net_7473), .A2(net_5812) );
NAND2_X2 inst_8646 ( .A2(net_16574), .ZN(net_16567), .A1(net_16413) );
NAND2_X2 inst_9028 ( .ZN(net_19823), .A1(net_14075), .A2(net_11904) );
INV_X4 inst_16512 ( .A(net_4299), .ZN(net_4212) );
NAND2_X2 inst_10677 ( .ZN(net_9838), .A2(net_5952), .A1(net_143) );
NAND2_X2 inst_10327 ( .ZN(net_11720), .A1(net_9090), .A2(net_7837) );
NOR2_X2 inst_5027 ( .ZN(net_3208), .A1(net_3014), .A2(net_1155) );
NAND3_X2 inst_5883 ( .ZN(net_15243), .A1(net_14735), .A3(net_13429), .A2(net_10299) );
NOR2_X4 inst_3113 ( .ZN(net_6842), .A1(net_3977), .A2(net_3491) );
INV_X4 inst_13500 ( .ZN(net_9435), .A(net_9434) );
CLKBUF_X2 inst_22470 ( .A(net_22049), .Z(net_22342) );
INV_X2 inst_19074 ( .ZN(net_4611), .A(net_4610) );
INV_X2 inst_18775 ( .A(net_11388), .ZN(net_7547) );
NOR2_X2 inst_3695 ( .ZN(net_11191), .A2(net_7998), .A1(net_6814) );
INV_X8 inst_12309 ( .ZN(net_7153), .A(net_5658) );
NAND3_X2 inst_6687 ( .ZN(net_7709), .A3(net_7044), .A1(net_3705), .A2(net_3179) );
OAI211_X2 inst_2385 ( .C1(net_20872), .ZN(net_16549), .C2(net_16371), .B(net_16088), .A(net_5497) );
OAI21_X2 inst_2336 ( .ZN(net_4683), .B1(net_3513), .A(net_3457), .B2(net_2252) );
INV_X4 inst_18061 ( .A(net_21138), .ZN(net_745) );
INV_X4 inst_16044 ( .ZN(net_11465), .A(net_6999) );
NAND3_X2 inst_5927 ( .ZN(net_14976), .A3(net_14441), .A1(net_14028), .A2(net_2959) );
NAND2_X2 inst_8574 ( .ZN(net_16731), .A1(net_16443), .A2(net_16410) );
INV_X4 inst_13549 ( .A(net_16659), .ZN(net_9173) );
NAND2_X2 inst_9482 ( .A1(net_11645), .ZN(net_11453), .A2(net_10941) );
INV_X4 inst_17263 ( .ZN(net_1269), .A(net_167) );
XNOR2_X2 inst_223 ( .ZN(net_17506), .A(net_17072), .B(net_605) );
NAND3_X2 inst_6814 ( .ZN(net_8394), .A2(net_3134), .A1(net_2361), .A3(net_2348) );
INV_X2 inst_19360 ( .A(net_3225), .ZN(net_2297) );
NAND4_X2 inst_5278 ( .ZN(net_16014), .A1(net_15608), .A4(net_15085), .A3(net_12403), .A2(net_10693) );
NAND3_X2 inst_6042 ( .ZN(net_14277), .A1(net_14276), .A2(net_12304), .A3(net_9820) );
INV_X4 inst_15884 ( .ZN(net_2991), .A(net_2519) );
INV_X4 inst_13811 ( .ZN(net_11065), .A(net_7539) );
OAI211_X2 inst_2420 ( .ZN(net_15323), .A(net_14413), .B(net_13574), .C2(net_9305), .C1(net_4350) );
NOR2_X2 inst_3564 ( .ZN(net_20178), .A2(net_11267), .A1(net_8640) );
INV_X2 inst_19150 ( .A(net_7111), .ZN(net_4067) );
INV_X4 inst_15453 ( .ZN(net_2488), .A(net_1774) );
NOR2_X2 inst_4205 ( .ZN(net_13187), .A1(net_7858), .A2(net_6742) );
NAND2_X2 inst_11452 ( .ZN(net_9552), .A1(net_8543), .A2(net_3246) );
NAND2_X2 inst_9633 ( .ZN(net_13140), .A1(net_11366), .A2(net_10370) );
INV_X4 inst_17039 ( .ZN(net_14490), .A(net_11968) );
CLKBUF_X2 inst_22859 ( .A(net_22433), .Z(net_22731) );
INV_X4 inst_17465 ( .ZN(net_1330), .A(net_805) );
CLKBUF_X2 inst_22133 ( .A(net_22004), .Z(net_22005) );
AOI22_X2 inst_19989 ( .A1(net_20346), .ZN(net_14982), .B1(net_12053), .B2(net_6388), .A2(net_652) );
INV_X2 inst_18747 ( .A(net_13323), .ZN(net_7875) );
NAND2_X2 inst_12027 ( .ZN(net_1010), .A2(net_1009), .A1(net_103) );
INV_X4 inst_18265 ( .A(net_19437), .ZN(net_19436) );
INV_X2 inst_18495 ( .ZN(net_13378), .A(net_12313) );
NAND2_X2 inst_11063 ( .ZN(net_4527), .A1(net_4526), .A2(net_2641) );
NAND2_X2 inst_9408 ( .ZN(net_20106), .A1(net_11663), .A2(net_11094) );
NAND3_X2 inst_6156 ( .ZN(net_13668), .A3(net_12710), .A2(net_9810), .A1(net_5626) );
DFF_X1 inst_19819 ( .D(net_17781), .CK(net_22554), .Q(x16) );
INV_X4 inst_17999 ( .A(net_21012), .ZN(net_422) );
NOR2_X4 inst_3019 ( .ZN(net_7960), .A1(net_5445), .A2(net_3242) );
OAI21_X2 inst_2327 ( .ZN(net_5318), .A(net_5317), .B2(net_4026), .B1(net_401) );
INV_X4 inst_13430 ( .ZN(net_19148), .A(net_8441) );
NOR2_X2 inst_5078 ( .ZN(net_11389), .A1(net_86), .A2(net_72) );
NAND2_X4 inst_6866 ( .A2(net_20616), .A1(net_20615), .ZN(net_18353) );
INV_X4 inst_14976 ( .ZN(net_3420), .A(net_3419) );
NAND2_X2 inst_11579 ( .ZN(net_2730), .A2(net_2479), .A1(net_252) );
XNOR2_X2 inst_113 ( .ZN(net_18508), .A(net_18417), .B(net_17579) );
INV_X4 inst_17212 ( .ZN(net_701), .A(net_170) );
NAND2_X2 inst_10433 ( .A1(net_9666), .A2(net_8704), .ZN(net_7206) );
CLKBUF_X2 inst_21697 ( .A(net_21568), .Z(net_21569) );
CLKBUF_X2 inst_21669 ( .A(net_21540), .Z(net_21541) );
INV_X4 inst_17217 ( .ZN(net_6314), .A(net_693) );
INV_X4 inst_16751 ( .A(net_10536), .ZN(net_6415) );
INV_X4 inst_14023 ( .A(net_8131), .ZN(net_7633) );
NAND2_X2 inst_9680 ( .ZN(net_10266), .A1(net_10265), .A2(net_10264) );
NAND2_X2 inst_9106 ( .ZN(net_19024), .A2(net_11596), .A1(net_3398) );
NAND2_X2 inst_8479 ( .A2(net_20516), .ZN(net_19958), .A1(net_17006) );
NAND2_X2 inst_10849 ( .ZN(net_10012), .A1(net_6092), .A2(net_5467) );
AOI21_X2 inst_20630 ( .ZN(net_13417), .B1(net_13416), .A(net_11673), .B2(net_8940) );
INV_X2 inst_18633 ( .ZN(net_9429), .A(net_9428) );
NAND2_X4 inst_7298 ( .A2(net_20533), .ZN(net_8758), .A1(net_2282) );
NOR2_X2 inst_4063 ( .ZN(net_9333), .A2(net_7816), .A1(net_1133) );
INV_X2 inst_19655 ( .A(net_20215), .ZN(net_20214) );
NAND2_X2 inst_10069 ( .A1(net_14605), .ZN(net_8660), .A2(net_8659) );
NAND2_X2 inst_8340 ( .ZN(net_19640), .A1(net_17492), .A2(net_17330) );
CLKBUF_X2 inst_21678 ( .A(net_21549), .Z(net_21550) );
INV_X2 inst_19525 ( .ZN(net_9620), .A(net_1061) );
INV_X4 inst_16427 ( .ZN(net_3041), .A(net_146) );
AND2_X2 inst_21329 ( .ZN(net_14437), .A1(net_7230), .A2(net_5525) );
NAND2_X2 inst_9016 ( .ZN(net_20017), .A2(net_12613), .A1(net_238) );
NOR3_X4 inst_2625 ( .A3(net_20060), .A1(net_20059), .ZN(net_19928), .A2(net_11566) );
INV_X4 inst_14088 ( .A(net_6210), .ZN(net_6208) );
NAND3_X2 inst_6064 ( .ZN(net_20660), .A1(net_10760), .A2(net_10739), .A3(net_7899) );
INV_X2 inst_19156 ( .A(net_7090), .ZN(net_3993) );
INV_X4 inst_16081 ( .ZN(net_3083), .A(net_1177) );
INV_X4 inst_12652 ( .ZN(net_17856), .A(net_17855) );
NAND2_X2 inst_9244 ( .ZN(net_19751), .A2(net_13742), .A1(net_11962) );
NOR2_X4 inst_3329 ( .A1(net_317), .ZN(net_273), .A2(net_272) );
NAND3_X2 inst_5769 ( .A3(net_20091), .A1(net_20090), .ZN(net_15896), .A2(net_15404) );
INV_X4 inst_13844 ( .ZN(net_13174), .A(net_7477) );
NOR2_X4 inst_2847 ( .ZN(net_19185), .A2(net_13819), .A1(net_10153) );
OAI21_X4 inst_1442 ( .ZN(net_15784), .A(net_15659), .B2(net_14784), .B1(net_5192) );
XNOR2_X2 inst_332 ( .ZN(net_16997), .A(net_16641), .B(net_6459) );
AOI211_X2 inst_21033 ( .ZN(net_14351), .A(net_14350), .B(net_13789), .C2(net_8641), .C1(net_6536) );
AOI21_X2 inst_20891 ( .B1(net_10183), .ZN(net_7786), .B2(net_6362), .A(net_6353) );
CLKBUF_X2 inst_22099 ( .A(net_21970), .Z(net_21971) );
INV_X4 inst_14192 ( .ZN(net_10539), .A(net_5977) );
NOR2_X2 inst_4013 ( .ZN(net_19845), .A2(net_8070), .A1(net_4893) );
OAI21_X2 inst_2132 ( .ZN(net_9992), .B1(net_6289), .B2(net_4848), .A(net_761) );
OAI22_X2 inst_1289 ( .ZN(net_12882), .A1(net_12881), .B2(net_12880), .A2(net_12842), .B1(net_10031) );
NOR2_X2 inst_4979 ( .ZN(net_3194), .A1(net_1934), .A2(net_1509) );
NOR2_X2 inst_4686 ( .A2(net_5557), .ZN(net_3195), .A1(net_2750) );
NOR2_X2 inst_4869 ( .A1(net_5537), .ZN(net_4171), .A2(net_1123) );
OAI21_X2 inst_1951 ( .ZN(net_12556), .A(net_11550), .B2(net_7533), .B1(net_4442) );
XNOR2_X2 inst_378 ( .A(net_17763), .ZN(net_16834), .B(net_16833) );
INV_X4 inst_17831 ( .ZN(net_1438), .A(net_308) );
NAND2_X4 inst_7444 ( .ZN(net_3431), .A1(net_1064), .A2(net_448) );
NAND2_X2 inst_8151 ( .ZN(net_18013), .A2(net_17980), .A1(net_17973) );
NAND2_X2 inst_11302 ( .ZN(net_9033), .A2(net_3819), .A1(net_3812) );
INV_X4 inst_18205 ( .A(net_21120), .ZN(net_17522) );
NAND2_X2 inst_8750 ( .ZN(net_15963), .A2(net_15801), .A1(net_1951) );
OAI21_X2 inst_2200 ( .A(net_9037), .ZN(net_8562), .B1(net_6002), .B2(net_5252) );
AOI221_X2 inst_20084 ( .ZN(net_15965), .B1(net_15869), .C1(net_15369), .C2(net_15283), .B2(net_14350), .A(net_12777) );
NOR2_X2 inst_4937 ( .ZN(net_2452), .A1(net_1470), .A2(net_112) );
AOI22_X2 inst_19980 ( .ZN(net_15392), .B1(net_15270), .A2(net_13969), .B2(net_5666), .A1(net_1869) );
NAND2_X2 inst_10320 ( .ZN(net_7823), .A1(net_7822), .A2(net_4678) );
NAND2_X2 inst_8284 ( .A2(net_20461), .ZN(net_19605), .A1(net_17441) );
NAND2_X2 inst_8080 ( .A1(net_18153), .ZN(net_18151), .A2(net_16912) );
NAND2_X2 inst_9948 ( .A1(net_9082), .ZN(net_8943), .A2(net_8942) );
INV_X4 inst_14707 ( .ZN(net_18576), .A(net_18025) );
XNOR2_X2 inst_250 ( .ZN(net_17313), .A(net_17312), .B(net_12269) );
NAND2_X2 inst_9275 ( .ZN(net_15024), .A1(net_14363), .A2(net_12616) );
CLKBUF_X2 inst_22363 ( .A(net_22176), .Z(net_22235) );
NAND2_X2 inst_7708 ( .ZN(net_18860), .A2(net_18853), .A1(net_18841) );
NAND3_X2 inst_5762 ( .ZN(net_15941), .A3(net_15218), .A1(net_14880), .A2(net_12955) );
CLKBUF_X2 inst_22257 ( .A(net_22128), .Z(net_22129) );
NAND3_X2 inst_6595 ( .ZN(net_9912), .A3(net_9911), .A1(net_6852), .A2(net_6231) );
NAND2_X2 inst_9384 ( .ZN(net_11936), .A2(net_8925), .A1(net_7918) );
OAI21_X2 inst_1523 ( .A(net_18582), .ZN(net_18064), .B1(net_18033), .B2(net_18028) );
NAND2_X2 inst_9941 ( .ZN(net_9091), .A1(net_9090), .A2(net_5816) );
INV_X4 inst_17787 ( .A(net_703), .ZN(net_409) );
SDFF_X2 inst_1048 ( .QN(net_20996), .D(net_1859), .SE(net_253), .CK(net_21820), .SI(x3090) );
NAND2_X4 inst_7120 ( .ZN(net_12636), .A1(net_10974), .A2(net_5632) );
INV_X4 inst_16822 ( .ZN(net_1312), .A(net_769) );
DFF_X1 inst_19902 ( .D(net_16995), .CK(net_22349), .Q(x856) );
INV_X2 inst_18429 ( .ZN(net_19734), .A(net_14323) );
INV_X4 inst_13537 ( .A(net_9209), .ZN(net_9208) );
AOI21_X2 inst_20333 ( .ZN(net_15819), .B1(net_15818), .B2(net_14919), .A(net_11835) );
OAI21_X2 inst_2270 ( .A(net_10142), .ZN(net_7142), .B1(net_5553), .B2(net_3473) );
INV_X4 inst_16050 ( .ZN(net_4482), .A(net_2317) );
NAND2_X2 inst_11624 ( .ZN(net_11292), .A1(net_2539), .A2(net_1537) );
OAI211_X2 inst_2401 ( .ZN(net_15935), .B(net_15208), .C1(net_15198), .C2(net_11323), .A(net_9898) );
AOI21_X4 inst_20202 ( .ZN(net_14814), .B1(net_14813), .B2(net_14241), .A(net_11341) );
INV_X4 inst_12979 ( .A(net_18214), .ZN(net_16882) );
NAND2_X2 inst_10092 ( .ZN(net_8621), .A2(net_6385), .A1(net_1894) );
INV_X4 inst_14723 ( .ZN(net_4149), .A(net_4148) );
INV_X4 inst_12649 ( .ZN(net_20704), .A(net_17870) );
NAND2_X2 inst_9356 ( .A1(net_13984), .ZN(net_12154), .A2(net_8805) );
NAND2_X2 inst_8367 ( .ZN(net_19932), .A2(net_17348), .A1(net_17126) );
INV_X2 inst_19548 ( .A(net_7230), .ZN(net_918) );
NAND2_X2 inst_8015 ( .ZN(net_18289), .A2(net_18239), .A1(net_17193) );
INV_X4 inst_15564 ( .ZN(net_3753), .A(net_2442) );
NAND2_X2 inst_8196 ( .ZN(net_17891), .A1(net_17890), .A2(net_17889) );
AND2_X4 inst_21196 ( .ZN(net_19582), .A1(net_10182), .A2(net_10181) );
NAND3_X2 inst_6050 ( .ZN(net_14239), .A3(net_13560), .A1(net_12602), .A2(net_9711) );
INV_X4 inst_14287 ( .ZN(net_7321), .A(net_5607) );
NAND3_X2 inst_6204 ( .ZN(net_13300), .A1(net_13164), .A3(net_10295), .A2(net_9921) );
INV_X4 inst_17351 ( .ZN(net_15452), .A(net_1471) );
NAND2_X2 inst_8618 ( .ZN(net_16610), .A2(net_16437), .A1(net_543) );
CLKBUF_X2 inst_21748 ( .A(net_21619), .Z(net_21620) );
NAND2_X2 inst_9710 ( .ZN(net_15413), .A1(net_10191), .A2(net_10190) );
XNOR2_X2 inst_420 ( .ZN(net_16531), .A(net_16530), .B(net_5237) );
NOR2_X2 inst_3992 ( .ZN(net_11667), .A1(net_8722), .A2(net_4993) );
INV_X4 inst_12522 ( .ZN(net_18491), .A(net_18490) );
NOR2_X4 inst_3265 ( .ZN(net_2078), .A1(net_2077), .A2(net_2076) );
CLKBUF_X2 inst_22071 ( .A(net_21561), .Z(net_21943) );
INV_X4 inst_15669 ( .ZN(net_4016), .A(net_2054) );
NAND2_X4 inst_7558 ( .ZN(net_3177), .A1(net_1608), .A2(net_61) );
OAI22_X2 inst_1305 ( .ZN(net_10448), .A1(net_10447), .A2(net_10446), .B1(net_10445), .B2(net_10444) );
NAND2_X2 inst_7997 ( .ZN(net_20718), .A2(net_18201), .A1(net_17234) );
CLKBUF_X2 inst_21858 ( .A(net_21729), .Z(net_21730) );
AND2_X4 inst_21254 ( .A1(net_20851), .A2(net_4030), .ZN(net_2449) );
XNOR2_X2 inst_314 ( .ZN(net_20377), .B(net_16698), .A(net_16679) );
INV_X4 inst_14813 ( .ZN(net_5255), .A(net_3948) );
NAND2_X2 inst_8713 ( .A1(net_21212), .ZN(net_16233), .A2(net_16052) );
NOR2_X4 inst_3225 ( .ZN(net_2586), .A2(net_2391), .A1(net_1697) );
INV_X4 inst_13367 ( .ZN(net_12324), .A(net_10909) );
INV_X4 inst_15342 ( .ZN(net_11366), .A(net_10389) );
XNOR2_X2 inst_597 ( .A(net_21129), .ZN(net_9240), .B(net_615) );
NAND3_X2 inst_6161 ( .ZN(net_13643), .A2(net_13580), .A3(net_13304), .A1(net_12397) );
NAND3_X4 inst_5524 ( .A3(net_20421), .A1(net_20420), .ZN(net_18192), .A2(net_13100) );
NAND2_X4 inst_7257 ( .ZN(net_7919), .A1(net_6633), .A2(net_5875) );
NAND2_X2 inst_11859 ( .ZN(net_12050), .A1(net_8596), .A2(net_7432) );
NAND2_X4 inst_6927 ( .A2(net_19010), .A1(net_19009), .ZN(net_17738) );
INV_X4 inst_15115 ( .ZN(net_13177), .A(net_7128) );
INV_X8 inst_12272 ( .ZN(net_2641), .A(net_1310) );
INV_X4 inst_16985 ( .ZN(net_883), .A(net_882) );
CLKBUF_X2 inst_21406 ( .A(net_21268), .Z(net_21278) );
XNOR2_X2 inst_472 ( .A(net_13655), .ZN(net_11890), .B(net_2507) );
XNOR2_X2 inst_447 ( .ZN(net_14916), .B(net_14915), .A(net_12873) );
NOR2_X2 inst_4533 ( .ZN(net_6860), .A2(net_3963), .A1(net_85) );
NAND3_X2 inst_5987 ( .ZN(net_18986), .A2(net_14537), .A1(net_13346), .A3(net_12013) );
INV_X4 inst_12872 ( .ZN(net_17275), .A(net_16950) );
INV_X4 inst_16940 ( .ZN(net_921), .A(net_920) );
NOR3_X4 inst_2623 ( .A3(net_20119), .A1(net_20118), .ZN(net_19967), .A2(net_10877) );
OAI21_X4 inst_1391 ( .A(net_20968), .B2(net_19725), .B1(net_19724), .ZN(net_16306) );
XNOR2_X2 inst_665 ( .A(net_21199), .B(net_21135), .ZN(net_240) );
AOI22_X2 inst_19975 ( .B1(net_15506), .ZN(net_15489), .A1(net_14788), .A2(net_14571), .B2(net_9952) );
NOR2_X2 inst_4843 ( .A1(net_20530), .ZN(net_4167), .A2(net_1117) );
CLKBUF_X2 inst_22615 ( .A(net_22486), .Z(net_22487) );
AOI21_X4 inst_20112 ( .B2(net_20928), .B1(net_19504), .ZN(net_16320), .A(net_12119) );
INV_X4 inst_16831 ( .A(net_3818), .ZN(net_1147) );
INV_X4 inst_12929 ( .ZN(net_17022), .A(net_16655) );
NAND2_X2 inst_12014 ( .A2(net_3056), .ZN(net_1400), .A1(net_1099) );
NAND2_X2 inst_10219 ( .ZN(net_14387), .A2(net_7948), .A1(net_6947) );
NOR2_X2 inst_3538 ( .ZN(net_13415), .A1(net_11664), .A2(net_10628) );
CLKBUF_X2 inst_21670 ( .A(net_21541), .Z(net_21542) );
NOR2_X2 inst_3755 ( .ZN(net_10384), .A2(net_9448), .A1(net_8894) );
NAND2_X2 inst_8718 ( .ZN(net_16188), .A1(net_16187), .A2(net_15980) );
NAND2_X2 inst_9810 ( .A1(net_14022), .ZN(net_9679), .A2(net_7202) );
OR2_X2 inst_1196 ( .A1(net_4508), .ZN(net_3958), .A2(net_3957) );
INV_X4 inst_17899 ( .A(net_20859), .ZN(net_167) );
INV_X4 inst_13815 ( .ZN(net_11114), .A(net_7527) );
INV_X4 inst_18154 ( .A(net_21087), .ZN(net_370) );
NOR2_X2 inst_3428 ( .ZN(net_15424), .A2(net_15040), .A1(net_14167) );
NAND2_X2 inst_10510 ( .ZN(net_12787), .A2(net_11113), .A1(net_9966) );
CLKBUF_X2 inst_21513 ( .A(net_21384), .Z(net_21385) );
NOR2_X4 inst_3336 ( .ZN(net_913), .A1(net_459), .A2(net_121) );
NAND2_X2 inst_7963 ( .ZN(net_18370), .A2(net_18363), .A1(net_17866) );
CLKBUF_X2 inst_21910 ( .A(net_21781), .Z(net_21782) );
INV_X2 inst_19043 ( .ZN(net_4761), .A(net_4760) );
NAND2_X2 inst_9034 ( .ZN(net_14067), .A2(net_12090), .A1(net_3376) );
INV_X4 inst_16625 ( .ZN(net_1478), .A(net_1229) );
NOR2_X4 inst_2837 ( .ZN(net_19194), .A2(net_14199), .A1(net_13409) );
NAND2_X4 inst_7115 ( .ZN(net_11051), .A1(net_11020), .A2(net_9396) );
INV_X2 inst_19580 ( .ZN(net_870), .A(net_298) );
OAI21_X2 inst_1845 ( .ZN(net_14018), .A(net_10891), .B2(net_10333), .B1(net_9092) );
INV_X4 inst_17847 ( .A(net_308), .ZN(net_97) );
INV_X4 inst_14681 ( .A(net_9569), .ZN(net_4300) );
NAND2_X2 inst_9296 ( .ZN(net_13439), .A1(net_10914), .A2(net_9211) );
INV_X4 inst_15598 ( .ZN(net_3452), .A(net_2887) );
NAND2_X4 inst_6905 ( .ZN(net_17919), .A1(net_17750), .A2(net_17656) );
OAI21_X4 inst_1429 ( .A(net_16210), .ZN(net_16023), .B2(net_15418), .B1(net_15201) );
NAND2_X2 inst_8439 ( .ZN(net_17270), .A2(net_16828), .A1(net_16673) );
INV_X16 inst_19739 ( .ZN(net_1192), .A(net_181) );
INV_X4 inst_12919 ( .A(net_16665), .ZN(net_16664) );
XNOR2_X2 inst_586 ( .B(net_9235), .ZN(net_577), .A(net_576) );
NAND4_X4 inst_5220 ( .ZN(net_17290), .A4(net_16181), .A1(net_16083), .A3(net_15993), .A2(net_10821) );
AOI21_X2 inst_20310 ( .ZN(net_16034), .B1(net_15842), .A(net_15575), .B2(net_15517) );
NAND2_X2 inst_9828 ( .ZN(net_9622), .A1(net_8759), .A2(net_8504) );
NAND2_X4 inst_7176 ( .ZN(net_14844), .A2(net_8334), .A1(net_7475) );
NAND2_X2 inst_10563 ( .A1(net_9109), .ZN(net_8772), .A2(net_6842) );
OAI211_X2 inst_2591 ( .ZN(net_5296), .B(net_5295), .A(net_2679), .C2(net_1405), .C1(net_1242) );
INV_X4 inst_15317 ( .A(net_3850), .ZN(net_2638) );
NOR3_X2 inst_2652 ( .A3(net_19679), .A1(net_19678), .ZN(net_19076), .A2(net_12655) );
NAND4_X4 inst_5221 ( .A3(net_18876), .A1(net_18875), .ZN(net_16602), .A4(net_16183), .A2(net_16116) );
OR2_X2 inst_1203 ( .ZN(net_3598), .A1(net_3452), .A2(net_2886) );
AND2_X4 inst_21171 ( .ZN(net_19829), .A1(net_14547), .A2(net_7236) );
SDFF_X2 inst_802 ( .Q(net_21241), .SI(net_17975), .SE(net_125), .CK(net_21570), .D(x6680) );
XNOR2_X2 inst_296 ( .B(net_21164), .ZN(net_17124), .A(net_17123) );
INV_X4 inst_16229 ( .ZN(net_9997), .A(net_6635) );
INV_X4 inst_14626 ( .ZN(net_18865), .A(net_18025) );
NOR2_X2 inst_4370 ( .ZN(net_20403), .A1(net_5487), .A2(net_3902) );
NAND2_X2 inst_11218 ( .ZN(net_5051), .A1(net_4918), .A2(net_4315) );
NAND2_X2 inst_9185 ( .A1(net_15706), .ZN(net_13133), .A2(net_13132) );
NAND2_X2 inst_11047 ( .ZN(net_7795), .A1(net_4715), .A2(net_3533) );
CLKBUF_X2 inst_22452 ( .A(net_22323), .Z(net_22324) );
NOR2_X2 inst_3943 ( .ZN(net_8643), .A1(net_8642), .A2(net_8641) );
INV_X4 inst_14280 ( .ZN(net_6261), .A(net_5651) );
OAI211_X2 inst_2532 ( .C1(net_13938), .ZN(net_11265), .A(net_11264), .C2(net_11263), .B(net_5197) );
INV_X4 inst_13263 ( .ZN(net_12678), .A(net_12677) );
OAI211_X2 inst_2463 ( .ZN(net_14146), .B(net_14145), .A(net_10144), .C2(net_9202), .C1(net_3274) );
INV_X4 inst_17267 ( .A(net_14678), .ZN(net_11404) );
NAND2_X2 inst_11206 ( .ZN(net_10355), .A1(net_9925), .A2(net_3129) );
NAND2_X2 inst_10907 ( .ZN(net_12221), .A1(net_5374), .A2(net_5373) );
NAND3_X4 inst_5610 ( .A3(net_19779), .A1(net_19778), .ZN(net_14117), .A2(net_7953) );
AOI211_X2 inst_21057 ( .C1(net_12852), .ZN(net_11210), .A(net_11209), .B(net_11208), .C2(net_11207) );
OAI21_X4 inst_1464 ( .ZN(net_15179), .B1(net_15178), .B2(net_13903), .A(net_13022) );
INV_X4 inst_15536 ( .ZN(net_3199), .A(net_2374) );
INV_X4 inst_12778 ( .ZN(net_17561), .A(net_17490) );
NAND2_X2 inst_8490 ( .A1(net_16959), .ZN(net_16957), .A2(net_16560) );
INV_X2 inst_19573 ( .A(net_3482), .ZN(net_702) );
NOR2_X2 inst_5031 ( .ZN(net_1763), .A2(net_1270), .A1(net_907) );
INV_X2 inst_19002 ( .A(net_9956), .ZN(net_5048) );
INV_X4 inst_17656 ( .ZN(net_14568), .A(net_14029) );
AND2_X2 inst_21284 ( .ZN(net_13104), .A1(net_13103), .A2(net_13102) );
INV_X4 inst_13498 ( .A(net_10117), .ZN(net_9439) );
INV_X4 inst_13215 ( .ZN(net_13638), .A(net_12815) );
AOI21_X2 inst_20424 ( .ZN(net_15212), .B1(net_14684), .B2(net_13894), .A(net_12649) );
NAND3_X2 inst_6441 ( .A2(net_12036), .ZN(net_11810), .A3(net_9061), .A1(net_5531) );
OAI22_X2 inst_1308 ( .A1(net_13752), .B1(net_12339), .ZN(net_9009), .B2(net_9008), .A2(net_8975) );
NOR2_X4 inst_3070 ( .ZN(net_8071), .A2(net_4784), .A1(net_411) );
XNOR2_X2 inst_85 ( .ZN(net_18569), .A(net_18506), .B(net_17757) );
NOR2_X2 inst_4733 ( .A1(net_5459), .ZN(net_3964), .A2(net_3070) );
AOI21_X2 inst_20973 ( .ZN(net_4667), .A(net_4666), .B2(net_4615), .B1(net_1170) );
INV_X4 inst_16949 ( .ZN(net_1395), .A(net_940) );
AOI21_X2 inst_20453 ( .ZN(net_15062), .B1(net_13416), .B2(net_13008), .A(net_7699) );
NAND3_X2 inst_5963 ( .ZN(net_14804), .A3(net_13492), .A1(net_10692), .A2(net_6865) );
AOI21_X2 inst_20771 ( .B1(net_19954), .ZN(net_10677), .A(net_10676), .B2(net_6624) );
DFF_X1 inst_19892 ( .D(net_16877), .CK(net_22080), .Q(x353) );
CLKBUF_X2 inst_22723 ( .A(net_21273), .Z(net_22595) );
INV_X4 inst_14693 ( .ZN(net_4278), .A(net_4277) );
NAND2_X2 inst_9681 ( .ZN(net_10262), .A1(net_10261), .A2(net_10260) );
INV_X4 inst_16310 ( .ZN(net_2299), .A(net_1456) );
NAND2_X2 inst_11850 ( .ZN(net_7743), .A1(net_1698), .A2(net_913) );
INV_X4 inst_12598 ( .ZN(net_18171), .A(net_18142) );
NAND2_X2 inst_11314 ( .A1(net_4074), .ZN(net_3772), .A2(net_3771) );
NOR2_X2 inst_4022 ( .ZN(net_12259), .A1(net_8748), .A2(net_6247) );
AOI21_X2 inst_20721 ( .ZN(net_11985), .B1(net_11442), .B2(net_7722), .A(net_3305) );
OAI21_X2 inst_1978 ( .A(net_13089), .ZN(net_12145), .B2(net_8234), .B1(net_5713) );
XNOR2_X2 inst_290 ( .B(net_21128), .A(net_19452), .ZN(net_17135) );
INV_X4 inst_15285 ( .A(net_3872), .ZN(net_2722) );
DFF_X1 inst_19827 ( .D(net_17593), .CK(net_21617), .Q(x648) );
INV_X4 inst_16346 ( .A(net_15697), .ZN(net_1296) );
INV_X4 inst_14122 ( .ZN(net_8154), .A(net_5529) );
OAI21_X2 inst_2112 ( .ZN(net_10038), .A(net_10037), .B2(net_8372), .B1(net_5001) );
NAND2_X2 inst_7743 ( .ZN(net_18797), .A2(net_18764), .A1(net_17721) );
INV_X4 inst_16610 ( .ZN(net_19826), .A(net_1314) );
INV_X4 inst_15431 ( .A(net_14493), .ZN(net_14051) );
NOR2_X4 inst_3036 ( .ZN(net_6269), .A1(net_5131), .A2(net_2431) );
SDFF_X2 inst_814 ( .Q(net_21239), .SI(net_17794), .SE(net_945), .CK(net_21566), .D(x6710) );
AND2_X4 inst_21208 ( .ZN(net_7055), .A1(net_7054), .A2(net_6558) );
INV_X4 inst_13441 ( .ZN(net_9805), .A(net_9804) );
NAND2_X2 inst_9465 ( .A2(net_20764), .ZN(net_13770), .A1(net_10898) );
INV_X2 inst_19007 ( .ZN(net_5022), .A(net_5021) );
NAND4_X4 inst_5203 ( .A2(net_18947), .A1(net_18946), .A3(net_18940), .ZN(net_16439), .A4(net_16325) );
NAND2_X2 inst_8973 ( .ZN(net_14517), .A2(net_13013), .A1(net_2355) );
NOR2_X2 inst_3471 ( .ZN(net_14457), .A1(net_14456), .A2(net_12773) );
OAI21_X4 inst_1458 ( .ZN(net_20745), .B2(net_19401), .B1(net_19400), .A(net_15119) );
INV_X4 inst_15933 ( .A(net_11376), .ZN(net_8983) );
NAND2_X2 inst_11332 ( .ZN(net_9951), .A1(net_9581), .A2(net_3751) );
OAI21_X2 inst_2275 ( .ZN(net_7134), .B2(net_7133), .A(net_6471), .B1(net_5677) );
INV_X4 inst_16650 ( .A(net_4305), .ZN(net_2909) );
INV_X4 inst_15727 ( .ZN(net_3872), .A(net_1460) );
NAND2_X2 inst_10212 ( .ZN(net_19236), .A1(net_8094), .A2(net_8093) );
INV_X4 inst_16567 ( .A(net_11407), .ZN(net_10891) );
SDFF_X2 inst_822 ( .Q(net_21181), .SI(net_17647), .SE(net_125), .CK(net_22331), .D(x6585) );
NAND2_X2 inst_12053 ( .A2(net_20876), .ZN(net_1205), .A1(net_973) );
OR2_X4 inst_1125 ( .ZN(net_6002), .A2(net_1790), .A1(net_77) );
NOR2_X2 inst_4341 ( .ZN(net_5686), .A1(net_4289), .A2(net_4223) );
NAND3_X2 inst_5996 ( .ZN(net_14440), .A2(net_14439), .A1(net_12786), .A3(net_11262) );
NAND2_X2 inst_10984 ( .ZN(net_8095), .A1(net_6598), .A2(net_3532) );
XNOR2_X2 inst_609 ( .B(net_17426), .ZN(net_510), .A(net_509) );
NAND2_X2 inst_11521 ( .ZN(net_4987), .A2(net_2980), .A1(net_170) );
NAND2_X2 inst_8261 ( .A2(net_19654), .ZN(net_17687), .A1(net_17686) );
SDFF_X2 inst_795 ( .Q(net_20887), .SE(net_18859), .SI(net_18008), .D(net_559), .CK(net_22770) );
OAI211_X2 inst_2491 ( .ZN(net_13162), .B(net_13161), .A(net_12809), .C2(net_11281), .C1(net_4437) );
NAND3_X2 inst_6668 ( .ZN(net_7918), .A1(net_7917), .A2(net_6854), .A3(net_5910) );
AOI21_X2 inst_20781 ( .B1(net_13080), .A(net_11317), .ZN(net_10559), .B2(net_6419) );
INV_X4 inst_14127 ( .ZN(net_9690), .A(net_6114) );
NAND2_X2 inst_11179 ( .ZN(net_8399), .A1(net_6611), .A2(net_4123) );
INV_X4 inst_12848 ( .ZN(net_17076), .A(net_17075) );
NAND2_X2 inst_8215 ( .ZN(net_17844), .A2(net_17843), .A1(net_6375) );
XNOR2_X2 inst_619 ( .ZN(net_14917), .A(net_670), .B(net_481) );
CLKBUF_X2 inst_21420 ( .A(net_21291), .Z(net_21292) );
INV_X4 inst_14481 ( .ZN(net_5847), .A(net_4871) );
NAND2_X1 inst_12139 ( .A1(net_19454), .ZN(net_17349), .A2(net_17348) );
OAI21_X2 inst_1654 ( .ZN(net_19934), .A(net_15451), .B1(net_15224), .B2(net_12579) );
CLKBUF_X2 inst_21966 ( .A(net_21837), .Z(net_21838) );
NOR2_X2 inst_4547 ( .ZN(net_6920), .A1(net_4052), .A2(net_3977) );
NAND2_X2 inst_7831 ( .ZN(net_19164), .A2(net_18649), .A1(net_17372) );
NAND2_X2 inst_10545 ( .ZN(net_12140), .A1(net_7246), .A2(net_3860) );
CLKBUF_X2 inst_21751 ( .A(net_21490), .Z(net_21623) );
NAND2_X2 inst_10553 ( .ZN(net_15425), .A2(net_6730), .A1(net_5415) );
CLKBUF_X2 inst_21476 ( .A(net_21347), .Z(net_21348) );
AOI22_X2 inst_20035 ( .B1(net_10989), .ZN(net_8459), .A2(net_6995), .B2(net_3670), .A1(net_761) );
CLKBUF_X2 inst_21956 ( .A(net_21827), .Z(net_21828) );
NAND2_X2 inst_10265 ( .ZN(net_7986), .A1(net_7985), .A2(net_7984) );
NAND3_X2 inst_6486 ( .ZN(net_11196), .A2(net_11195), .A3(net_11194), .A1(net_4234) );
OAI21_X2 inst_2076 ( .ZN(net_10586), .A(net_9076), .B2(net_6390), .B1(net_5449) );
INV_X2 inst_18896 ( .ZN(net_20427), .A(net_7960) );
NAND3_X2 inst_5879 ( .ZN(net_15283), .A1(net_14225), .A3(net_11210), .A2(net_9545) );
INV_X4 inst_16835 ( .ZN(net_14994), .A(net_13089) );
OAI211_X2 inst_2481 ( .ZN(net_13487), .B(net_13486), .C2(net_12569), .A(net_7502), .C1(net_2616) );
CLKBUF_X2 inst_21782 ( .A(net_21653), .Z(net_21654) );
NAND2_X2 inst_7824 ( .ZN(net_18646), .A1(net_18645), .A2(net_17435) );
NAND2_X2 inst_11474 ( .ZN(net_4077), .A2(net_2237), .A1(net_693) );
INV_X4 inst_13385 ( .ZN(net_20752), .A(net_10764) );
NOR2_X2 inst_4285 ( .ZN(net_6051), .A1(net_5455), .A2(net_4293) );
INV_X4 inst_15386 ( .ZN(net_7133), .A(net_2551) );
OR2_X2 inst_1162 ( .A2(net_10012), .ZN(net_8661), .A1(net_81) );
INV_X2 inst_18829 ( .ZN(net_6787), .A(net_6786) );
NAND2_X4 inst_7485 ( .ZN(net_4136), .A1(net_2490), .A2(net_2489) );
INV_X4 inst_14384 ( .A(net_7008), .ZN(net_5163) );
NAND3_X2 inst_6108 ( .ZN(net_19179), .A3(net_13764), .A1(net_11413), .A2(net_6103) );
NAND3_X2 inst_6572 ( .ZN(net_10464), .A2(net_9072), .A3(net_8782), .A1(net_5395) );
INV_X4 inst_13123 ( .ZN(net_15404), .A(net_15147) );
NAND2_X4 inst_7449 ( .A1(net_19669), .ZN(net_3918), .A2(net_2456) );
NOR2_X4 inst_2973 ( .ZN(net_9806), .A1(net_3308), .A2(net_1725) );
CLKBUF_X2 inst_22493 ( .A(net_21912), .Z(net_22365) );
NAND2_X2 inst_11454 ( .A1(net_10714), .ZN(net_3806), .A2(net_2669) );
INV_X4 inst_17297 ( .ZN(net_1133), .A(net_612) );
OAI21_X4 inst_1433 ( .B2(net_19597), .B1(net_19596), .A(net_16347), .ZN(net_15992) );
SDFF_X2 inst_793 ( .Q(net_20886), .SE(net_18862), .SI(net_18015), .D(net_747), .CK(net_22774) );
INV_X2 inst_18923 ( .ZN(net_5921), .A(net_5920) );
CLKBUF_X2 inst_21823 ( .A(net_21694), .Z(net_21695) );
NOR2_X2 inst_4815 ( .A2(net_3326), .ZN(net_2577), .A1(net_2576) );
OAI21_X2 inst_1999 ( .ZN(net_11850), .B2(net_11849), .A(net_8367), .B1(net_2212) );
NOR3_X2 inst_2733 ( .ZN(net_12823), .A2(net_12805), .A3(net_11574), .A1(net_7215) );
INV_X8 inst_12405 ( .ZN(net_20702), .A(net_322) );
NAND2_X2 inst_11750 ( .ZN(net_3286), .A2(net_2117), .A1(net_1848) );
CLKBUF_X2 inst_22193 ( .A(net_22064), .Z(net_22065) );
INV_X4 inst_15429 ( .A(net_11494), .ZN(net_8981) );
NAND2_X2 inst_8808 ( .ZN(net_15621), .A1(net_14963), .A2(net_14696) );
INV_X4 inst_17225 ( .ZN(net_904), .A(net_690) );
XNOR2_X2 inst_475 ( .ZN(net_11883), .A(net_11882), .B(net_2030) );
INV_X4 inst_13253 ( .ZN(net_12760), .A(net_11745) );
NAND2_X2 inst_9436 ( .ZN(net_11588), .A2(net_11587), .A1(net_10735) );
INV_X2 inst_19020 ( .A(net_8504), .ZN(net_4957) );
INV_X4 inst_17958 ( .A(net_20996), .ZN(net_1859) );
NOR2_X2 inst_4738 ( .ZN(net_3920), .A2(net_3065), .A1(net_1259) );
NAND2_X2 inst_9412 ( .A2(net_12995), .ZN(net_11657), .A1(net_11656) );
INV_X4 inst_17917 ( .ZN(net_10514), .A(net_60) );
NOR2_X2 inst_4412 ( .ZN(net_6187), .A1(net_5652), .A2(net_3890) );
INV_X4 inst_12595 ( .A(net_18098), .ZN(net_18097) );
AND3_X2 inst_21148 ( .A2(net_14684), .A3(net_12884), .A1(net_9834), .ZN(net_5323) );
AOI21_X2 inst_20323 ( .ZN(net_15859), .B1(net_15858), .B2(net_15311), .A(net_5446) );
NAND2_X2 inst_9564 ( .ZN(net_12657), .A1(net_9183), .A2(net_7373) );
INV_X4 inst_12804 ( .A(net_18478), .ZN(net_18451) );
INV_X4 inst_15573 ( .ZN(net_10229), .A(net_9260) );
NAND3_X2 inst_5724 ( .ZN(net_20138), .A3(net_15668), .A1(net_14026), .A2(net_12686) );
NAND2_X2 inst_8276 ( .ZN(net_17635), .A2(net_17462), .A1(net_17342) );
NOR2_X2 inst_4331 ( .ZN(net_5782), .A1(net_5781), .A2(net_3041) );
NAND2_X2 inst_11054 ( .ZN(net_4678), .A2(net_4677), .A1(net_3190) );
NAND2_X2 inst_8049 ( .ZN(net_18227), .A2(net_18226), .A1(net_17431) );
DFF_X1 inst_19846 ( .D(net_17218), .CK(net_22378), .Q(x683) );
NOR2_X2 inst_4705 ( .A1(net_5748), .ZN(net_3972), .A2(net_3168) );
NAND2_X2 inst_10940 ( .ZN(net_8378), .A2(net_5170), .A1(net_2976) );
AOI21_X2 inst_20591 ( .ZN(net_13937), .B2(net_11197), .B1(net_10920), .A(net_8803) );
NAND2_X2 inst_11543 ( .ZN(net_2911), .A1(net_1668), .A2(net_1201) );
INV_X4 inst_16178 ( .ZN(net_11678), .A(net_1777) );
INV_X4 inst_16320 ( .A(net_2841), .ZN(net_1431) );
NOR2_X2 inst_3580 ( .ZN(net_12686), .A2(net_12659), .A1(net_9704) );
INV_X8 inst_12321 ( .ZN(net_1237), .A(net_709) );
NAND2_X2 inst_11531 ( .ZN(net_3683), .A1(net_2934), .A2(net_2581) );
NAND2_X2 inst_10004 ( .A1(net_9751), .ZN(net_8816), .A2(net_5464) );
NOR2_X4 inst_3080 ( .ZN(net_6045), .A1(net_1877), .A2(net_925) );
NAND2_X4 inst_6857 ( .ZN(net_18423), .A2(net_18364), .A1(net_18305) );
INV_X2 inst_19181 ( .ZN(net_8377), .A(net_3775) );
OAI211_X2 inst_2434 ( .ZN(net_15013), .C1(net_15012), .C2(net_13876), .B(net_12772), .A(net_11003) );
NAND2_X4 inst_7432 ( .ZN(net_6243), .A1(net_3409), .A2(net_1365) );
OR2_X4 inst_1107 ( .A2(net_1886), .ZN(net_1530), .A1(net_1529) );
NAND2_X2 inst_10039 ( .ZN(net_13128), .A1(net_8720), .A2(net_8134) );
INV_X4 inst_15335 ( .ZN(net_4821), .A(net_2808) );
INV_X4 inst_12909 ( .A(net_16698), .ZN(net_16697) );
NAND3_X2 inst_5930 ( .ZN(net_14930), .A2(net_14929), .A1(net_13636), .A3(net_13510) );
AOI21_X2 inst_20724 ( .ZN(net_11967), .B2(net_10155), .B1(net_9824), .A(net_178) );
NAND2_X2 inst_9916 ( .ZN(net_12744), .A2(net_9348), .A1(net_9309) );
AOI211_X2 inst_21016 ( .ZN(net_15554), .C1(net_15553), .C2(net_14583), .B(net_13042), .A(net_8754) );
INV_X4 inst_18288 ( .A(net_20213), .ZN(net_20212) );
NOR2_X2 inst_4253 ( .A1(net_7450), .ZN(net_6337), .A2(net_6336) );
NOR3_X2 inst_2776 ( .A2(net_14675), .A3(net_8981), .A1(net_8378), .ZN(net_7765) );
INV_X2 inst_19474 ( .A(net_5265), .ZN(net_3960) );
NAND2_X2 inst_9646 ( .ZN(net_19390), .A1(net_10376), .A2(net_10375) );
AOI21_X2 inst_20754 ( .ZN(net_11232), .B1(net_10386), .B2(net_9683), .A(net_6232) );
NAND2_X2 inst_8612 ( .ZN(net_16617), .A2(net_16441), .A1(net_595) );
SDFF_X2 inst_746 ( .Q(net_20871), .SE(net_18856), .SI(net_18541), .D(net_462), .CK(net_22177) );
INV_X4 inst_13016 ( .ZN(net_18960), .A(net_16398) );
NAND3_X2 inst_6553 ( .ZN(net_10528), .A1(net_7662), .A3(net_7261), .A2(net_6837) );
INV_X4 inst_17618 ( .ZN(net_6838), .A(net_1815) );
NAND2_X2 inst_8660 ( .ZN(net_19668), .A2(net_16526), .A1(net_670) );
OAI21_X2 inst_2267 ( .A(net_9148), .ZN(net_7152), .B1(net_7151), .B2(net_3954) );
INV_X2 inst_18722 ( .A(net_8708), .ZN(net_8124) );
NAND2_X4 inst_7127 ( .ZN(net_20079), .A2(net_11270), .A1(net_10888) );
INV_X4 inst_18019 ( .A(net_21048), .ZN(net_581) );
INV_X4 inst_17664 ( .ZN(net_795), .A(net_289) );
NAND3_X2 inst_5662 ( .ZN(net_16419), .A1(net_16356), .A2(net_14844), .A3(net_12240) );
NAND2_X2 inst_7893 ( .ZN(net_18495), .A2(net_18490), .A1(net_17873) );
INV_X4 inst_16299 ( .A(net_11297), .ZN(net_10206) );
NAND2_X2 inst_10050 ( .A1(net_14552), .ZN(net_12184), .A2(net_8694) );
NAND3_X2 inst_5820 ( .ZN(net_15593), .A1(net_14888), .A3(net_13458), .A2(net_10768) );
NAND2_X2 inst_8721 ( .A1(net_20968), .ZN(net_16151), .A2(net_15895) );
OAI21_X2 inst_1577 ( .A(net_20872), .B2(net_19562), .B1(net_19561), .ZN(net_16316) );
NAND2_X2 inst_7722 ( .ZN(net_18836), .A2(net_18813), .A1(net_18797) );
OR2_X4 inst_1110 ( .ZN(net_8559), .A2(net_90), .A1(net_81) );
NAND3_X2 inst_5778 ( .ZN(net_15854), .A1(net_15344), .A3(net_15304), .A2(net_9026) );
INV_X2 inst_18607 ( .ZN(net_9725), .A(net_9724) );
INV_X4 inst_14870 ( .ZN(net_18859), .A(net_18025) );
NOR2_X4 inst_2873 ( .ZN(net_12305), .A2(net_10873), .A1(net_4702) );
NAND2_X2 inst_8468 ( .ZN(net_17033), .A1(net_16699), .A2(net_16545) );
OAI211_X2 inst_2442 ( .ZN(net_14821), .C1(net_13926), .C2(net_13728), .B(net_13426), .A(net_11374) );
DFF_X1 inst_19798 ( .D(net_18191), .CK(net_22401), .Q(x826) );
INV_X2 inst_19691 ( .A(net_20544), .ZN(net_20543) );
NAND2_X2 inst_9676 ( .ZN(net_10275), .A1(net_10274), .A2(net_7736) );
OAI21_X2 inst_2066 ( .ZN(net_10674), .A(net_10191), .B1(net_7811), .B2(net_6984) );
NAND2_X2 inst_12126 ( .A2(net_1848), .A1(net_703), .ZN(net_546) );
OAI21_X2 inst_1742 ( .ZN(net_20264), .A(net_15026), .B2(net_12748), .B1(net_7717) );
NAND2_X2 inst_12085 ( .ZN(net_1543), .A1(net_327), .A2(net_245) );
INV_X4 inst_13603 ( .ZN(net_8585), .A(net_7171) );
NAND2_X2 inst_12091 ( .ZN(net_660), .A1(net_337), .A2(net_229) );
AOI211_X2 inst_21035 ( .C1(net_14315), .ZN(net_14240), .B(net_13378), .A(net_5148), .C2(net_3203) );
INV_X4 inst_18282 ( .A(net_20075), .ZN(net_20074) );
NAND3_X2 inst_6236 ( .ZN(net_13212), .A3(net_13211), .A2(net_11927), .A1(net_6932) );
INV_X2 inst_18843 ( .A(net_12245), .ZN(net_6689) );
INV_X2 inst_18903 ( .ZN(net_6063), .A(net_6062) );
NOR2_X2 inst_4779 ( .A1(net_3456), .ZN(net_2896), .A2(net_1426) );
NAND2_X2 inst_9522 ( .ZN(net_11128), .A1(net_10654), .A2(net_7585) );
INV_X2 inst_19010 ( .ZN(net_5016), .A(net_5015) );
AOI21_X2 inst_20558 ( .ZN(net_14269), .B2(net_12418), .B1(net_3179), .A(net_1326) );
NOR2_X4 inst_3175 ( .ZN(net_7151), .A1(net_3122), .A2(net_1697) );
OAI21_X2 inst_2302 ( .ZN(net_5880), .B1(net_5547), .B2(net_3195), .A(net_1292) );
NAND2_X2 inst_11021 ( .ZN(net_10465), .A2(net_5443), .A1(net_4794) );
INV_X4 inst_16289 ( .ZN(net_6112), .A(net_86) );
NAND2_X2 inst_9967 ( .ZN(net_19251), .A1(net_11443), .A2(net_8894) );
NAND2_X4 inst_7181 ( .ZN(net_12854), .A2(net_9342), .A1(net_9341) );
OAI211_X2 inst_2447 ( .B(net_14867), .ZN(net_14660), .C2(net_14183), .A(net_13878), .C1(net_5477) );
INV_X2 inst_19700 ( .A(net_20562), .ZN(net_20561) );
NAND2_X2 inst_12043 ( .ZN(net_1542), .A2(net_103), .A1(net_59) );
INV_X4 inst_17377 ( .ZN(net_2389), .A(net_2371) );
INV_X2 inst_18393 ( .A(net_16576), .ZN(net_16536) );
NAND2_X2 inst_11648 ( .ZN(net_2465), .A2(net_2303), .A1(net_28) );
AOI21_X2 inst_20707 ( .B1(net_19860), .ZN(net_12107), .B2(net_6407), .A(net_2615) );
AOI21_X2 inst_20658 ( .ZN(net_13031), .B1(net_13030), .B2(net_12927), .A(net_11999) );
INV_X4 inst_15408 ( .ZN(net_3811), .A(net_2530) );
NAND2_X2 inst_11151 ( .ZN(net_7711), .A1(net_4205), .A2(net_2117) );
NAND2_X2 inst_10914 ( .A2(net_5393), .ZN(net_5350), .A1(net_115) );
NAND2_X2 inst_9695 ( .A1(net_14554), .A2(net_10720), .ZN(net_10226) );
NAND2_X4 inst_7622 ( .ZN(net_1745), .A1(net_1330), .A2(net_834) );
DFF_X1 inst_19814 ( .QN(net_21145), .D(net_17977), .CK(net_21698) );
NAND3_X2 inst_6141 ( .ZN(net_13714), .A2(net_13713), .A3(net_10146), .A1(net_4427) );
CLKBUF_X2 inst_21593 ( .A(net_21464), .Z(net_21465) );
NAND2_X2 inst_7921 ( .ZN(net_18453), .A2(net_18375), .A1(net_17727) );
INV_X4 inst_13303 ( .ZN(net_12271), .A(net_10808) );
NAND2_X4 inst_7163 ( .ZN(net_10949), .A2(net_9478), .A1(net_9397) );
NOR2_X2 inst_4803 ( .ZN(net_4928), .A2(net_2720), .A1(net_701) );
SDFF_X2 inst_935 ( .QN(net_20986), .SE(net_17277), .D(net_2507), .CK(net_22683), .SI(x3220) );
CLKBUF_X2 inst_21664 ( .A(net_21535), .Z(net_21536) );
CLKBUF_X2 inst_21720 ( .A(net_21553), .Z(net_21592) );
INV_X4 inst_17860 ( .ZN(net_92), .A(net_91) );
NAND3_X2 inst_6619 ( .ZN(net_9060), .A2(net_7984), .A3(net_7229), .A1(net_6497) );
NAND3_X2 inst_5699 ( .ZN(net_16227), .A3(net_15918), .A1(net_15598), .A2(net_15254) );
NOR2_X2 inst_4772 ( .ZN(net_2941), .A2(net_2494), .A1(net_1659) );
INV_X4 inst_12781 ( .ZN(net_19654), .A(net_17305) );
NOR2_X2 inst_4634 ( .ZN(net_4545), .A2(net_3514), .A1(net_809) );
AND4_X4 inst_21084 ( .ZN(net_16515), .A3(net_16309), .A4(net_16233), .A1(net_15972), .A2(net_14349) );
INV_X4 inst_16655 ( .ZN(net_7878), .A(net_6081) );
NAND2_X2 inst_11255 ( .ZN(net_19862), .A1(net_6951), .A2(net_3914) );
INV_X4 inst_15997 ( .ZN(net_2759), .A(net_1667) );
NAND2_X2 inst_9284 ( .A1(net_14363), .ZN(net_12545), .A2(net_9662) );
INV_X2 inst_19619 ( .A(net_20877), .ZN(net_39) );
NAND2_X2 inst_11587 ( .ZN(net_4389), .A2(net_2701), .A1(net_154) );
NOR2_X4 inst_2944 ( .A1(net_19575), .ZN(net_11670), .A2(net_10274) );
NOR2_X2 inst_5011 ( .ZN(net_1480), .A1(net_1270), .A2(net_1237) );
AOI21_X2 inst_20665 ( .B1(net_19923), .ZN(net_12922), .B2(net_12004), .A(net_8066) );
INV_X4 inst_15830 ( .ZN(net_11612), .A(net_1864) );
INV_X4 inst_15186 ( .ZN(net_3589), .A(net_2316) );
INV_X4 inst_13690 ( .ZN(net_9480), .A(net_7945) );
INV_X2 inst_19355 ( .ZN(net_9267), .A(net_2362) );
INV_X2 inst_18972 ( .ZN(net_5224), .A(net_5223) );
NAND2_X2 inst_8314 ( .A2(net_20520), .ZN(net_17581), .A1(net_17580) );
NOR2_X4 inst_2862 ( .ZN(net_14444), .A1(net_11552), .A2(net_11439) );
NAND2_X2 inst_7949 ( .ZN(net_18403), .A2(net_18277), .A1(net_18236) );
NAND2_X2 inst_8391 ( .ZN(net_17544), .A2(net_17004), .A1(net_16858) );
DFF_X1 inst_19880 ( .D(net_17134), .CK(net_22088), .Q(x473) );
INV_X4 inst_13397 ( .ZN(net_19990), .A(net_10652) );
INV_X4 inst_15109 ( .A(net_7097), .ZN(net_4296) );
NAND3_X2 inst_6510 ( .ZN(net_10788), .A3(net_10736), .A2(net_6640), .A1(net_5630) );
CLKBUF_X2 inst_22475 ( .A(net_22346), .Z(net_22347) );
NAND3_X2 inst_5808 ( .ZN(net_15656), .A3(net_14871), .A2(net_10121), .A1(net_8584) );
INV_X2 inst_19612 ( .A(net_20855), .ZN(net_49) );
INV_X4 inst_16132 ( .A(net_9450), .ZN(net_7004) );
INV_X8 inst_12181 ( .ZN(net_17441), .A(net_17100) );
INV_X4 inst_13390 ( .ZN(net_13367), .A(net_10726) );
CLKBUF_X2 inst_22000 ( .A(net_21871), .Z(net_21872) );
NAND2_X2 inst_11268 ( .A1(net_20568), .ZN(net_3893), .A2(net_2069) );
NAND2_X4 inst_6859 ( .ZN(net_18387), .A2(net_18318), .A1(net_18269) );
NAND2_X4 inst_7439 ( .A2(net_20559), .ZN(net_4063), .A1(net_3091) );
NOR2_X2 inst_4454 ( .A1(net_8836), .ZN(net_4713), .A2(net_4712) );
INV_X4 inst_17342 ( .ZN(net_4324), .A(net_1922) );
INV_X4 inst_12813 ( .ZN(net_17201), .A(net_17200) );
CLKBUF_X2 inst_22626 ( .A(net_22497), .Z(net_22498) );
NAND2_X2 inst_8709 ( .A1(net_21212), .ZN(net_16275), .A2(net_16105) );
NOR2_X2 inst_4315 ( .ZN(net_9400), .A2(net_5896), .A1(net_70) );
XNOR2_X2 inst_365 ( .A(net_19429), .ZN(net_16852), .B(net_16599) );
XNOR2_X2 inst_67 ( .ZN(net_18805), .A(net_18749), .B(net_17258) );
SDFF_X2 inst_954 ( .QN(net_21087), .D(net_370), .SE(net_263), .CK(net_22601), .SI(x1623) );
AOI21_X2 inst_20552 ( .ZN(net_14305), .A(net_13362), .B2(net_12371), .B1(net_2904) );
INV_X4 inst_16436 ( .ZN(net_6354), .A(net_761) );
INV_X4 inst_13162 ( .ZN(net_14812), .A(net_14231) );
INV_X4 inst_16844 ( .ZN(net_10000), .A(net_7487) );
AND3_X2 inst_21141 ( .ZN(net_9936), .A2(net_9935), .A3(net_3407), .A1(net_2478) );
INV_X4 inst_14186 ( .ZN(net_12137), .A(net_5982) );
NAND2_X2 inst_11216 ( .ZN(net_6885), .A1(net_4207), .A2(net_2086) );
NAND2_X2 inst_8569 ( .ZN(net_16738), .A2(net_16602), .A1(net_16511) );
INV_X4 inst_17729 ( .ZN(net_700), .A(net_185) );
NAND2_X2 inst_11685 ( .ZN(net_2338), .A2(net_2337), .A1(net_90) );
CLKBUF_X2 inst_22425 ( .A(net_22296), .Z(net_22297) );
OAI21_X2 inst_1823 ( .ZN(net_14152), .A(net_14151), .B2(net_10522), .B1(net_7249) );
NOR2_X2 inst_5084 ( .ZN(net_13310), .A1(net_855), .A2(net_60) );
XNOR2_X2 inst_202 ( .ZN(net_17647), .A(net_17295), .B(net_254) );
INV_X4 inst_16249 ( .ZN(net_1405), .A(net_1359) );
NAND2_X4 inst_7359 ( .ZN(net_7459), .A2(net_2641), .A1(net_260) );
CLKBUF_X2 inst_22797 ( .A(net_22668), .Z(net_22669) );
NAND2_X2 inst_9154 ( .ZN(net_13390), .A1(net_12070), .A2(net_10581) );
OAI21_X2 inst_2212 ( .A(net_13922), .ZN(net_8527), .B2(net_8526), .B1(net_5443) );
INV_X4 inst_13786 ( .ZN(net_9206), .A(net_7571) );
OAI21_X4 inst_1401 ( .A(net_20872), .B2(net_19116), .B1(net_19115), .ZN(net_16235) );
NOR2_X2 inst_4830 ( .A1(net_14378), .ZN(net_2455), .A2(net_2454) );
INV_X4 inst_13444 ( .ZN(net_9773), .A(net_9772) );
OAI21_X2 inst_2030 ( .ZN(net_11312), .A(net_11311), .B1(net_9578), .B2(net_3813) );
NAND2_X2 inst_8254 ( .A2(net_17718), .ZN(net_17707), .A1(net_17196) );
NAND2_X2 inst_11172 ( .ZN(net_12883), .A1(net_10962), .A2(net_4138) );
CLKBUF_X2 inst_22919 ( .A(net_21646), .Z(net_22791) );
XOR2_X2 inst_30 ( .A(net_17422), .Z(net_943), .B(net_942) );
XNOR2_X2 inst_610 ( .B(net_17262), .ZN(net_506), .A(net_505) );
NAND3_X2 inst_6271 ( .A3(net_13001), .ZN(net_12947), .A2(net_6691), .A1(net_5800) );
INV_X4 inst_16107 ( .ZN(net_2607), .A(net_1500) );
XNOR2_X2 inst_233 ( .ZN(net_17434), .A(net_17046), .B(net_11624) );
NAND2_X2 inst_9704 ( .A1(net_11721), .ZN(net_10205), .A2(net_10204) );
NAND2_X2 inst_8639 ( .ZN(net_16580), .A2(net_16579), .A1(net_16383) );
AND2_X4 inst_21246 ( .ZN(net_4280), .A1(net_2292), .A2(net_2291) );
NAND2_X2 inst_8595 ( .ZN(net_16690), .A1(net_16689), .A2(net_16688) );
INV_X4 inst_17852 ( .A(net_2744), .ZN(net_218) );
INV_X8 inst_12296 ( .ZN(net_1797), .A(net_1014) );
NAND2_X2 inst_9527 ( .ZN(net_19307), .A1(net_11767), .A2(net_5588) );
NAND2_X2 inst_9127 ( .ZN(net_13531), .A2(net_10793), .A1(net_816) );
INV_X2 inst_18822 ( .ZN(net_6950), .A(net_6949) );
XNOR2_X2 inst_60 ( .ZN(net_18825), .A(net_18773), .B(net_18718) );
NAND2_X2 inst_8939 ( .ZN(net_20165), .A2(net_14095), .A1(net_11676) );
NAND3_X2 inst_6651 ( .ZN(net_8548), .A3(net_7090), .A2(net_6632), .A1(net_5171) );
INV_X4 inst_13540 ( .ZN(net_12960), .A(net_10958) );
NAND2_X2 inst_7752 ( .ZN(net_18774), .A1(net_18760), .A2(net_17563) );
INV_X4 inst_13285 ( .ZN(net_12423), .A(net_12422) );
INV_X4 inst_12862 ( .ZN(net_17143), .A(net_17003) );
NAND2_X4 inst_7339 ( .ZN(net_7816), .A2(net_3359), .A1(net_2230) );
INV_X8 inst_12189 ( .ZN(net_16675), .A(net_16526) );
NAND2_X2 inst_10392 ( .A1(net_10595), .ZN(net_7306), .A2(net_7305) );
NAND2_X2 inst_8389 ( .A1(net_19974), .ZN(net_19268), .A2(net_17290) );
INV_X4 inst_14397 ( .ZN(net_6256), .A(net_5660) );
NOR2_X2 inst_3478 ( .ZN(net_14397), .A1(net_14378), .A2(net_13031) );
INV_X2 inst_18727 ( .ZN(net_14893), .A(net_8099) );
NAND2_X2 inst_11252 ( .A2(net_7144), .ZN(net_3916), .A1(net_3915) );
NAND2_X2 inst_10181 ( .ZN(net_19378), .A1(net_13673), .A2(net_8187) );
INV_X4 inst_17238 ( .ZN(net_1747), .A(net_661) );
NAND2_X4 inst_7147 ( .ZN(net_11593), .A1(net_10454), .A2(net_4994) );
INV_X4 inst_15505 ( .ZN(net_9748), .A(net_2269) );
NOR3_X2 inst_2782 ( .A3(net_14630), .A2(net_14319), .A1(net_9964), .ZN(net_6516) );
NAND2_X4 inst_7248 ( .ZN(net_8780), .A1(net_8068), .A2(net_6842) );
AOI21_X2 inst_20525 ( .ZN(net_14556), .A(net_12110), .B1(net_12067), .B2(net_12009) );
NAND4_X2 inst_5475 ( .A3(net_12958), .ZN(net_12914), .A2(net_10796), .A4(net_9663), .A1(net_3841) );
INV_X4 inst_13887 ( .ZN(net_16659), .A(net_7323) );
NAND2_X2 inst_11191 ( .ZN(net_5391), .A1(net_4090), .A2(net_4009) );
NOR2_X2 inst_3720 ( .A2(net_13490), .ZN(net_12659), .A1(net_8007) );
INV_X4 inst_14672 ( .A(net_6497), .ZN(net_5964) );
NAND2_X2 inst_11964 ( .A2(net_1789), .ZN(net_1377), .A1(net_1376) );
INV_X8 inst_12444 ( .ZN(net_20501), .A(net_16440) );
OAI21_X2 inst_2005 ( .B2(net_12734), .ZN(net_11411), .B1(net_3189), .A(net_843) );
NAND2_X2 inst_11988 ( .ZN(net_2886), .A1(net_2585), .A2(net_1991) );
INV_X4 inst_13377 ( .ZN(net_13605), .A(net_10872) );
SDFF_X2 inst_736 ( .Q(net_20967), .SE(net_18584), .SI(net_18555), .D(net_537), .CK(net_22706) );
XNOR2_X2 inst_544 ( .ZN(net_744), .A(net_743), .B(net_742) );
NAND3_X2 inst_5865 ( .ZN(net_15337), .A3(net_13730), .A1(net_11308), .A2(net_10367) );
NAND2_X2 inst_8021 ( .ZN(net_18276), .A2(net_18224), .A1(net_17561) );
NAND4_X2 inst_5465 ( .ZN(net_13259), .A1(net_12249), .A4(net_8790), .A2(net_5878), .A3(net_4278) );
NAND2_X2 inst_8232 ( .ZN(net_17787), .A2(net_17705), .A1(net_17641) );
AND4_X2 inst_21100 ( .A3(net_12807), .ZN(net_12754), .A2(net_11820), .A4(net_11819), .A1(net_9954) );
CLKBUF_X2 inst_22029 ( .A(net_21370), .Z(net_21901) );
INV_X4 inst_17290 ( .A(net_6867), .ZN(net_4702) );
NOR2_X2 inst_4402 ( .ZN(net_5897), .A2(net_5139), .A1(net_5077) );
SDFF_X2 inst_734 ( .Q(net_20969), .SE(net_18585), .SI(net_18559), .D(net_9001), .CK(net_21678) );
INV_X2 inst_19530 ( .ZN(net_3457), .A(net_1998) );
NAND2_X4 inst_7352 ( .A1(net_20807), .ZN(net_7695), .A2(net_1262) );
CLKBUF_X2 inst_21897 ( .A(net_21619), .Z(net_21769) );
OAI22_X2 inst_1282 ( .B1(net_15955), .ZN(net_15215), .A1(net_15214), .A2(net_14098), .B2(net_9950) );
NAND2_X2 inst_8528 ( .A2(net_20517), .ZN(net_20232), .A1(net_16982) );
INV_X4 inst_16125 ( .ZN(net_2584), .A(net_1526) );
INV_X4 inst_14818 ( .A(net_5400), .ZN(net_4937) );
INV_X4 inst_15673 ( .A(net_2674), .ZN(net_2051) );
INV_X4 inst_17715 ( .ZN(net_15301), .A(net_238) );
NAND2_X4 inst_7661 ( .ZN(net_1038), .A1(net_916), .A2(net_915) );
NAND2_X2 inst_10425 ( .A1(net_7253), .ZN(net_7222), .A2(net_5500) );
NAND2_X2 inst_8898 ( .A1(net_15366), .ZN(net_15103), .A2(net_13882) );
AND3_X2 inst_21150 ( .A3(net_11443), .A2(net_10216), .A1(net_8389), .ZN(net_4238) );
INV_X2 inst_19033 ( .A(net_5029), .ZN(net_4867) );
NAND3_X2 inst_5634 ( .ZN(net_20523), .A3(net_18600), .A1(net_16229), .A2(net_10823) );
CLKBUF_X2 inst_22567 ( .A(net_22438), .Z(net_22439) );
NAND2_X2 inst_9597 ( .ZN(net_10836), .A2(net_7595), .A1(net_2744) );
NOR2_X2 inst_3587 ( .ZN(net_19289), .A1(net_10973), .A2(net_9782) );
NAND2_X2 inst_8777 ( .ZN(net_19406), .A2(net_15359), .A1(net_14061) );
NAND2_X2 inst_10139 ( .A1(net_14458), .ZN(net_8319), .A2(net_8318) );
INV_X4 inst_13003 ( .A(net_16902), .ZN(net_16444) );
NAND2_X2 inst_10147 ( .A1(net_10676), .ZN(net_8296), .A2(net_8295) );
INV_X4 inst_18053 ( .A(net_21149), .ZN(net_17294) );
NAND3_X4 inst_5543 ( .A3(net_19547), .A1(net_19546), .ZN(net_17100), .A2(net_15579) );
AOI21_X2 inst_20799 ( .ZN(net_10400), .A(net_10037), .B2(net_9594), .B1(net_3615) );
NAND3_X2 inst_6392 ( .ZN(net_20458), .A3(net_9523), .A2(net_8949), .A1(net_8492) );
INV_X4 inst_17706 ( .ZN(net_2183), .A(net_508) );
NAND3_X4 inst_5588 ( .ZN(net_15309), .A3(net_13628), .A2(net_10263), .A1(net_8339) );
INV_X4 inst_15465 ( .ZN(net_8877), .A(net_573) );
NAND2_X2 inst_11427 ( .A1(net_6207), .ZN(net_4903), .A2(net_3866) );
INV_X4 inst_16203 ( .ZN(net_1410), .A(net_1409) );
CLKBUF_X2 inst_22286 ( .A(net_22157), .Z(net_22158) );
NAND3_X2 inst_6183 ( .ZN(net_13491), .A3(net_13490), .A1(net_10758), .A2(net_7483) );
CLKBUF_X2 inst_21582 ( .A(net_21453), .Z(net_21454) );
AOI211_X2 inst_21004 ( .ZN(net_18953), .C2(net_15338), .B(net_13924), .A(net_13386), .C1(net_2548) );
INV_X4 inst_17800 ( .A(net_703), .ZN(net_262) );
NAND2_X2 inst_11529 ( .ZN(net_2954), .A1(net_2953), .A2(net_2952) );
NAND2_X2 inst_8542 ( .A2(net_17752), .ZN(net_16819), .A1(net_1814) );
INV_X4 inst_17745 ( .ZN(net_5448), .A(net_226) );
INV_X4 inst_16445 ( .ZN(net_11776), .A(net_11511) );
INV_X2 inst_19640 ( .A(net_19432), .ZN(net_19431) );
NOR2_X2 inst_3701 ( .ZN(net_11105), .A2(net_11104), .A1(net_3523) );
NOR2_X2 inst_3357 ( .ZN(net_17650), .A1(net_17482), .A2(net_17367) );
NAND2_X4 inst_7082 ( .A1(net_19532), .ZN(net_15711), .A2(net_14276) );
NAND2_X2 inst_11822 ( .ZN(net_1800), .A2(net_1064), .A1(net_962) );
XOR2_X2 inst_8 ( .A(net_21125), .B(net_17166), .Z(net_17150) );
AND2_X4 inst_21260 ( .ZN(net_2842), .A1(net_809), .A2(net_85) );
INV_X4 inst_15559 ( .ZN(net_2741), .A(net_1448) );
INV_X4 inst_15456 ( .ZN(net_13504), .A(net_10395) );
AOI211_X2 inst_21019 ( .ZN(net_15043), .C1(net_14365), .C2(net_13499), .A(net_10968), .B(net_5929) );
NAND2_X2 inst_8925 ( .A1(net_15582), .ZN(net_14942), .A2(net_13604) );
NAND2_X4 inst_6984 ( .ZN(net_17651), .A1(net_16907), .A2(net_16719) );
INV_X4 inst_17420 ( .ZN(net_502), .A(net_493) );
OAI21_X2 inst_2090 ( .ZN(net_10299), .A(net_10298), .B2(net_5978), .B1(net_4582) );
SDFF_X2 inst_965 ( .QN(net_21100), .D(net_632), .SE(net_263), .CK(net_21778), .SI(x1401) );
NAND2_X2 inst_8228 ( .ZN(net_17794), .A2(net_17606), .A1(net_17545) );
INV_X4 inst_14583 ( .ZN(net_7899), .A(net_4021) );
INV_X8 inst_12267 ( .ZN(net_14038), .A(net_8199) );
NAND2_X2 inst_8677 ( .A1(net_20766), .A2(net_16465), .ZN(net_16457) );
NAND2_X2 inst_11991 ( .ZN(net_5248), .A2(net_4357), .A1(net_222) );
AOI211_X2 inst_21065 ( .ZN(net_9012), .C2(net_6211), .C1(net_3754), .A(net_3527), .B(net_3043) );
INV_X8 inst_12284 ( .ZN(net_4293), .A(net_3852) );
NAND2_X2 inst_11976 ( .ZN(net_3908), .A1(net_388), .A2(net_50) );
NAND4_X2 inst_5392 ( .ZN(net_20706), .A3(net_13323), .A4(net_13322), .A1(net_12598), .A2(net_11202) );
NAND3_X2 inst_6179 ( .ZN(net_13501), .A1(net_11052), .A3(net_8985), .A2(net_6229) );
INV_X4 inst_15520 ( .ZN(net_3051), .A(net_1616) );
AOI21_X2 inst_20500 ( .ZN(net_14654), .B1(net_14653), .A(net_12695), .B2(net_12097) );
INV_X4 inst_18073 ( .A(net_20866), .ZN(net_156) );
CLKBUF_X2 inst_22307 ( .A(net_22178), .Z(net_22179) );
CLKBUF_X2 inst_21598 ( .A(net_21469), .Z(net_21470) );
AOI21_X4 inst_20146 ( .ZN(net_20652), .B1(net_19125), .A(net_10751), .B2(net_588) );
CLKBUF_X2 inst_21787 ( .A(net_21658), .Z(net_21659) );
INV_X4 inst_16003 ( .ZN(net_11681), .A(net_1663) );
NAND2_X2 inst_7913 ( .ZN(net_18460), .A2(net_18346), .A1(net_18294) );
CLKBUF_X2 inst_22890 ( .A(net_22761), .Z(net_22762) );
INV_X4 inst_16097 ( .ZN(net_2491), .A(net_2193) );
INV_X4 inst_13288 ( .ZN(net_12412), .A(net_12411) );
INV_X4 inst_14013 ( .ZN(net_13213), .A(net_6305) );
AOI211_X4 inst_20993 ( .C1(net_19624), .ZN(net_14180), .C2(net_14179), .A(net_6800), .B(net_6746) );
OAI21_X2 inst_1934 ( .ZN(net_12931), .B1(net_10723), .B2(net_9431), .A(net_8293) );
NAND3_X2 inst_6759 ( .A1(net_8241), .ZN(net_5631), .A3(net_5209), .A2(net_3297) );
INV_X4 inst_16022 ( .A(net_10504), .ZN(net_1641) );
NAND2_X2 inst_9429 ( .ZN(net_11613), .A1(net_11612), .A2(net_11039) );
INV_X4 inst_18207 ( .A(net_21148), .ZN(net_16646) );
NOR2_X2 inst_3916 ( .ZN(net_8817), .A2(net_8166), .A1(net_8062) );
NAND3_X2 inst_5739 ( .ZN(net_16048), .A3(net_15469), .A1(net_14025), .A2(net_12685) );
NAND4_X2 inst_5401 ( .ZN(net_14776), .A2(net_13345), .A1(net_12700), .A4(net_10626), .A3(net_8282) );
INV_X2 inst_18752 ( .ZN(net_7794), .A(net_7793) );
NAND2_X2 inst_9970 ( .ZN(net_18949), .A1(net_11018), .A2(net_8891) );
INV_X4 inst_17007 ( .ZN(net_865), .A(net_849) );
NAND2_X2 inst_8319 ( .ZN(net_19557), .A2(net_19396), .A1(net_19395) );
NAND2_X2 inst_8539 ( .A1(net_21208), .A2(net_16994), .ZN(net_16828) );
INV_X2 inst_19136 ( .ZN(net_4144), .A(net_4143) );
INV_X4 inst_13359 ( .ZN(net_12355), .A(net_10949) );
CLKBUF_X2 inst_22676 ( .A(net_22547), .Z(net_22548) );
NAND2_X2 inst_8464 ( .A1(net_20788), .A2(net_20069), .ZN(net_19656) );
NAND2_X2 inst_10968 ( .ZN(net_6175), .A2(net_5109), .A1(net_1103) );
OAI21_X2 inst_2097 ( .A(net_10164), .ZN(net_10073), .B2(net_10072), .B1(net_3980) );
INV_X4 inst_12943 ( .A(net_16789), .ZN(net_16634) );
NOR2_X2 inst_4484 ( .A1(net_6876), .ZN(net_5562), .A2(net_4295) );
CLKBUF_X2 inst_21401 ( .A(net_21272), .Z(net_21273) );
INV_X4 inst_14948 ( .ZN(net_5893), .A(net_3515) );
NAND2_X2 inst_8053 ( .ZN(net_18215), .A1(net_18214), .A2(net_18213) );
NAND3_X2 inst_6215 ( .ZN(net_13263), .A2(net_11746), .A3(net_10530), .A1(net_10513) );
INV_X2 inst_18798 ( .ZN(net_11138), .A(net_7424) );
INV_X4 inst_16350 ( .A(net_8521), .ZN(net_1777) );
INV_X4 inst_16700 ( .ZN(net_7196), .A(net_1066) );
CLKBUF_X2 inst_21792 ( .A(net_21663), .Z(net_21664) );
INV_X8 inst_12225 ( .A(net_5934), .ZN(net_5834) );
SDFF_X2 inst_1050 ( .QN(net_21027), .D(net_648), .SE(net_263), .CK(net_21945), .SI(x2547) );
NAND3_X2 inst_6476 ( .ZN(net_11284), .A2(net_11273), .A3(net_3081), .A1(net_1700) );
DFF_X1 inst_19864 ( .D(net_17065), .CK(net_22102), .Q(x503) );
INV_X4 inst_17546 ( .A(net_14104), .ZN(net_11968) );
INV_X4 inst_17195 ( .ZN(net_20424), .A(net_987) );
NOR2_X2 inst_4661 ( .ZN(net_8090), .A2(net_3287), .A1(net_1423) );
OAI21_X2 inst_1852 ( .A(net_15020), .ZN(net_14003), .B2(net_10341), .B1(net_8561) );
NAND3_X2 inst_6809 ( .A2(net_2996), .ZN(net_2498), .A3(net_2497), .A1(net_112) );
NAND3_X2 inst_6273 ( .ZN(net_12943), .A2(net_11974), .A3(net_9406), .A1(net_5359) );
CLKBUF_X2 inst_22826 ( .A(net_21818), .Z(net_22698) );
CLKBUF_X2 inst_21869 ( .A(net_21379), .Z(net_21741) );
NOR2_X4 inst_3282 ( .ZN(net_2460), .A1(net_1614), .A2(net_1556) );
INV_X4 inst_12667 ( .ZN(net_20634), .A(net_17799) );
NOR2_X2 inst_4074 ( .ZN(net_7531), .A2(net_7530), .A1(net_1076) );
NOR2_X2 inst_3783 ( .ZN(net_20731), .A1(net_10124), .A2(net_9446) );
INV_X4 inst_13613 ( .ZN(net_12762), .A(net_8419) );
OAI21_X2 inst_1557 ( .ZN(net_17565), .B2(net_17498), .A(net_17248), .B1(net_17247) );
OAI211_X2 inst_2399 ( .ZN(net_16010), .A(net_16009), .B(net_15650), .C2(net_15155), .C1(net_15020) );
INV_X2 inst_18498 ( .ZN(net_13364), .A(net_12305) );
INV_X2 inst_18430 ( .ZN(net_14861), .A(net_14322) );
INV_X8 inst_12207 ( .ZN(net_13324), .A(net_7568) );
NOR2_X2 inst_3412 ( .A2(net_20362), .A1(net_20361), .ZN(net_19402) );
NOR2_X2 inst_4698 ( .ZN(net_4146), .A2(net_3174), .A1(net_3146) );
NAND2_X2 inst_9620 ( .ZN(net_10689), .A1(net_10688), .A2(net_8496) );
NAND2_X2 inst_8485 ( .ZN(net_20189), .A1(net_16985), .A2(net_16973) );
INV_X4 inst_17431 ( .ZN(net_959), .A(net_482) );
CLKBUF_X2 inst_21660 ( .A(net_21531), .Z(net_21532) );
INV_X4 inst_17247 ( .ZN(net_4890), .A(net_993) );
NAND2_X2 inst_11326 ( .ZN(net_5319), .A1(net_4299), .A2(net_3339) );
CLKBUF_X2 inst_22449 ( .A(net_22320), .Z(net_22321) );
OAI21_X2 inst_1616 ( .A(net_20952), .ZN(net_16087), .B2(net_15555), .B1(net_12186) );
INV_X4 inst_14090 ( .ZN(net_11198), .A(net_7753) );
NAND2_X2 inst_8813 ( .ZN(net_15606), .A2(net_14946), .A1(net_13024) );
NAND3_X2 inst_5646 ( .A3(net_19062), .A1(net_19061), .ZN(net_16897), .A2(net_16249) );
INV_X4 inst_13167 ( .ZN(net_14799), .A(net_14206) );
NAND2_X2 inst_11295 ( .ZN(net_6225), .A1(net_3509), .A2(net_759) );
NAND2_X2 inst_11403 ( .ZN(net_3455), .A2(net_2439), .A1(net_1232) );
DFF_X1 inst_19861 ( .D(net_17133), .CK(net_22544), .Q(x140) );
NAND4_X2 inst_5356 ( .ZN(net_15410), .A1(net_14667), .A3(net_14303), .A4(net_10884), .A2(net_8680) );
INV_X4 inst_13110 ( .ZN(net_15651), .A(net_15419) );
INV_X2 inst_19551 ( .ZN(net_1184), .A(net_899) );
NAND2_X2 inst_8690 ( .ZN(net_18997), .A1(net_16385), .A2(net_16271) );
NAND2_X2 inst_11786 ( .ZN(net_2631), .A1(net_1376), .A2(net_1136) );
NAND2_X2 inst_11621 ( .A2(net_2685), .ZN(net_2556), .A1(net_1751) );
INV_X4 inst_17410 ( .ZN(net_15450), .A(net_14563) );
INV_X4 inst_15303 ( .A(net_3946), .ZN(net_2665) );
INV_X4 inst_16536 ( .ZN(net_15607), .A(net_14793) );
NOR2_X4 inst_3186 ( .ZN(net_9525), .A1(net_3111), .A2(net_1099) );
INV_X4 inst_15266 ( .ZN(net_6445), .A(net_3838) );
NOR2_X2 inst_3762 ( .A2(net_14900), .ZN(net_12965), .A1(net_10309) );
NAND3_X2 inst_5653 ( .ZN(net_16550), .A3(net_16403), .A2(net_16174), .A1(net_15427) );
CLKBUF_X2 inst_22445 ( .A(net_22262), .Z(net_22317) );
NAND2_X2 inst_10925 ( .ZN(net_9935), .A2(net_6541), .A1(net_3745) );
NOR2_X4 inst_3259 ( .ZN(net_5689), .A1(net_1788), .A2(net_1404) );
SDFF_X2 inst_854 ( .Q(net_21186), .SI(net_17210), .SE(net_125), .CK(net_22234), .D(x6461) );
INV_X4 inst_12464 ( .ZN(net_18803), .A(net_18802) );
INV_X4 inst_13293 ( .A(net_12614), .ZN(net_12377) );
AOI222_X2 inst_20066 ( .ZN(net_9015), .A1(net_9014), .A2(net_6665), .C2(net_3353), .B2(net_2097), .B1(net_494), .C1(net_81) );
INV_X4 inst_13796 ( .ZN(net_13330), .A(net_7559) );
INV_X4 inst_15369 ( .ZN(net_4045), .A(net_2572) );
INV_X4 inst_16600 ( .ZN(net_2229), .A(net_1602) );
NOR2_X2 inst_3678 ( .ZN(net_20610), .A1(net_11432), .A2(net_9246) );
NOR2_X2 inst_3979 ( .ZN(net_8390), .A1(net_8389), .A2(net_4788) );
NAND3_X2 inst_6297 ( .ZN(net_12817), .A3(net_12816), .A2(net_9346), .A1(net_8119) );
INV_X4 inst_15578 ( .ZN(net_7219), .A(net_7004) );
NAND2_X2 inst_7865 ( .ZN(net_18556), .A2(net_18502), .A1(net_18395) );
NAND2_X2 inst_10478 ( .A2(net_10629), .ZN(net_6977), .A1(net_6976) );
NAND2_X2 inst_12006 ( .ZN(net_7002), .A2(net_1697), .A1(net_1158) );
NAND2_X2 inst_8008 ( .ZN(net_18355), .A2(net_18217), .A1(net_18189) );
INV_X4 inst_13401 ( .ZN(net_13962), .A(net_8943) );
AOI21_X2 inst_20983 ( .B1(net_4340), .ZN(net_2538), .B2(net_2283), .A(net_1824) );
NAND2_X2 inst_10861 ( .ZN(net_13697), .A1(net_5438), .A2(net_5384) );
NAND2_X2 inst_9464 ( .ZN(net_11486), .A2(net_9277), .A1(net_828) );
OAI21_X2 inst_1749 ( .ZN(net_14839), .A(net_14838), .B1(net_14837), .B2(net_13883) );
INV_X4 inst_16508 ( .ZN(net_1647), .A(net_1190) );
NAND2_X2 inst_9717 ( .ZN(net_10165), .A1(net_10164), .A2(net_7707) );
NAND3_X2 inst_6519 ( .ZN(net_10645), .A2(net_10644), .A3(net_10643), .A1(net_7547) );
INV_X4 inst_14105 ( .ZN(net_11243), .A(net_6169) );
NAND4_X2 inst_5514 ( .ZN(net_10541), .A2(net_10540), .A3(net_10539), .A4(net_9719), .A1(net_4541) );
INV_X4 inst_12518 ( .ZN(net_20703), .A(net_18562) );
NAND2_X2 inst_9071 ( .ZN(net_13975), .A2(net_12198), .A1(net_10069) );
NAND2_X2 inst_11872 ( .ZN(net_2467), .A2(net_1636), .A1(net_1385) );
NAND2_X2 inst_9017 ( .ZN(net_14202), .A2(net_14201), .A1(net_588) );
AOI21_X2 inst_20493 ( .ZN(net_14753), .B1(net_12669), .B2(net_12285), .A(net_11098) );
SDFF_X2 inst_840 ( .Q(net_21117), .SI(net_17296), .SE(net_125), .CK(net_21553), .D(x4481) );
INV_X4 inst_16555 ( .ZN(net_1170), .A(net_1169) );
INV_X4 inst_17073 ( .ZN(net_4037), .A(net_3187) );
NAND2_X2 inst_11900 ( .A2(net_6563), .ZN(net_1576), .A1(net_1394) );
INV_X4 inst_13523 ( .ZN(net_13621), .A(net_9343) );
INV_X4 inst_12498 ( .ZN(net_18680), .A(net_18663) );
NAND3_X2 inst_6117 ( .ZN(net_13865), .A3(net_13864), .A2(net_12266), .A1(net_4271) );
NAND2_X2 inst_10736 ( .A1(net_7028), .ZN(net_5769), .A2(net_5768) );
CLKBUF_X2 inst_22771 ( .A(net_22642), .Z(net_22643) );
NAND3_X2 inst_5876 ( .ZN(net_20591), .A1(net_14505), .A3(net_10425), .A2(net_4686) );
NAND2_X4 inst_7497 ( .ZN(net_4290), .A2(net_2331), .A1(net_225) );
NOR2_X2 inst_4294 ( .ZN(net_11209), .A2(net_3354), .A1(net_1809) );
INV_X2 inst_18512 ( .A(net_14536), .ZN(net_11579) );
NAND2_X4 inst_7589 ( .ZN(net_2026), .A2(net_807), .A1(net_129) );
INV_X16 inst_19741 ( .ZN(net_973), .A(net_179) );
INV_X4 inst_14302 ( .A(net_15582), .ZN(net_8411) );
CLKBUF_X2 inst_22046 ( .A(net_21917), .Z(net_21918) );
NAND2_X2 inst_10799 ( .ZN(net_5974), .A1(net_4862), .A2(net_3478) );
NAND3_X2 inst_5710 ( .A3(net_19988), .A1(net_19987), .ZN(net_19623), .A2(net_9773) );
INV_X2 inst_19347 ( .ZN(net_2417), .A(net_2416) );
AOI21_X2 inst_20880 ( .ZN(net_8280), .B1(net_6488), .B2(net_3651), .A(net_3251) );
NAND2_X2 inst_9536 ( .ZN(net_12694), .A2(net_11067), .A1(net_9459) );
NAND3_X2 inst_5939 ( .A3(net_20197), .A1(net_20196), .ZN(net_19090), .A2(net_11537) );
AOI21_X2 inst_20535 ( .ZN(net_14502), .A(net_12930), .B1(net_12880), .B2(net_11519) );
INV_X4 inst_15966 ( .ZN(net_10930), .A(net_1688) );
NAND2_X2 inst_11846 ( .A1(net_20495), .ZN(net_3150), .A2(net_247) );
NAND3_X2 inst_5679 ( .A3(net_19799), .A1(net_19798), .ZN(net_16332), .A2(net_12758) );
NAND2_X4 inst_7272 ( .ZN(net_9633), .A1(net_5945), .A2(net_2585) );
NAND2_X2 inst_11141 ( .A1(net_7659), .ZN(net_4237), .A2(net_4236) );
AND2_X2 inst_21312 ( .A2(net_11338), .ZN(net_8385), .A1(net_8384) );
NAND2_X2 inst_9200 ( .A1(net_15183), .ZN(net_13085), .A2(net_11360) );
INV_X4 inst_16527 ( .ZN(net_10445), .A(net_9378) );
XNOR2_X2 inst_617 ( .B(net_5788), .ZN(net_486), .A(net_485) );
INV_X4 inst_14897 ( .A(net_5109), .ZN(net_4634) );
NAND2_X2 inst_9167 ( .A2(net_19991), .A1(net_19990), .ZN(net_13368) );
NAND3_X2 inst_5734 ( .ZN(net_16062), .A3(net_15505), .A1(net_15045), .A2(net_14169) );
NAND2_X2 inst_10823 ( .ZN(net_6803), .A1(net_5499), .A2(net_5468) );
INV_X4 inst_18089 ( .A(net_21077), .ZN(net_589) );
INV_X4 inst_16634 ( .ZN(net_3045), .A(net_1109) );
NAND2_X2 inst_8123 ( .A2(net_18067), .ZN(net_18057), .A1(net_15510) );
NAND3_X2 inst_6614 ( .ZN(net_9074), .A1(net_9073), .A2(net_9072), .A3(net_7014) );
INV_X2 inst_18457 ( .ZN(net_13370), .A(net_13369) );
INV_X4 inst_15749 ( .ZN(net_3866), .A(net_1944) );
NAND3_X2 inst_6029 ( .ZN(net_14370), .A3(net_13766), .A1(net_8591), .A2(net_6104) );
CLKBUF_X2 inst_22300 ( .A(net_22171), .Z(net_22172) );
INV_X2 inst_19089 ( .ZN(net_4561), .A(net_4560) );
NAND2_X2 inst_11956 ( .ZN(net_1396), .A1(net_1395), .A2(net_216) );
NAND4_X2 inst_5482 ( .ZN(net_12489), .A3(net_12488), .A4(net_12487), .A2(net_12063), .A1(net_4382) );
NAND2_X4 inst_7159 ( .ZN(net_11607), .A1(net_9618), .A2(net_9537) );
CLKBUF_X2 inst_21682 ( .A(net_21536), .Z(net_21554) );
NAND3_X2 inst_6739 ( .ZN(net_6462), .A1(net_6461), .A3(net_4273), .A2(net_3585) );
INV_X4 inst_17494 ( .ZN(net_14160), .A(net_816) );
INV_X4 inst_18045 ( .A(net_21123), .ZN(net_543) );
NAND2_X2 inst_8916 ( .ZN(net_14963), .A1(net_14962), .A2(net_13647) );
INV_X4 inst_14487 ( .ZN(net_9954), .A(net_6561) );
NAND2_X2 inst_9818 ( .A2(net_12738), .ZN(net_9651), .A1(net_9650) );
NAND2_X2 inst_8798 ( .ZN(net_15672), .A2(net_15157), .A1(net_13075) );
INV_X4 inst_15064 ( .ZN(net_5480), .A(net_2501) );
NOR2_X4 inst_2909 ( .ZN(net_19183), .A2(net_8429), .A1(net_8421) );
INV_X4 inst_12636 ( .ZN(net_17916), .A(net_17915) );
AOI21_X4 inst_20161 ( .B1(net_20190), .ZN(net_15696), .A(net_13835), .B2(net_9191) );
NOR2_X4 inst_3135 ( .ZN(net_6998), .A1(net_4022), .A2(net_3800) );
SDFF_X2 inst_701 ( .Q(net_20924), .SE(net_18864), .SI(net_18838), .D(net_737), .CK(net_22038) );
OAI211_X4 inst_2380 ( .C1(net_19367), .ZN(net_15713), .B(net_9744), .C2(net_9080), .A(net_8528) );
INV_X4 inst_16780 ( .ZN(net_12496), .A(net_1019) );
INV_X8 inst_12337 ( .ZN(net_3056), .A(net_3026) );
NAND2_X4 inst_7583 ( .A1(net_20581), .ZN(net_1571), .A2(net_1442) );
NAND4_X2 inst_5261 ( .A4(net_20173), .A1(net_20172), .ZN(net_16225), .A2(net_15267), .A3(net_12949) );
CLKBUF_X2 inst_22587 ( .A(net_22458), .Z(net_22459) );
CLKBUF_X2 inst_21862 ( .A(net_21733), .Z(net_21734) );
INV_X4 inst_15998 ( .ZN(net_20741), .A(net_1666) );
INV_X4 inst_17356 ( .ZN(net_15616), .A(net_178) );
NAND2_X2 inst_7739 ( .ZN(net_18801), .A2(net_18771), .A1(net_17856) );
AOI211_X2 inst_21040 ( .ZN(net_13493), .B(net_12771), .C2(net_10767), .A(net_3440), .C1(net_81) );
CLKBUF_X2 inst_22260 ( .A(net_21618), .Z(net_22132) );
NAND2_X4 inst_6933 ( .A2(net_18933), .A1(net_18932), .ZN(net_17629) );
SDFF_X2 inst_1007 ( .QN(net_21096), .D(net_389), .SE(net_263), .CK(net_22581), .SI(x1457) );
NAND2_X2 inst_11011 ( .ZN(net_4873), .A1(net_4872), .A2(net_2690) );
INV_X2 inst_19348 ( .A(net_2940), .ZN(net_2415) );
INV_X4 inst_15989 ( .ZN(net_13274), .A(net_10134) );
CLKBUF_X2 inst_22948 ( .A(net_22819), .Z(net_22820) );
NAND2_X2 inst_11674 ( .ZN(net_6392), .A2(net_2093), .A1(net_165) );
CLKBUF_X2 inst_22734 ( .A(net_21817), .Z(net_22606) );
NAND2_X2 inst_11932 ( .ZN(net_3241), .A1(net_1529), .A2(net_1486) );
NOR2_X2 inst_5066 ( .ZN(net_11997), .A1(net_788), .A2(net_70) );
NAND2_X2 inst_11998 ( .ZN(net_4378), .A1(net_1186), .A2(net_90) );
INV_X4 inst_16160 ( .ZN(net_2847), .A(net_2060) );
NOR2_X4 inst_2883 ( .A1(net_18920), .ZN(net_11675), .A2(net_9745) );
NAND2_X2 inst_11313 ( .ZN(net_11843), .A1(net_8877), .A2(net_3776) );
CLKBUF_X2 inst_22562 ( .A(net_22433), .Z(net_22434) );
CLKBUF_X2 inst_21536 ( .A(net_21406), .Z(net_21408) );
NAND2_X2 inst_11108 ( .ZN(net_4935), .A2(net_2837), .A1(net_2712) );
INV_X2 inst_18733 ( .A(net_8651), .ZN(net_7999) );
NAND2_X2 inst_10083 ( .A2(net_8681), .ZN(net_8634), .A1(net_7394) );
INV_X2 inst_19726 ( .A(net_20796), .ZN(net_20795) );
NOR2_X2 inst_3685 ( .A1(net_14791), .ZN(net_11416), .A2(net_9300) );
NAND2_X2 inst_10527 ( .A2(net_13203), .ZN(net_6836), .A1(net_6835) );
INV_X4 inst_16407 ( .ZN(net_15088), .A(net_14684) );
NAND2_X4 inst_6891 ( .ZN(net_19493), .A2(net_18070), .A1(net_16375) );
AOI22_X2 inst_20019 ( .ZN(net_11229), .B1(net_10962), .A1(net_10096), .A2(net_7497), .B2(net_4499) );
NAND2_X2 inst_11301 ( .A2(net_20801), .ZN(net_5047), .A1(net_3792) );
INV_X2 inst_19140 ( .ZN(net_4129), .A(net_4128) );
OAI21_X4 inst_1472 ( .B2(net_19134), .B1(net_19133), .ZN(net_14792), .A(net_1070) );
INV_X2 inst_19161 ( .ZN(net_5015), .A(net_3934) );
INV_X4 inst_17633 ( .ZN(net_285), .A(net_284) );
NOR2_X2 inst_4261 ( .ZN(net_7594), .A1(net_6089), .A2(net_4623) );
NAND2_X4 inst_7616 ( .ZN(net_2328), .A2(net_1344), .A1(net_1142) );
INV_X4 inst_12511 ( .A(net_18626), .ZN(net_18605) );
INV_X4 inst_14784 ( .ZN(net_9695), .A(net_5547) );
NOR2_X2 inst_3784 ( .ZN(net_14908), .A2(net_10156), .A1(net_9083) );
OR2_X2 inst_1183 ( .A2(net_4837), .ZN(net_4748), .A1(net_4747) );
NAND2_X2 inst_9577 ( .ZN(net_10938), .A1(net_10937), .A2(net_9096) );
OAI21_X4 inst_1489 ( .B2(net_19122), .B1(net_19121), .ZN(net_13394), .A(net_10225) );
OAI211_X2 inst_2415 ( .ZN(net_20389), .C1(net_15506), .B(net_14629), .C2(net_13907), .A(net_11923) );
INV_X8 inst_12353 ( .ZN(net_2431), .A(net_260) );
INV_X4 inst_14498 ( .ZN(net_6006), .A(net_4841) );
NOR2_X2 inst_4981 ( .ZN(net_2998), .A1(net_1485), .A2(net_1354) );
NAND2_X2 inst_8352 ( .A2(net_17493), .ZN(net_17467), .A1(net_17466) );
NAND4_X2 inst_5506 ( .ZN(net_11280), .A2(net_11279), .A4(net_11278), .A1(net_6116), .A3(net_6005) );
NAND2_X4 inst_7102 ( .ZN(net_12367), .A2(net_12366), .A1(net_10742) );
OAI21_X2 inst_1808 ( .A(net_14634), .ZN(net_14467), .B2(net_11631), .B1(net_6084) );
INV_X4 inst_17896 ( .ZN(net_307), .A(net_62) );
NAND2_X2 inst_8440 ( .ZN(net_17266), .A2(net_16819), .A1(net_16661) );
SDFF_X2 inst_988 ( .QN(net_20978), .D(net_2277), .SE(net_263), .CK(net_22669), .SI(x3339) );
INV_X4 inst_16988 ( .ZN(net_2348), .A(net_878) );
NAND2_X2 inst_10288 ( .ZN(net_9469), .A2(net_4922), .A1(net_4288) );
INV_X4 inst_15668 ( .ZN(net_12881), .A(net_9330) );
INV_X4 inst_14941 ( .ZN(net_4879), .A(net_3531) );
NAND2_X2 inst_9333 ( .ZN(net_12299), .A1(net_12298), .A2(net_9054) );
NOR2_X2 inst_4954 ( .ZN(net_2261), .A1(net_1848), .A2(net_1250) );
NOR2_X2 inst_4308 ( .ZN(net_7420), .A2(net_5914), .A1(net_399) );
NAND2_X2 inst_11026 ( .ZN(net_5946), .A1(net_4783), .A2(net_3365) );
INV_X2 inst_18460 ( .ZN(net_19180), .A(net_12042) );
NAND2_X4 inst_7569 ( .A1(net_20495), .ZN(net_2399), .A2(net_1640) );
INV_X4 inst_18100 ( .A(net_21030), .ZN(net_586) );
CLKBUF_X2 inst_22667 ( .A(net_21708), .Z(net_22539) );
INV_X2 inst_18654 ( .ZN(net_9217), .A(net_9216) );
NAND2_X2 inst_10049 ( .A2(net_10534), .ZN(net_8695), .A1(net_7441) );
INV_X4 inst_15249 ( .A(net_3797), .ZN(net_3560) );
AOI21_X2 inst_20364 ( .B1(net_15731), .ZN(net_15639), .B2(net_14433), .A(net_10494) );
AOI21_X4 inst_20207 ( .B1(net_20663), .ZN(net_14638), .B2(net_13350), .A(net_7694) );
INV_X1 inst_19750 ( .ZN(net_14254), .A(net_12374) );
NAND2_X2 inst_9808 ( .ZN(net_12131), .A2(net_7814), .A1(net_5776) );
AND2_X2 inst_21333 ( .ZN(net_4617), .A1(net_4616), .A2(net_4615) );
NAND3_X4 inst_5527 ( .A1(net_20787), .A3(net_19817), .ZN(net_17876), .A2(net_15927) );
NAND2_X4 inst_7007 ( .A1(net_17239), .ZN(net_17053), .A2(net_17052) );
NAND3_X2 inst_6718 ( .ZN(net_7929), .A3(net_6648), .A1(net_4109), .A2(net_2585) );
INV_X4 inst_12562 ( .ZN(net_18240), .A(net_18239) );
NAND3_X2 inst_5919 ( .ZN(net_15005), .A3(net_13077), .A2(net_11314), .A1(net_8850) );
AOI21_X2 inst_20788 ( .ZN(net_20847), .A(net_10688), .B1(net_10546), .B2(net_8727) );
INV_X4 inst_13471 ( .ZN(net_11027), .A(net_9646) );
CLKBUF_X2 inst_21708 ( .A(net_21523), .Z(net_21580) );
DFF_X1 inst_19885 ( .D(net_17117), .CK(net_21596), .Q(x629) );
INV_X4 inst_17910 ( .A(net_824), .ZN(net_182) );
INV_X2 inst_18939 ( .ZN(net_5821), .A(net_5820) );
NOR2_X2 inst_4618 ( .A1(net_6812), .ZN(net_6556), .A2(net_4328) );
NAND2_X4 inst_6827 ( .ZN(net_18850), .A2(net_18833), .A1(net_18819) );
OAI21_X2 inst_1922 ( .ZN(net_13024), .A(net_13023), .B2(net_11501), .B1(net_5221) );
NOR2_X2 inst_3361 ( .ZN(net_17367), .A1(net_17366), .A2(net_17365) );
NOR2_X4 inst_3170 ( .A2(net_20568), .ZN(net_3671), .A1(net_3177) );
NOR2_X4 inst_3232 ( .ZN(net_3127), .A1(net_2456), .A2(net_1795) );
NAND2_X2 inst_8335 ( .A2(net_20508), .ZN(net_17516), .A1(net_17515) );
INV_X4 inst_13062 ( .ZN(net_16351), .A(net_16295) );
NAND2_X2 inst_10524 ( .ZN(net_6847), .A2(net_3978), .A1(net_3310) );
NAND2_X2 inst_10444 ( .ZN(net_7184), .A1(net_7183), .A2(net_7182) );
NAND3_X2 inst_5973 ( .ZN(net_14762), .A3(net_13366), .A1(net_12385), .A2(net_10469) );
NAND2_X4 inst_6942 ( .A1(net_20584), .ZN(net_19047), .A2(net_17483) );
AOI21_X2 inst_20627 ( .B1(net_19005), .ZN(net_13433), .B2(net_10206), .A(net_4185) );
INV_X4 inst_16731 ( .ZN(net_15636), .A(net_15468) );
OAI21_X4 inst_1350 ( .ZN(net_18665), .B2(net_18640), .A(net_18623), .B1(net_17123) );
AND2_X2 inst_21307 ( .A2(net_9759), .ZN(net_9304), .A1(net_2182) );
NAND2_X1 inst_12156 ( .A1(net_11505), .ZN(net_6768), .A2(net_5521) );
INV_X4 inst_16489 ( .ZN(net_12231), .A(net_11297) );
NOR2_X4 inst_3012 ( .ZN(net_6270), .A2(net_3890), .A1(net_3563) );
NAND2_X2 inst_11369 ( .ZN(net_3579), .A1(net_3297), .A2(net_2387) );
NOR3_X2 inst_2635 ( .ZN(net_16198), .A1(net_16002), .A2(net_11192), .A3(net_10218) );
INV_X4 inst_16502 ( .ZN(net_10490), .A(net_1790) );
INV_X4 inst_14014 ( .A(net_6305), .ZN(net_6304) );
NAND2_X2 inst_8673 ( .A2(net_16721), .ZN(net_16461), .A1(net_5731) );
CLKBUF_X2 inst_22897 ( .A(net_22768), .Z(net_22769) );
NOR2_X2 inst_3363 ( .A2(net_17239), .ZN(net_17238), .A1(net_17237) );
NOR3_X2 inst_2666 ( .ZN(net_14984), .A1(net_14036), .A2(net_13184), .A3(net_12937) );
AOI21_X2 inst_20274 ( .B1(net_19066), .ZN(net_16342), .B2(net_16214), .A(net_15615) );
NAND2_X4 inst_7188 ( .ZN(net_10152), .A2(net_8706), .A1(net_4995) );
INV_X2 inst_19217 ( .ZN(net_3475), .A(net_3474) );
OAI21_X4 inst_1357 ( .ZN(net_18260), .B2(net_18192), .A(net_18164), .B1(net_17244) );
INV_X2 inst_18969 ( .ZN(net_8583), .A(net_5229) );
NAND2_X2 inst_10938 ( .A2(net_20785), .ZN(net_9985), .A1(net_5205) );
NAND2_X2 inst_9547 ( .A1(net_14657), .ZN(net_11036), .A2(net_10924) );
AND2_X2 inst_21361 ( .A2(net_3780), .ZN(net_2424), .A1(net_154) );
NAND4_X2 inst_5302 ( .ZN(net_15898), .A4(net_15262), .A2(net_15190), .A1(net_14929), .A3(net_13084) );
NOR2_X2 inst_4476 ( .A2(net_20851), .ZN(net_5121), .A1(net_3024) );
NAND2_X2 inst_11307 ( .ZN(net_8236), .A1(net_6636), .A2(net_4035) );
NAND2_X4 inst_6861 ( .ZN(net_18372), .A2(net_18302), .A1(net_18264) );
OAI21_X2 inst_2288 ( .B1(net_6589), .ZN(net_6523), .A(net_6480), .B2(net_3303) );
INV_X4 inst_13644 ( .ZN(net_9122), .A(net_8162) );
AOI211_X2 inst_21020 ( .ZN(net_15042), .C1(net_14743), .C2(net_13498), .A(net_4830), .B(net_4755) );
NAND2_X2 inst_11505 ( .ZN(net_5665), .A2(net_3053), .A1(net_1617) );
NOR2_X2 inst_4841 ( .ZN(net_7128), .A2(net_7002), .A1(net_3187) );
NAND2_X2 inst_9368 ( .ZN(net_12119), .A1(net_12118), .A2(net_12117) );
OAI21_X2 inst_1834 ( .B1(net_20730), .ZN(net_14050), .A(net_8611), .B2(net_4201) );
INV_X2 inst_18870 ( .ZN(net_9306), .A(net_6276) );
INV_X4 inst_17989 ( .A(net_21057), .ZN(net_544) );
NOR2_X2 inst_3574 ( .ZN(net_12721), .A1(net_12720), .A2(net_10905) );
OAI21_X2 inst_2228 ( .ZN(net_19401), .B1(net_9940), .B2(net_8442), .A(net_2658) );
INV_X2 inst_18864 ( .A(net_9999), .ZN(net_6291) );
SDFF_X2 inst_768 ( .Q(net_20939), .SE(net_18859), .SI(net_18497), .D(net_14826), .CK(net_22744) );
OAI21_X2 inst_2121 ( .ZN(net_20056), .A(net_11442), .B2(net_7958), .B1(net_3782) );
NOR2_X2 inst_4850 ( .ZN(net_9611), .A2(net_2974), .A1(net_816) );
NAND2_X2 inst_12067 ( .A1(net_20881), .ZN(net_1061), .A2(net_761) );
NAND3_X2 inst_6639 ( .ZN(net_8956), .A2(net_8093), .A1(net_4941), .A3(net_4445) );
INV_X4 inst_16450 ( .A(net_10521), .ZN(net_8722) );
NAND2_X2 inst_11001 ( .ZN(net_4889), .A2(net_3951), .A1(net_2274) );
INV_X4 inst_13225 ( .ZN(net_13599), .A(net_13598) );
AOI21_X2 inst_20759 ( .ZN(net_11180), .B2(net_11179), .A(net_7884), .B1(net_3404) );
INV_X2 inst_19272 ( .A(net_4280), .ZN(net_3022) );
NAND3_X2 inst_6774 ( .ZN(net_4980), .A1(net_4681), .A2(net_4088), .A3(net_2942) );
NOR2_X2 inst_3494 ( .A1(net_14820), .ZN(net_14198), .A2(net_14197) );
INV_X2 inst_18960 ( .A(net_12994), .ZN(net_5440) );
INV_X4 inst_17172 ( .ZN(net_19205), .A(net_2585) );
OAI21_X2 inst_1867 ( .ZN(net_13735), .A(net_13734), .B1(net_12734), .B2(net_10980) );
INV_X2 inst_18997 ( .ZN(net_6163), .A(net_5066) );
INV_X4 inst_17165 ( .ZN(net_5472), .A(net_2585) );
INV_X4 inst_13627 ( .A(net_10437), .ZN(net_9782) );
NAND3_X2 inst_6314 ( .ZN(net_12739), .A2(net_12738), .A3(net_12737), .A1(net_5645) );
NAND2_X4 inst_7580 ( .ZN(net_3096), .A1(net_1584), .A2(net_1583) );
INV_X2 inst_18882 ( .A(net_8288), .ZN(net_6181) );
NAND2_X4 inst_7046 ( .A2(net_19847), .A1(net_19846), .ZN(net_19444) );
AOI21_X2 inst_20577 ( .B1(net_14166), .ZN(net_14102), .B2(net_10645), .A(net_10362) );
CLKBUF_X2 inst_22700 ( .A(net_22571), .Z(net_22572) );
AOI21_X2 inst_20382 ( .ZN(net_15541), .A(net_15156), .B2(net_14609), .B1(net_7429) );
INV_X4 inst_13782 ( .ZN(net_9209), .A(net_7574) );
NAND2_X2 inst_7909 ( .ZN(net_18466), .A1(net_18415), .A2(net_17823) );
NAND3_X2 inst_5670 ( .A3(net_19635), .A1(net_19634), .ZN(net_16375), .A2(net_14809) );
INV_X4 inst_15222 ( .A(net_2868), .ZN(net_2867) );
NAND3_X2 inst_6791 ( .ZN(net_11126), .A1(net_9542), .A2(net_4039), .A3(net_4038) );
INV_X4 inst_15862 ( .ZN(net_1809), .A(net_1808) );
CLKBUF_X2 inst_22806 ( .A(net_22677), .Z(net_22678) );
INV_X4 inst_13695 ( .ZN(net_11021), .A(net_9572) );
INV_X4 inst_12575 ( .ZN(net_18180), .A(net_18179) );
INV_X4 inst_14143 ( .A(net_9954), .ZN(net_6066) );
NOR2_X2 inst_4912 ( .A2(net_7002), .ZN(net_4244), .A1(net_193) );
NOR2_X2 inst_3342 ( .ZN(net_18148), .A2(net_18147), .A1(net_18086) );
NOR2_X2 inst_4825 ( .ZN(net_3607), .A1(net_1848), .A2(net_1816) );
NAND2_X2 inst_9832 ( .ZN(net_9602), .A2(net_9601), .A1(net_9345) );
AOI21_X2 inst_20290 ( .ZN(net_16193), .B2(net_15871), .A(net_14683), .B1(net_1052) );
INV_X4 inst_14666 ( .ZN(net_11729), .A(net_5071) );
NAND2_X2 inst_8175 ( .A2(net_18715), .ZN(net_17940), .A1(net_17924) );
NOR2_X2 inst_3895 ( .ZN(net_9153), .A1(net_9152), .A2(net_9151) );
CLKBUF_X2 inst_21888 ( .A(net_21523), .Z(net_21760) );
XNOR2_X2 inst_303 ( .B(net_21197), .ZN(net_17105), .A(net_17104) );
INV_X4 inst_13518 ( .ZN(net_12836), .A(net_9391) );
INV_X4 inst_14324 ( .ZN(net_7192), .A(net_5442) );
OAI22_X2 inst_1275 ( .B1(net_21141), .ZN(net_16929), .A2(net_16622), .B2(net_16554), .A1(net_726) );
INV_X2 inst_18362 ( .ZN(net_18116), .A(net_18098) );
XOR2_X2 inst_26 ( .B(net_21124), .A(net_16501), .Z(net_16500) );
AOI21_X2 inst_20583 ( .ZN(net_14039), .B1(net_14038), .B2(net_10143), .A(net_9980) );
INV_X4 inst_15326 ( .ZN(net_4859), .A(net_1967) );
INV_X4 inst_13052 ( .ZN(net_16716), .A(net_16556) );
NAND2_X2 inst_10480 ( .A2(net_8546), .ZN(net_6972), .A1(net_6971) );
NAND2_X2 inst_8104 ( .ZN(net_18115), .A2(net_18112), .A1(net_17625) );
NAND2_X2 inst_10198 ( .A2(net_9801), .ZN(net_8133), .A1(net_7962) );
INV_X4 inst_17096 ( .A(net_6849), .ZN(net_6177) );
INV_X4 inst_12731 ( .A(net_17458), .ZN(net_17457) );
INV_X4 inst_14038 ( .ZN(net_9594), .A(net_6270) );
NAND2_X2 inst_10001 ( .A2(net_12109), .ZN(net_8819), .A1(net_8478) );
NAND3_X2 inst_6530 ( .ZN(net_10603), .A2(net_10449), .A1(net_9632), .A3(net_7302) );
CLKBUF_X2 inst_22331 ( .A(net_22202), .Z(net_22203) );
NAND2_X4 inst_7490 ( .A1(net_18965), .ZN(net_3212), .A2(net_818) );
INV_X4 inst_12895 ( .A(net_16864), .ZN(net_16788) );
CLKBUF_X2 inst_21529 ( .A(net_21255), .Z(net_21401) );
AND2_X4 inst_21226 ( .A1(net_14865), .A2(net_11211), .ZN(net_5151) );
NOR2_X2 inst_4864 ( .A1(net_6606), .ZN(net_4172), .A2(net_1285) );
INV_X4 inst_15900 ( .ZN(net_2663), .A(net_1770) );
INV_X4 inst_16211 ( .A(net_8674), .ZN(net_2302) );
NOR2_X2 inst_3765 ( .ZN(net_10302), .A1(net_9201), .A2(net_6775) );
CLKBUF_X2 inst_21689 ( .A(net_21560), .Z(net_21561) );
INV_X4 inst_15924 ( .A(net_9968), .ZN(net_2903) );
INV_X4 inst_17056 ( .ZN(net_15602), .A(net_14014) );
NOR2_X2 inst_4218 ( .A1(net_7610), .ZN(net_6630), .A2(net_6629) );
NAND2_X2 inst_7718 ( .ZN(net_18844), .A1(net_18810), .A2(net_18793) );
AOI21_X4 inst_20235 ( .B1(net_19787), .ZN(net_12297), .A(net_8836), .B2(net_6902) );
INV_X4 inst_15808 ( .ZN(net_3181), .A(net_1382) );
NAND2_X2 inst_10062 ( .A1(net_13703), .ZN(net_8679), .A2(net_8678) );
NAND3_X2 inst_6456 ( .ZN(net_19859), .A3(net_10573), .A1(net_9505), .A2(net_5827) );
INV_X4 inst_16689 ( .ZN(net_7962), .A(net_3760) );
INV_X4 inst_17511 ( .A(net_493), .ZN(net_411) );
INV_X4 inst_16720 ( .ZN(net_10831), .A(net_2311) );
NAND2_X4 inst_7064 ( .A2(net_20896), .A1(net_19101), .ZN(net_16248) );
INV_X4 inst_18020 ( .A(net_20857), .ZN(net_72) );
NAND2_X2 inst_11636 ( .ZN(net_3318), .A1(net_1060), .A2(net_809) );
INV_X4 inst_13702 ( .ZN(net_13914), .A(net_7880) );
NAND2_X4 inst_7623 ( .ZN(net_2485), .A1(net_1299), .A2(net_781) );
NAND2_X2 inst_11469 ( .A1(net_10309), .ZN(net_3154), .A2(net_3153) );
NOR2_X2 inst_5053 ( .ZN(net_1465), .A1(net_1044), .A2(net_1043) );
INV_X4 inst_15137 ( .ZN(net_4055), .A(net_2334) );
INV_X2 inst_18373 ( .A(net_17515), .ZN(net_17456) );
INV_X4 inst_17484 ( .ZN(net_3984), .A(net_539) );
OAI21_X4 inst_1438 ( .B2(net_18922), .B1(net_18921), .A(net_16347), .ZN(net_15916) );
CLKBUF_X2 inst_22581 ( .A(net_21469), .Z(net_22453) );
NAND2_X2 inst_10454 ( .ZN(net_12175), .A2(net_6860), .A1(net_1298) );
NAND3_X2 inst_6373 ( .A2(net_13941), .ZN(net_12055), .A1(net_11854), .A3(net_9381) );
INV_X4 inst_17795 ( .ZN(net_6078), .A(net_308) );
INV_X4 inst_18005 ( .A(net_21153), .ZN(net_742) );
INV_X4 inst_12681 ( .ZN(net_17727), .A(net_17726) );
SDFF_X2 inst_880 ( .Q(net_21188), .SI(net_16889), .SE(net_125), .CK(net_22291), .D(x6404) );
INV_X8 inst_12241 ( .ZN(net_5136), .A(net_1924) );
NAND2_X2 inst_11437 ( .ZN(net_3327), .A2(net_1414), .A1(net_1339) );
INV_X4 inst_16596 ( .ZN(net_2597), .A(net_131) );
NOR3_X2 inst_2681 ( .ZN(net_14569), .A3(net_11760), .A1(net_8861), .A2(net_8479) );
NOR2_X2 inst_3445 ( .A1(net_16035), .ZN(net_14952), .A2(net_13609) );
CLKBUF_X2 inst_22654 ( .A(net_22525), .Z(net_22526) );
NAND2_X2 inst_9118 ( .ZN(net_14838), .A1(net_13565), .A2(net_13564) );
INV_X8 inst_12370 ( .ZN(net_990), .A(net_205) );
CLKBUF_X2 inst_22519 ( .A(net_21517), .Z(net_22391) );
INV_X4 inst_16023 ( .ZN(net_4530), .A(net_1638) );
NAND2_X2 inst_9044 ( .ZN(net_14048), .A1(net_13999), .A2(net_12034) );
NOR2_X2 inst_3972 ( .ZN(net_8406), .A1(net_4565), .A2(net_4096) );
NAND3_X2 inst_6670 ( .A2(net_14643), .A3(net_14078), .ZN(net_7770), .A1(net_7769) );
NAND2_X2 inst_11633 ( .ZN(net_3907), .A2(net_2523), .A1(net_1582) );
INV_X4 inst_17186 ( .ZN(net_15353), .A(net_278) );
OAI21_X4 inst_1388 ( .A(net_20968), .B2(net_19995), .B1(net_19994), .ZN(net_19356) );
AOI21_X2 inst_20936 ( .A(net_6884), .ZN(net_6498), .B2(net_6497), .B1(net_4241) );
NOR3_X2 inst_2699 ( .ZN(net_14093), .A2(net_11255), .A3(net_10483), .A1(net_8863) );
NOR2_X2 inst_3517 ( .ZN(net_13782), .A1(net_13781), .A2(net_12465) );
NAND2_X2 inst_9291 ( .ZN(net_14242), .A2(net_10764), .A1(net_9018) );
INV_X4 inst_14927 ( .A(net_4109), .ZN(net_3556) );
NAND2_X2 inst_8506 ( .ZN(net_16925), .A2(net_16540), .A1(net_8089) );
NOR2_X2 inst_3396 ( .ZN(net_15973), .A2(net_15660), .A1(net_15041) );
OAI21_X4 inst_1372 ( .ZN(net_20356), .B2(net_20228), .B1(net_20227), .A(net_16260) );
NAND2_X4 inst_7332 ( .ZN(net_6079), .A1(net_3589), .A2(net_1848) );
AOI21_X2 inst_20767 ( .ZN(net_10722), .A(net_9984), .B1(net_6913), .B2(net_6671) );
AOI21_X2 inst_20356 ( .ZN(net_19760), .B2(net_15011), .A(net_13334), .B1(net_869) );
NAND2_X2 inst_12109 ( .ZN(net_313), .A2(net_312), .A1(net_291) );
CLKBUF_X2 inst_21929 ( .A(net_21771), .Z(net_21801) );
NAND2_X2 inst_10631 ( .A1(net_12409), .ZN(net_6454), .A2(net_2698) );
NAND2_X2 inst_9759 ( .ZN(net_13149), .A1(net_9966), .A2(net_6234) );
NAND3_X2 inst_6081 ( .ZN(net_13967), .A1(net_13966), .A3(net_13965), .A2(net_12079) );
NOR3_X2 inst_2761 ( .ZN(net_10578), .A3(net_7973), .A2(net_7937), .A1(net_4084) );
CLKBUF_X2 inst_22044 ( .A(net_21915), .Z(net_21916) );
SDFF_X2 inst_989 ( .QN(net_21060), .SE(net_17277), .D(net_653), .CK(net_21250), .SI(x2042) );
INV_X4 inst_15087 ( .A(net_4468), .ZN(net_4325) );
OAI21_X2 inst_2283 ( .A(net_13996), .ZN(net_6577), .B2(net_3261), .B1(net_2792) );
CLKBUF_X2 inst_21565 ( .A(net_21436), .Z(net_21437) );
SDFF_X2 inst_858 ( .Q(net_21165), .SE(net_17277), .D(net_17174), .CK(net_21400), .SI(x5099) );
INV_X2 inst_19080 ( .A(net_6040), .ZN(net_4593) );
CLKBUF_X2 inst_22112 ( .A(net_21608), .Z(net_21984) );
NAND2_X2 inst_9111 ( .A1(net_14216), .ZN(net_13583), .A2(net_13582) );
INV_X4 inst_13779 ( .ZN(net_7578), .A(net_7577) );
NAND2_X2 inst_12060 ( .ZN(net_1320), .A2(net_897), .A1(net_834) );
NOR2_X4 inst_2936 ( .A2(net_13734), .A1(net_10247), .ZN(net_8777) );
OAI211_X2 inst_2468 ( .ZN(net_13911), .B(net_13910), .A(net_12058), .C2(net_7735), .C1(net_1145) );
XOR2_X1 inst_54 ( .B(net_21153), .Z(net_17778), .A(net_17777) );
INV_X4 inst_12610 ( .ZN(net_19192), .A(net_18078) );
NAND2_X2 inst_10556 ( .ZN(net_12109), .A1(net_8190), .A2(net_4954) );
OAI21_X4 inst_1482 ( .B1(net_20636), .ZN(net_14464), .A(net_14463), .B2(net_13025) );
OAI21_X4 inst_1420 ( .B2(net_18968), .B1(net_18967), .A(net_16390), .ZN(net_16116) );
INV_X2 inst_18678 ( .A(net_12105), .ZN(net_8813) );
CLKBUF_X2 inst_21758 ( .A(net_21629), .Z(net_21630) );
INV_X8 inst_12177 ( .ZN(net_17590), .A(net_17109) );
INV_X4 inst_12988 ( .ZN(net_16637), .A(net_16494) );
CLKBUF_X2 inst_22310 ( .A(net_21817), .Z(net_22182) );
NAND4_X2 inst_5337 ( .ZN(net_15517), .A1(net_14520), .A2(net_13855), .A4(net_13405), .A3(net_8778) );
NOR2_X2 inst_4062 ( .A1(net_10405), .ZN(net_7820), .A2(net_7819) );
NAND3_X2 inst_5730 ( .ZN(net_20161), .A1(net_15853), .A3(net_15140), .A2(net_11328) );
INV_X4 inst_16819 ( .ZN(net_9972), .A(net_2280) );
INV_X4 inst_15775 ( .ZN(net_16046), .A(net_15917) );
INV_X4 inst_15685 ( .ZN(net_3492), .A(net_2037) );
NOR2_X2 inst_4108 ( .ZN(net_7172), .A2(net_5298), .A1(net_4729) );
NOR2_X2 inst_4626 ( .ZN(net_3603), .A1(net_3105), .A2(net_2681) );
NAND2_X2 inst_8780 ( .ZN(net_15803), .A2(net_15293), .A1(net_10858) );
NAND2_X2 inst_9491 ( .ZN(net_11438), .A2(net_11437), .A1(net_9409) );
NAND2_X2 inst_11595 ( .A1(net_7844), .ZN(net_7840), .A2(net_2672) );
INV_X4 inst_15496 ( .ZN(net_6993), .A(net_1670) );
INV_X4 inst_15272 ( .ZN(net_5082), .A(net_2761) );
XNOR2_X2 inst_497 ( .A(net_16546), .ZN(net_9004), .B(net_1874) );
INV_X4 inst_13826 ( .ZN(net_10888), .A(net_7506) );
NAND2_X4 inst_7517 ( .ZN(net_4256), .A1(net_2071), .A2(net_1819) );
INV_X4 inst_18320 ( .A(net_20534), .ZN(net_20533) );
INV_X2 inst_19414 ( .A(net_3146), .ZN(net_1932) );
INV_X4 inst_15919 ( .ZN(net_11494), .A(net_10134) );
OAI21_X2 inst_2195 ( .ZN(net_8582), .B2(net_8581), .B1(net_4509), .A(net_1471) );
NAND2_X2 inst_8787 ( .ZN(net_15752), .A1(net_15628), .A2(net_15161) );
OAI221_X2 inst_1335 ( .ZN(net_15367), .A(net_14347), .B2(net_12798), .C2(net_12293), .C1(net_5166), .B1(net_3180) );
AND2_X4 inst_21221 ( .ZN(net_12805), .A1(net_5450), .A2(net_4448) );
INV_X4 inst_15197 ( .ZN(net_4675), .A(net_2306) );
NAND2_X2 inst_9924 ( .A1(net_14689), .ZN(net_9233), .A2(net_6435) );
NOR2_X2 inst_3845 ( .ZN(net_10991), .A1(net_8502), .A2(net_7548) );
NAND2_X4 inst_7173 ( .ZN(net_12999), .A2(net_9396), .A1(net_9338) );
NAND2_X2 inst_10124 ( .A1(net_10383), .ZN(net_8365), .A2(net_8364) );
NAND4_X4 inst_5168 ( .A4(net_18887), .A1(net_18886), .ZN(net_17110), .A2(net_16342), .A3(net_8106) );
NOR2_X4 inst_3128 ( .ZN(net_4435), .A2(net_3904), .A1(net_3566) );
DFF_X1 inst_19824 ( .D(net_17778), .CK(net_21620), .Q(x598) );
NAND2_X2 inst_10715 ( .ZN(net_11629), .A2(net_5933), .A1(net_4907) );
INV_X4 inst_17749 ( .A(net_4850), .ZN(net_4718) );
INV_X4 inst_14653 ( .ZN(net_13956), .A(net_4368) );
OAI211_X2 inst_2517 ( .ZN(net_11899), .B(net_11898), .C1(net_11897), .A(net_6291), .C2(net_3717) );
NOR2_X2 inst_4183 ( .ZN(net_6793), .A1(net_6792), .A2(net_4431) );
NAND2_X2 inst_10806 ( .A1(net_8334), .ZN(net_5541), .A2(net_3395) );
CLKBUF_X2 inst_22821 ( .A(net_22692), .Z(net_22693) );
SDFF_X2 inst_714 ( .Q(net_20856), .SE(net_18847), .SI(net_18796), .D(net_531), .CK(net_22019) );
INV_X4 inst_15735 ( .ZN(net_15708), .A(net_14500) );
INV_X4 inst_15518 ( .A(net_11682), .ZN(net_11617) );
NOR2_X4 inst_3005 ( .ZN(net_7574), .A1(net_4588), .A2(net_3332) );
NOR2_X4 inst_2895 ( .ZN(net_12847), .A1(net_9410), .A2(net_9401) );
NAND2_X2 inst_9005 ( .ZN(net_19953), .A2(net_13491), .A1(net_9260) );
INV_X4 inst_16199 ( .A(net_12203), .ZN(net_2408) );
OR3_X2 inst_1061 ( .A3(net_13206), .A1(net_8969), .ZN(net_8968), .A2(net_8967) );
NAND2_X2 inst_11201 ( .ZN(net_5202), .A2(net_4065), .A1(net_2585) );
CLKBUF_X2 inst_22083 ( .A(net_21551), .Z(net_21955) );
OAI21_X2 inst_2326 ( .ZN(net_5542), .A(net_2696), .B1(net_2340), .B2(net_1976) );
NAND3_X2 inst_6657 ( .ZN(net_8470), .A3(net_8469), .A2(net_6034), .A1(net_3928) );
INV_X4 inst_18183 ( .A(net_21229), .ZN(net_855) );
XNOR2_X2 inst_72 ( .ZN(net_18760), .B(net_18683), .A(net_17631) );
NAND2_X4 inst_6967 ( .ZN(net_17414), .A1(net_17012), .A2(net_16865) );
AOI21_X2 inst_20284 ( .B2(net_19004), .B1(net_19003), .A(net_16394), .ZN(net_16252) );
NAND2_X2 inst_11703 ( .ZN(net_2301), .A2(net_1313), .A1(net_168) );
INV_X4 inst_17920 ( .A(net_21092), .ZN(net_491) );
OAI21_X2 inst_1634 ( .ZN(net_15984), .B2(net_15609), .A(net_12252), .B1(net_1930) );
INV_X4 inst_15961 ( .ZN(net_3581), .A(net_1701) );
NAND2_X2 inst_8998 ( .ZN(net_14299), .A2(net_14298), .A1(net_13238) );
NAND2_X2 inst_7980 ( .ZN(net_18340), .A2(net_18339), .A1(net_18137) );
CLKBUF_X2 inst_22107 ( .A(net_21486), .Z(net_21979) );
NAND2_X2 inst_10619 ( .ZN(net_7842), .A1(net_6580), .A2(net_6579) );
NAND3_X2 inst_6729 ( .ZN(net_19756), .A2(net_6487), .A1(net_5665), .A3(net_1615) );
INV_X2 inst_19278 ( .ZN(net_2946), .A(net_2945) );
NAND3_X2 inst_6650 ( .ZN(net_8551), .A1(net_8550), .A3(net_7093), .A2(net_6646) );
AOI21_X2 inst_20427 ( .B1(net_19179), .ZN(net_15206), .B2(net_15205), .A(net_8731) );
CLKBUF_X2 inst_22559 ( .A(net_22430), .Z(net_22431) );
INV_X2 inst_19114 ( .A(net_14075), .ZN(net_8416) );
INV_X4 inst_15609 ( .ZN(net_19861), .A(net_2189) );
NAND2_X2 inst_9485 ( .ZN(net_14342), .A1(net_11451), .A2(net_11450) );
AOI21_X4 inst_20182 ( .ZN(net_15335), .B1(net_15334), .B2(net_13684), .A(net_12101) );
INV_X8 inst_12415 ( .A(net_20909), .ZN(net_879) );
INV_X8 inst_12357 ( .ZN(net_1662), .A(net_1347) );
NOR2_X2 inst_4638 ( .ZN(net_5958), .A2(net_3904), .A1(net_3481) );
AOI22_X2 inst_19998 ( .ZN(net_14176), .A1(net_14175), .B1(net_14174), .A2(net_10775), .B2(net_9965) );
NAND2_X2 inst_11487 ( .A1(net_8160), .ZN(net_4007), .A2(net_3094) );
INV_X4 inst_13426 ( .ZN(net_13199), .A(net_8503) );
OAI21_X2 inst_1582 ( .A(net_16743), .ZN(net_16309), .B2(net_15996), .B1(net_7841) );
INV_X4 inst_16122 ( .ZN(net_11182), .A(net_6112) );
INV_X4 inst_13202 ( .ZN(net_13859), .A(net_13178) );
AOI21_X2 inst_20846 ( .ZN(net_20134), .A(net_9254), .B2(net_4417), .B1(net_2159) );
INV_X4 inst_17585 ( .ZN(net_2646), .A(net_1660) );
NAND3_X2 inst_6334 ( .ZN(net_12448), .A2(net_12447), .A3(net_12446), .A1(net_4886) );
INV_X4 inst_13905 ( .ZN(net_7622), .A(net_7057) );
NAND3_X2 inst_5846 ( .ZN(net_15442), .A1(net_15385), .A3(net_14499), .A2(net_13822) );
INV_X2 inst_18858 ( .ZN(net_6331), .A(net_6330) );
OAI21_X2 inst_1840 ( .A(net_15452), .ZN(net_14026), .B2(net_10273), .B1(net_3739) );
NAND3_X2 inst_6345 ( .ZN(net_12244), .A3(net_12243), .A1(net_9848), .A2(net_6645) );
AOI222_X2 inst_20061 ( .A1(net_20389), .A2(net_16402), .ZN(net_16162), .B1(net_15976), .C2(net_14660), .B2(net_13119), .C1(net_10048) );
XNOR2_X2 inst_133 ( .ZN(net_18225), .A(net_18187), .B(net_18141) );
INV_X4 inst_17805 ( .A(net_131), .ZN(net_122) );
CLKBUF_X2 inst_22731 ( .A(net_22602), .Z(net_22603) );
INV_X4 inst_14734 ( .ZN(net_7772), .A(net_4114) );
INV_X4 inst_13847 ( .ZN(net_13483), .A(net_10337) );
CLKBUF_X2 inst_21384 ( .A(net_21253), .Z(net_21256) );
INV_X4 inst_16587 ( .ZN(net_9745), .A(net_4990) );
INV_X2 inst_18955 ( .ZN(net_5533), .A(net_5532) );
NAND2_X2 inst_9988 ( .ZN(net_10332), .A2(net_8308), .A1(net_8260) );
INV_X2 inst_18552 ( .A(net_12944), .ZN(net_10905) );
INV_X4 inst_14688 ( .ZN(net_5952), .A(net_2730) );
OAI21_X2 inst_1721 ( .ZN(net_15115), .B2(net_12919), .B1(net_7042), .A(net_1030) );
AOI221_X2 inst_20078 ( .ZN(net_19556), .C1(net_16037), .B1(net_15955), .C2(net_15599), .B2(net_13694), .A(net_6516) );
NAND2_X2 inst_9744 ( .ZN(net_10094), .A1(net_10093), .A2(net_7674) );
NAND2_X2 inst_10884 ( .A2(net_12954), .A1(net_8330), .ZN(net_5412) );
INV_X2 inst_18930 ( .ZN(net_9181), .A(net_5856) );
INV_X4 inst_12854 ( .ZN(net_17064), .A(net_17063) );
XNOR2_X2 inst_126 ( .ZN(net_18373), .A(net_18203), .B(net_17046) );
INV_X2 inst_19454 ( .A(net_1761), .ZN(net_1532) );
INV_X2 inst_18413 ( .ZN(net_15989), .A(net_15877) );
CLKBUF_X2 inst_22825 ( .A(net_22696), .Z(net_22697) );
NOR2_X2 inst_3887 ( .ZN(net_9245), .A1(net_6371), .A2(net_5939) );
CLKBUF_X2 inst_21846 ( .A(net_21639), .Z(net_21718) );
INV_X4 inst_14163 ( .ZN(net_9320), .A(net_6015) );
OAI21_X2 inst_1631 ( .ZN(net_16020), .A(net_15974), .B2(net_15458), .B1(net_6300) );
INV_X2 inst_19292 ( .ZN(net_2850), .A(net_2849) );
INV_X4 inst_12651 ( .ZN(net_17860), .A(net_17859) );
NAND2_X4 inst_7510 ( .ZN(net_3986), .A2(net_1753), .A1(net_1220) );
INV_X4 inst_13106 ( .ZN(net_15736), .A(net_15530) );
OR2_X4 inst_1086 ( .A1(net_9490), .ZN(net_8410), .A2(net_5211) );
AOI21_X2 inst_20343 ( .B1(net_20145), .ZN(net_19393), .B2(net_15343), .A(net_15189) );
INV_X4 inst_14360 ( .ZN(net_9945), .A(net_5233) );
NOR3_X2 inst_2643 ( .ZN(net_15900), .A3(net_15389), .A1(net_15215), .A2(net_10005) );
NAND2_X2 inst_12088 ( .ZN(net_704), .A2(net_703), .A1(net_124) );
INV_X2 inst_18354 ( .ZN(net_19489), .A(net_18626) );
INV_X4 inst_13950 ( .A(net_8727), .ZN(net_8637) );
INV_X4 inst_12615 ( .ZN(net_18066), .A(net_18058) );
CLKBUF_X2 inst_22087 ( .A(net_21834), .Z(net_21959) );
INV_X4 inst_12713 ( .A(net_17762), .ZN(net_17551) );
OAI21_X2 inst_1688 ( .B1(net_19824), .ZN(net_15395), .A(net_13658), .B2(net_588) );
INV_X4 inst_15621 ( .A(net_11451), .ZN(net_5486) );
INV_X4 inst_13651 ( .ZN(net_13266), .A(net_8151) );
INV_X4 inst_13732 ( .ZN(net_19773), .A(net_6481) );
INV_X4 inst_17481 ( .A(net_8304), .ZN(net_8241) );
NAND2_X1 inst_12146 ( .A2(net_17815), .ZN(net_16661), .A1(net_1895) );
AOI21_X4 inst_20242 ( .ZN(net_19349), .B1(net_19110), .A(net_5099), .B2(net_86) );
INV_X4 inst_14836 ( .ZN(net_14331), .A(net_7125) );
INV_X4 inst_17580 ( .A(net_1529), .ZN(net_340) );
INV_X4 inst_13084 ( .ZN(net_19486), .A(net_15967) );
SDFF_X2 inst_914 ( .Q(net_21116), .D(net_16649), .SE(net_263), .CK(net_22275), .SI(x4496) );
CLKBUF_X2 inst_22872 ( .A(net_22743), .Z(net_22744) );
CLKBUF_X2 inst_21713 ( .A(net_21584), .Z(net_21585) );
AOI21_X4 inst_20225 ( .ZN(net_14030), .A(net_14029), .B2(net_11400), .B1(net_10382) );
NAND3_X2 inst_6364 ( .ZN(net_12080), .A3(net_12079), .A2(net_9676), .A1(net_5222) );
NAND4_X4 inst_5170 ( .A3(net_18998), .A1(net_18997), .ZN(net_17031), .A4(net_16306), .A2(net_13195) );
NAND4_X4 inst_5182 ( .ZN(net_16631), .A1(net_16355), .A2(net_16188), .A3(net_16092), .A4(net_16019) );
INV_X8 inst_12198 ( .ZN(net_16562), .A(net_16336) );
INV_X4 inst_14962 ( .ZN(net_5455), .A(net_2668) );
NAND2_X2 inst_11588 ( .ZN(net_2698), .A1(net_2697), .A2(net_2696) );
XNOR2_X2 inst_384 ( .ZN(net_16800), .A(net_16799), .B(net_16743) );
OAI22_X2 inst_1252 ( .ZN(net_18446), .A2(net_18339), .B2(net_18283), .A1(net_17819), .B1(net_17818) );
INV_X4 inst_12773 ( .ZN(net_17329), .A(net_17328) );
NOR2_X2 inst_3800 ( .ZN(net_9858), .A2(net_9460), .A1(net_6326) );
INV_X4 inst_17568 ( .ZN(net_358), .A(net_170) );
INV_X4 inst_17458 ( .ZN(net_8041), .A(net_522) );
NAND3_X2 inst_6086 ( .ZN(net_13954), .A1(net_12435), .A3(net_11321), .A2(net_11118) );
CLKBUF_X2 inst_22695 ( .A(net_22566), .Z(net_22567) );
INV_X4 inst_12989 ( .ZN(net_19411), .A(net_16426) );
NAND2_X2 inst_10271 ( .ZN(net_9520), .A1(net_7975), .A2(net_7947) );
OAI21_X2 inst_2209 ( .A(net_14460), .ZN(net_8532), .B2(net_3475), .B1(net_3058) );
NOR3_X2 inst_2722 ( .ZN(net_13254), .A1(net_10532), .A3(net_9603), .A2(net_7542) );
INV_X4 inst_13034 ( .A(net_16716), .ZN(net_16590) );
INV_X4 inst_17738 ( .ZN(net_4918), .A(net_1655) );
INV_X2 inst_19093 ( .ZN(net_8287), .A(net_4549) );
INV_X4 inst_16817 ( .ZN(net_3505), .A(net_999) );
OR2_X2 inst_1238 ( .ZN(net_10074), .A2(net_993), .A1(net_816) );
NAND2_X4 inst_7361 ( .ZN(net_4458), .A1(net_4073), .A2(net_3586) );
OAI21_X2 inst_2171 ( .ZN(net_8927), .A(net_8644), .B2(net_6143), .B1(net_1430) );
INV_X4 inst_15385 ( .ZN(net_3568), .A(net_3384) );
NAND2_X2 inst_9031 ( .ZN(net_14072), .A1(net_13091), .A2(net_11887) );
NAND2_X2 inst_7941 ( .ZN(net_18461), .A2(net_18362), .A1(net_18304) );
NAND2_X2 inst_8527 ( .ZN(net_16871), .A2(net_16870), .A1(net_430) );
CLKBUF_X2 inst_22922 ( .A(net_21367), .Z(net_22794) );
CLKBUF_X2 inst_22717 ( .A(net_22588), .Z(net_22589) );
NOR2_X2 inst_3402 ( .A2(net_18873), .ZN(net_15822), .A1(net_15109) );
INV_X2 inst_18616 ( .ZN(net_9606), .A(net_9605) );
INV_X4 inst_14318 ( .ZN(net_5463), .A(net_5462) );
SDFF_X2 inst_1011 ( .QN(net_21043), .D(net_613), .SE(net_263), .CK(net_22499), .SI(x2272) );
XNOR2_X2 inst_404 ( .ZN(net_16652), .A(net_16650), .B(net_1676) );
NAND3_X2 inst_5838 ( .ZN(net_15509), .A1(net_14637), .A3(net_14573), .A2(net_13524) );
NOR2_X2 inst_3615 ( .ZN(net_19573), .A1(net_10652), .A2(net_6239) );
NAND2_X2 inst_9628 ( .ZN(net_10547), .A2(net_7201), .A1(net_171) );
NOR2_X4 inst_3216 ( .ZN(net_6512), .A2(net_3225), .A1(net_2855) );
NAND2_X2 inst_8748 ( .ZN(net_15981), .A2(net_15822), .A1(net_15059) );
INV_X4 inst_15093 ( .ZN(net_14315), .A(net_8991) );
INV_X2 inst_19499 ( .ZN(net_1267), .A(net_1266) );
INV_X4 inst_18228 ( .ZN(net_32), .A(net_26) );
INV_X4 inst_15489 ( .A(net_11550), .ZN(net_11440) );
INV_X2 inst_19428 ( .A(net_2299), .ZN(net_1782) );
NOR2_X2 inst_3540 ( .ZN(net_13401), .A1(net_11217), .A2(net_10473) );
CLKBUF_X2 inst_22921 ( .A(net_22792), .Z(net_22793) );
INV_X4 inst_15277 ( .ZN(net_8539), .A(net_2742) );
NAND2_X4 inst_7701 ( .ZN(net_932), .A2(net_386), .A1(net_289) );
INV_X4 inst_17723 ( .ZN(net_1529), .A(net_880) );
INV_X4 inst_14005 ( .ZN(net_6345), .A(net_6344) );
NAND2_X2 inst_10904 ( .ZN(net_12126), .A1(net_7975), .A2(net_5371) );
INV_X2 inst_18541 ( .ZN(net_19062), .A(net_11009) );
OAI211_X2 inst_2413 ( .ZN(net_15520), .C1(net_15519), .B(net_14652), .A(net_14321), .C2(net_12857) );
OAI21_X2 inst_1574 ( .A(net_20864), .ZN(net_16343), .B1(net_16100), .B2(net_15824) );
INV_X1 inst_19762 ( .ZN(net_3875), .A(net_3101) );
INV_X2 inst_18755 ( .ZN(net_7671), .A(net_6393) );
INV_X4 inst_16549 ( .ZN(net_2332), .A(net_1172) );
NAND2_X4 inst_7528 ( .ZN(net_3850), .A2(net_1990), .A1(net_1847) );
INV_X4 inst_14518 ( .ZN(net_4797), .A(net_4796) );
XNOR2_X2 inst_228 ( .ZN(net_17499), .A(net_17250), .B(net_16931) );
CLKBUF_X2 inst_22729 ( .A(net_22600), .Z(net_22601) );
AOI21_X4 inst_20198 ( .ZN(net_20432), .B1(net_18911), .B2(net_13383), .A(net_7697) );
INV_X4 inst_14034 ( .ZN(net_9813), .A(net_5154) );
NAND2_X4 inst_6872 ( .ZN(net_18271), .A1(net_18146), .A2(net_18123) );
NAND2_X2 inst_12008 ( .ZN(net_6387), .A1(net_4918), .A2(net_3675) );
INV_X2 inst_19019 ( .ZN(net_4970), .A(net_4969) );
INV_X8 inst_12279 ( .ZN(net_2168), .A(net_815) );
NAND2_X2 inst_8759 ( .ZN(net_18993), .A2(net_15527), .A1(net_12861) );
XNOR2_X2 inst_244 ( .B(net_21112), .ZN(net_17319), .A(net_16980) );
INV_X2 inst_18801 ( .A(net_9512), .ZN(net_7417) );
INV_X4 inst_17881 ( .ZN(net_79), .A(net_78) );
INV_X4 inst_13514 ( .A(net_11824), .ZN(net_11450) );
NAND4_X2 inst_5262 ( .A2(net_20345), .A1(net_20344), .ZN(net_16200), .A4(net_15392), .A3(net_8527) );
NAND2_X2 inst_11472 ( .ZN(net_8550), .A2(net_2595), .A1(net_1790) );
INV_X4 inst_13464 ( .ZN(net_13596), .A(net_8223) );
NAND2_X1 inst_12136 ( .A1(net_20066), .ZN(net_17477), .A2(net_17236) );
NAND2_X2 inst_11794 ( .ZN(net_9278), .A1(net_5009), .A2(net_1959) );
NAND3_X4 inst_5537 ( .ZN(net_17334), .A3(net_16707), .A2(net_15925), .A1(net_10748) );
AND2_X2 inst_21275 ( .A1(net_14751), .ZN(net_14069), .A2(net_11879) );
INV_X2 inst_18887 ( .ZN(net_18920), .A(net_6143) );
NAND2_X2 inst_11339 ( .A2(net_4615), .ZN(net_4522), .A1(net_3641) );
NOR2_X4 inst_3079 ( .ZN(net_6395), .A2(net_4438), .A1(net_547) );
AOI21_X2 inst_20683 ( .ZN(net_12293), .A(net_9225), .B2(net_5272), .B1(net_4377) );
INV_X4 inst_16951 ( .ZN(net_6856), .A(net_911) );
NAND2_X2 inst_10143 ( .ZN(net_8309), .A1(net_7004), .A2(net_6227) );
INV_X4 inst_12529 ( .ZN(net_18415), .A(net_18414) );
NAND4_X2 inst_5487 ( .ZN(net_12289), .A2(net_12076), .A4(net_11822), .A3(net_10627), .A1(net_6716) );
NAND2_X4 inst_7599 ( .ZN(net_2483), .A2(net_807), .A1(net_445) );
NAND2_X2 inst_11789 ( .ZN(net_5288), .A1(net_1163), .A2(net_840) );
NAND2_X2 inst_10303 ( .ZN(net_11836), .A1(net_7872), .A2(net_7871) );
INV_X2 inst_18949 ( .ZN(net_5648), .A(net_4032) );
NOR2_X2 inst_3606 ( .ZN(net_12429), .A2(net_12428), .A1(net_9834) );
XNOR2_X2 inst_93 ( .ZN(net_18551), .B(net_18493), .A(net_18492) );
INV_X4 inst_17192 ( .ZN(net_771), .A(net_322) );
NOR2_X2 inst_4832 ( .ZN(net_20579), .A1(net_3505), .A2(net_2422) );
NAND2_X4 inst_7026 ( .ZN(net_17234), .A1(net_16585), .A2(net_16457) );
INV_X4 inst_14631 ( .A(net_15369), .ZN(net_5567) );
INV_X4 inst_17632 ( .A(net_1080), .ZN(net_286) );
NAND2_X2 inst_12105 ( .ZN(net_7156), .A1(net_3745), .A2(net_790) );
NAND2_X2 inst_7784 ( .A1(net_20473), .ZN(net_18905), .A2(net_18626) );
NOR2_X2 inst_4595 ( .A1(net_6854), .ZN(net_4752), .A2(net_1700) );
OAI21_X2 inst_1675 ( .ZN(net_15546), .B2(net_14626), .B1(net_8612), .A(net_1046) );
CLKBUF_X2 inst_22866 ( .A(net_22737), .Z(net_22738) );
NAND2_X2 inst_11086 ( .ZN(net_9961), .A1(net_7121), .A2(net_4402) );
NOR2_X2 inst_3433 ( .ZN(net_15279), .A1(net_15278), .A2(net_14269) );
INV_X2 inst_19727 ( .A(net_20799), .ZN(net_20798) );
NAND2_X2 inst_11274 ( .A1(net_5120), .ZN(net_4883), .A2(net_2443) );
NOR2_X1 inst_5149 ( .ZN(net_10138), .A1(net_10137), .A2(net_6820) );
NAND2_X2 inst_8958 ( .ZN(net_14715), .A1(net_13530), .A2(net_13208) );
INV_X4 inst_13713 ( .ZN(net_10160), .A(net_7845) );
NOR2_X2 inst_4237 ( .ZN(net_7825), .A1(net_6612), .A2(net_6571) );
NAND2_X2 inst_10709 ( .ZN(net_9386), .A2(net_6153), .A1(net_170) );
XNOR2_X2 inst_148 ( .ZN(net_18039), .A(net_18006), .B(net_17381) );
XNOR2_X2 inst_554 ( .B(net_16921), .ZN(net_708), .A(net_707) );
INV_X4 inst_13675 ( .A(net_9795), .ZN(net_8004) );
INV_X4 inst_13621 ( .ZN(net_9804), .A(net_8356) );
OR2_X2 inst_1187 ( .ZN(net_4550), .A2(net_4336), .A1(net_2202) );
NAND3_X2 inst_6000 ( .ZN(net_14433), .A3(net_13054), .A1(net_12790), .A2(net_11699) );
NAND4_X2 inst_5499 ( .ZN(net_11901), .A4(net_11900), .A3(net_10834), .A2(net_9317), .A1(net_6327) );
INV_X2 inst_19147 ( .ZN(net_4095), .A(net_4094) );
CLKBUF_X2 inst_21652 ( .A(net_21522), .Z(net_21524) );
INV_X4 inst_17963 ( .A(net_21091), .ZN(net_584) );
NAND2_X2 inst_10740 ( .ZN(net_20402), .A1(net_5727), .A2(net_4233) );
NAND2_X2 inst_8951 ( .ZN(net_14724), .A2(net_13315), .A1(net_13058) );
OAI21_X2 inst_1917 ( .ZN(net_13044), .A(net_10831), .B2(net_9551), .B1(net_4035) );
INV_X4 inst_14764 ( .ZN(net_9035), .A(net_5480) );
INV_X2 inst_19060 ( .ZN(net_4697), .A(net_4696) );
AOI21_X2 inst_20317 ( .B1(net_20920), .ZN(net_19558), .A(net_15532), .B2(net_15286) );
INV_X4 inst_15302 ( .A(net_3986), .ZN(net_3601) );
INV_X4 inst_15753 ( .ZN(net_1936), .A(net_1935) );
INV_X4 inst_12695 ( .ZN(net_17639), .A(net_17638) );
NOR2_X2 inst_4955 ( .A2(net_2204), .ZN(net_2184), .A1(net_2050) );
NAND2_X2 inst_11553 ( .ZN(net_2848), .A1(net_2847), .A2(net_2846) );
INV_X8 inst_12386 ( .A(net_272), .ZN(net_205) );
CLKBUF_X2 inst_22313 ( .A(net_22184), .Z(net_22185) );
INV_X4 inst_16292 ( .ZN(net_8822), .A(net_8568) );
CLKBUF_X2 inst_21685 ( .A(net_21556), .Z(net_21557) );
INV_X4 inst_17909 ( .A(net_459), .ZN(net_58) );
OAI21_X2 inst_2087 ( .ZN(net_10378), .A(net_10377), .B2(net_6238), .B1(net_4275) );
AOI21_X2 inst_20971 ( .ZN(net_4671), .A(net_4670), .B2(net_4669), .B1(net_1018) );
INV_X4 inst_16215 ( .ZN(net_3165), .A(net_1393) );
INV_X4 inst_13891 ( .ZN(net_9164), .A(net_7308) );
INV_X4 inst_15671 ( .ZN(net_11907), .A(net_9260) );
INV_X2 inst_19058 ( .ZN(net_4706), .A(net_4705) );
NAND2_X2 inst_9881 ( .A1(net_12542), .ZN(net_9440), .A2(net_5838) );
NAND2_X2 inst_8571 ( .ZN(net_16736), .A2(net_16729), .A1(net_16544) );
AOI21_X2 inst_20912 ( .B2(net_12994), .A(net_7968), .ZN(net_7342), .B1(net_3432) );
INV_X4 inst_16858 ( .A(net_2569), .ZN(net_2264) );
NAND3_X2 inst_6501 ( .ZN(net_19497), .A3(net_5832), .A1(net_4658), .A2(net_3687) );
SDFF_X2 inst_819 ( .Q(net_21137), .SI(net_17677), .SE(net_125), .CK(net_21413), .D(x3732) );
NOR2_X2 inst_4464 ( .ZN(net_5804), .A1(net_4530), .A2(net_4529) );
NOR2_X4 inst_3320 ( .ZN(net_1420), .A2(net_211), .A1(net_123) );
OAI21_X4 inst_1468 ( .B2(net_20132), .B1(net_20131), .ZN(net_15078), .A(net_15077) );
NAND2_X2 inst_9663 ( .ZN(net_13099), .A2(net_8332), .A1(net_1889) );
INV_X4 inst_18068 ( .A(net_21236), .ZN(net_16644) );
NOR2_X2 inst_3776 ( .A1(net_15612), .ZN(net_10173), .A2(net_10172) );
INV_X4 inst_18244 ( .A(net_21243), .ZN(net_1009) );
INV_X4 inst_14046 ( .ZN(net_7614), .A(net_6257) );
AOI21_X2 inst_20469 ( .B1(net_15366), .ZN(net_14993), .B2(net_12920), .A(net_7175) );
INV_X4 inst_16992 ( .ZN(net_1190), .A(net_873) );
NAND2_X2 inst_8857 ( .A1(net_15666), .ZN(net_15351), .A2(net_14425) );
NAND3_X2 inst_5859 ( .ZN(net_15386), .A2(net_15385), .A3(net_14048), .A1(net_11119) );
INV_X4 inst_17641 ( .ZN(net_448), .A(net_143) );
NOR3_X4 inst_2617 ( .A3(net_19699), .A1(net_19698), .ZN(net_15527), .A2(net_10879) );
CLKBUF_X2 inst_21765 ( .A(net_21636), .Z(net_21637) );
DFF_X1 inst_19897 ( .D(net_16942), .CK(net_21318), .Q(x288) );
INV_X2 inst_19515 ( .ZN(net_2109), .A(net_1139) );
NOR2_X2 inst_3942 ( .A2(net_8772), .ZN(net_8647), .A1(net_4892) );
NAND2_X2 inst_9459 ( .ZN(net_11498), .A2(net_11497), .A1(net_10690) );
NOR2_X4 inst_3068 ( .ZN(net_7921), .A1(net_5042), .A2(net_4810) );
CLKBUF_X2 inst_22403 ( .A(net_21428), .Z(net_22275) );
NAND3_X2 inst_5850 ( .ZN(net_15426), .A2(net_15425), .A1(net_14989), .A3(net_12411) );
INV_X2 inst_18716 ( .A(net_11763), .ZN(net_8174) );
OAI21_X2 inst_2277 ( .ZN(net_7131), .B1(net_5573), .A(net_3293), .B2(net_2565) );
NAND2_X2 inst_9518 ( .ZN(net_11143), .A2(net_7412), .A1(net_4129) );
INV_X4 inst_18335 ( .A(net_20582), .ZN(net_20580) );
NAND2_X2 inst_8245 ( .A1(net_17760), .ZN(net_17719), .A2(net_17718) );
AOI21_X2 inst_20896 ( .B1(net_8181), .ZN(net_7766), .B2(net_6119), .A(net_4643) );
INV_X2 inst_19626 ( .A(net_20894), .ZN(net_35) );
NOR2_X4 inst_2962 ( .ZN(net_7864), .A2(net_6951), .A1(net_6629) );
INV_X4 inst_16455 ( .ZN(net_1680), .A(net_1225) );
CLKBUF_X2 inst_22394 ( .A(net_22265), .Z(net_22266) );
INV_X2 inst_18940 ( .ZN(net_5813), .A(net_5812) );
INV_X4 inst_13973 ( .ZN(net_8793), .A(net_6656) );
NAND2_X2 inst_10605 ( .ZN(net_12118), .A2(net_6555), .A1(net_703) );
NAND2_X2 inst_9973 ( .A2(net_10643), .ZN(net_8882), .A1(net_8881) );
XNOR2_X2 inst_208 ( .ZN(net_17644), .B(net_17208), .A(net_17121) );
CLKBUF_X2 inst_21946 ( .A(net_21817), .Z(net_21818) );
INV_X4 inst_13756 ( .ZN(net_10557), .A(net_7614) );
INV_X4 inst_16477 ( .ZN(net_12298), .A(net_1209) );
INV_X4 inst_14272 ( .A(net_5670), .ZN(net_5668) );
INV_X4 inst_15247 ( .ZN(net_2807), .A(net_2806) );
NOR2_X2 inst_4202 ( .ZN(net_8703), .A2(net_4966), .A1(net_952) );
NOR2_X2 inst_3774 ( .A2(net_14387), .ZN(net_12937), .A1(net_3156) );
NAND2_X4 inst_7101 ( .ZN(net_13595), .A1(net_12694), .A2(net_4780) );
INV_X2 inst_19445 ( .A(net_2275), .ZN(net_1626) );
NAND4_X2 inst_5282 ( .ZN(net_15982), .A1(net_15581), .A4(net_14521), .A3(net_12185), .A2(net_3840) );
CLKBUF_X2 inst_21439 ( .A(net_21310), .Z(net_21311) );
INV_X4 inst_12751 ( .ZN(net_17889), .A(net_17413) );
NAND2_X2 inst_11935 ( .ZN(net_3175), .A1(net_1461), .A2(net_1309) );
NAND2_X2 inst_10294 ( .ZN(net_7913), .A1(net_7912), .A2(net_5904) );
AND2_X2 inst_21326 ( .A2(net_5733), .ZN(net_5717), .A1(net_5716) );
XNOR2_X2 inst_636 ( .ZN(net_432), .A(net_431), .B(net_430) );
INV_X4 inst_15823 ( .A(net_14636), .ZN(net_1869) );
INV_X2 inst_18868 ( .A(net_8372), .ZN(net_6280) );
CLKBUF_X2 inst_21675 ( .A(net_21546), .Z(net_21547) );
INV_X4 inst_12499 ( .ZN(net_18639), .A(net_18624) );
NAND2_X2 inst_11777 ( .ZN(net_2036), .A2(net_253), .A1(x3463) );
INV_X4 inst_17208 ( .A(net_897), .ZN(net_751) );
OAI21_X2 inst_1907 ( .ZN(net_13110), .A(net_11007), .B1(net_9742), .B2(net_9494) );
CLKBUF_X2 inst_22322 ( .A(net_22193), .Z(net_22194) );
NAND2_X4 inst_7015 ( .A1(net_19450), .A2(net_16973), .ZN(net_16968) );
NAND2_X2 inst_8384 ( .ZN(net_17435), .A2(net_17055), .A1(net_16920) );
INV_X4 inst_16672 ( .ZN(net_6610), .A(net_154) );
INV_X4 inst_17859 ( .A(net_1790), .ZN(net_93) );
NAND2_X2 inst_10313 ( .ZN(net_9376), .A1(net_7858), .A2(net_7847) );
INV_X4 inst_17169 ( .ZN(net_3035), .A(net_85) );
NOR2_X2 inst_3836 ( .ZN(net_12851), .A2(net_9690), .A1(net_1233) );
NAND2_X4 inst_6999 ( .ZN(net_17365), .A1(net_16730), .A2(net_16575) );
INV_X4 inst_13461 ( .ZN(net_11497), .A(net_10237) );
NAND2_X2 inst_8472 ( .A1(net_21146), .A2(net_20514), .ZN(net_20231) );
OAI21_X2 inst_2192 ( .ZN(net_19118), .B2(net_8587), .B1(net_4510), .A(net_278) );
NAND3_X2 inst_5980 ( .ZN(net_14597), .A2(net_14596), .A1(net_13035), .A3(net_10671) );
NAND2_X2 inst_7806 ( .ZN(net_18688), .A1(net_18687), .A2(net_18667) );
CLKBUF_X2 inst_22484 ( .A(net_22355), .Z(net_22356) );
INV_X4 inst_14675 ( .ZN(net_5513), .A(net_4310) );
NOR2_X2 inst_4216 ( .ZN(net_8689), .A1(net_6325), .A2(net_4851) );
XNOR2_X2 inst_106 ( .ZN(net_18526), .A(net_18459), .B(net_17718) );
OAI211_X2 inst_2583 ( .ZN(net_7668), .C1(net_7667), .B(net_7428), .A(net_6018), .C2(net_2853) );
AOI21_X2 inst_20883 ( .A(net_10229), .ZN(net_8267), .B1(net_5302), .B2(net_3599) );
NAND2_X2 inst_10753 ( .ZN(net_13843), .A1(net_11311), .A2(net_5383) );
NOR2_X2 inst_3997 ( .A1(net_9768), .ZN(net_8234), .A2(net_8233) );
NAND2_X2 inst_11344 ( .ZN(net_3659), .A2(net_3658), .A1(net_2590) );
INV_X4 inst_16685 ( .A(net_6131), .ZN(net_1072) );
NAND4_X4 inst_5241 ( .ZN(net_15433), .A1(net_14550), .A2(net_13490), .A4(net_13069), .A3(net_11367) );
NAND2_X2 inst_9903 ( .ZN(net_12163), .A1(net_9360), .A2(net_9341) );
NOR2_X2 inst_4383 ( .ZN(net_6128), .A1(net_5277), .A2(net_5006) );
INV_X4 inst_14507 ( .ZN(net_14314), .A(net_6573) );
NAND2_X2 inst_9208 ( .ZN(net_13055), .A1(net_13054), .A2(net_13053) );
NAND4_X2 inst_5434 ( .ZN(net_13972), .A4(net_12923), .A3(net_11702), .A1(net_11194), .A2(net_10900) );
NAND2_X2 inst_10418 ( .ZN(net_7238), .A1(net_7237), .A2(net_5672) );
NOR2_X2 inst_3756 ( .ZN(net_10371), .A1(net_10370), .A2(net_9407) );
NOR2_X2 inst_4991 ( .A1(net_3836), .ZN(net_3462), .A2(net_3368) );
INV_X4 inst_16939 ( .ZN(net_12004), .A(net_4995) );
INV_X2 inst_18965 ( .A(net_6794), .ZN(net_6115) );
INV_X4 inst_14993 ( .ZN(net_10137), .A(net_3398) );
INV_X4 inst_16997 ( .ZN(net_8361), .A(net_3297) );
NAND2_X2 inst_10811 ( .ZN(net_6828), .A1(net_5845), .A2(net_5526) );
OAI21_X2 inst_1733 ( .B2(net_19908), .B1(net_19907), .ZN(net_15075), .A(net_421) );
NAND2_X2 inst_9489 ( .ZN(net_14330), .A1(net_11443), .A2(net_9417) );
NAND2_X2 inst_8832 ( .A1(net_16037), .ZN(net_15536), .A2(net_15118) );
INV_X4 inst_17139 ( .ZN(net_1321), .A(net_763) );
NAND2_X2 inst_11714 ( .ZN(net_6790), .A2(net_2271), .A1(net_1940) );
NAND2_X2 inst_8911 ( .ZN(net_14971), .A2(net_13745), .A1(net_13194) );
NOR2_X2 inst_3900 ( .A1(net_11526), .ZN(net_9093), .A2(net_5659) );
INV_X4 inst_18059 ( .A(net_20881), .ZN(net_44) );
OAI21_X2 inst_2199 ( .A(net_9039), .ZN(net_8564), .B1(net_8563), .B2(net_5248) );
SDFF_X2 inst_918 ( .Q(net_21139), .D(net_16484), .SE(net_263), .CK(net_21639), .SI(x3667) );
NOR2_X2 inst_4751 ( .A1(net_3842), .ZN(net_3018), .A2(net_2377) );
CLKBUF_X2 inst_22349 ( .A(net_21705), .Z(net_22221) );
NAND3_X2 inst_6588 ( .ZN(net_13849), .A3(net_10139), .A2(net_9541), .A1(net_9466) );
NAND2_X4 inst_7678 ( .ZN(net_1217), .A1(net_1134), .A2(net_699) );
INV_X4 inst_16146 ( .A(net_1825), .ZN(net_1466) );
INV_X4 inst_13921 ( .ZN(net_8659), .A(net_7261) );
NAND2_X2 inst_9177 ( .ZN(net_13341), .A1(net_10714), .A2(net_10453) );
INV_X4 inst_17846 ( .ZN(net_508), .A(net_98) );
NOR2_X2 inst_4035 ( .A1(net_11376), .ZN(net_7940), .A2(net_7939) );
OAI21_X2 inst_1862 ( .ZN(net_13792), .B2(net_11066), .B1(net_8429), .A(net_1125) );
INV_X4 inst_14108 ( .A(net_11285), .ZN(net_6162) );
INV_X4 inst_12928 ( .ZN(net_16867), .A(net_16656) );
INV_X4 inst_15973 ( .ZN(net_13734), .A(net_8889) );
NAND2_X4 inst_7466 ( .ZN(net_4789), .A1(net_2727), .A2(net_225) );
AOI21_X4 inst_20172 ( .B2(net_20144), .B1(net_20143), .ZN(net_15549), .A(net_15468) );
OAI211_X2 inst_2429 ( .ZN(net_15154), .B(net_13930), .C1(net_10810), .A(net_8963), .C2(net_6439) );
INV_X4 inst_15292 ( .ZN(net_6466), .A(net_2716) );
INV_X2 inst_18571 ( .ZN(net_10743), .A(net_10742) );
INV_X4 inst_17027 ( .ZN(net_1568), .A(net_236) );
NAND2_X2 inst_10596 ( .ZN(net_7909), .A1(net_6631), .A2(net_3853) );
NAND2_X2 inst_10463 ( .ZN(net_10609), .A2(net_7008), .A1(net_3356) );
SDFF_X2 inst_754 ( .Q(net_20943), .SE(net_18577), .SI(net_18529), .D(net_8990), .CK(net_22748) );
NAND2_X2 inst_10531 ( .ZN(net_8788), .A1(net_6863), .A2(net_6860) );
NAND2_X2 inst_10030 ( .ZN(net_19917), .A1(net_10683), .A2(net_8735) );
INV_X2 inst_18696 ( .A(net_10604), .ZN(net_8337) );
CLKBUF_X2 inst_22592 ( .A(net_22463), .Z(net_22464) );
INV_X4 inst_18165 ( .A(net_21033), .ZN(net_463) );
NAND2_X2 inst_10332 ( .ZN(net_7595), .A1(net_4471), .A2(net_3479) );
NOR2_X4 inst_2913 ( .ZN(net_9758), .A2(net_6155), .A1(net_2431) );
NAND2_X4 inst_7647 ( .A1(net_20901), .ZN(net_1240), .A2(net_163) );
AOI21_X4 inst_20216 ( .ZN(net_19039), .B1(net_13514), .B2(net_12404), .A(net_10677) );
NAND2_X2 inst_8783 ( .A1(net_16259), .ZN(net_15788), .A2(net_15226) );
NOR2_X4 inst_3295 ( .ZN(net_2331), .A1(net_1261), .A2(net_570) );
AOI21_X2 inst_20926 ( .ZN(net_7123), .A(net_7122), .B1(net_7121), .B2(net_2567) );
NAND2_X2 inst_8792 ( .A1(net_19915), .ZN(net_18940), .A2(net_15744) );
NOR2_X2 inst_5057 ( .ZN(net_10569), .A1(net_1021), .A2(net_1020) );
INV_X4 inst_16368 ( .ZN(net_14709), .A(net_60) );
CLKBUF_X2 inst_21606 ( .A(net_21477), .Z(net_21478) );
NAND2_X2 inst_8828 ( .A1(net_15690), .ZN(net_15539), .A2(net_14771) );
CLKBUF_X2 inst_21814 ( .A(net_21274), .Z(net_21686) );
NAND2_X4 inst_7394 ( .A2(net_20875), .A1(net_19861), .ZN(net_12409) );
INV_X4 inst_13997 ( .ZN(net_7404), .A(net_6395) );
INV_X4 inst_13140 ( .ZN(net_15084), .A(net_14688) );
INV_X4 inst_12998 ( .ZN(net_17115), .A(net_16799) );
INV_X4 inst_16383 ( .ZN(net_6905), .A(net_5766) );
NOR2_X4 inst_2923 ( .ZN(net_9446), .A2(net_7906), .A1(net_761) );
NAND2_X2 inst_7957 ( .ZN(net_18392), .A1(net_18355), .A2(net_18251) );
NOR3_X2 inst_2707 ( .ZN(net_20635), .A3(net_13904), .A1(net_11942), .A2(net_8295) );
NOR2_X2 inst_3958 ( .ZN(net_19818), .A1(net_6707), .A2(net_6486) );
AND4_X2 inst_21109 ( .A1(net_13156), .A3(net_11744), .ZN(net_11726), .A2(net_11725), .A4(net_11724) );
CLKBUF_X2 inst_22366 ( .A(net_22237), .Z(net_22238) );
AOI21_X2 inst_20567 ( .ZN(net_14207), .B2(net_12400), .A(net_12113), .B1(net_11407) );
INV_X4 inst_17543 ( .ZN(net_17277), .A(net_375) );
NAND2_X2 inst_10465 ( .ZN(net_7005), .A1(net_7004), .A2(net_4258) );
NAND2_X2 inst_10166 ( .ZN(net_9723), .A2(net_8241), .A1(net_8131) );
NOR2_X2 inst_4620 ( .ZN(net_3620), .A2(net_3391), .A1(net_1407) );
INV_X4 inst_12674 ( .ZN(net_17741), .A(net_17740) );
INV_X4 inst_15719 ( .ZN(net_3591), .A(net_2797) );
NAND2_X2 inst_9277 ( .A1(net_13023), .ZN(net_12595), .A2(net_10913) );
NOR2_X2 inst_3707 ( .ZN(net_11058), .A2(net_11057), .A1(net_7636) );
NAND2_X2 inst_11869 ( .ZN(net_1642), .A2(net_1224), .A1(net_691) );
INV_X4 inst_14243 ( .ZN(net_5779), .A(net_5778) );
CLKBUF_X2 inst_22509 ( .A(net_22380), .Z(net_22381) );
CLKBUF_X2 inst_22056 ( .A(net_21927), .Z(net_21928) );
INV_X8 inst_12431 ( .A(net_19459), .ZN(net_19455) );
NAND2_X2 inst_10158 ( .ZN(net_8262), .A1(net_8261), .A2(net_8095) );
NAND2_X2 inst_8131 ( .ZN(net_18042), .A2(net_18030), .A1(net_18023) );
AND2_X2 inst_21370 ( .A1(net_20495), .A2(net_1271), .ZN(net_438) );
INV_X4 inst_14767 ( .ZN(net_7018), .A(net_5483) );
NAND4_X2 inst_5388 ( .ZN(net_19545), .A2(net_13476), .A4(net_9992), .A1(net_9831), .A3(net_9216) );
INV_X2 inst_19436 ( .A(net_3451), .ZN(net_1731) );
NOR2_X2 inst_4492 ( .ZN(net_7351), .A2(net_4355), .A1(net_4299) );
INV_X4 inst_13551 ( .ZN(net_9166), .A(net_9165) );
NAND2_X2 inst_9773 ( .ZN(net_11647), .A2(net_9793), .A1(net_7850) );
INV_X4 inst_14553 ( .ZN(net_18903), .A(net_4590) );
NOR2_X4 inst_3056 ( .A1(net_20825), .ZN(net_7937), .A2(net_1163) );
INV_X4 inst_14550 ( .ZN(net_6205), .A(net_4592) );
INV_X8 inst_12214 ( .ZN(net_9540), .A(net_5059) );
CLKBUF_X2 inst_21616 ( .A(net_21487), .Z(net_21488) );
CLKBUF_X2 inst_22837 ( .A(net_22708), .Z(net_22709) );
NOR3_X4 inst_2609 ( .A3(net_18983), .A1(net_18982), .ZN(net_16133), .A2(net_15503) );
CLKBUF_X2 inst_22818 ( .A(net_21506), .Z(net_22690) );
OAI211_X2 inst_2556 ( .C1(net_13495), .A(net_11293), .ZN(net_9952), .B(net_9951), .C2(net_2872) );
INV_X2 inst_19716 ( .A(net_20773), .ZN(net_20770) );
INV_X4 inst_15022 ( .A(net_6548), .ZN(net_3375) );
NAND4_X2 inst_5371 ( .ZN(net_15233), .A4(net_14031), .A3(net_11773), .A2(net_11490), .A1(net_9783) );
OAI21_X2 inst_1704 ( .ZN(net_15287), .A(net_15046), .B2(net_13563), .B1(net_11187) );
NOR2_X2 inst_4604 ( .ZN(net_11207), .A1(net_3750), .A2(net_3749) );
INV_X2 inst_19459 ( .A(net_2076), .ZN(net_1912) );
INV_X4 inst_15156 ( .ZN(net_3486), .A(net_3055) );
INV_X4 inst_15766 ( .ZN(net_3766), .A(net_1416) );
XNOR2_X2 inst_161 ( .B(net_20462), .ZN(net_17935), .A(net_17800) );
CLKBUF_X2 inst_22832 ( .A(net_22703), .Z(net_22704) );
NAND2_X2 inst_10956 ( .A1(net_10105), .A2(net_5373), .ZN(net_5084) );
NAND3_X2 inst_6118 ( .A2(net_14669), .ZN(net_13863), .A3(net_13862), .A1(net_8692) );
NAND2_X2 inst_11287 ( .ZN(net_6646), .A1(net_4093), .A2(net_2763) );
NAND2_X2 inst_9624 ( .ZN(net_10665), .A1(net_10664), .A2(net_7366) );
NAND2_X2 inst_11764 ( .ZN(net_4024), .A1(net_2828), .A2(net_2066) );
INV_X4 inst_17389 ( .ZN(net_1259), .A(net_146) );
OAI211_X2 inst_2408 ( .B(net_20838), .A(net_20837), .C1(net_19227), .ZN(net_15533), .C2(net_14759) );
NAND2_X2 inst_10519 ( .A1(net_9339), .ZN(net_6873), .A2(net_6781) );
CLKBUF_X2 inst_21503 ( .A(net_21374), .Z(net_21375) );
NAND2_X2 inst_9778 ( .ZN(net_20813), .A1(net_15573), .A2(net_6271) );
OAI222_X2 inst_1324 ( .ZN(net_11919), .A2(net_11918), .C1(net_10514), .A1(net_10490), .C2(net_7094), .B1(net_6524), .B2(net_2052) );
INV_X4 inst_15585 ( .ZN(net_2837), .A(net_2265) );
AOI21_X2 inst_20822 ( .ZN(net_9990), .A(net_9989), .B1(net_9988), .B2(net_5691) );
NAND2_X2 inst_11848 ( .ZN(net_1950), .A1(net_1584), .A2(net_754) );
NAND2_X2 inst_10646 ( .ZN(net_11708), .A1(net_6611), .A2(net_6369) );
XNOR2_X2 inst_342 ( .B(net_20708), .ZN(net_17119), .A(net_16451) );
XNOR2_X2 inst_463 ( .ZN(net_13285), .A(net_13284), .B(net_8994) );
CLKBUF_X2 inst_22914 ( .A(net_21584), .Z(net_22786) );
CLKBUF_X2 inst_22014 ( .A(net_21885), .Z(net_21886) );
NAND2_X2 inst_10667 ( .ZN(net_6266), .A1(net_6265), .A2(net_6264) );
INV_X2 inst_18648 ( .ZN(net_9231), .A(net_9230) );
INV_X4 inst_13571 ( .ZN(net_9130), .A(net_9129) );
NOR2_X2 inst_3820 ( .ZN(net_19091), .A1(net_10031), .A2(net_9795) );
NOR2_X2 inst_4667 ( .ZN(net_4356), .A1(net_3138), .A2(net_703) );
CLKBUF_X2 inst_22457 ( .A(net_22328), .Z(net_22329) );
INV_X4 inst_12762 ( .ZN(net_17387), .A(net_17386) );
NAND2_X4 inst_6992 ( .ZN(net_17215), .A1(net_16720), .A2(net_16559) );
NAND3_X2 inst_5923 ( .ZN(net_19827), .A1(net_14057), .A3(net_12735), .A2(net_7384) );
INV_X4 inst_15857 ( .A(net_6840), .ZN(net_1916) );
OAI21_X2 inst_2158 ( .ZN(net_19811), .A(net_7396), .B1(net_4601), .B2(net_3914) );
INV_X4 inst_15702 ( .A(net_2739), .ZN(net_2004) );
NAND3_X4 inst_5560 ( .ZN(net_19470), .A2(net_15447), .A3(net_15247), .A1(net_14592) );
OAI21_X2 inst_1711 ( .A(net_15876), .ZN(net_15196), .B1(net_14056), .B2(net_10755) );
NAND2_X2 inst_10660 ( .ZN(net_7637), .A2(net_3621), .A1(net_1182) );
NOR2_X2 inst_3426 ( .ZN(net_15429), .A2(net_14978), .A1(net_7285) );
INV_X4 inst_16063 ( .ZN(net_2444), .A(net_2291) );
INV_X4 inst_16118 ( .ZN(net_1901), .A(net_1492) );
OAI21_X2 inst_2052 ( .B1(net_10976), .A(net_10975), .ZN(net_10845), .B2(net_10844) );
SDFF_X2 inst_995 ( .QN(net_20999), .D(net_2132), .SE(net_263), .CK(net_21840), .SI(x3052) );
NAND2_X2 inst_8850 ( .ZN(net_15388), .A2(net_14559), .A1(net_11672) );
NAND2_X2 inst_7726 ( .ZN(net_18830), .A2(net_18786), .A1(net_17703) );
INV_X4 inst_13948 ( .ZN(net_6769), .A(net_6768) );
NAND2_X2 inst_10697 ( .A1(net_6840), .ZN(net_6069), .A2(net_4586) );
OAI211_X2 inst_2470 ( .C2(net_20781), .ZN(net_13850), .B(net_13849), .C1(net_13848), .A(net_12802) );
NAND3_X2 inst_6049 ( .ZN(net_14245), .A3(net_13562), .A2(net_12483), .A1(net_6361) );
CLKBUF_X2 inst_22216 ( .A(net_22087), .Z(net_22088) );
NOR2_X2 inst_3857 ( .A2(net_9472), .ZN(net_9471), .A1(net_7470) );
INV_X2 inst_18384 ( .A(net_16901), .ZN(net_16696) );
OR3_X2 inst_1060 ( .A3(net_13206), .ZN(net_8970), .A1(net_8969), .A2(net_277) );
NAND3_X2 inst_5920 ( .ZN(net_20105), .A3(net_12840), .A2(net_11257), .A1(net_8860) );
SDFF_X2 inst_900 ( .Q(net_21150), .D(net_16771), .SE(net_253), .CK(net_22215), .SI(x5685) );
NAND2_X4 inst_6950 ( .A2(net_20051), .A1(net_20050), .ZN(net_17529) );
NAND2_X2 inst_10568 ( .A1(net_7298), .ZN(net_6708), .A2(net_6707) );
INV_X4 inst_18172 ( .A(net_20989), .ZN(net_1867) );
INV_X4 inst_18123 ( .A(net_21029), .ZN(net_853) );
INV_X4 inst_14511 ( .ZN(net_4819), .A(net_4818) );
NOR2_X2 inst_4949 ( .A1(net_20530), .ZN(net_8389), .A2(net_1664) );
INV_X2 inst_18835 ( .ZN(net_6759), .A(net_6758) );
INV_X2 inst_19104 ( .ZN(net_7530), .A(net_4498) );
INV_X4 inst_12677 ( .ZN(net_20129), .A(net_17734) );
NOR2_X4 inst_2807 ( .A2(net_20317), .A1(net_20316), .ZN(net_17912) );
INV_X4 inst_13608 ( .ZN(net_8791), .A(net_8573) );
NAND4_X2 inst_5327 ( .A4(net_19173), .A1(net_19172), .ZN(net_15653), .A2(net_12447), .A3(net_10255) );
NAND4_X2 inst_5423 ( .ZN(net_14208), .A2(net_13497), .A1(net_12351), .A4(net_12260), .A3(net_7107) );
NAND2_X2 inst_9995 ( .ZN(net_8838), .A2(net_8837), .A1(net_8618) );
NAND2_X2 inst_8803 ( .ZN(net_19496), .A2(net_15348), .A1(net_14265) );
CLKBUF_X2 inst_22880 ( .A(net_22024), .Z(net_22752) );
NAND2_X2 inst_8651 ( .A2(net_20068), .ZN(net_16559), .A1(net_16520) );
AOI21_X2 inst_20866 ( .B1(net_19332), .ZN(net_8600), .B2(net_6484), .A(net_57) );
INV_X4 inst_15948 ( .ZN(net_11087), .A(net_4694) );
INV_X2 inst_18683 ( .A(net_14537), .ZN(net_8756) );
NAND2_X2 inst_10470 ( .ZN(net_8356), .A1(net_6996), .A2(net_4737) );
NAND2_X2 inst_7882 ( .ZN(net_18519), .A1(net_18457), .A2(net_18407) );
NAND2_X2 inst_11617 ( .A2(net_9310), .ZN(net_6478), .A1(net_2581) );
AOI21_X2 inst_20373 ( .ZN(net_15605), .B1(net_15375), .B2(net_14263), .A(net_5262) );
NAND2_X1 inst_12161 ( .A1(net_2590), .A2(net_2192), .ZN(net_1408) );
NAND3_X2 inst_6767 ( .ZN(net_5303), .A3(net_5302), .A1(net_3160), .A2(net_1580) );
CLKBUF_X2 inst_21497 ( .A(net_21253), .Z(net_21369) );
INV_X2 inst_19287 ( .ZN(net_4393), .A(net_4022) );
NAND2_X2 inst_8084 ( .A2(net_20505), .ZN(net_18145), .A1(net_17137) );
OR2_X2 inst_1225 ( .ZN(net_3815), .A2(net_1686), .A1(net_170) );
INV_X2 inst_19029 ( .A(net_6740), .ZN(net_4904) );
CLKBUF_X2 inst_22006 ( .A(net_21877), .Z(net_21878) );
NAND2_X4 inst_7535 ( .A2(net_19661), .A1(net_19660), .ZN(net_1952) );
INV_X8 inst_12411 ( .A(net_20907), .ZN(net_896) );
INV_X4 inst_14256 ( .A(net_10608), .ZN(net_8837) );
NAND4_X2 inst_5316 ( .ZN(net_15777), .A4(net_15053), .A2(net_13994), .A1(net_11583), .A3(net_8314) );
INV_X2 inst_19686 ( .ZN(net_20530), .A(net_20529) );
NAND3_X4 inst_5530 ( .A3(net_19531), .A1(net_19530), .ZN(net_17775), .A2(net_16036) );
INV_X4 inst_14427 ( .A(net_6705), .ZN(net_6178) );
INV_X4 inst_14215 ( .ZN(net_5879), .A(net_5878) );
NOR2_X2 inst_4551 ( .ZN(net_4992), .A2(net_3963), .A1(net_809) );
NAND2_X2 inst_11397 ( .ZN(net_5460), .A2(net_3472), .A1(net_2697) );
NOR2_X2 inst_4313 ( .ZN(net_7409), .A2(net_6893), .A1(net_6610) );
INV_X4 inst_13153 ( .ZN(net_14880), .A(net_14343) );
NOR2_X2 inst_4714 ( .A2(net_7745), .A1(net_5153), .ZN(net_4094) );
INV_X4 inst_12898 ( .ZN(net_17007), .A(net_16786) );
INV_X4 inst_16114 ( .ZN(net_12440), .A(net_8138) );
CLKBUF_X2 inst_22101 ( .A(net_21972), .Z(net_21973) );
NOR2_X4 inst_2956 ( .ZN(net_8706), .A1(net_5175), .A2(net_955) );
NOR2_X2 inst_4713 ( .A2(net_5845), .ZN(net_4116), .A1(net_3146) );
INV_X4 inst_16071 ( .ZN(net_8184), .A(net_1566) );
XNOR2_X2 inst_412 ( .B(net_21150), .A(net_16619), .ZN(net_16618) );
NAND4_X2 inst_5463 ( .ZN(net_13325), .A1(net_13324), .A2(net_13323), .A4(net_13322), .A3(net_7644) );
INV_X4 inst_14721 ( .ZN(net_4161), .A(net_3962) );
INV_X2 inst_19693 ( .A(net_20547), .ZN(net_20546) );
INV_X4 inst_13022 ( .A(net_16619), .ZN(net_16605) );
NAND2_X2 inst_8295 ( .A1(net_20318), .ZN(net_19919), .A2(net_17194) );
INV_X4 inst_13969 ( .A(net_10442), .ZN(net_8604) );
INV_X2 inst_19358 ( .ZN(net_2347), .A(net_2346) );
NOR2_X4 inst_3163 ( .ZN(net_5629), .A1(net_3196), .A2(net_2539) );
INV_X2 inst_19228 ( .A(net_16125), .ZN(net_3390) );
OAI211_X2 inst_2504 ( .ZN(net_12775), .B(net_12774), .C2(net_12091), .A(net_5235), .C1(net_60) );
INV_X4 inst_17132 ( .ZN(net_6081), .A(net_925) );
INV_X4 inst_13511 ( .ZN(net_13010), .A(net_9405) );
INV_X4 inst_14076 ( .A(net_6224), .ZN(net_6223) );
INV_X4 inst_14824 ( .ZN(net_5780), .A(net_4387) );
INV_X4 inst_15469 ( .ZN(net_15628), .A(net_14687) );
NOR2_X2 inst_3374 ( .ZN(net_16498), .A2(net_16497), .A1(net_552) );
NOR2_X2 inst_4354 ( .ZN(net_5962), .A2(net_5614), .A1(net_4288) );
INV_X4 inst_18049 ( .A(net_21143), .ZN(net_430) );
NOR2_X2 inst_3438 ( .A1(net_16076), .ZN(net_15251), .A2(net_14732) );
INV_X4 inst_12541 ( .ZN(net_18352), .A(net_18351) );
INV_X4 inst_14614 ( .ZN(net_7443), .A(net_4204) );
INV_X2 inst_18781 ( .ZN(net_7515), .A(net_7514) );
NOR2_X2 inst_3811 ( .ZN(net_19089), .A2(net_10089), .A1(net_7033) );
NOR2_X2 inst_3653 ( .ZN(net_11668), .A2(net_11667), .A1(net_9609) );
CLKBUF_X2 inst_22184 ( .A(net_22055), .Z(net_22056) );
INV_X2 inst_18694 ( .A(net_11659), .ZN(net_8358) );
NAND2_X4 inst_6959 ( .ZN(net_17952), .A2(net_17102), .A1(net_16944) );
CLKBUF_X2 inst_21877 ( .A(net_21748), .Z(net_21749) );
INV_X4 inst_15652 ( .ZN(net_8537), .A(net_2111) );
NAND2_X2 inst_8213 ( .ZN(net_17847), .A1(net_17782), .A2(net_17594) );
NAND2_X2 inst_10700 ( .ZN(net_6043), .A2(net_6042), .A1(net_5506) );
INV_X4 inst_16187 ( .ZN(net_7659), .A(net_3187) );
INV_X4 inst_15438 ( .ZN(net_3105), .A(net_2502) );
OR2_X2 inst_1241 ( .A1(net_790), .ZN(net_499), .A2(net_104) );
SDFF_X2 inst_1038 ( .QN(net_20989), .SE(net_17277), .D(net_1867), .CK(net_22651), .SI(x3178) );
INV_X4 inst_15418 ( .ZN(net_4581), .A(net_2779) );
SDFF_X2 inst_940 ( .QN(net_21015), .D(net_536), .SE(net_263), .CK(net_22679), .SI(x2784) );
AND2_X4 inst_21193 ( .ZN(net_20013), .A1(net_14782), .A2(net_7247) );
INV_X2 inst_19307 ( .ZN(net_5614), .A(net_2728) );
NAND2_X2 inst_9417 ( .ZN(net_14359), .A2(net_9796), .A1(net_9681) );
NAND2_X2 inst_11705 ( .A1(net_3919), .ZN(net_2582), .A2(net_1878) );
NAND2_X2 inst_11641 ( .A1(net_3542), .ZN(net_3279), .A2(net_1422) );
NOR2_X2 inst_3595 ( .A1(net_14055), .A2(net_13644), .ZN(net_12599) );
NAND2_X2 inst_11830 ( .ZN(net_3030), .A2(net_1331), .A1(net_61) );
NOR2_X2 inst_4876 ( .ZN(net_2203), .A2(net_2202), .A1(net_1018) );
NAND2_X2 inst_8103 ( .ZN(net_18117), .A2(net_18094), .A1(net_16815) );
NAND2_X2 inst_7732 ( .ZN(net_18817), .A2(net_18787), .A1(net_17729) );
NAND2_X2 inst_9008 ( .ZN(net_14271), .A2(net_14270), .A1(net_10637) );
NOR2_X2 inst_4362 ( .ZN(net_6844), .A1(net_5537), .A2(net_3981) );
NAND2_X2 inst_9581 ( .ZN(net_12605), .A1(net_7610), .A2(net_7605) );
INV_X4 inst_15761 ( .ZN(net_4230), .A(net_1417) );
INV_X4 inst_12608 ( .ZN(net_18081), .A(net_18080) );
NOR2_X2 inst_4369 ( .ZN(net_5489), .A2(net_5488), .A1(net_3690) );
INV_X4 inst_17869 ( .ZN(net_798), .A(net_95) );
NAND2_X2 inst_11899 ( .A2(net_9309), .ZN(net_1579), .A1(net_913) );
CLKBUF_X2 inst_22357 ( .A(net_21568), .Z(net_22229) );
NAND2_X2 inst_11236 ( .A1(net_20482), .ZN(net_3942), .A2(net_3941) );
INV_X4 inst_13076 ( .ZN(net_16223), .A(net_16164) );
NOR2_X2 inst_4007 ( .ZN(net_11754), .A1(net_10447), .A2(net_8095) );
SDFF_X2 inst_879 ( .Q(net_21231), .SI(net_16886), .SE(net_125), .CK(net_21452), .D(x6966) );
INV_X4 inst_17325 ( .ZN(net_4163), .A(net_572) );
INV_X4 inst_17105 ( .ZN(net_9191), .A(net_333) );
NOR2_X2 inst_4291 ( .ZN(net_11365), .A1(net_6034), .A2(net_3703) );
NAND3_X2 inst_5692 ( .ZN(net_16270), .A2(net_15977), .A3(net_15838), .A1(net_5377) );
INV_X4 inst_17603 ( .ZN(net_1471), .A(net_320) );
XNOR2_X2 inst_629 ( .B(net_17422), .ZN(net_453), .A(net_452) );
NOR2_X2 inst_4903 ( .ZN(net_1976), .A2(net_1205), .A1(net_1142) );
OR2_X4 inst_1100 ( .ZN(net_7074), .A1(net_3867), .A2(net_2986) );
NAND2_X2 inst_10872 ( .A2(net_5526), .ZN(net_5429), .A1(net_143) );
INV_X4 inst_18037 ( .A(net_20962), .ZN(net_824) );
INV_X4 inst_15105 ( .ZN(net_6801), .A(net_4229) );
INV_X2 inst_18372 ( .ZN(net_17369), .A(net_17240) );
NOR2_X2 inst_3383 ( .ZN(net_16367), .A2(net_16218), .A1(net_15679) );
AOI221_X2 inst_20091 ( .ZN(net_15235), .B1(net_14734), .C1(net_14600), .B2(net_13875), .C2(net_13227), .A(net_9044) );
INV_X4 inst_15682 ( .ZN(net_3249), .A(net_2039) );
OR2_X2 inst_1191 ( .ZN(net_19710), .A1(net_11045), .A2(net_10635) );
INV_X4 inst_18307 ( .A(net_20495), .ZN(net_20493) );
XNOR2_X2 inst_533 ( .ZN(net_1897), .A(net_1896), .B(net_1895) );
OAI211_X2 inst_2478 ( .ZN(net_13506), .C1(net_11441), .C2(net_10730), .B(net_6065), .A(net_5035) );
NOR2_X2 inst_4972 ( .ZN(net_2973), .A1(net_2204), .A2(net_1349) );
NOR3_X2 inst_2751 ( .ZN(net_12087), .A3(net_11813), .A1(net_9827), .A2(net_7524) );
AOI21_X2 inst_20694 ( .ZN(net_12181), .A(net_10323), .B1(net_8272), .B2(net_6685) );
INV_X4 inst_16928 ( .ZN(net_1640), .A(net_932) );
OAI21_X2 inst_1760 ( .ZN(net_14723), .A(net_14657), .B2(net_11963), .B1(net_5622) );
OAI21_X2 inst_1874 ( .B1(net_15374), .ZN(net_13698), .B2(net_13697), .A(net_12618) );
OAI21_X2 inst_2022 ( .ZN(net_11330), .A(net_10105), .B2(net_9793), .B1(net_3949) );
AOI21_X2 inst_20646 ( .ZN(net_13142), .B2(net_9535), .B1(net_2920), .A(net_968) );
NOR2_X2 inst_3960 ( .ZN(net_20226), .A1(net_6740), .A2(net_6475) );
NOR2_X4 inst_2821 ( .ZN(net_16292), .A1(net_16114), .A2(net_16045) );
OR2_X4 inst_1095 ( .ZN(net_8480), .A2(net_8446), .A1(net_4711) );
NAND2_X2 inst_8042 ( .ZN(net_18238), .A1(net_18237), .A2(net_18222) );
INV_X4 inst_16738 ( .ZN(net_12522), .A(net_9994) );
NAND2_X2 inst_10516 ( .ZN(net_10406), .A1(net_8330), .A2(net_4999) );
NAND2_X2 inst_10096 ( .ZN(net_13176), .A1(net_10022), .A2(net_7876) );
NAND2_X2 inst_9052 ( .ZN(net_20330), .A2(net_11957), .A1(net_8596) );
OAI211_X2 inst_2439 ( .ZN(net_14868), .A(net_14867), .B(net_14866), .C1(net_14865), .C2(net_11959) );
XNOR2_X2 inst_176 ( .ZN(net_17779), .A(net_17551), .B(net_201) );
NOR2_X4 inst_2826 ( .A2(net_20426), .A1(net_20425), .ZN(net_19290) );
NAND2_X2 inst_9069 ( .ZN(net_13978), .A2(net_12200), .A1(net_8577) );
NAND2_X2 inst_10894 ( .A1(net_20571), .ZN(net_5399), .A2(net_3731) );
AOI22_X2 inst_20027 ( .A1(net_11472), .ZN(net_9928), .A2(net_8204), .B1(net_7867), .B2(net_3442) );
OAI221_X2 inst_1336 ( .ZN(net_15175), .C1(net_15174), .B1(net_15174), .A(net_14311), .B2(net_9828), .C2(net_7730) );
NAND4_X2 inst_5472 ( .ZN(net_13204), .A1(net_13203), .A2(net_10315), .A4(net_7734), .A3(net_4248) );
NAND2_X2 inst_10387 ( .A1(net_10141), .ZN(net_8913), .A2(net_7321) );
OAI21_X2 inst_1665 ( .B1(net_20142), .ZN(net_18982), .B2(net_15753), .A(net_13836) );
NOR2_X2 inst_4500 ( .ZN(net_4255), .A2(net_3051), .A1(net_1813) );
INV_X4 inst_13962 ( .ZN(net_6724), .A(net_6723) );
NOR2_X2 inst_4763 ( .ZN(net_3895), .A2(net_3095), .A1(net_955) );
INV_X4 inst_17224 ( .A(net_3297), .ZN(net_749) );
SDFF_X2 inst_780 ( .Q(net_20935), .SE(net_18576), .SI(net_18341), .D(net_486), .CK(net_21424) );
NAND3_X4 inst_5626 ( .ZN(net_7757), .A2(net_5208), .A3(net_4535), .A1(net_2900) );
NAND3_X2 inst_6783 ( .A1(net_6402), .ZN(net_4233), .A2(net_3172), .A3(net_2561) );
NAND2_X2 inst_8255 ( .A2(net_17851), .ZN(net_17700), .A1(net_17699) );
NAND2_X2 inst_12016 ( .ZN(net_2369), .A2(net_937), .A1(net_741) );
NOR2_X2 inst_3967 ( .ZN(net_8417), .A1(net_8416), .A2(net_8415) );
INV_X2 inst_19099 ( .ZN(net_4539), .A(net_4538) );
INV_X4 inst_16769 ( .ZN(net_13514), .A(net_1028) );
NAND2_X2 inst_8722 ( .A1(net_21228), .ZN(net_16149), .A2(net_15894) );
NOR2_X2 inst_3669 ( .ZN(net_12631), .A2(net_11528), .A1(net_60) );
OAI21_X2 inst_1767 ( .ZN(net_14701), .A(net_14700), .B2(net_12060), .B1(net_9825) );
CLKBUF_X2 inst_22145 ( .A(net_22016), .Z(net_22017) );
CLKBUF_X2 inst_21727 ( .A(net_21598), .Z(net_21599) );
INV_X4 inst_13564 ( .ZN(net_9141), .A(net_9140) );
INV_X4 inst_16087 ( .A(net_1703), .ZN(net_1531) );
OAI21_X1 inst_2361 ( .ZN(net_12543), .A(net_12542), .B1(net_11067), .B2(net_5804) );
CLKBUF_X2 inst_22140 ( .A(net_21526), .Z(net_22012) );
NAND2_X2 inst_11497 ( .ZN(net_7099), .A2(net_3402), .A1(net_2500) );
NAND2_X2 inst_10237 ( .ZN(net_8040), .A1(net_8039), .A2(net_6978) );
NAND3_X2 inst_6006 ( .ZN(net_14424), .A3(net_12453), .A1(net_10887), .A2(net_2661) );
INV_X4 inst_14652 ( .ZN(net_5719), .A(net_4369) );
AOI21_X2 inst_20691 ( .ZN(net_19034), .B1(net_12137), .B2(net_8387), .A(net_7116) );
NAND3_X2 inst_6802 ( .A3(net_19418), .ZN(net_13920), .A2(net_4481), .A1(net_761) );
INV_X4 inst_16797 ( .ZN(net_10091), .A(net_1007) );
SDFF_X2 inst_694 ( .Q(net_20955), .SE(net_18856), .SI(net_18854), .D(net_614), .CK(net_21502) );
INV_X4 inst_17025 ( .ZN(net_11442), .A(net_3729) );
INV_X4 inst_15689 ( .ZN(net_4029), .A(net_2026) );
NAND3_X4 inst_5574 ( .ZN(net_19874), .A3(net_14768), .A1(net_12878), .A2(net_4165) );
NAND3_X2 inst_6382 ( .ZN(net_12024), .A3(net_11807), .A2(net_9137), .A1(net_6888) );
CLKBUF_X2 inst_22515 ( .A(net_22225), .Z(net_22387) );
OAI211_X2 inst_2498 ( .ZN(net_12865), .C1(net_12864), .B(net_11642), .A(net_6808), .C2(net_4653) );
INV_X4 inst_17274 ( .ZN(net_1007), .A(net_70) );
INV_X8 inst_12402 ( .ZN(net_223), .A(net_83) );
NOR2_X4 inst_3154 ( .A1(net_20544), .ZN(net_4054), .A2(net_1230) );
AOI21_X2 inst_20480 ( .B1(net_20204), .ZN(net_14906), .A(net_11540), .B2(net_1244) );
NAND4_X2 inst_5396 ( .ZN(net_19912), .A2(net_19737), .A1(net_19736), .A4(net_10117), .A3(net_8124) );
NAND2_X2 inst_9394 ( .ZN(net_11706), .A2(net_11705), .A1(net_9829) );
INV_X4 inst_15531 ( .A(net_3351), .ZN(net_2376) );
AOI21_X2 inst_20688 ( .B1(net_13709), .ZN(net_12224), .B2(net_7265), .A(net_6559) );
NAND2_X2 inst_7814 ( .ZN(net_18671), .A2(net_18670), .A1(net_16874) );
INV_X4 inst_17390 ( .ZN(net_529), .A(net_167) );
INV_X4 inst_16767 ( .ZN(net_15217), .A(net_14720) );
INV_X4 inst_16271 ( .ZN(net_7912), .A(net_5727) );
NAND2_X2 inst_12071 ( .A1(net_3745), .ZN(net_1325), .A2(net_168) );
SDFF_X2 inst_787 ( .Q(net_20948), .SE(net_18584), .SI(net_18037), .D(net_666), .CK(net_21277) );
NOR2_X2 inst_4396 ( .ZN(net_20060), .A1(net_5479), .A2(net_5193) );
NAND2_X2 inst_11211 ( .ZN(net_5069), .A2(net_4157), .A1(net_2274) );
INV_X4 inst_12958 ( .ZN(net_16684), .A(net_16537) );
INV_X4 inst_18214 ( .A(net_20977), .ZN(net_1843) );
INV_X4 inst_15541 ( .A(net_11443), .ZN(net_9636) );
INV_X4 inst_14439 ( .A(net_6683), .ZN(net_6278) );
SDFF_X2 inst_825 ( .Q(net_21237), .SI(net_17574), .SE(net_125), .CK(net_21564), .D(x6764) );
OAI211_X2 inst_2586 ( .ZN(net_6483), .C2(net_6482), .B(net_5317), .A(net_3167), .C1(net_1203) );
NAND2_X2 inst_7928 ( .ZN(net_18443), .A1(net_18356), .A2(net_18204) );
INV_X4 inst_17684 ( .ZN(net_10676), .A(net_232) );
INV_X2 inst_19661 ( .ZN(net_20444), .A(net_20443) );
INV_X4 inst_15310 ( .ZN(net_2656), .A(net_2655) );
INV_X4 inst_12886 ( .ZN(net_17162), .A(net_17031) );
OAI21_X2 inst_1892 ( .ZN(net_13391), .A(net_12179), .B2(net_8816), .B1(net_2392) );
NAND2_X2 inst_7860 ( .ZN(net_18564), .A1(net_18544), .A2(net_18516) );
NAND2_X2 inst_11404 ( .ZN(net_3454), .A2(net_2285), .A1(net_772) );
SDFF_X2 inst_726 ( .Q(net_20973), .SE(net_18585), .SI(net_18569), .D(net_8998), .CK(net_21923) );
DFF_X1 inst_19913 ( .D(net_16834), .CK(net_21576), .Q(x592) );
INV_X4 inst_18112 ( .A(net_20913), .ZN(net_816) );
INV_X2 inst_18436 ( .ZN(net_14341), .A(net_13863) );
NAND2_X2 inst_10583 ( .A1(net_6861), .ZN(net_6673), .A2(net_6672) );
DFF_X1 inst_19851 ( .D(net_17219), .CK(net_22372), .Q(x887) );
INV_X2 inst_18988 ( .A(net_6960), .ZN(net_5110) );
NOR2_X2 inst_4726 ( .A2(net_4865), .ZN(net_4013), .A1(net_3138) );
NAND2_X2 inst_8073 ( .ZN(net_18163), .A2(net_18162), .A1(net_17458) );
CLKBUF_X2 inst_22068 ( .A(net_21939), .Z(net_21940) );
CLKBUF_X2 inst_21738 ( .A(net_21609), .Z(net_21610) );
INV_X2 inst_18623 ( .ZN(net_9566), .A(net_9565) );
XNOR2_X2 inst_320 ( .ZN(net_17041), .A(net_17040), .B(net_13947) );
INV_X4 inst_16861 ( .ZN(net_1752), .A(net_962) );
XOR2_X2 inst_1 ( .A(net_21194), .Z(net_18195), .B(net_18158) );
INV_X4 inst_16327 ( .ZN(net_2950), .A(net_1095) );
OAI21_X2 inst_1891 ( .ZN(net_19167), .B2(net_8755), .B1(net_8423), .A(net_3828) );
CLKBUF_X2 inst_22234 ( .A(net_21778), .Z(net_22106) );
INV_X4 inst_12794 ( .A(net_17894), .ZN(net_17845) );
AOI22_X2 inst_20051 ( .A1(net_8007), .ZN(net_3705), .B1(net_3704), .B2(net_3703), .A2(net_2384) );
NOR2_X2 inst_4558 ( .A1(net_5677), .ZN(net_3926), .A2(net_2883) );
INV_X4 inst_14862 ( .ZN(net_7256), .A(net_3765) );
INV_X4 inst_14525 ( .ZN(net_11781), .A(net_10580) );
INV_X2 inst_19175 ( .ZN(net_3807), .A(net_3806) );
INV_X4 inst_17411 ( .ZN(net_19583), .A(net_493) );
NOR2_X4 inst_3063 ( .ZN(net_6080), .A2(net_4934), .A1(net_3322) );
INV_X4 inst_13881 ( .ZN(net_7356), .A(net_7355) );
INV_X4 inst_17770 ( .ZN(net_4770), .A(net_226) );
INV_X4 inst_17691 ( .ZN(net_958), .A(net_223) );
OAI21_X2 inst_1812 ( .ZN(net_14181), .A(net_12306), .B1(net_10682), .B2(net_6124) );
DFF_X2 inst_19769 ( .QN(net_20875), .D(net_18597), .CK(net_21936) );
NAND2_X4 inst_7608 ( .ZN(net_2650), .A2(net_1669), .A1(net_1384) );
CLKBUF_X2 inst_22767 ( .A(net_22638), .Z(net_22639) );
CLKBUF_X2 inst_21822 ( .A(net_21390), .Z(net_21694) );
AOI21_X2 inst_20908 ( .ZN(net_7379), .B2(net_7378), .A(net_4858), .B1(net_1691) );
CLKBUF_X2 inst_22347 ( .A(net_22218), .Z(net_22219) );
INV_X4 inst_15036 ( .A(net_9529), .ZN(net_3358) );
INV_X4 inst_14608 ( .ZN(net_9955), .A(net_4433) );
AND2_X2 inst_21342 ( .A2(net_4669), .ZN(net_2856), .A1(net_2847) );
INV_X4 inst_17258 ( .A(net_2183), .ZN(net_952) );
INV_X4 inst_12726 ( .ZN(net_20428), .A(net_17507) );
INV_X4 inst_13066 ( .ZN(net_20199), .A(net_16228) );
NOR2_X2 inst_4721 ( .ZN(net_10006), .A2(net_4378), .A1(net_1977) );
INV_X2 inst_19668 ( .A(net_20495), .ZN(net_20481) );
INV_X4 inst_13601 ( .ZN(net_20738), .A(net_8613) );
NAND3_X2 inst_6638 ( .A3(net_10620), .ZN(net_8957), .A1(net_6087), .A2(net_4898) );
INV_X4 inst_13019 ( .ZN(net_16643), .A(net_16423) );
OAI21_X2 inst_2207 ( .A(net_12609), .B1(net_11212), .ZN(net_8535), .B2(net_4331) );
CLKBUF_X2 inst_22887 ( .A(net_21543), .Z(net_22759) );
NAND2_X2 inst_7841 ( .A1(net_21155), .ZN(net_18621), .A2(net_18620) );
INV_X4 inst_16254 ( .ZN(net_3648), .A(net_1038) );
NAND2_X2 inst_10088 ( .A1(net_10279), .ZN(net_8626), .A2(net_8625) );
INV_X4 inst_17086 ( .ZN(net_810), .A(net_532) );
INV_X4 inst_15692 ( .ZN(net_15810), .A(net_10182) );
NAND3_X2 inst_5902 ( .ZN(net_15135), .A3(net_13385), .A2(net_12661), .A1(net_9770) );
NAND2_X4 inst_7322 ( .ZN(net_8022), .A1(net_5109), .A2(net_955) );
NOR2_X2 inst_3892 ( .A2(net_20776), .ZN(net_9229), .A1(net_1502) );
INV_X4 inst_16265 ( .ZN(net_1350), .A(net_1349) );
INV_X4 inst_14906 ( .A(net_3589), .ZN(net_3588) );
NAND2_X2 inst_8829 ( .ZN(net_19628), .A2(net_14840), .A1(net_10082) );
AOI21_X2 inst_20829 ( .ZN(net_9860), .B1(net_5976), .B2(net_3297), .A(net_3100) );
NOR2_X2 inst_3930 ( .A1(net_13734), .ZN(net_12187), .A2(net_8736) );
NOR2_X4 inst_2867 ( .ZN(net_19257), .A2(net_9357), .A1(net_7589) );
INV_X4 inst_16388 ( .ZN(net_2477), .A(net_1276) );
CLKBUF_X2 inst_22894 ( .A(net_22574), .Z(net_22766) );
NAND2_X2 inst_9768 ( .ZN(net_11699), .A2(net_9812), .A1(net_8639) );
AND2_X4 inst_21153 ( .ZN(net_17092), .A2(net_16431), .A1(net_15538) );
AOI221_X4 inst_20070 ( .B1(net_20661), .C1(net_16644), .ZN(net_16290), .C2(net_15981), .A(net_15962), .B2(net_15936) );
NAND2_X2 inst_7953 ( .ZN(net_18398), .A2(net_18393), .A1(net_17648) );
INV_X4 inst_17147 ( .ZN(net_6589), .A(net_5454) );
INV_X4 inst_14235 ( .ZN(net_7568), .A(net_5078) );
CLKBUF_X2 inst_21938 ( .A(net_21809), .Z(net_21810) );
NOR2_X4 inst_3305 ( .ZN(net_2358), .A1(net_886), .A2(net_225) );
INV_X4 inst_14637 ( .A(net_4785), .ZN(net_4382) );
CLKBUF_X2 inst_21971 ( .A(net_21687), .Z(net_21843) );
AOI21_X4 inst_20136 ( .ZN(net_19790), .B1(net_19370), .B2(net_15607), .A(net_14486) );
NAND2_X2 inst_10153 ( .ZN(net_14900), .A1(net_8273), .A2(net_6114) );
DFF_X1 inst_19926 ( .Q(net_21109), .D(net_12106), .CK(net_22468) );
SDFF_X2 inst_710 ( .Q(net_20895), .SE(net_18858), .SI(net_18806), .D(net_521), .CK(net_21308) );
SDFF_X2 inst_941 ( .QN(net_21040), .D(net_610), .SE(net_263), .CK(net_22529), .SI(x2333) );
NOR2_X2 inst_3350 ( .ZN(net_17957), .A1(net_17946), .A2(net_17916) );
NAND2_X2 inst_8398 ( .A1(net_21122), .ZN(net_19153), .A2(net_17146) );
XOR2_X1 inst_56 ( .A(net_21124), .Z(net_441), .B(net_440) );
NAND2_X4 inst_6835 ( .A2(net_20811), .A1(net_20810), .ZN(net_18769) );
XNOR2_X2 inst_308 ( .ZN(net_17090), .A(net_16676), .B(net_680) );
OAI21_X2 inst_1546 ( .ZN(net_17866), .A(net_17617), .B1(net_17616), .B2(net_17615) );
NAND2_X4 inst_7208 ( .ZN(net_7959), .A1(net_7958), .A2(net_3729) );
NAND2_X2 inst_11224 ( .ZN(net_3961), .A1(net_3960), .A2(net_3959) );
XNOR2_X2 inst_455 ( .ZN(net_13663), .A(net_11623), .B(net_2277) );
NAND2_X2 inst_8449 ( .ZN(net_19221), .A1(net_17101), .A2(net_17100) );
NAND2_X2 inst_10015 ( .ZN(net_10270), .A1(net_9926), .A2(net_8157) );
OAI21_X2 inst_1694 ( .ZN(net_15357), .A(net_15356), .B1(net_13635), .B2(net_12141) );
AOI22_X2 inst_20000 ( .ZN(net_14097), .B1(net_14027), .A1(net_12006), .B2(net_10854), .A2(net_9078) );
INV_X4 inst_17153 ( .A(net_821), .ZN(net_754) );
INV_X4 inst_17158 ( .ZN(net_2671), .A(net_1848) );
OAI211_X2 inst_2540 ( .ZN(net_10830), .A(net_10829), .C2(net_10818), .B(net_9366), .C1(net_4221) );
NAND2_X4 inst_6833 ( .A2(net_18905), .A1(net_18904), .ZN(net_18789) );
AOI21_X2 inst_20700 ( .ZN(net_12138), .B1(net_12137), .A(net_8751), .B2(net_8018) );
AOI21_X2 inst_20601 ( .B2(net_19258), .B1(net_19257), .ZN(net_13835), .A(net_296) );
INV_X4 inst_13298 ( .ZN(net_13562), .A(net_12336) );
INV_X4 inst_17231 ( .ZN(net_674), .A(net_673) );
NAND2_X4 inst_7052 ( .A2(net_20288), .A1(net_20287), .ZN(net_16677) );
NAND3_X2 inst_6602 ( .A3(net_11363), .ZN(net_9884), .A1(net_6013), .A2(net_3346) );
NAND2_X2 inst_8114 ( .A2(net_20076), .ZN(net_19341), .A1(net_18084) );
NOR2_X4 inst_3024 ( .A2(net_20755), .ZN(net_6615), .A1(net_4291) );
AOI21_X4 inst_20137 ( .ZN(net_16078), .B1(net_15926), .B2(net_15557), .A(net_15459) );
INV_X2 inst_18406 ( .ZN(net_16804), .A(net_16560) );
NAND2_X2 inst_8454 ( .ZN(net_17192), .A2(net_16745), .A1(net_16608) );
AND2_X2 inst_21293 ( .A2(net_11518), .ZN(net_11496), .A1(net_761) );
INV_X4 inst_17942 ( .A(net_21209), .ZN(net_15957) );
NAND2_X2 inst_11860 ( .ZN(net_2463), .A1(net_1660), .A2(net_1291) );
INV_X4 inst_16370 ( .ZN(net_2070), .A(net_1040) );
NOR2_X2 inst_3951 ( .ZN(net_8605), .A2(net_8604), .A1(net_6618) );
NAND2_X2 inst_8240 ( .ZN(net_17813), .A2(net_17562), .A1(net_17491) );
INV_X4 inst_16337 ( .ZN(net_10812), .A(net_1300) );
NOR2_X2 inst_4282 ( .ZN(net_12380), .A1(net_7357), .A2(net_4604) );
NAND4_X2 inst_5428 ( .ZN(net_14116), .A4(net_13849), .A3(net_9528), .A1(net_8726), .A2(net_8614) );
AOI21_X2 inst_20360 ( .ZN(net_15667), .A(net_15666), .B2(net_14939), .B1(net_13985) );
INV_X4 inst_18197 ( .A(net_21156), .ZN(net_580) );
NOR2_X4 inst_2943 ( .ZN(net_6925), .A1(net_5527), .A2(net_4161) );
AOI21_X4 inst_20127 ( .ZN(net_19634), .B1(net_19099), .A(net_14082), .B2(net_1171) );
OAI21_X2 inst_1593 ( .A(net_20920), .B2(net_20137), .B1(net_20136), .ZN(net_19539) );
INV_X2 inst_19479 ( .A(net_10398), .ZN(net_1399) );
INV_X2 inst_18595 ( .ZN(net_10039), .A(net_8548) );
SDFF_X2 inst_724 ( .Q(net_20878), .SE(net_18584), .SI(net_18572), .D(net_5707), .CK(net_21926) );
CLKBUF_X2 inst_22176 ( .A(net_22047), .Z(net_22048) );
INV_X4 inst_17526 ( .ZN(net_1823), .A(net_279) );
INV_X4 inst_14869 ( .ZN(net_4779), .A(net_3727) );
SDFF_X2 inst_975 ( .QN(net_21049), .D(net_697), .SE(net_253), .CK(net_21730), .SI(x2197) );
INV_X4 inst_15546 ( .ZN(net_3467), .A(net_2357) );
AOI22_X2 inst_19959 ( .ZN(net_16269), .A2(net_15982), .A1(net_15666), .B2(net_13162), .B1(net_1906) );
INV_X4 inst_16677 ( .A(net_1563), .ZN(net_1462) );
INV_X4 inst_13683 ( .ZN(net_10200), .A(net_7977) );
NOR2_X4 inst_3191 ( .A1(net_20487), .ZN(net_3421), .A2(net_3102) );
NOR3_X2 inst_2789 ( .A2(net_15202), .A3(net_12852), .A1(net_9959), .ZN(net_5287) );
NAND2_X2 inst_7792 ( .ZN(net_18711), .A2(net_18668), .A1(net_17919) );
NAND2_X2 inst_9504 ( .ZN(net_11337), .A2(net_10480), .A1(net_8263) );
CLKBUF_X2 inst_22727 ( .A(net_22598), .Z(net_22599) );
NAND3_X2 inst_5714 ( .ZN(net_16161), .A3(net_15785), .A2(net_14282), .A1(net_13133) );
NAND2_X2 inst_10110 ( .ZN(net_8428), .A2(net_7731), .A1(net_4144) );
NAND2_X2 inst_10783 ( .ZN(net_20414), .A1(net_8865), .A2(net_5593) );
OAI21_X2 inst_1804 ( .ZN(net_14477), .A(net_14476), .B2(net_12524), .B1(net_8430) );
AOI21_X2 inst_20470 ( .ZN(net_19852), .A(net_13559), .B2(net_12837), .B1(net_238) );
NAND3_X2 inst_6418 ( .ZN(net_11945), .A3(net_10213), .A1(net_7654), .A2(net_6186) );
INV_X2 inst_18778 ( .ZN(net_11076), .A(net_7537) );
NAND2_X2 inst_11037 ( .ZN(net_7807), .A1(net_4762), .A2(net_4741) );
OAI21_X2 inst_2183 ( .A(net_8959), .ZN(net_8835), .B2(net_5481), .B1(net_4496) );
AOI21_X2 inst_20489 ( .ZN(net_14766), .B1(net_14600), .B2(net_13202), .A(net_11481) );
NAND2_X2 inst_11981 ( .ZN(net_5866), .A2(net_4329), .A1(net_359) );
NOR2_X2 inst_5068 ( .ZN(net_13699), .A2(net_10676), .A1(net_710) );
NOR3_X2 inst_2659 ( .ZN(net_15151), .A3(net_14023), .A2(net_12759), .A1(net_11496) );
NAND3_X2 inst_6545 ( .ZN(net_10563), .A3(net_10562), .A1(net_7614), .A2(net_5911) );
INV_X4 inst_13878 ( .ZN(net_10757), .A(net_7367) );
CLKBUF_X2 inst_21627 ( .A(net_21338), .Z(net_21499) );
NOR2_X2 inst_5018 ( .A1(net_1339), .ZN(net_1239), .A2(net_1101) );
NAND2_X2 inst_11609 ( .A2(net_6951), .ZN(net_4529), .A1(net_3459) );
INV_X4 inst_18144 ( .A(net_20863), .ZN(net_272) );
NAND3_X2 inst_5641 ( .ZN(net_17988), .A2(net_17979), .A3(net_17978), .A1(net_17874) );
INV_X2 inst_19511 ( .ZN(net_1185), .A(net_1184) );
NAND2_X2 inst_11134 ( .A2(net_6437), .ZN(net_5410), .A1(net_4264) );
INV_X2 inst_18708 ( .A(net_8657), .ZN(net_8240) );
INV_X2 inst_18814 ( .A(net_7433), .ZN(net_7288) );
OR2_X2 inst_1155 ( .ZN(net_19683), .A2(net_8765), .A1(net_6917) );
XNOR2_X2 inst_207 ( .ZN(net_17577), .A(net_17576), .B(net_10496) );
INV_X4 inst_16169 ( .ZN(net_2726), .A(net_1413) );
NAND2_X2 inst_8886 ( .ZN(net_15147), .A2(net_14099), .A1(net_5745) );
INV_X4 inst_14467 ( .ZN(net_4913), .A(net_4912) );
AOI21_X2 inst_20618 ( .ZN(net_13536), .B1(net_12160), .A(net_5783), .B2(net_5026) );
INV_X4 inst_18096 ( .A(net_21085), .ZN(net_591) );
NAND2_X2 inst_10490 ( .ZN(net_19403), .A1(net_10930), .A2(net_6931) );
NAND2_X2 inst_9615 ( .ZN(net_10707), .A2(net_8445), .A1(net_8097) );
CLKBUF_X2 inst_22094 ( .A(net_21965), .Z(net_21966) );
NAND2_X2 inst_9912 ( .A2(net_12795), .ZN(net_11513), .A1(net_9313) );
OR2_X2 inst_1215 ( .ZN(net_8091), .A1(net_1624), .A2(net_1118) );
NAND2_X2 inst_9303 ( .ZN(net_13427), .A2(net_9218), .A1(net_7253) );
XNOR2_X2 inst_131 ( .B(net_21228), .ZN(net_18246), .A(net_18134) );
INV_X4 inst_15353 ( .A(net_9085), .ZN(net_2589) );
CLKBUF_X2 inst_22768 ( .A(net_22626), .Z(net_22640) );
NAND3_X2 inst_6104 ( .ZN(net_13899), .A3(net_13898), .A2(net_11352), .A1(net_5688) );
CLKBUF_X2 inst_22563 ( .A(net_22434), .Z(net_22435) );
INV_X4 inst_16412 ( .ZN(net_9733), .A(net_749) );
XOR2_X2 inst_47 ( .A(net_21207), .Z(net_470), .B(net_469) );
INV_X8 inst_12360 ( .A(net_20860), .ZN(net_3919) );
INV_X4 inst_14958 ( .ZN(net_3495), .A(net_3494) );
AOI21_X4 inst_20231 ( .ZN(net_19736), .B1(net_12884), .A(net_11069), .B2(net_8948) );
OAI21_X2 inst_1984 ( .ZN(net_12065), .A(net_11468), .B1(net_11406), .B2(net_10720) );
NAND4_X4 inst_5231 ( .A2(net_19877), .A1(net_19876), .A4(net_19098), .ZN(net_16008), .A3(net_11969) );
INV_X4 inst_14567 ( .ZN(net_20409), .A(net_4559) );
NAND2_X2 inst_9458 ( .A1(net_13703), .ZN(net_11500), .A2(net_11499) );
INV_X4 inst_15563 ( .ZN(net_5402), .A(net_955) );
NAND3_X2 inst_6520 ( .ZN(net_10640), .A1(net_10639), .A2(net_10638), .A3(net_10637) );
INV_X4 inst_14356 ( .ZN(net_5830), .A(net_5255) );
INV_X8 inst_12397 ( .A(net_301), .ZN(net_248) );
NOR2_X2 inst_4101 ( .ZN(net_19809), .A2(net_9099), .A1(net_8460) );
NAND2_X2 inst_10316 ( .ZN(net_12798), .A2(net_7846), .A1(net_7844) );
INV_X2 inst_19507 ( .A(net_1637), .ZN(net_1223) );
NAND2_X2 inst_9469 ( .A1(net_12763), .ZN(net_12618), .A2(net_11480) );
NOR2_X2 inst_4792 ( .ZN(net_2780), .A1(net_2779), .A2(net_1325) );
INV_X4 inst_14027 ( .ZN(net_12471), .A(net_6289) );
CLKBUF_X2 inst_22842 ( .A(net_22713), .Z(net_22714) );
INV_X4 inst_18249 ( .A(net_20861), .ZN(net_318) );
INV_X4 inst_17078 ( .ZN(net_7432), .A(net_6788) );
INV_X4 inst_12738 ( .ZN(net_17613), .A(net_17552) );
XNOR2_X2 inst_434 ( .ZN(net_16268), .A(net_16267), .B(net_16090) );
NOR2_X2 inst_3455 ( .ZN(net_14853), .A2(net_14147), .A1(net_1306) );
INV_X4 inst_14099 ( .ZN(net_9021), .A(net_8013) );
OAI21_X4 inst_1392 ( .A(net_20864), .B2(net_19072), .B1(net_19071), .ZN(net_16280) );
NAND2_X4 inst_7376 ( .A1(net_19647), .ZN(net_11090), .A2(net_4288) );
NAND2_X2 inst_11816 ( .ZN(net_2987), .A1(net_1568), .A2(net_711) );
NOR2_X2 inst_4044 ( .ZN(net_11739), .A2(net_6020), .A1(net_1441) );
INV_X2 inst_18926 ( .ZN(net_5907), .A(net_5906) );
INV_X4 inst_17116 ( .A(net_898), .ZN(net_782) );
INV_X4 inst_16971 ( .A(net_7917), .ZN(net_7822) );
AOI21_X2 inst_20812 ( .ZN(net_10088), .A(net_10087), .B1(net_6776), .B2(net_6023) );
INV_X4 inst_16282 ( .ZN(net_15202), .A(net_15158) );
INV_X4 inst_16697 ( .A(net_6321), .ZN(net_1067) );
OAI21_X4 inst_1476 ( .B2(net_18907), .B1(net_18906), .ZN(net_18891), .A(net_239) );
NAND2_X2 inst_8265 ( .A1(net_20709), .ZN(net_17661), .A2(net_17660) );
OAI21_X2 inst_2249 ( .A(net_11440), .ZN(net_7301), .B2(net_5521), .B1(net_3401) );
INV_X4 inst_18187 ( .A(net_21158), .ZN(net_16680) );
INV_X4 inst_13773 ( .ZN(net_9215), .A(net_7591) );
NAND2_X2 inst_8995 ( .ZN(net_14446), .A2(net_13135), .A1(net_10070) );
NAND4_X2 inst_5404 ( .ZN(net_14682), .A2(net_12520), .A4(net_12317), .A1(net_12195), .A3(net_5025) );
OAI211_X2 inst_2390 ( .ZN(net_16166), .C1(net_16011), .B(net_15766), .A(net_11978), .C2(net_11326) );
INV_X2 inst_19581 ( .ZN(net_779), .A(net_281) );
INV_X4 inst_17315 ( .ZN(net_2942), .A(net_596) );
NAND3_X2 inst_6033 ( .ZN(net_14343), .A3(net_14342), .A1(net_8693), .A2(net_3840) );
INV_X4 inst_17592 ( .A(net_808), .ZN(net_507) );
INV_X4 inst_15149 ( .ZN(net_4028), .A(net_3076) );
INV_X4 inst_14305 ( .ZN(net_6817), .A(net_5519) );
NAND2_X2 inst_8424 ( .A2(net_19455), .ZN(net_17182), .A1(net_16675) );
NOR2_X2 inst_3871 ( .ZN(net_9369), .A1(net_7492), .A2(net_6670) );
AND3_X4 inst_21112 ( .ZN(net_15683), .A3(net_15092), .A2(net_12816), .A1(net_10115) );
NAND2_X2 inst_9268 ( .A1(net_15012), .ZN(net_14863), .A2(net_10908) );
NOR2_X2 inst_4449 ( .ZN(net_5932), .A1(net_4770), .A2(net_2764) );
NAND3_X2 inst_6077 ( .ZN(net_14090), .A1(net_12323), .A3(net_8935), .A2(net_2962) );
NAND2_X4 inst_7637 ( .ZN(net_1969), .A2(net_1662), .A1(net_597) );
OAI21_X2 inst_2045 ( .ZN(net_11183), .B1(net_11182), .B2(net_11181), .A(net_7863) );
INV_X2 inst_19289 ( .A(net_11208), .ZN(net_2873) );
INV_X4 inst_17807 ( .ZN(net_6692), .A(net_146) );
NAND2_X2 inst_11746 ( .ZN(net_5292), .A1(net_4907), .A2(net_2129) );
OAI22_X2 inst_1311 ( .A2(net_9623), .ZN(net_8474), .B1(net_8473), .B2(net_8472), .A1(net_4296) );
NAND2_X2 inst_9307 ( .ZN(net_12369), .A1(net_10550), .A2(net_9208) );
NAND2_X4 inst_7185 ( .ZN(net_12193), .A2(net_9330), .A1(net_8903) );
NOR2_X2 inst_3415 ( .ZN(net_15610), .A2(net_14895), .A1(net_1822) );
INV_X2 inst_19417 ( .ZN(net_4138), .A(net_1884) );
NAND2_X2 inst_9534 ( .ZN(net_11078), .A1(net_11077), .A2(net_11076) );
INV_X4 inst_16667 ( .ZN(net_1796), .A(net_813) );
NAND2_X2 inst_10780 ( .A1(net_11442), .ZN(net_5601), .A2(net_4411) );
NOR2_X2 inst_4654 ( .ZN(net_3506), .A1(net_2702), .A2(net_940) );
OAI21_X2 inst_1640 ( .ZN(net_20301), .A(net_16259), .B1(net_15336), .B2(net_14804) );
AOI21_X2 inst_20622 ( .ZN(net_20426), .A(net_15039), .B1(net_9377), .B2(net_9013) );
NAND2_X2 inst_11359 ( .ZN(net_3615), .A2(net_3614), .A1(net_1925) );
INV_X4 inst_13928 ( .A(net_6870), .ZN(net_6869) );
AND4_X4 inst_21090 ( .ZN(net_19198), .A2(net_12981), .A4(net_10057), .A3(net_8156), .A1(net_5880) );
INV_X4 inst_15127 ( .ZN(net_5571), .A(net_3144) );
NOR2_X2 inst_4747 ( .ZN(net_4003), .A1(net_3184), .A2(net_3029) );
NAND2_X4 inst_7682 ( .ZN(net_1303), .A2(net_646), .A1(net_234) );
AOI21_X2 inst_20637 ( .ZN(net_13276), .B1(net_10947), .B2(net_9888), .A(net_6870) );
NAND2_X4 inst_7571 ( .A1(net_19016), .ZN(net_1635), .A2(net_445) );
NOR2_X2 inst_4630 ( .ZN(net_3593), .A1(net_3592), .A2(net_3591) );
OAI211_X2 inst_2509 ( .ZN(net_12498), .A(net_12497), .C1(net_12496), .C2(net_12495), .B(net_5193) );
NAND3_X2 inst_5971 ( .ZN(net_14771), .A3(net_13411), .A1(net_11671), .A2(net_10338) );
NOR2_X4 inst_3091 ( .ZN(net_5462), .A1(net_4383), .A2(net_4290) );
NOR2_X2 inst_4197 ( .ZN(net_7973), .A1(net_6706), .A2(net_6705) );
INV_X4 inst_15784 ( .ZN(net_13781), .A(net_13448) );
INV_X4 inst_16151 ( .ZN(net_10182), .A(net_9656) );
INV_X4 inst_15914 ( .ZN(net_13512), .A(net_8278) );
INV_X4 inst_15354 ( .ZN(net_19414), .A(net_15991) );
NAND2_X4 inst_7400 ( .ZN(net_4418), .A1(net_3299), .A2(net_2490) );
INV_X4 inst_13745 ( .A(net_12483), .ZN(net_7632) );
INV_X4 inst_17176 ( .ZN(net_6951), .A(net_733) );
NOR2_X2 inst_4524 ( .ZN(net_7006), .A2(net_3381), .A1(net_3371) );
NOR2_X2 inst_4871 ( .ZN(net_2226), .A2(net_1723), .A1(net_85) );
INV_X4 inst_16030 ( .ZN(net_2108), .A(net_1143) );
NAND4_X2 inst_5520 ( .ZN(net_4421), .A2(net_4420), .A3(net_2524), .A4(net_1098), .A1(x7654) );
AOI21_X2 inst_20924 ( .ZN(net_7174), .A(net_7173), .B1(net_6476), .B2(net_3897) );
NOR2_X2 inst_4257 ( .ZN(net_6283), .A2(net_6076), .A1(net_4209) );
NOR2_X2 inst_4586 ( .A1(net_8273), .ZN(net_7207), .A2(net_3815) );
INV_X4 inst_18342 ( .A(net_20762), .ZN(net_20761) );
INV_X4 inst_13722 ( .ZN(net_12647), .A(net_7806) );
OAI22_X2 inst_1317 ( .A1(net_6719), .ZN(net_5245), .B1(net_5244), .B2(net_5243), .A2(net_3219) );
NAND3_X1 inst_6820 ( .ZN(net_18795), .A2(net_18783), .A3(net_18782), .A1(net_17736) );
AOI211_X2 inst_21078 ( .C2(net_7428), .ZN(net_6450), .B(net_6449), .A(net_3236), .C1(net_187) );
NAND2_X2 inst_9623 ( .ZN(net_10668), .A1(net_10667), .A2(net_8555) );
INV_X4 inst_12603 ( .ZN(net_18128), .A(net_18085) );
INV_X2 inst_19321 ( .A(net_3355), .ZN(net_2605) );
XNOR2_X2 inst_624 ( .A(net_21145), .ZN(net_16265), .B(net_466) );
NAND3_X2 inst_6284 ( .ZN(net_12868), .A3(net_12528), .A2(net_12471), .A1(net_6364) );
INV_X4 inst_17767 ( .A(net_275), .ZN(net_155) );
NAND3_X2 inst_5728 ( .ZN(net_19380), .A3(net_15815), .A2(net_15580), .A1(net_11585) );
AND2_X4 inst_21234 ( .ZN(net_19699), .A1(net_9350), .A2(net_4166) );
NAND3_X2 inst_6404 ( .ZN(net_11975), .A2(net_11974), .A3(net_9469), .A1(net_2614) );
CLKBUF_X2 inst_21436 ( .A(net_21307), .Z(net_21308) );
NAND3_X2 inst_6419 ( .A2(net_12516), .ZN(net_11944), .A3(net_10245), .A1(net_6383) );
NAND2_X2 inst_9886 ( .ZN(net_12844), .A1(net_9421), .A2(net_9388) );
INV_X4 inst_18327 ( .A(net_20923), .ZN(net_20545) );
NAND2_X2 inst_11247 ( .ZN(net_8985), .A2(net_4242), .A1(net_117) );
NAND2_X2 inst_9375 ( .ZN(net_11987), .A2(net_10128), .A1(net_4476) );
AOI21_X2 inst_20836 ( .B1(net_12330), .ZN(net_9300), .A(net_5849), .B2(net_3955) );
NOR2_X2 inst_3624 ( .A1(net_14430), .ZN(net_13578), .A2(net_12408) );
INV_X4 inst_17048 ( .ZN(net_5785), .A(net_5476) );
INV_X4 inst_13207 ( .ZN(net_13727), .A(net_12986) );
INV_X4 inst_14598 ( .ZN(net_13922), .A(net_11779) );
NAND2_X2 inst_11440 ( .ZN(net_3727), .A1(net_3310), .A2(net_2981) );
CLKBUF_X2 inst_22905 ( .A(net_22776), .Z(net_22777) );
INV_X8 inst_12389 ( .ZN(net_275), .A(net_137) );
INV_X4 inst_16495 ( .ZN(net_1712), .A(net_1194) );
INV_X4 inst_13262 ( .ZN(net_20196), .A(net_11599) );
INV_X4 inst_14805 ( .ZN(net_5018), .A(net_3981) );
NOR2_X2 inst_4532 ( .ZN(net_6946), .A2(net_4041), .A1(net_1163) );
NAND3_X2 inst_6277 ( .ZN(net_20233), .A3(net_12854), .A2(net_11886), .A1(net_11185) );
INV_X4 inst_12962 ( .ZN(net_18886), .A(net_16435) );
NAND3_X4 inst_5600 ( .ZN(net_14532), .A3(net_12189), .A2(net_11941), .A1(net_9489) );
NOR2_X2 inst_3508 ( .ZN(net_13964), .A2(net_12107), .A1(net_8613) );
CLKBUF_X2 inst_22831 ( .A(net_22654), .Z(net_22703) );
NOR2_X2 inst_5132 ( .ZN(net_216), .A2(net_116), .A1(net_87) );
NAND3_X2 inst_6327 ( .ZN(net_12509), .A2(net_12508), .A3(net_12507), .A1(net_2924) );
INV_X4 inst_14955 ( .A(net_4109), .ZN(net_3500) );
INV_X2 inst_18519 ( .ZN(net_11523), .A(net_11522) );
OR2_X2 inst_1133 ( .ZN(net_13073), .A2(net_13072), .A1(net_8981) );
NOR2_X2 inst_4580 ( .ZN(net_3839), .A2(net_3838), .A1(net_170) );
NAND2_X2 inst_9990 ( .ZN(net_12169), .A2(net_8846), .A1(net_8169) );
OAI21_X2 inst_2103 ( .ZN(net_10062), .A(net_10061), .B1(net_8404), .B2(net_6281) );
INV_X4 inst_16577 ( .A(net_11296), .ZN(net_5344) );
NAND2_X2 inst_8710 ( .A1(net_21212), .ZN(net_16250), .A2(net_16053) );
INV_X4 inst_14040 ( .ZN(net_11307), .A(net_7084) );
INV_X4 inst_16234 ( .ZN(net_2750), .A(net_1375) );
XNOR2_X2 inst_339 ( .B(net_21196), .ZN(net_16966), .A(net_16965) );
NOR2_X2 inst_4750 ( .ZN(net_5423), .A2(net_3019), .A1(net_1689) );
INV_X4 inst_17551 ( .ZN(net_5951), .A(net_1165) );
INV_X4 inst_13995 ( .ZN(net_6413), .A(net_5271) );
XNOR2_X2 inst_351 ( .ZN(net_16937), .A(net_16527), .B(net_342) );
INV_X4 inst_17379 ( .ZN(net_5120), .A(net_170) );
NAND3_X2 inst_6615 ( .A3(net_19374), .ZN(net_9069), .A1(net_6970), .A2(net_5312) );
NAND2_X2 inst_10257 ( .ZN(net_7996), .A2(net_6086), .A1(net_5016) );
NAND2_X2 inst_9557 ( .A1(net_11550), .ZN(net_11005), .A2(net_11004) );
NAND2_X2 inst_7852 ( .ZN(net_18587), .A2(net_18579), .A1(net_18574) );
INV_X4 inst_12507 ( .ZN(net_18615), .A(net_18608) );
INV_X2 inst_19650 ( .A(net_19465), .ZN(net_19464) );
CLKBUF_X2 inst_22854 ( .A(net_22056), .Z(net_22726) );
NAND2_X4 inst_7651 ( .ZN(net_1075), .A2(net_897), .A1(net_161) );
AND3_X2 inst_21144 ( .ZN(net_7744), .A2(net_7743), .A3(net_7380), .A1(net_4328) );
OAI21_X2 inst_1560 ( .ZN(net_17442), .B1(net_17441), .A(net_17176), .B2(net_17175) );
NAND2_X2 inst_11463 ( .A2(net_4358), .ZN(net_3186), .A1(net_1508) );
CLKBUF_X2 inst_22669 ( .A(net_22540), .Z(net_22541) );
INV_X4 inst_12622 ( .ZN(net_17994), .A(net_17993) );
NAND2_X2 inst_10868 ( .ZN(net_6709), .A1(net_5632), .A2(net_5401) );
AOI21_X4 inst_20250 ( .B1(net_8442), .ZN(net_8129), .A(net_8128), .B2(net_2635) );
NAND2_X2 inst_10994 ( .ZN(net_9923), .A1(net_8369), .A2(net_4859) );
INV_X4 inst_13915 ( .A(net_8734), .ZN(net_7318) );
CLKBUF_X2 inst_22021 ( .A(net_21266), .Z(net_21893) );
NAND2_X2 inst_10203 ( .A1(net_8709), .ZN(net_8121), .A2(net_8120) );
NAND2_X4 inst_7035 ( .A2(net_19636), .A1(net_16588), .ZN(net_16587) );
NAND2_X2 inst_9224 ( .ZN(net_19893), .A2(net_10841), .A1(net_1244) );
INV_X4 inst_15205 ( .ZN(net_3524), .A(net_2905) );
AOI211_X2 inst_20998 ( .ZN(net_15970), .C1(net_15969), .C2(net_15570), .B(net_10385), .A(net_8647) );
NAND2_X2 inst_11164 ( .A1(net_8226), .ZN(net_4178), .A2(net_4177) );
NAND2_X2 inst_10161 ( .ZN(net_8257), .A1(net_8256), .A2(net_8100) );
SDFF_X2 inst_847 ( .Q(net_21213), .SI(net_17313), .SE(net_125), .CK(net_22306), .D(x7584) );
NOR3_X2 inst_2720 ( .ZN(net_13302), .A2(net_11382), .A3(net_9864), .A1(net_7001) );
NAND3_X2 inst_6577 ( .A3(net_12038), .ZN(net_10451), .A2(net_7495), .A1(net_6082) );
OAI21_X2 inst_1716 ( .ZN(net_15188), .B2(net_13954), .A(net_11407), .B1(net_7038) );
OAI21_X2 inst_1942 ( .ZN(net_12768), .B1(net_12708), .A(net_10220), .B2(net_8467) );
NAND2_X2 inst_10857 ( .ZN(net_12644), .A1(net_11189), .A2(net_5451) );
INV_X4 inst_18271 ( .A(net_19452), .ZN(net_19451) );
NAND2_X2 inst_9788 ( .A1(net_11297), .ZN(net_11094), .A2(net_9743) );
NAND3_X2 inst_5950 ( .ZN(net_14885), .A3(net_14798), .A2(net_9693), .A1(net_8294) );
INV_X4 inst_13573 ( .ZN(net_9127), .A(net_9126) );
NAND2_X2 inst_9136 ( .ZN(net_13453), .A1(net_13452), .A2(net_10839) );
NOR3_X2 inst_2648 ( .A3(net_20847), .A1(net_20846), .ZN(net_15715), .A2(net_12713) );
NAND2_X4 inst_7055 ( .A2(net_19539), .A1(net_19538), .ZN(net_16393) );
AOI21_X2 inst_20406 ( .B1(net_19620), .ZN(net_15333), .B2(net_10709), .A(net_5263) );
INV_X4 inst_15470 ( .ZN(net_15522), .A(net_14986) );
NAND2_X2 inst_7919 ( .ZN(net_18455), .A1(net_18380), .A2(net_18332) );
NAND2_X2 inst_8372 ( .ZN(net_19043), .A1(net_17355), .A2(net_16859) );
OR2_X2 inst_1146 ( .A1(net_12339), .ZN(net_10107), .A2(net_10106) );
INV_X2 inst_18503 ( .ZN(net_12000), .A(net_11999) );
INV_X4 inst_12947 ( .A(net_16628), .ZN(net_16627) );
NOR2_X2 inst_3708 ( .ZN(net_11043), .A2(net_11042), .A1(net_9158) );
AOI21_X2 inst_20405 ( .ZN(net_15341), .B1(net_15340), .B2(net_13748), .A(net_10294) );
INV_X2 inst_18570 ( .ZN(net_10745), .A(net_10744) );
NOR2_X2 inst_4023 ( .ZN(net_9563), .A1(net_8021), .A2(net_6248) );
NOR2_X2 inst_3673 ( .A2(net_11607), .ZN(net_11477), .A1(net_11476) );
NOR2_X4 inst_3105 ( .A2(net_20868), .ZN(net_7009), .A1(net_4081) );
NAND4_X4 inst_5162 ( .ZN(net_18093), .A4(net_18071), .A1(net_18062), .A2(net_15843), .A3(net_13139) );
CLKBUF_X2 inst_21948 ( .A(net_21386), .Z(net_21820) );
INV_X2 inst_18422 ( .ZN(net_15304), .A(net_15005) );
NOR2_X2 inst_4519 ( .ZN(net_4137), .A2(net_4136), .A1(net_832) );
NAND4_X2 inst_5349 ( .ZN(net_15418), .A1(net_14664), .A3(net_14537), .A4(net_13802), .A2(net_7212) );
NAND3_X2 inst_6210 ( .ZN(net_13272), .A2(net_11898), .A3(net_9882), .A1(net_9340) );
NAND2_X2 inst_9899 ( .ZN(net_12165), .A1(net_9365), .A2(net_6555) );
NOR2_X2 inst_3539 ( .A1(net_19650), .ZN(net_13411), .A2(net_9819) );
OAI211_X2 inst_2457 ( .ZN(net_14217), .A(net_14216), .B(net_14215), .C2(net_14214), .C1(net_6360) );
INV_X4 inst_16442 ( .ZN(net_2846), .A(net_1234) );
NAND2_X2 inst_8307 ( .ZN(net_19295), .A2(net_17653), .A1(net_219) );
NAND2_X2 inst_10188 ( .ZN(net_8170), .A1(net_8169), .A2(net_8168) );
XNOR2_X2 inst_274 ( .B(net_21141), .A(net_17441), .ZN(net_17191) );
INV_X4 inst_15076 ( .ZN(net_16127), .A(net_15542) );
INV_X4 inst_14543 ( .ZN(net_10818), .A(net_4637) );
NAND2_X4 inst_7329 ( .ZN(net_6173), .A1(net_5009), .A2(net_4393) );
NOR2_X4 inst_2817 ( .A2(net_19209), .A1(net_19208), .ZN(net_16544) );
INV_X4 inst_13135 ( .ZN(net_19743), .A(net_14749) );
INV_X4 inst_13436 ( .ZN(net_12582), .A(net_9818) );
NOR2_X4 inst_3207 ( .A1(net_20564), .ZN(net_7125), .A2(net_3030) );
NOR2_X4 inst_3143 ( .ZN(net_6550), .A2(net_4026), .A1(net_85) );
NAND2_X4 inst_7112 ( .ZN(net_12726), .A2(net_11135), .A1(net_6626) );
DFF_X2 inst_19781 ( .QN(net_21104), .D(net_1993), .CK(net_22187) );
NAND2_X2 inst_11387 ( .A2(net_3641), .ZN(net_3526), .A1(net_923) );
NOR3_X2 inst_2696 ( .ZN(net_14096), .A3(net_10482), .A2(net_9931), .A1(net_7303) );
INV_X4 inst_14063 ( .A(net_7979), .ZN(net_7601) );
NAND2_X4 inst_7136 ( .A1(net_20380), .ZN(net_14301), .A2(net_10188) );
NOR2_X4 inst_2880 ( .ZN(net_20640), .A1(net_9455), .A2(net_6690) );
OAI21_X2 inst_1771 ( .A(net_15468), .ZN(net_14693), .B2(net_11939), .B1(net_10408) );
INV_X4 inst_14402 ( .ZN(net_5112), .A(net_5111) );
NOR3_X2 inst_2660 ( .ZN(net_20142), .A3(net_12821), .A2(net_12590), .A1(net_8890) );
NAND2_X2 inst_7859 ( .ZN(net_18568), .A1(net_18547), .A2(net_18517) );
CLKBUF_X2 inst_22956 ( .A(net_22827), .Z(net_22828) );
INV_X4 inst_13729 ( .ZN(net_11891), .A(net_7774) );
OAI211_X2 inst_2389 ( .ZN(net_16196), .A(net_15975), .B(net_15837), .C2(net_13648), .C1(net_4452) );
INV_X4 inst_17967 ( .A(net_20985), .ZN(net_2030) );
NAND3_X2 inst_5912 ( .ZN(net_15014), .A3(net_12823), .A2(net_12672), .A1(net_6929) );
NAND2_X2 inst_10802 ( .ZN(net_5548), .A2(net_5547), .A1(net_1037) );
INV_X4 inst_16906 ( .ZN(net_6201), .A(net_1813) );
NAND3_X2 inst_6199 ( .ZN(net_19944), .A3(net_13168), .A2(net_12829), .A1(net_7154) );
AOI21_X2 inst_20369 ( .B1(net_19103), .ZN(net_15629), .B2(net_15628), .A(net_11848) );
INV_X4 inst_16406 ( .A(net_10105), .ZN(net_8685) );
NOR2_X2 inst_4946 ( .ZN(net_1683), .A1(net_1682), .A2(net_1681) );
OAI21_X2 inst_2148 ( .ZN(net_9621), .A(net_9620), .B2(net_9619), .B1(net_2577) );
AOI21_X2 inst_20301 ( .B2(net_19733), .B1(net_19732), .ZN(net_16102), .A(net_15833) );
NAND3_X2 inst_5784 ( .ZN(net_19507), .A3(net_14767), .A1(net_12910), .A2(net_4176) );
INV_X4 inst_17947 ( .A(net_21026), .ZN(net_688) );
INV_X4 inst_13488 ( .ZN(net_11540), .A(net_9522) );
NOR2_X4 inst_2900 ( .ZN(net_20764), .A1(net_8220), .A2(net_7486) );
CLKBUF_X2 inst_22595 ( .A(net_22466), .Z(net_22467) );
NOR2_X4 inst_3247 ( .ZN(net_4316), .A1(net_2293), .A2(net_61) );
INV_X4 inst_13544 ( .A(net_12467), .ZN(net_9196) );
XNOR2_X2 inst_379 ( .B(net_21170), .A(net_17763), .ZN(net_16832) );
SDFF_X2 inst_926 ( .Q(net_21234), .SI(net_16531), .SE(net_125), .CK(net_22406), .D(x6870) );
INV_X8 inst_12348 ( .ZN(net_1682), .A(net_328) );
NAND2_X2 inst_10997 ( .ZN(net_10999), .A1(net_4915), .A2(net_4914) );
CLKBUF_X2 inst_21836 ( .A(net_21372), .Z(net_21708) );
NOR2_X2 inst_4153 ( .ZN(net_6900), .A1(net_6899), .A2(net_6898) );
INV_X4 inst_13586 ( .A(net_10749), .ZN(net_8911) );
NAND2_X2 inst_8684 ( .A2(net_16622), .ZN(net_16446), .A1(net_16445) );
NAND2_X2 inst_10624 ( .ZN(net_19733), .A1(net_6563), .A2(net_3507) );
INV_X4 inst_15741 ( .ZN(net_1951), .A(net_588) );
INV_X4 inst_16884 ( .A(net_7173), .ZN(net_1244) );
NOR2_X2 inst_3646 ( .ZN(net_13820), .A2(net_11699), .A1(net_11691) );
SDFF_X2 inst_891 ( .Q(net_21120), .D(net_16989), .SE(net_263), .CK(net_22287), .SI(x4384) );
NAND2_X2 inst_9479 ( .ZN(net_20001), .A1(net_11459), .A2(net_8995) );
NAND3_X2 inst_5682 ( .A3(net_19273), .A1(net_19272), .ZN(net_16329), .A2(net_14219) );
XNOR2_X2 inst_288 ( .A(net_17170), .ZN(net_17151), .B(net_16464) );
INV_X2 inst_19233 ( .A(net_5044), .ZN(net_3357) );
INV_X4 inst_14414 ( .ZN(net_11285), .A(net_5083) );
CLKBUF_X2 inst_22019 ( .A(net_21251), .Z(net_21891) );
NAND2_X2 inst_11729 ( .ZN(net_5243), .A2(net_2224), .A1(net_1632) );
NAND2_X4 inst_7263 ( .ZN(net_7646), .A2(net_6968), .A1(net_6366) );
OAI22_X2 inst_1298 ( .B1(net_20551), .ZN(net_20417), .B2(net_13497), .A1(net_10320), .A2(net_4668) );
INV_X4 inst_15059 ( .ZN(net_5483), .A(net_2333) );
INV_X4 inst_14636 ( .A(net_5789), .ZN(net_5274) );
NAND2_X2 inst_9147 ( .ZN(net_13404), .A1(net_10709), .A2(net_10498) );
INV_X4 inst_14856 ( .A(net_4801), .ZN(net_3808) );
NAND2_X2 inst_12032 ( .A2(net_2744), .ZN(net_1355), .A1(net_992) );
NAND2_X2 inst_8241 ( .ZN(net_17735), .A1(net_17558), .A2(net_17475) );
NAND3_X2 inst_6499 ( .ZN(net_10848), .A2(net_10847), .A3(net_6004), .A1(net_6001) );
INV_X2 inst_18484 ( .A(net_12726), .ZN(net_12427) );
XNOR2_X2 inst_372 ( .ZN(net_16992), .A(net_16843), .B(net_16842) );
NAND2_X4 inst_7388 ( .A2(net_20851), .ZN(net_6825), .A1(net_4201) );
NAND2_X2 inst_8031 ( .ZN(net_20378), .A1(net_18185), .A2(net_18160) );
AOI21_X2 inst_20297 ( .ZN(net_16128), .B1(net_16127), .B2(net_15729), .A(net_14692) );
INV_X4 inst_15142 ( .ZN(net_4366), .A(net_3112) );
INV_X4 inst_14623 ( .ZN(net_4557), .A(net_4405) );
NAND2_X2 inst_9218 ( .ZN(net_12985), .A1(net_12408), .A2(net_10336) );
NAND2_X2 inst_8512 ( .ZN(net_16917), .A1(net_16901), .A2(net_16409) );
NAND3_X2 inst_5835 ( .ZN(net_15512), .A3(net_14625), .A2(net_11759), .A1(net_5185) );
NAND2_X2 inst_11128 ( .ZN(net_4276), .A2(net_4275), .A1(net_2274) );
OAI21_X2 inst_1775 ( .B2(net_20175), .B1(net_20174), .A(net_15366), .ZN(net_14681) );
NAND3_X2 inst_6223 ( .ZN(net_13239), .A3(net_13238), .A1(net_8426), .A2(net_6660) );
AND2_X2 inst_21278 ( .ZN(net_18937), .A2(net_13770), .A1(net_13001) );
OR2_X2 inst_1172 ( .ZN(net_6005), .A2(net_6004), .A1(net_4843) );
NOR2_X2 inst_3903 ( .ZN(net_12196), .A1(net_9728), .A2(net_8356) );
INV_X4 inst_17606 ( .A(net_900), .ZN(net_601) );
NAND2_X4 inst_7467 ( .ZN(net_3490), .A2(net_2712), .A1(net_1312) );
INV_X4 inst_13454 ( .ZN(net_13018), .A(net_10213) );
CLKBUF_X2 inst_22104 ( .A(net_21345), .Z(net_21976) );
INV_X4 inst_17400 ( .ZN(net_1186), .A(net_170) );
OR2_X2 inst_1239 ( .ZN(net_2311), .A2(net_154), .A1(net_70) );
INV_X2 inst_18583 ( .ZN(net_10296), .A(net_10295) );
NAND2_X2 inst_8991 ( .A1(net_14962), .ZN(net_14462), .A2(net_12947) );
INV_X4 inst_13832 ( .ZN(net_11053), .A(net_7495) );
INV_X4 inst_14068 ( .ZN(net_7586), .A(net_6239) );
CLKBUF_X2 inst_22151 ( .A(net_21950), .Z(net_22023) );
AOI21_X2 inst_20716 ( .A(net_13184), .ZN(net_12005), .B2(net_6413), .B1(net_4154) );
NAND2_X4 inst_7094 ( .A1(net_19554), .ZN(net_14722), .A2(net_238) );
INV_X4 inst_17468 ( .ZN(net_3818), .A(net_112) );
NAND2_X2 inst_11319 ( .ZN(net_3763), .A2(net_2058), .A1(net_1243) );
NAND2_X2 inst_8556 ( .A1(net_21205), .A2(net_20501), .ZN(net_16753) );
CLKBUF_X2 inst_22269 ( .A(net_22140), .Z(net_22141) );
AOI21_X2 inst_20261 ( .A(net_20936), .B2(net_19185), .B1(net_19184), .ZN(net_18590) );
CLKBUF_X2 inst_21701 ( .A(net_21572), .Z(net_21573) );
INV_X4 inst_17427 ( .A(net_5415), .ZN(net_4707) );
INV_X4 inst_14445 ( .ZN(net_5833), .A(net_4978) );
NAND2_X2 inst_8300 ( .ZN(net_17599), .A2(net_17598), .A1(net_17588) );
INV_X4 inst_18199 ( .A(net_21235), .ZN(net_229) );
INV_X4 inst_13235 ( .ZN(net_13473), .A(net_12432) );
NAND2_X2 inst_10580 ( .ZN(net_6678), .A2(net_4921), .A1(net_4028) );
NAND2_X2 inst_8907 ( .ZN(net_14992), .A2(net_14035), .A1(net_12592) );
NOR2_X2 inst_5088 ( .A2(net_3493), .A1(net_1214), .ZN(net_850) );
INV_X4 inst_16938 ( .A(net_3862), .ZN(net_1363) );
NOR2_X2 inst_4193 ( .ZN(net_9791), .A1(net_6720), .A2(net_1931) );
INV_X4 inst_17287 ( .A(net_816), .ZN(net_630) );
INV_X4 inst_13316 ( .ZN(net_11609), .A(net_10268) );
NAND2_X4 inst_7074 ( .ZN(net_20608), .A1(net_20256), .A2(net_16395) );
INV_X4 inst_14200 ( .ZN(net_14867), .A(net_5966) );
INV_X4 inst_12858 ( .ZN(net_19404), .A(net_16897) );
XNOR2_X1 inst_686 ( .B(net_21118), .A(net_17082), .ZN(net_17070) );
NAND2_X2 inst_9871 ( .ZN(net_9473), .A2(net_9472), .A1(net_8889) );
CLKBUF_X2 inst_22545 ( .A(net_22416), .Z(net_22417) );
INV_X4 inst_14777 ( .A(net_9529), .ZN(net_4046) );
CLKBUF_X2 inst_22633 ( .A(net_22504), .Z(net_22505) );
NOR2_X2 inst_4892 ( .ZN(net_11002), .A2(net_6537), .A1(net_1542) );
NOR2_X2 inst_3643 ( .ZN(net_12019), .A2(net_8812), .A1(net_4494) );
NAND2_X2 inst_10635 ( .A1(net_6705), .ZN(net_6428), .A2(net_3910) );
NAND2_X2 inst_9075 ( .ZN(net_13836), .A2(net_12509), .A1(net_11968) );
OAI21_X2 inst_2119 ( .ZN(net_19769), .A(net_10022), .B2(net_7954), .B1(net_4752) );
OAI21_X2 inst_1929 ( .ZN(net_12949), .B1(net_9854), .B2(net_9706), .A(net_9656) );
NOR2_X2 inst_3391 ( .A2(net_19518), .A1(net_19517), .ZN(net_18914) );
NAND2_X2 inst_9422 ( .A2(net_12061), .ZN(net_11631), .A1(net_9167) );
NAND2_X2 inst_8519 ( .A1(net_20708), .ZN(net_16910), .A2(net_16909) );
NAND2_X2 inst_9025 ( .ZN(net_19635), .A1(net_14086), .A2(net_11916) );
INV_X4 inst_12472 ( .ZN(net_18761), .A(net_18760) );
OAI21_X2 inst_1794 ( .ZN(net_14595), .A(net_13255), .B2(net_6425), .B1(net_1919) );
INV_X2 inst_19404 ( .ZN(net_1997), .A(net_1996) );
INV_X4 inst_15023 ( .ZN(net_3373), .A(net_3372) );
NAND2_X2 inst_8126 ( .A2(net_20880), .ZN(net_19499), .A1(net_15770) );
CLKBUF_X2 inst_22548 ( .A(net_22419), .Z(net_22420) );
INV_X4 inst_16010 ( .ZN(net_9345), .A(net_6896) );
NOR2_X4 inst_3047 ( .ZN(net_8245), .A1(net_4916), .A2(net_131) );
NAND3_X2 inst_5957 ( .ZN(net_14846), .A2(net_13446), .A3(net_12605), .A1(net_8415) );
INV_X2 inst_19339 ( .A(net_3172), .ZN(net_2459) );
NOR2_X2 inst_3847 ( .ZN(net_9559), .A1(net_9558), .A2(net_7458) );
INV_X2 inst_18464 ( .ZN(net_12733), .A(net_11701) );
INV_X4 inst_14494 ( .ZN(net_6010), .A(net_4844) );
INV_X4 inst_18192 ( .A(net_21215), .ZN(net_165) );
NAND3_X2 inst_5756 ( .ZN(net_19700), .A1(net_15700), .A3(net_14754), .A2(net_7141) );
NAND2_X2 inst_11376 ( .ZN(net_4604), .A2(net_3554), .A1(net_606) );
INV_X4 inst_14369 ( .A(net_6895), .ZN(net_6298) );
NAND2_X2 inst_9748 ( .ZN(net_19735), .A1(net_9518), .A2(net_8382) );
OAI21_X2 inst_1660 ( .A(net_16743), .ZN(net_15785), .B2(net_14779), .B1(net_14676) );
NAND2_X2 inst_10113 ( .A1(net_9490), .ZN(net_8425), .A2(net_6319) );
CLKBUF_X2 inst_22647 ( .A(net_21591), .Z(net_22519) );
NOR2_X2 inst_4375 ( .ZN(net_11737), .A1(net_5635), .A2(net_5403) );
CLKBUF_X2 inst_22415 ( .A(net_22286), .Z(net_22287) );
INV_X4 inst_13416 ( .ZN(net_10278), .A(net_8789) );
XNOR2_X2 inst_517 ( .ZN(net_5707), .B(net_5706), .A(net_1865) );
AOI21_X2 inst_20544 ( .ZN(net_19978), .B1(net_14634), .A(net_13428), .B2(net_12534) );
OAI22_X2 inst_1261 ( .B1(net_21152), .ZN(net_17405), .A1(net_17404), .A2(net_16949), .B2(net_16948) );
NAND4_X2 inst_5368 ( .ZN(net_19509), .A4(net_14010), .A1(net_12423), .A3(net_11736), .A2(net_11498) );
AOI22_X2 inst_19987 ( .ZN(net_15140), .B1(net_14622), .A2(net_13331), .A1(net_12675), .B2(net_7377) );
NAND2_X2 inst_8967 ( .ZN(net_14610), .A2(net_13268), .A1(net_12813) );
NAND2_X2 inst_10220 ( .ZN(net_9599), .A1(net_6318), .A2(net_6262) );
NAND3_X2 inst_6130 ( .ZN(net_19277), .A1(net_13676), .A3(net_6342), .A2(net_3783) );
NAND4_X2 inst_5382 ( .ZN(net_15050), .A3(net_13920), .A2(net_12979), .A4(net_12507), .A1(net_9697) );
INV_X4 inst_14661 ( .ZN(net_5627), .A(net_4353) );
XNOR2_X2 inst_310 ( .ZN(net_17088), .A(net_16870), .B(net_16268) );
INV_X2 inst_18875 ( .ZN(net_6212), .A(net_6211) );
INV_X4 inst_17982 ( .A(net_20884), .ZN(net_1719) );
NAND2_X2 inst_8900 ( .ZN(net_15100), .A1(net_15099), .A2(net_13948) );
AOI21_X4 inst_20119 ( .B2(net_19526), .B1(net_19525), .A(net_16359), .ZN(net_16241) );
NOR3_X2 inst_2688 ( .ZN(net_14354), .A3(net_14291), .A1(net_12606), .A2(net_9791) );
NAND3_X2 inst_6172 ( .ZN(net_13604), .A1(net_12338), .A3(net_10534), .A2(net_10174) );
NAND3_X4 inst_5592 ( .ZN(net_15134), .A2(net_14783), .A3(net_13381), .A1(net_6935) );
INV_X4 inst_18091 ( .A(net_21037), .ZN(net_456) );
AND2_X4 inst_21210 ( .A1(net_14962), .A2(net_7065), .ZN(net_6731) );
OAI21_X2 inst_2351 ( .B1(net_7075), .A(net_5252), .ZN(net_3718), .B2(net_2410) );
NAND2_X2 inst_8067 ( .ZN(net_18184), .A2(net_18183), .A1(net_18182) );
INV_X8 inst_12302 ( .ZN(net_1071), .A(net_503) );
NOR2_X2 inst_5125 ( .A1(net_879), .A2(net_646), .ZN(net_274) );
OAI21_X2 inst_1853 ( .ZN(net_13998), .B1(net_12954), .B2(net_11283), .A(net_10325) );
AOI22_X2 inst_19968 ( .ZN(net_20812), .A1(net_19786), .B1(net_18900), .B2(net_14264), .A2(net_1402) );
NAND2_X4 inst_7576 ( .ZN(net_2559), .A1(net_1607), .A2(net_63) );
CLKBUF_X2 inst_22754 ( .A(net_22625), .Z(net_22626) );
NAND2_X2 inst_11101 ( .ZN(net_4335), .A2(net_4334), .A1(net_154) );
XNOR2_X2 inst_264 ( .A(net_19420), .ZN(net_17256), .B(net_16644) );
CLKBUF_X2 inst_22928 ( .A(net_22799), .Z(net_22800) );
INV_X4 inst_15834 ( .ZN(net_2869), .A(net_1858) );
NOR2_X2 inst_3710 ( .A1(net_13495), .ZN(net_11026), .A2(net_11025) );
CLKBUF_X2 inst_22523 ( .A(net_22394), .Z(net_22395) );
OAI22_X2 inst_1260 ( .ZN(net_17417), .A2(net_17416), .B2(net_17415), .A1(net_14825), .B1(net_13594) );
NAND3_X2 inst_6490 ( .ZN(net_11169), .A2(net_11168), .A3(net_11167), .A1(net_6033) );
CLKBUF_X2 inst_22435 ( .A(net_22287), .Z(net_22307) );
NAND2_X2 inst_10190 ( .ZN(net_10343), .A1(net_6736), .A2(net_5515) );
NOR2_X4 inst_3332 ( .ZN(net_841), .A2(net_646), .A1(net_234) );
NAND2_X2 inst_7885 ( .ZN(net_18515), .A2(net_18447), .A1(net_17950) );
NOR2_X2 inst_4898 ( .ZN(net_2015), .A1(net_1241), .A2(net_621) );
INV_X4 inst_17126 ( .ZN(net_2171), .A(net_773) );
NOR3_X2 inst_2717 ( .ZN(net_13425), .A2(net_11220), .A1(net_10307), .A3(net_8964) );
AND2_X4 inst_21219 ( .ZN(net_6870), .A2(net_5305), .A1(net_573) );
INV_X4 inst_13836 ( .ZN(net_10929), .A(net_8759) );
NOR2_X2 inst_4176 ( .A1(net_12620), .ZN(net_6824), .A2(net_6823) );
XNOR2_X2 inst_129 ( .A(net_18299), .ZN(net_18262), .B(net_1873) );
NOR3_X2 inst_2740 ( .ZN(net_12756), .A1(net_10203), .A3(net_8075), .A2(net_4823) );
OAI21_X2 inst_1754 ( .ZN(net_14794), .A(net_14793), .B2(net_13281), .B1(net_6964) );
INV_X4 inst_16777 ( .ZN(net_1024), .A(net_1023) );
NAND2_X4 inst_6974 ( .A1(net_19454), .ZN(net_19243), .A2(net_17242) );
INV_X4 inst_12955 ( .A(net_16748), .ZN(net_16539) );
NAND2_X2 inst_7789 ( .A2(net_20209), .ZN(net_18717), .A1(net_17498) );
NOR3_X2 inst_2727 ( .ZN(net_13247), .A2(net_13246), .A1(net_10596), .A3(net_5172) );
NAND2_X2 inst_7974 ( .ZN(net_18438), .A1(net_18254), .A2(net_18207) );
INV_X16 inst_19734 ( .A(net_1730), .ZN(net_1022) );
NAND2_X2 inst_8848 ( .A2(net_20035), .A1(net_20034), .ZN(net_15396) );
NAND3_X2 inst_6305 ( .ZN(net_12792), .A3(net_12791), .A2(net_10867), .A1(net_5523) );
INV_X2 inst_18664 ( .ZN(net_9179), .A(net_9178) );
SDFF_X2 inst_777 ( .Q(net_20930), .SE(net_18862), .SI(net_18402), .D(net_575), .CK(net_21426) );
NAND3_X2 inst_6164 ( .A3(net_20698), .ZN(net_20449), .A2(net_12968), .A1(net_12694) );
INV_X4 inst_14175 ( .ZN(net_7469), .A(net_5994) );
NOR2_X2 inst_5016 ( .A2(net_4030), .ZN(net_1243), .A1(net_846) );
INV_X4 inst_17872 ( .ZN(net_19897), .A(net_1733) );
INV_X4 inst_17199 ( .ZN(net_3418), .A(net_110) );
NAND2_X2 inst_10276 ( .ZN(net_19887), .A2(net_7957), .A1(net_5951) );
NAND2_X4 inst_7000 ( .ZN(net_17500), .A1(net_16725), .A2(net_16570) );
AOI21_X2 inst_20852 ( .B1(net_10108), .ZN(net_9071), .A(net_7484), .B2(net_5303) );
INV_X4 inst_15975 ( .ZN(net_14463), .A(net_12522) );
NAND2_X2 inst_9983 ( .ZN(net_8855), .A1(net_8854), .A2(net_6493) );
NOR2_X2 inst_3724 ( .A1(net_13353), .ZN(net_10923), .A2(net_10922) );
AOI21_X4 inst_20249 ( .ZN(net_9977), .A(net_6692), .B2(net_4740), .B1(net_3768) );
INV_X4 inst_14393 ( .ZN(net_10716), .A(net_7313) );
INV_X4 inst_14138 ( .ZN(net_9384), .A(net_6085) );
INV_X2 inst_19731 ( .A(net_20807), .ZN(net_20806) );
INV_X4 inst_15943 ( .ZN(net_2020), .A(net_783) );
INV_X4 inst_16930 ( .ZN(net_11751), .A(net_8676) );
NAND2_X2 inst_10509 ( .ZN(net_11790), .A1(net_11296), .A2(net_5046) );
NAND3_X2 inst_6146 ( .ZN(net_13684), .A2(net_12322), .A1(net_7088), .A3(net_5354) );
INV_X4 inst_13978 ( .ZN(net_6623), .A(net_6622) );
NAND2_X2 inst_11909 ( .ZN(net_2428), .A1(net_2283), .A2(net_1697) );
NOR2_X2 inst_4965 ( .A1(net_2744), .ZN(net_1598), .A2(net_1311) );
INV_X4 inst_13039 ( .A(net_16576), .ZN(net_16410) );
NAND2_X2 inst_11158 ( .ZN(net_7021), .A2(net_4123), .A1(net_809) );
OAI21_X2 inst_2354 ( .ZN(net_2963), .B1(net_2769), .B2(net_2489), .A(net_2389) );
NAND2_X2 inst_9447 ( .A1(net_12160), .ZN(net_11531), .A2(net_11530) );
NAND2_X2 inst_8735 ( .A1(net_19871), .A2(net_16368), .ZN(net_16027) );
NAND2_X2 inst_10729 ( .ZN(net_5828), .A2(net_4482), .A1(net_4392) );
INV_X4 inst_13315 ( .ZN(net_11611), .A(net_11610) );
INV_X4 inst_15514 ( .A(net_3334), .ZN(net_2406) );
INV_X4 inst_15872 ( .ZN(net_16051), .A(net_15706) );
INV_X4 inst_14965 ( .ZN(net_3434), .A(net_3433) );
INV_X8 inst_12316 ( .ZN(net_2497), .A(net_752) );
NAND2_X2 inst_10883 ( .ZN(net_11794), .A1(net_6318), .A2(net_5278) );
NOR2_X2 inst_3869 ( .A1(net_11368), .ZN(net_9371), .A2(net_7871) );
NOR2_X2 inst_3488 ( .ZN(net_14275), .A1(net_14274), .A2(net_12623) );
INV_X4 inst_15801 ( .A(net_13512), .ZN(net_12888) );
INV_X4 inst_12689 ( .ZN(net_17669), .A(net_17668) );
NOR2_X2 inst_4563 ( .ZN(net_5021), .A1(net_3308), .A2(net_1848) );
CLKBUF_X2 inst_22053 ( .A(net_21924), .Z(net_21925) );
INV_X2 inst_19401 ( .A(net_2970), .ZN(net_2024) );
INV_X4 inst_17813 ( .A(net_265), .ZN(net_159) );
AOI21_X2 inst_20371 ( .ZN(net_15615), .A(net_15463), .B2(net_14275), .B1(net_12358) );
NAND4_X2 inst_5504 ( .ZN(net_11791), .A4(net_11790), .A2(net_11725), .A3(net_11724), .A1(net_9878) );
CLKBUF_X2 inst_21429 ( .A(net_21300), .Z(net_21301) );
INV_X2 inst_19422 ( .ZN(net_1832), .A(net_1831) );
INV_X2 inst_19134 ( .ZN(net_4160), .A(net_4159) );
NAND2_X4 inst_7453 ( .ZN(net_4381), .A1(net_4158), .A2(net_1626) );
CLKBUF_X2 inst_21657 ( .A(net_21270), .Z(net_21529) );
OAI21_X2 inst_1519 ( .ZN(net_18429), .A(net_18314), .B1(net_18313), .B2(net_18312) );
NAND2_X4 inst_7243 ( .ZN(net_10452), .A1(net_6997), .A2(net_874) );
AND2_X2 inst_21358 ( .ZN(net_2595), .A1(net_1376), .A2(net_187) );
NAND2_X2 inst_9936 ( .ZN(net_9147), .A1(net_9146), .A2(net_7102) );
NAND2_X2 inst_8461 ( .A1(net_17162), .ZN(net_17051), .A2(net_16614) );
NOR2_X2 inst_4989 ( .A1(net_2388), .ZN(net_1430), .A2(net_1429) );
CLKBUF_X2 inst_22228 ( .A(net_22071), .Z(net_22100) );
INV_X4 inst_16617 ( .ZN(net_2606), .A(net_1118) );
CLKBUF_X2 inst_22531 ( .A(net_22402), .Z(net_22403) );
INV_X2 inst_18601 ( .ZN(net_9816), .A(net_9815) );
NOR2_X2 inst_4324 ( .ZN(net_5861), .A1(net_3635), .A2(net_3608) );
NAND3_X2 inst_5746 ( .ZN(net_16016), .A3(net_15429), .A1(net_14156), .A2(net_12917) );
NAND3_X4 inst_5597 ( .ZN(net_14746), .A2(net_14745), .A3(net_12327), .A1(net_9643) );
INV_X4 inst_12705 ( .ZN(net_17592), .A(net_17591) );
CLKBUF_X2 inst_21413 ( .A(net_21264), .Z(net_21285) );
NAND2_X2 inst_8531 ( .A1(net_17006), .ZN(net_16865), .A2(net_16864) );
INV_X8 inst_12244 ( .ZN(net_5042), .A(net_2800) );
OAI21_X4 inst_1491 ( .ZN(net_19075), .B1(net_11504), .B2(net_10928), .A(net_368) );
NAND2_X2 inst_8070 ( .ZN(net_18167), .A2(net_18166), .A1(net_16792) );
CLKBUF_X2 inst_21619 ( .A(net_21490), .Z(net_21491) );
INV_X4 inst_12747 ( .ZN(net_17420), .A(net_17419) );
INV_X4 inst_15446 ( .ZN(net_9487), .A(net_9458) );
AOI21_X2 inst_20945 ( .ZN(net_6389), .A(net_4119), .B2(net_3673), .B1(net_2788) );
NOR3_X2 inst_2676 ( .ZN(net_14773), .A3(net_13151), .A1(net_11402), .A2(net_7217) );
CLKBUF_X2 inst_21998 ( .A(net_21772), .Z(net_21870) );
NAND2_X2 inst_8566 ( .ZN(net_20405), .A1(net_16743), .A2(net_16742) );
XNOR2_X2 inst_154 ( .ZN(net_17974), .B(net_17973), .A(net_17850) );
AOI21_X2 inst_20435 ( .ZN(net_15159), .B1(net_15158), .B2(net_13877), .A(net_13564) );
NAND2_X2 inst_9794 ( .A1(net_14493), .ZN(net_11073), .A2(net_9709) );
NAND3_X2 inst_6057 ( .ZN(net_14218), .A3(net_13427), .A2(net_10194), .A1(net_9598) );
INV_X8 inst_12325 ( .A(net_2629), .ZN(net_1056) );
NAND2_X2 inst_10078 ( .A1(net_8793), .ZN(net_8646), .A2(net_8645) );
INV_X4 inst_13427 ( .ZN(net_9899), .A(net_8468) );
NAND2_X2 inst_10368 ( .A1(net_11482), .ZN(net_7403), .A2(net_5830) );
INV_X2 inst_19441 ( .A(net_15790), .ZN(net_1693) );
CLKBUF_X2 inst_21541 ( .A(net_21412), .Z(net_21413) );
NOR2_X2 inst_4240 ( .A1(net_11045), .ZN(net_6559), .A2(net_6558) );
NAND2_X2 inst_10813 ( .A1(net_11148), .A2(net_5575), .ZN(net_5523) );
AND2_X4 inst_21160 ( .ZN(net_13804), .A1(net_13803), .A2(net_13802) );
INV_X2 inst_19705 ( .ZN(net_20572), .A(net_20568) );
INV_X4 inst_12570 ( .ZN(net_18301), .A(net_18263) );
OAI21_X2 inst_1790 ( .ZN(net_14644), .A(net_14643), .B1(net_12481), .B2(net_11758) );
NAND3_X2 inst_6621 ( .A2(net_14145), .ZN(net_9057), .A1(net_9056), .A3(net_9055) );
CLKBUF_X2 inst_22161 ( .A(net_21707), .Z(net_22033) );
NAND2_X2 inst_10989 ( .ZN(net_9911), .A1(net_5291), .A2(net_1214) );
NAND3_X2 inst_6355 ( .ZN(net_12094), .A3(net_12093), .A1(net_10595), .A2(net_8256) );
CLKBUF_X2 inst_21467 ( .A(net_21338), .Z(net_21339) );
INV_X4 inst_13982 ( .ZN(net_14456), .A(net_6607) );
INV_X4 inst_18155 ( .A(net_20944), .ZN(net_16260) );
XNOR2_X2 inst_243 ( .B(net_21210), .ZN(net_17325), .A(net_16854) );
OAI21_X4 inst_1378 ( .B1(net_19989), .ZN(net_16650), .B2(net_16644), .A(net_16290) );
INV_X4 inst_14156 ( .ZN(net_11195), .A(net_3874) );
INV_X4 inst_14049 ( .ZN(net_7613), .A(net_6253) );
INV_X2 inst_18521 ( .ZN(net_19226), .A(net_10081) );
INV_X4 inst_16894 ( .ZN(net_2841), .A(net_1044) );
INV_X2 inst_19245 ( .ZN(net_6698), .A(net_4032) );
INV_X4 inst_15738 ( .ZN(net_12877), .A(net_11182) );
NAND2_X2 inst_8189 ( .ZN(net_17946), .A1(net_17792), .A2(net_17691) );
CLKBUF_X2 inst_21551 ( .A(net_21422), .Z(net_21423) );
NAND2_X4 inst_7281 ( .ZN(net_13323), .A2(net_5097), .A1(net_4435) );
INV_X4 inst_16491 ( .ZN(net_10188), .A(net_1197) );
NAND3_X2 inst_6704 ( .ZN(net_7347), .A3(net_7346), .A2(net_6829), .A1(net_4365) );
CLKBUF_X2 inst_22120 ( .A(net_21991), .Z(net_21992) );
NAND2_X2 inst_9501 ( .A1(net_11682), .ZN(net_11351), .A2(net_8237) );
CLKBUF_X2 inst_22709 ( .A(net_22580), .Z(net_22581) );
INV_X4 inst_16709 ( .ZN(net_4952), .A(net_1786) );
NAND2_X2 inst_8799 ( .ZN(net_15671), .A2(net_15159), .A1(net_13786) );
CLKBUF_X2 inst_21377 ( .A(net_21248), .Z(net_21249) );
NOR2_X4 inst_3229 ( .A2(net_20494), .ZN(net_7149), .A1(net_4014) );
NOR2_X2 inst_4135 ( .ZN(net_6943), .A2(net_6942), .A1(net_4005) );
INV_X4 inst_14459 ( .ZN(net_8204), .A(net_4944) );
OAI21_X4 inst_1369 ( .ZN(net_17121), .A(net_16795), .B1(net_16794), .B2(net_16451) );
NOR2_X2 inst_3988 ( .ZN(net_20383), .A1(net_8311), .A2(net_8310) );
NAND3_X2 inst_6548 ( .ZN(net_10535), .A3(net_10534), .A2(net_8225), .A1(net_5998) );
INV_X2 inst_18548 ( .ZN(net_10940), .A(net_10939) );
INV_X4 inst_15172 ( .ZN(net_3979), .A(net_3012) );
INV_X4 inst_15280 ( .A(net_3759), .ZN(net_2740) );
OAI211_X2 inst_2561 ( .ZN(net_9910), .C1(net_9909), .A(net_7530), .C2(net_7313), .B(net_3923) );
NAND2_X2 inst_7767 ( .ZN(net_18747), .A2(net_18741), .A1(net_17068) );
NAND2_X2 inst_8495 ( .ZN(net_16943), .A1(net_16597), .A2(net_16461) );
NAND2_X2 inst_8974 ( .ZN(net_14516), .A1(net_14515), .A2(net_13004) );
NAND2_X2 inst_8163 ( .ZN(net_17971), .A1(net_17970), .A2(net_17969) );
INV_X4 inst_13669 ( .ZN(net_9593), .A(net_8060) );
INV_X4 inst_13257 ( .ZN(net_12717), .A(net_11658) );
NAND2_X2 inst_9583 ( .ZN(net_10925), .A2(net_10924), .A1(net_10141) );
NOR2_X2 inst_4226 ( .ZN(net_6605), .A1(net_6604), .A2(net_6603) );
INV_X4 inst_16011 ( .ZN(net_3192), .A(net_1666) );
INV_X4 inst_15847 ( .ZN(net_3719), .A(net_1834) );
NAND2_X2 inst_9222 ( .ZN(net_12971), .A2(net_12970), .A1(net_7403) );
INV_X4 inst_12843 ( .ZN(net_17084), .A(net_17083) );
NAND3_X2 inst_5795 ( .ZN(net_15723), .A1(net_15333), .A2(net_15115), .A3(net_14993) );
NAND2_X2 inst_12112 ( .A1(net_20938), .A2(net_955), .ZN(net_549) );
OAI21_X2 inst_2238 ( .A(net_13198), .ZN(net_7720), .B1(net_6376), .B2(net_6153) );
NAND4_X4 inst_5207 ( .A4(net_20729), .A1(net_20728), .A3(net_19494), .ZN(net_16569), .A2(net_13872) );
NOR2_X2 inst_4543 ( .ZN(net_5046), .A2(net_3986), .A1(net_526) );
NOR2_X2 inst_5072 ( .ZN(net_1282), .A2(net_926), .A1(net_63) );
INV_X4 inst_14347 ( .ZN(net_5812), .A(net_5329) );
NOR2_X4 inst_3151 ( .ZN(net_6641), .A1(net_4293), .A2(net_1544) );
INV_X4 inst_15312 ( .ZN(net_3419), .A(net_2648) );
AND3_X4 inst_21123 ( .ZN(net_12515), .A3(net_11971), .A2(net_8399), .A1(net_7789) );
INV_X4 inst_13073 ( .ZN(net_16247), .A(net_16177) );
NAND2_X2 inst_10764 ( .A1(net_9541), .ZN(net_5645), .A2(net_5644) );
NOR2_X2 inst_4436 ( .ZN(net_12771), .A1(net_4850), .A2(net_4849) );
NAND2_X2 inst_8180 ( .ZN(net_17932), .A1(net_17926), .A2(net_17914) );
INV_X4 inst_16307 ( .ZN(net_4259), .A(net_2050) );
INV_X4 inst_13042 ( .ZN(net_16401), .A(net_16377) );
INV_X4 inst_14732 ( .ZN(net_12406), .A(net_4116) );
NAND3_X2 inst_5801 ( .ZN(net_20425), .A3(net_19514), .A1(net_19513), .A2(net_8834) );
NAND2_X2 inst_9363 ( .ZN(net_12136), .A1(net_11430), .A2(net_9904) );
NAND3_X2 inst_6674 ( .ZN(net_7759), .A1(net_7743), .A2(net_5908), .A3(net_5054) );
OAI21_X2 inst_2259 ( .ZN(net_18931), .A(net_12041), .B2(net_11194), .B1(net_2604) );
INV_X4 inst_12935 ( .ZN(net_17242), .A(net_17126) );
NAND3_X2 inst_6196 ( .ZN(net_13313), .A1(net_10895), .A3(net_9877), .A2(net_2752) );
INV_X4 inst_14314 ( .A(net_7849), .ZN(net_5477) );
AOI21_X2 inst_20805 ( .B2(net_11124), .ZN(net_10342), .A(net_4931), .B1(net_3631) );
NAND3_X2 inst_6462 ( .ZN(net_11371), .A3(net_9798), .A2(net_7474), .A1(net_7111) );
INV_X4 inst_14101 ( .A(net_12908), .ZN(net_9474) );
INV_X4 inst_12824 ( .ZN(net_17164), .A(net_17163) );
NAND2_X2 inst_11915 ( .ZN(net_3029), .A2(net_1787), .A1(net_765) );
INV_X4 inst_18232 ( .A(net_20924), .ZN(net_61) );
INV_X8 inst_12280 ( .A(net_1764), .ZN(net_1586) );
NAND2_X2 inst_11072 ( .ZN(net_4483), .A1(net_4482), .A2(net_3119) );
NAND3_X2 inst_6428 ( .ZN(net_11926), .A2(net_11925), .A3(net_11924), .A1(net_3655) );
CLKBUF_X2 inst_21395 ( .A(net_21266), .Z(net_21267) );
INV_X4 inst_14221 ( .A(net_6197), .ZN(net_5846) );
NAND2_X4 inst_7312 ( .A1(net_20534), .ZN(net_8995), .A2(net_5370) );
INV_X2 inst_19049 ( .ZN(net_4743), .A(net_4742) );
INV_X4 inst_17731 ( .ZN(net_6207), .A(net_184) );
INV_X4 inst_17409 ( .ZN(net_15087), .A(net_512) );
CLKBUF_X2 inst_21460 ( .A(net_21303), .Z(net_21332) );
NAND2_X2 inst_10749 ( .ZN(net_5708), .A2(net_5462), .A1(net_1229) );
INV_X2 inst_18479 ( .ZN(net_12619), .A(net_12618) );
INV_X4 inst_12737 ( .ZN(net_17541), .A(net_17446) );
CLKBUF_X2 inst_22272 ( .A(net_22143), .Z(net_22144) );
INV_X4 inst_17499 ( .ZN(net_2872), .A(net_250) );
XNOR2_X2 inst_524 ( .B(net_16700), .ZN(net_3755), .A(net_2472) );
INV_X4 inst_15568 ( .A(net_3235), .ZN(net_2288) );
INV_X4 inst_13027 ( .ZN(net_16584), .A(net_16465) );
XNOR2_X2 inst_104 ( .ZN(net_18529), .B(net_18470), .A(net_18422) );
INV_X4 inst_14986 ( .A(net_12339), .ZN(net_8169) );
OAI21_X2 inst_2331 ( .ZN(net_5247), .B1(net_5246), .B2(net_3879), .A(net_3078) );
NAND3_X2 inst_6096 ( .ZN(net_19126), .A3(net_13919), .A1(net_11424), .A2(net_9524) );
NAND2_X2 inst_9752 ( .ZN(net_10049), .A1(net_10048), .A2(net_6933) );
OAI211_X4 inst_2377 ( .A(net_19214), .C2(net_19195), .C1(net_19194), .ZN(net_16170), .B(net_14596) );
OAI211_X2 inst_2522 ( .B(net_11959), .ZN(net_11862), .A(net_11861), .C1(net_11860), .C2(net_1561) );
INV_X4 inst_13793 ( .ZN(net_13494), .A(net_7562) );
NAND2_X2 inst_11910 ( .ZN(net_3294), .A2(net_1636), .A1(net_222) );
NAND2_X2 inst_10673 ( .ZN(net_10582), .A2(net_2537), .A1(net_842) );
INV_X2 inst_18530 ( .A(net_11487), .ZN(net_11085) );
NAND2_X2 inst_7967 ( .ZN(net_18366), .A2(net_18365), .A1(net_17386) );
NAND4_X4 inst_5216 ( .A2(net_20623), .A1(net_20622), .A3(net_20278), .A4(net_19176), .ZN(net_16379) );
NAND4_X2 inst_5257 ( .A4(net_19503), .A1(net_19502), .ZN(net_16337), .A2(net_16113), .A3(net_15985) );
NAND2_X2 inst_8011 ( .ZN(net_18296), .A2(net_18295), .A1(net_17271) );
NAND2_X2 inst_11226 ( .ZN(net_10629), .A2(net_3954), .A1(net_3187) );
SDFF_X2 inst_708 ( .Q(net_20956), .SE(net_18858), .SI(net_18826), .D(net_468), .CK(net_22069) );
OAI221_X2 inst_1346 ( .C1(net_14865), .ZN(net_13148), .A(net_13147), .B2(net_13146), .B1(net_12763), .C2(net_7721) );
NOR2_X2 inst_3523 ( .ZN(net_13722), .A2(net_11573), .A1(net_8756) );
INV_X2 inst_19673 ( .A(net_20495), .ZN(net_20491) );
NAND3_X2 inst_5811 ( .ZN(net_15647), .A3(net_14516), .A1(net_11646), .A2(net_10397) );
NOR2_X2 inst_3510 ( .ZN(net_13902), .A2(net_12026), .A1(net_9427) );
NOR2_X2 inst_5108 ( .A2(net_915), .ZN(net_755), .A1(net_606) );
NAND3_X2 inst_6723 ( .ZN(net_6506), .A2(net_6489), .A1(net_5652), .A3(net_5556) );
OR2_X4 inst_1071 ( .A1(net_13544), .ZN(net_12174), .A2(net_10565) );
NOR2_X2 inst_4277 ( .A1(net_9667), .A2(net_6229), .ZN(net_6117) );
NAND3_X2 inst_6421 ( .ZN(net_11942), .A3(net_10237), .A1(net_7658), .A2(net_6160) );
NAND4_X2 inst_5291 ( .A4(net_19240), .A1(net_19239), .ZN(net_15934), .A2(net_13932), .A3(net_8024) );
DFF_X1 inst_19801 ( .D(net_18194), .CK(net_21998), .Q(x1044) );
INV_X4 inst_17476 ( .ZN(net_3830), .A(net_1327) );
NAND2_X2 inst_11352 ( .ZN(net_3642), .A1(net_3641), .A2(net_3640) );
INV_X4 inst_17783 ( .ZN(net_365), .A(net_242) );
INV_X4 inst_13211 ( .ZN(net_13665), .A(net_12882) );
CLKBUF_X2 inst_21483 ( .A(net_21264), .Z(net_21355) );
OAI21_X2 inst_1994 ( .ZN(net_11969), .A(net_11968), .B1(net_11535), .B2(net_8704) );
INV_X4 inst_13132 ( .ZN(net_15266), .A(net_14875) );
INV_X4 inst_15952 ( .A(net_7244), .ZN(net_2212) );
NAND2_X2 inst_9192 ( .ZN(net_13116), .A2(net_11227), .A1(net_10521) );
NAND4_X2 inst_5298 ( .A4(net_19261), .A1(net_19260), .ZN(net_19219), .A2(net_15287), .A3(net_13027) );
CLKBUF_X2 inst_21915 ( .A(net_21786), .Z(net_21787) );
INV_X4 inst_14436 ( .ZN(net_6165), .A(net_5005) );
NAND2_X2 inst_10108 ( .A1(net_11536), .ZN(net_8432), .A2(net_8431) );
INV_X4 inst_15179 ( .ZN(net_3798), .A(net_3362) );
INV_X4 inst_14935 ( .ZN(net_20446), .A(net_4967) );
INV_X4 inst_14744 ( .ZN(net_10630), .A(net_3137) );
INV_X4 inst_13191 ( .ZN(net_14170), .A(net_13513) );
NAND2_X2 inst_8940 ( .ZN(net_14761), .A2(net_14143), .A1(net_13191) );
OAI21_X2 inst_2162 ( .ZN(net_9089), .A(net_4642), .B2(net_4472), .B1(net_3429) );
CLKBUF_X2 inst_21691 ( .A(net_21562), .Z(net_21563) );
XNOR2_X2 inst_392 ( .B(net_21155), .A(net_16769), .ZN(net_16768) );
XNOR2_X2 inst_120 ( .ZN(net_18406), .B(net_18405), .A(net_18234) );
INV_X4 inst_14533 ( .ZN(net_7449), .A(net_3714) );
NAND2_X2 inst_7747 ( .ZN(net_18781), .A2(net_18733), .A1(net_18707) );
NAND2_X2 inst_10917 ( .ZN(net_13260), .A1(net_5342), .A2(net_3849) );
INV_X4 inst_17575 ( .ZN(net_14628), .A(net_855) );
OAI21_X2 inst_1514 ( .ZN(net_18570), .B2(net_18498), .B1(net_18025), .A(net_7391) );
NAND2_X2 inst_8361 ( .ZN(net_20411), .A2(net_17148), .A1(net_17016) );
XNOR2_X2 inst_567 ( .ZN(net_645), .A(net_644), .B(net_643) );
NOR2_X4 inst_3200 ( .ZN(net_5553), .A2(net_3056), .A1(net_3025) );
NAND2_X2 inst_9134 ( .ZN(net_20837), .A1(net_13514), .A2(net_10778) );
OAI21_X2 inst_1601 ( .A(net_21228), .ZN(net_16174), .B2(net_15775), .B1(net_14290) );
NOR2_X2 inst_3526 ( .ZN(net_18935), .A2(net_11551), .A1(net_11545) );
NAND2_X2 inst_9010 ( .ZN(net_14268), .A2(net_13540), .A1(net_4685) );
INV_X2 inst_18501 ( .A(net_14164), .ZN(net_12148) );
NAND2_X1 inst_12147 ( .A2(net_16619), .ZN(net_16463), .A1(net_16462) );
AOI21_X4 inst_20256 ( .ZN(net_20419), .A(net_4079), .B1(net_3681), .B2(net_2492) );
NAND2_X2 inst_10910 ( .ZN(net_10185), .A1(net_7121), .A2(net_5371) );
NAND2_X4 inst_6916 ( .A2(net_19189), .A1(net_19188), .ZN(net_17831) );
INV_X4 inst_13999 ( .ZN(net_6382), .A(net_5245) );
NAND2_X2 inst_9876 ( .ZN(net_9454), .A1(net_7801), .A2(net_7420) );
INV_X2 inst_18365 ( .ZN(net_17947), .A(net_17946) );
NOR2_X2 inst_4123 ( .ZN(net_7032), .A2(net_7031), .A1(net_4114) );
OAI21_X2 inst_1751 ( .A(net_15454), .ZN(net_14800), .B2(net_13336), .B1(net_5888) );
NAND2_X4 inst_6919 ( .A2(net_19313), .A1(net_19312), .ZN(net_17809) );
NAND2_X2 inst_7766 ( .ZN(net_18748), .A2(net_18745), .A1(net_18661) );
INV_X4 inst_14490 ( .A(net_4848), .ZN(net_4847) );
INV_X2 inst_19243 ( .ZN(net_3280), .A(net_3279) );
NAND2_X2 inst_8140 ( .A1(net_20651), .ZN(net_18027), .A2(net_17724) );
INV_X2 inst_18388 ( .A(net_16985), .ZN(net_16638) );
INV_X4 inst_17462 ( .ZN(net_1588), .A(net_157) );
OAI21_X2 inst_2235 ( .A(net_12640), .ZN(net_7763), .B1(net_3458), .B2(net_1907) );
SDFF_X2 inst_779 ( .Q(net_20911), .SE(net_18864), .SI(net_18403), .D(net_11864), .CK(net_22686) );
NAND2_X2 inst_11465 ( .ZN(net_3183), .A2(net_1474), .A1(net_1432) );
INV_X4 inst_16563 ( .ZN(net_5201), .A(net_4783) );
INV_X2 inst_18567 ( .A(net_12960), .ZN(net_10772) );
NAND2_X2 inst_10503 ( .ZN(net_13678), .A1(net_10031), .A2(net_6918) );
NOR2_X2 inst_4131 ( .ZN(net_20646), .A2(net_6931), .A1(net_2346) );
INV_X4 inst_17502 ( .ZN(net_3049), .A(net_117) );
NAND2_X2 inst_9805 ( .ZN(net_19134), .A1(net_10251), .A2(net_9692) );
INV_X4 inst_13591 ( .A(net_9165), .ZN(net_8841) );
INV_X2 inst_18860 ( .ZN(net_6327), .A(net_6326) );
INV_X4 inst_16184 ( .ZN(net_2102), .A(net_1424) );
AOI21_X2 inst_20294 ( .B1(net_19507), .ZN(net_16159), .A(net_14024), .B2(net_13089) );
CLKBUF_X2 inst_22185 ( .A(net_21744), .Z(net_22057) );
NOR2_X2 inst_4228 ( .ZN(net_13654), .A1(net_6592), .A2(net_6591) );
INV_X4 inst_15838 ( .ZN(net_9909), .A(net_8232) );
INV_X4 inst_16647 ( .ZN(net_1956), .A(net_1095) );
NAND2_X2 inst_10808 ( .ZN(net_5530), .A2(net_3895), .A1(net_1028) );
INV_X2 inst_19672 ( .A(net_20495), .ZN(net_20489) );
NAND2_X2 inst_12017 ( .ZN(net_5869), .A1(net_2361), .A2(net_308) );
NOR2_X2 inst_4647 ( .A1(net_6637), .ZN(net_4433), .A2(net_3371) );
AOI21_X2 inst_20923 ( .ZN(net_7175), .B1(net_4222), .B2(net_3876), .A(net_410) );
INV_X2 inst_18758 ( .ZN(net_7639), .A(net_7638) );
NAND2_X4 inst_7408 ( .A2(net_20805), .ZN(net_4851), .A1(net_3645) );
AOI21_X2 inst_20946 ( .B1(net_7975), .ZN(net_6381), .B2(net_4920), .A(net_3021) );
INV_X2 inst_19443 ( .ZN(net_1984), .A(net_1793) );
CLKBUF_X2 inst_21893 ( .A(net_21764), .Z(net_21765) );
NOR2_X2 inst_4709 ( .A1(net_20648), .A2(net_5570), .ZN(net_4114) );
CLKBUF_X2 inst_22380 ( .A(net_22022), .Z(net_22252) );
NAND2_X2 inst_10461 ( .ZN(net_10613), .A2(net_8541), .A1(net_4288) );
INV_X4 inst_15436 ( .ZN(net_3262), .A(net_2503) );
CLKBUF_X2 inst_22644 ( .A(net_22515), .Z(net_22516) );
NAND2_X2 inst_10820 ( .ZN(net_5878), .A1(net_5694), .A2(net_4864) );
CLKBUF_X2 inst_21424 ( .A(net_21295), .Z(net_21296) );
NAND2_X4 inst_7060 ( .ZN(net_20369), .A1(net_19623), .A2(net_16347) );
NOR2_X4 inst_3130 ( .ZN(net_8553), .A1(net_3898), .A2(net_3862) );
NOR2_X2 inst_3347 ( .ZN(net_18033), .A2(net_18012), .A1(net_17282) );
NAND2_X2 inst_9568 ( .ZN(net_19291), .A1(net_15297), .A2(net_7602) );
NAND2_X2 inst_11446 ( .ZN(net_4062), .A2(net_3093), .A1(net_193) );
NOR2_X2 inst_4136 ( .ZN(net_6941), .A2(net_6940), .A1(net_4000) );
NAND4_X2 inst_5341 ( .A4(net_19979), .A1(net_19978), .ZN(net_19197), .A2(net_13966), .A3(net_11216) );
INV_X4 inst_12585 ( .A(net_18138), .ZN(net_18137) );
INV_X4 inst_17573 ( .ZN(net_860), .A(net_180) );
NAND2_X2 inst_9372 ( .ZN(net_12052), .A1(net_10071), .A2(net_8878) );
NAND2_X2 inst_9653 ( .ZN(net_20054), .A1(net_9342), .A2(net_7686) );
NOR2_X2 inst_4985 ( .A2(net_10550), .ZN(net_10170), .A1(net_1471) );
NAND4_X4 inst_5164 ( .ZN(net_20442), .A3(net_18061), .A4(net_18046), .A1(net_16299), .A2(net_7678) );
NAND2_X2 inst_9461 ( .ZN(net_11491), .A2(net_9279), .A1(net_977) );
NAND2_X2 inst_9736 ( .ZN(net_11448), .A1(net_10521), .A2(net_9405) );
INV_X4 inst_15971 ( .ZN(net_13448), .A(net_12620) );
OAI21_X2 inst_1655 ( .ZN(net_15805), .B1(net_15804), .B2(net_14841), .A(net_6531) );
NAND2_X2 inst_10720 ( .A1(net_9309), .ZN(net_5883), .A2(net_3808) );
INV_X4 inst_15174 ( .ZN(net_19632), .A(net_3010) );
CLKBUF_X2 inst_22684 ( .A(net_22555), .Z(net_22556) );
NAND2_X4 inst_7415 ( .ZN(net_7665), .A2(net_3696), .A1(net_3695) );
INV_X4 inst_14165 ( .ZN(net_9368), .A(net_6010) );
NAND2_X2 inst_8731 ( .ZN(net_16058), .A2(net_15764), .A1(net_14045) );
INV_X4 inst_16200 ( .ZN(net_9458), .A(net_1903) );
INV_X4 inst_16594 ( .A(net_11186), .ZN(net_10398) );
NOR2_X2 inst_4847 ( .A1(net_4621), .ZN(net_2336), .A2(net_1538) );
NAND3_X2 inst_6010 ( .ZN(net_19103), .A3(net_12553), .A2(net_11615), .A1(net_10357) );
INV_X4 inst_16318 ( .ZN(net_1319), .A(net_1240) );
INV_X4 inst_15733 ( .ZN(net_4151), .A(net_4018) );
OR3_X2 inst_1066 ( .ZN(net_1534), .A1(net_838), .A2(net_602), .A3(net_225) );
NAND2_X2 inst_9978 ( .ZN(net_8866), .A1(net_8865), .A2(net_6511) );
NAND2_X2 inst_7977 ( .ZN(net_18347), .A2(net_18241), .A1(net_17270) );
INV_X4 inst_16542 ( .ZN(net_7676), .A(net_1005) );
NAND2_X2 inst_10377 ( .A1(net_18025), .ZN(net_7389), .A2(net_633) );
NAND2_X2 inst_12122 ( .A1(net_525), .A2(net_220), .ZN(net_191) );
NOR2_X2 inst_5063 ( .A1(net_10714), .ZN(net_10335), .A2(net_989) );
CLKBUF_X2 inst_22885 ( .A(net_22756), .Z(net_22757) );
INV_X4 inst_15707 ( .A(net_4530), .ZN(net_1992) );
NOR2_X2 inst_4608 ( .A1(net_10875), .A2(net_9024), .ZN(net_3739) );
OAI21_X2 inst_2294 ( .ZN(net_20447), .B2(net_6495), .A(net_4592), .B1(net_303) );
INV_X4 inst_16909 ( .ZN(net_7661), .A(net_4737) );
INV_X4 inst_14321 ( .ZN(net_7250), .A(net_5457) );
INV_X4 inst_12495 ( .ZN(net_18661), .A(net_18645) );
NOR2_X2 inst_4821 ( .A2(net_11845), .A1(net_7950), .ZN(net_3813) );
NAND2_X2 inst_8696 ( .A2(net_20848), .A1(net_19253), .ZN(net_16356) );
NOR2_X2 inst_3931 ( .ZN(net_8726), .A2(net_8681), .A1(net_6259) );
AND2_X2 inst_21302 ( .ZN(net_10095), .A2(net_7673), .A1(net_308) );
INV_X8 inst_12409 ( .ZN(net_329), .A(net_317) );
INV_X4 inst_12682 ( .ZN(net_18439), .A(net_17634) );
NAND2_X4 inst_7239 ( .ZN(net_8829), .A1(net_7008), .A2(net_6849) );
INV_X4 inst_13237 ( .A(net_13566), .ZN(net_13446) );
NAND2_X2 inst_11590 ( .A1(net_6599), .ZN(net_3470), .A2(net_1412) );
NAND2_X2 inst_10785 ( .ZN(net_7302), .A1(net_5611), .A2(net_5591) );
INV_X4 inst_13098 ( .ZN(net_15861), .A(net_15712) );
NAND2_X2 inst_8864 ( .ZN(net_18922), .A2(net_14464), .A1(net_10830) );
XNOR2_X2 inst_158 ( .ZN(net_17949), .B(net_17797), .A(net_17790) );
INV_X4 inst_13529 ( .ZN(net_10796), .A(net_9226) );
CLKBUF_X2 inst_22726 ( .A(net_22182), .Z(net_22598) );
XNOR2_X2 inst_507 ( .B(net_21181), .A(net_15537), .ZN(net_7652) );
AOI21_X2 inst_20806 ( .ZN(net_10321), .A(net_10320), .B2(net_6268), .B1(net_3241) );
NOR2_X2 inst_4289 ( .A2(net_7727), .A1(net_7473), .ZN(net_6036) );
NAND2_X2 inst_10566 ( .A1(net_6867), .A2(net_6740), .ZN(net_6711) );
INV_X4 inst_14365 ( .ZN(net_6309), .A(net_5203) );
SDFF_X2 inst_884 ( .Q(net_21202), .SI(net_16937), .SE(net_125), .CK(net_21652), .D(x6043) );
INV_X8 inst_12311 ( .ZN(net_3713), .A(net_818) );
SDFF_X2 inst_711 ( .Q(net_20920), .SI(net_18805), .SE(net_18585), .D(net_582), .CK(net_22026) );
NAND3_X2 inst_6542 ( .ZN(net_20839), .A2(net_10570), .A1(net_8945), .A3(net_7977) );
INV_X2 inst_19714 ( .A(net_20769), .ZN(net_20768) );
AND3_X4 inst_21124 ( .ZN(net_12502), .A2(net_12501), .A3(net_12500), .A1(net_6565) );
INV_X4 inst_14452 ( .ZN(net_9967), .A(net_4956) );
INV_X2 inst_18847 ( .ZN(net_6653), .A(net_6652) );
INV_X4 inst_14845 ( .ZN(net_11172), .A(net_3846) );
INV_X4 inst_17559 ( .ZN(net_15113), .A(net_14006) );
NAND2_X2 inst_8465 ( .A2(net_20435), .ZN(net_19885), .A1(net_19432) );
NAND2_X2 inst_11213 ( .A1(net_6930), .ZN(net_6888), .A2(net_4009) );
INV_X4 inst_16725 ( .A(net_8924), .ZN(net_1830) );
NOR2_X2 inst_4191 ( .A2(net_11746), .ZN(net_6737), .A1(net_172) );
NOR2_X2 inst_4269 ( .ZN(net_6138), .A2(net_6137), .A1(net_3372) );
INV_X4 inst_14171 ( .ZN(net_9353), .A(net_7790) );
INV_X2 inst_18581 ( .ZN(net_10316), .A(net_10315) );
INV_X2 inst_18486 ( .ZN(net_13568), .A(net_12373) );
NAND2_X2 inst_8559 ( .ZN(net_16749), .A2(net_16748), .A1(net_8098) );
INV_X4 inst_17936 ( .A(net_20945), .ZN(net_788) );
INV_X4 inst_15616 ( .ZN(net_5209), .A(net_2166) );
INV_X4 inst_14534 ( .ZN(net_8997), .A(net_4661) );
OAI21_X2 inst_2263 ( .ZN(net_7162), .B2(net_7161), .A(net_2452), .B1(net_1932) );
NAND3_X4 inst_5608 ( .A3(net_20040), .A1(net_20039), .ZN(net_14119), .A2(net_9066) );
NOR2_X2 inst_4796 ( .A2(net_3239), .ZN(net_2755), .A1(net_1429) );
NOR2_X2 inst_3549 ( .ZN(net_19943), .A1(net_13101), .A2(net_11307) );
CLKBUF_X2 inst_21936 ( .A(net_21807), .Z(net_21808) );
NOR2_X2 inst_3501 ( .A1(net_14986), .ZN(net_14064), .A2(net_11842) );
INV_X4 inst_12602 ( .ZN(net_18124), .A(net_18086) );
NAND2_X2 inst_10035 ( .ZN(net_13234), .A2(net_13065), .A1(net_7087) );
INV_X4 inst_13029 ( .ZN(net_16615), .A(net_16594) );
NOR2_X2 inst_4175 ( .ZN(net_6834), .A2(net_3930), .A1(net_3529) );
NAND2_X4 inst_7076 ( .A2(net_19599), .A1(net_19598), .ZN(net_19477) );
NAND2_X2 inst_8535 ( .A2(net_16870), .ZN(net_16858), .A1(net_16857) );
NAND2_X2 inst_9783 ( .ZN(net_9763), .A1(net_9762), .A2(net_9761) );
INV_X4 inst_14217 ( .A(net_7816), .ZN(net_7484) );
NAND2_X4 inst_6954 ( .A1(net_20438), .A2(net_20067), .ZN(net_17364) );
NAND2_X4 inst_7378 ( .ZN(net_11530), .A1(net_4280), .A2(net_2627) );
NAND2_X2 inst_9416 ( .ZN(net_11648), .A1(net_11647), .A2(net_9480) );
NOR2_X2 inst_4397 ( .A1(net_14622), .ZN(net_5190), .A2(net_5189) );
NOR2_X4 inst_3102 ( .ZN(net_6853), .A2(net_4042), .A1(net_1700) );
NAND2_X4 inst_7392 ( .ZN(net_8933), .A2(net_8304), .A1(net_4180) );
NAND2_X2 inst_10818 ( .ZN(net_5507), .A1(net_5506), .A2(net_2282) );
INV_X4 inst_12847 ( .ZN(net_17078), .A(net_17077) );
NOR2_X2 inst_3860 ( .ZN(net_10939), .A2(net_9824), .A1(net_9575) );
INV_X4 inst_12748 ( .A(net_17544), .ZN(net_17418) );
OAI21_X2 inst_2063 ( .ZN(net_10684), .A(net_10683), .B1(net_5923), .B2(net_4803) );
CLKBUF_X2 inst_21463 ( .A(net_21316), .Z(net_21335) );
INV_X4 inst_14659 ( .ZN(net_9913), .A(net_4356) );
CLKBUF_X2 inst_21924 ( .A(net_21705), .Z(net_21796) );
INV_X4 inst_14917 ( .ZN(net_19881), .A(net_3565) );
NOR2_X2 inst_4801 ( .ZN(net_2734), .A1(net_2733), .A2(net_2732) );
NOR2_X2 inst_3723 ( .ZN(net_12350), .A1(net_10091), .A2(net_9102) );
INV_X4 inst_15978 ( .ZN(net_3133), .A(net_956) );
CLKBUF_X2 inst_21609 ( .A(net_21480), .Z(net_21481) );
NAND2_X2 inst_9346 ( .ZN(net_12206), .A2(net_8910), .A1(net_2266) );
INV_X8 inst_12286 ( .ZN(net_1737), .A(net_914) );
INV_X4 inst_15282 ( .ZN(net_3976), .A(net_2736) );
OAI21_X2 inst_2036 ( .B1(net_11549), .ZN(net_11305), .A(net_10865), .B2(net_10211) );
NOR2_X2 inst_3985 ( .ZN(net_8346), .A1(net_8345), .A2(net_8318) );
NAND4_X2 inst_5386 ( .ZN(net_15017), .A2(net_13475), .A3(net_9955), .A1(net_8401), .A4(net_7132) );
INV_X4 inst_14350 ( .ZN(net_8131), .A(net_5311) );
NAND2_X2 inst_9853 ( .ZN(net_9517), .A1(net_9516), .A2(net_6209) );
NAND2_X2 inst_11107 ( .ZN(net_12829), .A1(net_7153), .A2(net_2572) );
SDFF_X2 inst_868 ( .Q(net_21163), .D(net_17093), .SE(net_263), .CK(net_21462), .SI(x5188) );
OAI21_X2 inst_2049 ( .ZN(net_10853), .A(net_7563), .B2(net_6537), .B1(net_933) );
NAND2_X2 inst_8187 ( .ZN(net_17909), .A2(net_17795), .A1(net_17709) );
NAND2_X2 inst_10747 ( .ZN(net_10792), .A1(net_6570), .A2(net_4311) );
NAND3_X2 inst_6625 ( .ZN(net_9048), .A3(net_6760), .A1(net_5620), .A2(net_3793) );
CLKBUF_X2 inst_22516 ( .A(net_22387), .Z(net_22388) );
XNOR2_X2 inst_201 ( .ZN(net_17663), .A(net_17662), .B(net_17586) );
NAND2_X2 inst_11240 ( .ZN(net_6518), .A2(net_3834), .A1(net_526) );
NOR2_X2 inst_3627 ( .ZN(net_12291), .A2(net_9048), .A1(net_8846) );
XNOR2_X2 inst_304 ( .ZN(net_17096), .A(net_16922), .B(net_7278) );
OR2_X4 inst_1084 ( .ZN(net_20306), .A1(net_14241), .A2(net_5584) );
CLKBUF_X2 inst_21525 ( .A(net_21396), .Z(net_21397) );
NOR2_X2 inst_4157 ( .A1(net_20552), .ZN(net_10493), .A2(net_6926) );
NAND3_X2 inst_5793 ( .ZN(net_15738), .A3(net_15105), .A1(net_13710), .A2(net_13528) );
OAI221_X2 inst_1345 ( .C1(net_13448), .ZN(net_13227), .C2(net_13226), .A(net_13112), .B1(net_11858), .B2(net_7023) );
NAND2_X2 inst_10670 ( .A2(net_8480), .ZN(net_6234), .A1(net_5319) );
INV_X4 inst_12823 ( .ZN(net_17293), .A(net_17184) );
AOI21_X2 inst_20886 ( .ZN(net_7813), .B1(net_4395), .B2(net_2916), .A(net_877) );
NOR2_X4 inst_2947 ( .ZN(net_11627), .A2(net_5450), .A1(net_4883) );
INV_X4 inst_17650 ( .ZN(net_1231), .A(net_270) );
CLKBUF_X2 inst_22925 ( .A(net_22796), .Z(net_22797) );
NOR2_X2 inst_5122 ( .ZN(net_281), .A1(net_91), .A2(net_45) );
INV_X4 inst_12951 ( .ZN(net_16899), .A(net_16544) );
INV_X4 inst_14225 ( .ZN(net_7367), .A(net_5839) );
NAND3_X2 inst_5638 ( .A3(net_19474), .A1(net_19473), .ZN(net_18080), .A2(net_18055) );
NOR2_X2 inst_3608 ( .ZN(net_12424), .A1(net_12315), .A2(net_10034) );
DFF_X1 inst_19877 ( .D(net_17032), .CK(net_21328), .Q(x315) );
NAND2_X4 inst_7306 ( .A1(net_5553), .ZN(net_5473), .A2(net_5472) );
NAND2_X2 inst_10724 ( .A2(net_5910), .ZN(net_5873), .A1(net_5872) );
INV_X4 inst_15235 ( .ZN(net_4632), .A(net_4091) );
SDFF_X2 inst_1016 ( .QN(net_21075), .SE(net_17277), .D(net_568), .CK(net_22172), .SI(x1808) );
INV_X4 inst_18195 ( .A(net_21058), .ZN(net_477) );
SDFF_X2 inst_848 ( .Q(net_21240), .SI(net_17311), .SE(net_125), .CK(net_21550), .D(x6697) );
INV_X4 inst_17480 ( .ZN(net_4079), .A(net_602) );
INV_X4 inst_13394 ( .ZN(net_14164), .A(net_10705) );
OAI211_X2 inst_2479 ( .ZN(net_13505), .C1(net_13504), .B(net_10999), .C2(net_7617), .A(net_5044) );
INV_X4 inst_14333 ( .A(net_6646), .ZN(net_5392) );
CLKBUF_X2 inst_21655 ( .A(net_21526), .Z(net_21527) );
INV_X2 inst_19153 ( .A(net_5437), .ZN(net_5101) );
INV_X4 inst_17814 ( .A(net_493), .ZN(net_196) );
OAI21_X2 inst_1554 ( .B1(net_20433), .B2(net_20067), .ZN(net_17686), .A(net_17364) );
INV_X2 inst_19162 ( .ZN(net_3932), .A(net_3931) );
OAI21_X2 inst_1542 ( .ZN(net_17887), .A(net_17687), .B2(net_17686), .B1(net_17306) );
NOR2_X2 inst_4511 ( .A2(net_20470), .ZN(net_6597), .A1(net_170) );
NAND2_X2 inst_7830 ( .ZN(net_20033), .A2(net_18617), .A1(net_17445) );
NAND2_X2 inst_8849 ( .ZN(net_20113), .A2(net_14716), .A1(net_14173) );
NAND2_X2 inst_11580 ( .A2(net_9247), .ZN(net_5564), .A1(net_3991) );
XNOR2_X2 inst_644 ( .A(net_21131), .ZN(net_10804), .B(net_636) );
AOI21_X2 inst_20478 ( .ZN(net_14944), .A(net_14151), .B2(net_13551), .B1(net_10392) );
INV_X4 inst_15946 ( .ZN(net_2876), .A(net_1713) );
INV_X2 inst_19263 ( .A(net_4330), .ZN(net_3128) );
NOR2_X2 inst_5015 ( .A1(net_5448), .ZN(net_2063), .A2(net_1155) );
CLKBUF_X2 inst_21491 ( .A(net_21362), .Z(net_21363) );
AOI211_X2 inst_21077 ( .C2(net_10812), .ZN(net_6452), .B(net_6451), .A(net_2675), .C1(net_2129) );
INV_X2 inst_19122 ( .A(net_5060), .ZN(net_4624) );
CLKBUF_X2 inst_22035 ( .A(net_21906), .Z(net_21907) );
INV_X4 inst_17229 ( .ZN(net_933), .A(net_103) );
AOI21_X2 inst_20519 ( .B1(net_20061), .ZN(net_14567), .A(net_10085), .B2(net_10082) );
NOR2_X4 inst_2806 ( .ZN(net_17964), .A1(net_17839), .A2(net_17788) );
AOI21_X2 inst_20851 ( .B2(net_13697), .ZN(net_9086), .B1(net_9085), .A(net_8685) );
NOR2_X2 inst_4008 ( .ZN(net_8079), .A2(net_7838), .A1(net_6062) );
NAND3_X2 inst_6736 ( .ZN(net_6473), .A1(net_6133), .A3(net_4793), .A2(net_2786) );
NAND3_X2 inst_6449 ( .ZN(net_11762), .A3(net_10254), .A2(net_8833), .A1(net_2670) );
NAND2_X2 inst_10652 ( .ZN(net_12880), .A1(net_6346), .A2(net_3680) );
CLKBUF_X2 inst_22537 ( .A(net_22408), .Z(net_22409) );
INV_X8 inst_12229 ( .ZN(net_6255), .A(net_3644) );
CLKBUF_X2 inst_22692 ( .A(net_21625), .Z(net_22564) );
NOR2_X2 inst_4896 ( .ZN(net_3362), .A2(net_2045), .A1(net_193) );
AND4_X4 inst_21092 ( .A1(net_20781), .A3(net_12802), .ZN(net_12753), .A4(net_12752), .A2(net_4982) );
INV_X4 inst_14800 ( .A(net_8264), .ZN(net_3985) );
AOI21_X2 inst_20597 ( .ZN(net_13872), .B1(net_13871), .A(net_12176), .B2(net_10646) );
XNOR2_X2 inst_432 ( .A(net_16482), .ZN(net_16478), .B(net_13297) );
XNOR2_X2 inst_282 ( .ZN(net_17167), .A(net_17166), .B(net_13295) );
INV_X4 inst_16827 ( .ZN(net_10947), .A(net_6743) );
INV_X4 inst_15829 ( .ZN(net_3781), .A(net_1440) );
NAND2_X2 inst_8906 ( .ZN(net_15031), .A2(net_14008), .A1(net_11933) );
NAND2_X2 inst_11584 ( .A2(net_4690), .A1(net_2745), .ZN(net_2711) );
NAND2_X2 inst_8428 ( .A1(net_17445), .ZN(net_17179), .A2(net_17178) );
NAND2_X2 inst_9605 ( .ZN(net_10734), .A1(net_10733), .A2(net_10732) );
INV_X4 inst_12533 ( .ZN(net_18383), .A(net_18382) );
NOR2_X4 inst_3171 ( .ZN(net_7059), .A1(net_5537), .A2(net_2206) );
NOR2_X4 inst_3266 ( .ZN(net_3076), .A2(net_2007), .A1(net_2006) );
NAND2_X4 inst_7694 ( .ZN(net_762), .A2(net_598), .A1(net_287) );
NAND2_X2 inst_8725 ( .ZN(net_16100), .A2(net_15835), .A1(net_10051) );
INV_X4 inst_14060 ( .ZN(net_12612), .A(net_7729) );
INV_X4 inst_14910 ( .ZN(net_19399), .A(net_3583) );
INV_X4 inst_12479 ( .ZN(net_18732), .A(net_18692) );
INV_X2 inst_18681 ( .ZN(net_8792), .A(net_7281) );
INV_X4 inst_18106 ( .A(net_21074), .ZN(net_671) );
NAND2_X2 inst_7887 ( .ZN(net_18511), .A2(net_18430), .A1(net_18378) );
NAND2_X2 inst_10296 ( .ZN(net_10116), .A2(net_7900), .A1(net_3678) );
CLKBUF_X2 inst_22413 ( .A(net_21594), .Z(net_22285) );
SDFF_X2 inst_774 ( .Q(net_20869), .SE(net_18847), .SI(net_18472), .D(net_457), .CK(net_21671) );
OAI21_X2 inst_2292 ( .A(net_6976), .ZN(net_6514), .B2(net_2187), .B1(net_1766) );
CLKBUF_X2 inst_22115 ( .A(net_21986), .Z(net_21987) );
CLKBUF_X2 inst_21711 ( .A(net_21427), .Z(net_21583) );
INV_X4 inst_16418 ( .ZN(net_8455), .A(net_2948) );
CLKBUF_X2 inst_22697 ( .A(net_21272), .Z(net_22569) );
INV_X4 inst_14826 ( .ZN(net_4896), .A(net_3902) );
CLKBUF_X2 inst_21398 ( .A(net_21269), .Z(net_21270) );
INV_X4 inst_16871 ( .ZN(net_15104), .A(net_13437) );
NAND4_X2 inst_5300 ( .ZN(net_20146), .A4(net_19853), .A1(net_19852), .A3(net_14904), .A2(net_14471) );
NOR3_X2 inst_2766 ( .ZN(net_9933), .A2(net_9932), .A3(net_9931), .A1(net_5347) );
INV_X8 inst_12340 ( .ZN(net_5875), .A(net_493) );
NOR2_X2 inst_4326 ( .A1(net_6884), .A2(net_6039), .ZN(net_5817) );
NAND2_X2 inst_7938 ( .ZN(net_18428), .A2(net_18369), .A1(net_18311) );
AOI21_X2 inst_20515 ( .A(net_15300), .ZN(net_14603), .B2(net_11802), .B1(net_7720) );
INV_X4 inst_13985 ( .ZN(net_13617), .A(net_6560) );
INV_X2 inst_18663 ( .A(net_12520), .ZN(net_9180) );
INV_X2 inst_18382 ( .ZN(net_19123), .A(net_16551) );
INV_X2 inst_19221 ( .ZN(net_3466), .A(net_3465) );
XNOR2_X2 inst_127 ( .ZN(net_18300), .B(net_18256), .A(net_16997) );
INV_X4 inst_14754 ( .ZN(net_6995), .A(net_3124) );
INV_X4 inst_17535 ( .ZN(net_7780), .A(net_224) );
NAND2_X2 inst_11279 ( .ZN(net_4566), .A1(net_2585), .A2(net_2439) );
NAND2_X2 inst_10657 ( .ZN(net_9842), .A1(net_6314), .A2(net_4647) );
INV_X4 inst_14562 ( .A(net_7705), .ZN(net_4565) );
XNOR2_X2 inst_122 ( .ZN(net_18435), .A(net_18250), .B(net_16853) );
OAI22_X2 inst_1268 ( .ZN(net_17202), .A1(net_17082), .B1(net_16732), .A2(net_16637), .B2(net_16494) );
NOR2_X4 inst_3029 ( .ZN(net_8421), .A2(net_5106), .A1(net_703) );
INV_X4 inst_14270 ( .A(net_7182), .ZN(net_6690) );
NAND2_X2 inst_8944 ( .A1(net_15217), .ZN(net_14730), .A2(net_13235) );
AND2_X4 inst_21167 ( .ZN(net_19193), .A1(net_14536), .A2(net_12193) );
AOI21_X2 inst_20436 ( .ZN(net_15157), .B1(net_15156), .B2(net_13881), .A(net_11480) );
INV_X4 inst_15053 ( .ZN(net_5649), .A(net_3318) );
NAND2_X2 inst_9740 ( .A1(net_13651), .ZN(net_10102), .A2(net_10101) );
CLKBUF_X2 inst_22336 ( .A(net_21649), .Z(net_22208) );
NAND3_X2 inst_6281 ( .ZN(net_12898), .A3(net_11587), .A1(net_10807), .A2(net_7550) );
NAND2_X4 inst_7540 ( .A1(net_20860), .ZN(net_3028), .A2(net_1878) );
INV_X4 inst_17657 ( .ZN(net_4205), .A(net_262) );
NOR2_X2 inst_3912 ( .A1(net_20419), .ZN(net_8857), .A2(net_5160) );
NAND2_X2 inst_10077 ( .ZN(net_12117), .A2(net_7810), .A1(net_6719) );
NAND2_X2 inst_8499 ( .ZN(net_16931), .A1(net_16610), .A2(net_16474) );
OAI21_X2 inst_2306 ( .ZN(net_5767), .A(net_5766), .B2(net_3964), .B1(net_2222) );
NAND2_X2 inst_9191 ( .ZN(net_13118), .A2(net_13117), .A1(net_8815) );
INV_X2 inst_19334 ( .ZN(net_3258), .A(net_2494) );
OAI21_X2 inst_1646 ( .A(net_16743), .ZN(net_15910), .B2(net_15406), .B1(net_15175) );
INV_X4 inst_14008 ( .ZN(net_10553), .A(net_6313) );
INV_X4 inst_14468 ( .ZN(net_7989), .A(net_4911) );
INV_X4 inst_15361 ( .A(net_5482), .ZN(net_3398) );
NAND3_X2 inst_6748 ( .A2(net_10415), .ZN(net_5798), .A1(net_5797), .A3(net_3624) );
NAND3_X2 inst_5773 ( .ZN(net_15893), .A3(net_15371), .A2(net_14757), .A1(net_11509) );
NAND2_X4 inst_7547 ( .ZN(net_3111), .A2(net_1687), .A1(net_938) );
INV_X4 inst_17167 ( .ZN(net_4158), .A(net_2274) );
NAND3_X2 inst_6294 ( .A3(net_19997), .ZN(net_12820), .A1(net_10936), .A2(net_9351) );
NAND3_X2 inst_6741 ( .ZN(net_6408), .A2(net_6407), .A3(net_6406), .A1(net_2943) );
INV_X4 inst_13664 ( .A(net_12286), .ZN(net_10189) );
CLKBUF_X2 inst_22522 ( .A(net_22393), .Z(net_22394) );
INV_X2 inst_18536 ( .ZN(net_11049), .A(net_11048) );
NAND3_X4 inst_5550 ( .ZN(net_16764), .A3(net_16327), .A1(net_15937), .A2(net_10813) );
OR2_X4 inst_1102 ( .ZN(net_5037), .A1(net_2992), .A2(net_823) );
NAND3_X2 inst_6368 ( .ZN(net_12075), .A2(net_8243), .A3(net_7189), .A1(net_7046) );
INV_X4 inst_13329 ( .ZN(net_11171), .A(net_9876) );
CLKBUF_X2 inst_22438 ( .A(net_21355), .Z(net_22310) );
SDFF_X2 inst_702 ( .Q(net_20953), .SE(net_18863), .SI(net_18844), .D(net_497), .CK(net_21500) );
NAND3_X2 inst_5860 ( .ZN(net_15384), .A3(net_14058), .A2(net_7767), .A1(net_6937) );
INV_X8 inst_12448 ( .A(net_20538), .ZN(net_20529) );
INV_X2 inst_18668 ( .ZN(net_9170), .A(net_9169) );
INV_X4 inst_15192 ( .A(net_10298), .ZN(net_4350) );
NAND2_X2 inst_9297 ( .ZN(net_12399), .A1(net_12398), .A2(net_9160) );
NAND2_X2 inst_9980 ( .A1(net_14669), .A2(net_10606), .ZN(net_8863) );
CLKBUF_X2 inst_22753 ( .A(net_22624), .Z(net_22625) );
INV_X8 inst_12233 ( .ZN(net_6200), .A(net_3553) );
INV_X4 inst_13912 ( .ZN(net_8846), .A(net_6967) );
NAND2_X2 inst_9049 ( .ZN(net_14020), .A1(net_13089), .A2(net_11955) );
CLKBUF_X2 inst_21992 ( .A(net_21863), .Z(net_21864) );
CLKBUF_X2 inst_21977 ( .A(net_21503), .Z(net_21849) );
INV_X2 inst_18533 ( .A(net_11497), .ZN(net_11079) );
INV_X8 inst_12365 ( .ZN(net_897), .A(net_174) );
NOR2_X4 inst_2928 ( .ZN(net_9405), .A2(net_4868), .A1(net_1298) );
INV_X4 inst_13335 ( .ZN(net_12707), .A(net_11647) );
XNOR2_X2 inst_400 ( .ZN(net_16682), .A(net_16677), .B(net_14415) );
NOR2_X2 inst_3813 ( .ZN(net_9828), .A2(net_9827), .A1(net_3352) );
NOR2_X4 inst_2991 ( .A1(net_19022), .ZN(net_9430), .A2(net_5169) );
NAND2_X2 inst_8895 ( .ZN(net_20630), .A1(net_15107), .A2(net_13890) );
NOR2_X2 inst_3513 ( .ZN(net_13825), .A1(net_13824), .A2(net_13823) );
NAND3_X2 inst_6309 ( .ZN(net_12776), .A1(net_11064), .A3(net_9701), .A2(net_8130) );
INV_X4 inst_16196 ( .ZN(net_16035), .A(net_1831) );
XNOR2_X2 inst_261 ( .A(net_20789), .ZN(net_17259), .B(net_16804) );
AOI21_X4 inst_20158 ( .ZN(net_15709), .B1(net_15708), .B2(net_14980), .A(net_9725) );
INV_X8 inst_12418 ( .A(net_20891), .ZN(net_874) );
CLKBUF_X2 inst_22007 ( .A(net_21878), .Z(net_21879) );
XNOR2_X2 inst_268 ( .B(net_21139), .ZN(net_17221), .A(net_17220) );
OAI21_X2 inst_1518 ( .ZN(net_18413), .A(net_18292), .B1(net_18291), .B2(net_18290) );
NAND2_X2 inst_8198 ( .A1(net_17926), .ZN(net_17885), .A2(net_17870) );
NAND2_X2 inst_10985 ( .ZN(net_8100), .A1(net_4711), .A2(net_3600) );
NAND2_X2 inst_8586 ( .A2(net_17526), .ZN(net_16714), .A1(net_16509) );
NAND2_X2 inst_9199 ( .ZN(net_13086), .A2(net_11361), .A1(net_1070) );
INV_X4 inst_18313 ( .ZN(net_20509), .A(net_20508) );
INV_X8 inst_12264 ( .ZN(net_3791), .A(net_2108) );
CLKBUF_X2 inst_21538 ( .A(net_21409), .Z(net_21410) );
INV_X4 inst_18092 ( .A(net_21090), .ZN(net_676) );
NAND2_X4 inst_7245 ( .ZN(net_13728), .A1(net_6599), .A2(net_5549) );
INV_X4 inst_14118 ( .ZN(net_6142), .A(net_6141) );
NOR2_X2 inst_3509 ( .ZN(net_20016), .A2(net_12181), .A1(net_11084) );
INV_X4 inst_13936 ( .ZN(net_8150), .A(net_6828) );
INV_X4 inst_17758 ( .ZN(net_526), .A(net_165) );
NAND2_X2 inst_7971 ( .A2(net_20392), .A1(net_20391), .ZN(net_18359) );
NAND2_X2 inst_10746 ( .ZN(net_10736), .A1(net_5712), .A2(net_5519) );
NAND2_X2 inst_11511 ( .ZN(net_10570), .A2(net_2971), .A1(net_308) );
NAND3_X2 inst_6348 ( .ZN(net_12227), .A2(net_12226), .A3(net_12225), .A1(net_8687) );
NOR2_X4 inst_3097 ( .ZN(net_20497), .A2(net_4208), .A1(net_3212) );
NAND2_X2 inst_8357 ( .ZN(net_17452), .A1(net_17451), .A2(net_17450) );
NAND2_X2 inst_9229 ( .ZN(net_12896), .A1(net_10938), .A2(net_5765) );
NAND2_X2 inst_9625 ( .ZN(net_20841), .A2(net_7334), .A1(net_7246) );
CLKBUF_X2 inst_21830 ( .A(x7698), .Z(net_21702) );
XNOR2_X2 inst_502 ( .ZN(net_8998), .B(net_8997), .A(net_2515) );
CLKBUF_X2 inst_21837 ( .A(net_21708), .Z(net_21709) );
INV_X4 inst_13976 ( .ZN(net_9572), .A(net_4955) );
NAND2_X2 inst_8745 ( .A1(net_19406), .ZN(net_15987), .A2(net_1046) );
INV_X4 inst_18212 ( .A(net_21055), .ZN(net_637) );
INV_X4 inst_17966 ( .A(net_20921), .ZN(net_10216) );
INV_X4 inst_14771 ( .ZN(net_6418), .A(net_4049) );
NOR2_X2 inst_3645 ( .ZN(net_11933), .A2(net_9944), .A1(net_7186) );
OAI21_X2 inst_1598 ( .A(net_20968), .B2(net_20605), .B1(net_20604), .ZN(net_19315) );
INV_X4 inst_15724 ( .A(net_9438), .ZN(net_1965) );
INV_X4 inst_17040 ( .ZN(net_11189), .A(net_6879) );
INV_X4 inst_17098 ( .A(net_2965), .ZN(net_1358) );
NAND2_X2 inst_10167 ( .ZN(net_8237), .A1(net_8236), .A2(net_8235) );
INV_X4 inst_15670 ( .ZN(net_3946), .A(net_1558) );
CLKBUF_X2 inst_21945 ( .A(net_21499), .Z(net_21817) );
NAND2_X2 inst_7880 ( .ZN(net_18524), .A1(net_18465), .A2(net_18437) );
NOR2_X4 inst_3152 ( .ZN(net_4049), .A1(net_3322), .A2(net_2213) );
INV_X4 inst_15073 ( .A(net_11770), .ZN(net_3399) );
NOR2_X2 inst_4161 ( .A1(net_8664), .ZN(net_8217), .A2(net_6526) );
INV_X4 inst_18166 ( .ZN(net_125), .A(x7642) );
NAND2_X2 inst_11678 ( .ZN(net_3135), .A2(net_2358), .A1(net_2329) );
NAND2_X2 inst_10117 ( .ZN(net_20259), .A1(net_8395), .A2(net_5915) );
NAND3_X2 inst_5869 ( .ZN(net_15311), .A1(net_14377), .A3(net_13456), .A2(net_6206) );
CLKBUF_X2 inst_21556 ( .A(net_21427), .Z(net_21428) );
NOR2_X4 inst_3196 ( .A1(net_20479), .ZN(net_5401), .A2(net_3102) );
CLKBUF_X2 inst_21831 ( .A(net_21702), .Z(net_21703) );
INV_X4 inst_14603 ( .ZN(net_9236), .A(net_4466) );
CLKBUF_X2 inst_21646 ( .A(net_21266), .Z(net_21518) );
NAND3_X2 inst_6525 ( .ZN(net_10621), .A1(net_10620), .A2(net_10619), .A3(net_10618) );
INV_X4 inst_15452 ( .ZN(net_4221), .A(net_1722) );
INV_X4 inst_18252 ( .A(net_21145), .ZN(net_101) );
NOR2_X2 inst_4025 ( .A1(net_15297), .ZN(net_8012), .A2(net_8011) );
XNOR2_X2 inst_322 ( .B(net_17494), .A(net_17040), .ZN(net_17035) );
NOR2_X2 inst_3516 ( .ZN(net_13790), .A1(net_13789), .A2(net_13788) );
NAND2_X2 inst_10070 ( .A1(net_14365), .ZN(net_8658), .A2(net_8657) );
CLKBUF_X2 inst_22051 ( .A(net_21922), .Z(net_21923) );
NOR2_X2 inst_4200 ( .A1(net_14378), .ZN(net_6688), .A2(net_5734) );
INV_X2 inst_19570 ( .ZN(net_19016), .A(net_762) );
NOR2_X2 inst_3902 ( .ZN(net_13205), .A2(net_8969), .A1(net_253) );
NAND3_X2 inst_6191 ( .ZN(net_13321), .A1(net_13320), .A3(net_13319), .A2(net_12987) );
NAND2_X2 inst_10858 ( .ZN(net_7280), .A2(net_5114), .A1(net_4401) );
CLKBUF_X2 inst_22220 ( .A(net_22091), .Z(net_22092) );
NAND2_X2 inst_10647 ( .A2(net_6366), .ZN(net_6361), .A1(net_6360) );
AOI22_X2 inst_19969 ( .ZN(net_15813), .B1(net_14986), .A2(net_14889), .A1(net_14548), .B2(net_11806) );
NAND3_X2 inst_6243 ( .ZN(net_13178), .A2(net_13177), .A3(net_13176), .A1(net_7224) );
NAND2_X4 inst_6908 ( .A2(net_19605), .A1(net_19604), .ZN(net_17907) );
NAND2_X2 inst_8302 ( .A1(net_20428), .ZN(net_20235), .A2(net_17391) );
NAND3_X2 inst_6289 ( .ZN(net_20346), .A3(net_12286), .A2(net_11249), .A1(net_10257) );
OAI21_X2 inst_2315 ( .ZN(net_5705), .A(net_5239), .B1(net_3292), .B2(net_3291) );
INV_X4 inst_12662 ( .ZN(net_17810), .A(net_17809) );
SDFF_X2 inst_962 ( .QN(net_21095), .D(net_558), .SE(net_263), .CK(net_21783), .SI(x1471) );
NAND3_X2 inst_6350 ( .ZN(net_12162), .A1(net_11532), .A2(net_8762), .A3(net_6859) );
INV_X2 inst_18789 ( .ZN(net_10915), .A(net_9739) );
NAND2_X2 inst_11489 ( .A1(net_4751), .ZN(net_4001), .A2(net_3092) );
NAND2_X2 inst_9673 ( .ZN(net_10281), .A2(net_10280), .A1(net_9547) );
DFF_X2 inst_19773 ( .QN(net_20852), .D(net_18053), .CK(net_21804) );
NAND2_X2 inst_7955 ( .ZN(net_18396), .A2(net_18395), .A1(net_17993) );
INV_X4 inst_17395 ( .ZN(net_524), .A(net_523) );
INV_X4 inst_14044 ( .A(net_6260), .ZN(net_6259) );
INV_X2 inst_19119 ( .ZN(net_4434), .A(net_3828) );
NAND2_X2 inst_9308 ( .ZN(net_12368), .A1(net_9339), .A2(net_7573) );
CLKBUF_X2 inst_21596 ( .A(net_21467), .Z(net_21468) );
NAND2_X2 inst_11876 ( .ZN(net_2101), .A2(net_1625), .A1(net_131) );
CLKBUF_X2 inst_21674 ( .A(net_21533), .Z(net_21546) );
AOI211_X4 inst_20990 ( .C1(net_19197), .ZN(net_16084), .C2(net_15681), .B(net_14836), .A(net_12597) );
XNOR2_X2 inst_350 ( .B(net_21179), .ZN(net_16938), .A(net_16442) );
NAND2_X2 inst_11322 ( .ZN(net_7037), .A2(net_3756), .A1(net_154) );
INV_X2 inst_19501 ( .ZN(net_1260), .A(net_200) );
NAND2_X2 inst_10403 ( .A1(net_10562), .ZN(net_7274), .A2(net_6738) );
INV_X4 inst_14437 ( .A(net_5066), .ZN(net_5003) );
NOR2_X2 inst_5104 ( .A2(net_20851), .ZN(net_1152), .A1(net_846) );
INV_X4 inst_16853 ( .ZN(net_10956), .A(net_1019) );
INV_X4 inst_18275 ( .A(net_19457), .ZN(net_19456) );
AOI21_X2 inst_20379 ( .B1(net_15684), .ZN(net_15559), .B2(net_14712), .A(net_13280) );
INV_X4 inst_12851 ( .ZN(net_17362), .A(net_17234) );
NAND2_X2 inst_8518 ( .ZN(net_20089), .A1(net_19447), .A2(net_16911) );
NAND2_X2 inst_11901 ( .ZN(net_2781), .A1(net_1574), .A2(net_216) );
NAND2_X4 inst_7506 ( .A2(net_19897), .ZN(net_3903), .A1(net_1956) );
OAI21_X4 inst_1452 ( .B2(net_19081), .B1(net_19080), .ZN(net_15446), .A(net_15353) );
NAND2_X2 inst_11867 ( .A2(net_5959), .A1(net_2744), .ZN(net_1648) );
INV_X4 inst_13740 ( .ZN(net_13515), .A(net_7643) );
NAND3_X2 inst_6549 ( .ZN(net_10533), .A2(net_10207), .A3(net_10185), .A1(net_8435) );
INV_X4 inst_16743 ( .ZN(net_1425), .A(net_1047) );
INV_X4 inst_18176 ( .A(net_21056), .ZN(net_394) );
INV_X4 inst_12967 ( .ZN(net_16662), .A(net_16520) );
CLKBUF_X2 inst_22529 ( .A(net_22238), .Z(net_22401) );
CLKBUF_X2 inst_22638 ( .A(net_22509), .Z(net_22510) );
AND2_X2 inst_21325 ( .ZN(net_6300), .A2(net_6299), .A1(net_3383) );
OAI21_X4 inst_1396 ( .ZN(net_19577), .B2(net_19256), .B1(net_19255), .A(net_16347) );
AOI21_X2 inst_20400 ( .ZN(net_15393), .B1(net_14496), .B2(net_13971), .A(net_9734) );
NAND2_X2 inst_8901 ( .ZN(net_15089), .A1(net_15088), .A2(net_13916) );
CLKBUF_X2 inst_22204 ( .A(net_22075), .Z(net_22076) );
INV_X4 inst_15768 ( .ZN(net_12382), .A(net_11087) );
INV_X4 inst_15311 ( .A(net_11858), .ZN(net_2649) );
INV_X4 inst_16774 ( .ZN(net_19150), .A(net_932) );
NOR2_X4 inst_3003 ( .ZN(net_7424), .A1(net_4537), .A2(net_167) );
NAND3_X4 inst_5579 ( .ZN(net_19758), .A3(net_14234), .A1(net_8897), .A2(net_8601) );
INV_X8 inst_12169 ( .ZN(net_18624), .A(net_18612) );
INV_X4 inst_16978 ( .ZN(net_15064), .A(net_449) );
INV_X4 inst_16641 ( .ZN(net_5077), .A(net_3929) );
OAI21_X2 inst_2185 ( .ZN(net_8823), .A(net_8822), .B2(net_4976), .B1(net_3905) );
NAND2_X2 inst_8550 ( .A1(net_21236), .ZN(net_16793), .A2(net_16792) );
NAND2_X2 inst_9165 ( .ZN(net_13374), .A2(net_10649), .A1(net_10158) );
INV_X4 inst_13134 ( .ZN(net_19032), .A(net_14778) );
NOR2_X2 inst_4050 ( .A2(net_7881), .ZN(net_7856), .A1(net_5982) );
INV_X4 inst_16604 ( .ZN(net_14548), .A(net_60) );
OAI211_X4 inst_2370 ( .C2(net_20896), .C1(net_18960), .ZN(net_16898), .B(net_16244), .A(net_8886) );
NOR2_X2 inst_3882 ( .ZN(net_10862), .A2(net_9467), .A1(net_4718) );
INV_X4 inst_14069 ( .ZN(net_9750), .A(net_8316) );
INV_X2 inst_19302 ( .ZN(net_4712), .A(net_2770) );
INV_X4 inst_16868 ( .ZN(net_10183), .A(net_4900) );
NOR2_X4 inst_2811 ( .ZN(net_17697), .A1(net_17279), .A2(net_17145) );
INV_X4 inst_17597 ( .ZN(net_1699), .A(net_327) );
XNOR2_X2 inst_137 ( .ZN(net_18218), .A(net_18093), .B(net_16694) );
NOR2_X2 inst_4615 ( .ZN(net_6348), .A1(net_4205), .A2(net_3249) );
NAND3_X2 inst_6120 ( .ZN(net_13856), .A2(net_13855), .A3(net_13854), .A1(net_8671) );
INV_X4 inst_18067 ( .A(net_20982), .ZN(net_1900) );
NAND2_X4 inst_6889 ( .ZN(net_18090), .A1(net_18089), .A2(net_5616) );
AOI21_X2 inst_20711 ( .ZN(net_12068), .A(net_12067), .B2(net_12066), .B1(net_9935) );
OAI211_X2 inst_2567 ( .B(net_20590), .A(net_20589), .ZN(net_9042), .C2(net_9041), .C1(net_8618) );
NAND2_X2 inst_11384 ( .ZN(net_4606), .A2(net_3538), .A1(net_338) );
NOR2_X4 inst_3206 ( .ZN(net_5526), .A1(net_3033), .A2(net_2979) );
NAND2_X2 inst_11742 ( .ZN(net_4328), .A1(net_1213), .A2(net_1130) );
NAND2_X2 inst_8591 ( .ZN(net_16699), .A2(net_16514), .A1(net_349) );
INV_X4 inst_17576 ( .ZN(net_832), .A(net_341) );
NOR2_X2 inst_4046 ( .A1(net_9571), .ZN(net_9428), .A2(net_7885) );
NAND2_X2 inst_10245 ( .ZN(net_8018), .A1(net_7097), .A2(net_5313) );
NAND2_X4 inst_7179 ( .ZN(net_10878), .A2(net_9430), .A1(net_9350) );
NAND2_X2 inst_11752 ( .ZN(net_4210), .A1(net_2955), .A2(net_1222) );
AOI21_X2 inst_20831 ( .ZN(net_9736), .A(net_9735), .B1(net_6491), .B2(net_4602) );
NAND2_X2 inst_8112 ( .ZN(net_18104), .A2(net_18101), .A1(net_17416) );
OAI21_X2 inst_1897 ( .ZN(net_13359), .B2(net_10330), .A(net_8596), .B1(net_5886) );
NAND2_X2 inst_8511 ( .ZN(net_16918), .A1(net_16899), .A2(net_16574) );
INV_X2 inst_18634 ( .ZN(net_9408), .A(net_9407) );
NAND2_X2 inst_10615 ( .A2(net_7037), .ZN(net_6590), .A1(net_4727) );
NAND2_X2 inst_11810 ( .A2(net_2073), .ZN(net_1853), .A1(net_1562) );
NOR2_X4 inst_3159 ( .A2(net_4394), .ZN(net_4080), .A1(net_2197) );
INV_X4 inst_15587 ( .ZN(net_3756), .A(net_1610) );
INV_X4 inst_15786 ( .ZN(net_3751), .A(net_3013) );
AOI21_X2 inst_20305 ( .B2(net_19795), .B1(net_19794), .A(net_16242), .ZN(net_16071) );
OAI21_X2 inst_1569 ( .ZN(net_16405), .A(net_16404), .B2(net_16257), .B1(net_14066) );
NAND2_X4 inst_7130 ( .ZN(net_14542), .A1(net_9672), .A2(net_8021) );
NAND2_X2 inst_11722 ( .A2(net_3654), .ZN(net_2916), .A1(net_225) );
INV_X4 inst_12990 ( .ZN(net_16636), .A(net_16492) );
OAI21_X2 inst_1772 ( .ZN(net_14691), .A(net_14643), .B2(net_11944), .B1(net_11684) );
NAND2_X4 inst_7080 ( .A1(net_19967), .ZN(net_19331), .A2(net_14242) );
NAND2_X4 inst_7314 ( .ZN(net_7906), .A1(net_5333), .A2(net_107) );
INV_X4 inst_13565 ( .ZN(net_9139), .A(net_9138) );
CLKBUF_X2 inst_22621 ( .A(net_22492), .Z(net_22493) );
INV_X4 inst_13725 ( .ZN(net_9316), .A(net_6551) );
INV_X4 inst_14738 ( .A(net_5574), .ZN(net_5181) );
OAI21_X2 inst_2143 ( .ZN(net_9939), .B1(net_7912), .A(net_5868), .B2(net_4676) );
OAI22_X2 inst_1291 ( .ZN(net_12503), .B1(net_7872), .B2(net_7625), .A1(net_6899), .A2(net_5864) );
INV_X4 inst_14233 ( .ZN(net_7486), .A(net_5823) );
NAND2_X4 inst_7671 ( .ZN(net_1095), .A1(net_244), .A2(net_155) );
XNOR2_X2 inst_359 ( .ZN(net_16888), .A(net_16887), .B(net_14911) );
NAND2_X2 inst_8239 ( .ZN(net_17748), .A1(net_17747), .A2(net_17746) );
INV_X4 inst_18030 ( .A(net_21195), .ZN(net_5788) );
CLKBUF_X2 inst_22005 ( .A(net_21876), .Z(net_21877) );
INV_X8 inst_12382 ( .A(net_325), .ZN(net_282) );
CLKBUF_X2 inst_22270 ( .A(net_21398), .Z(net_22142) );
AOI21_X2 inst_20718 ( .B1(net_20617), .ZN(net_19242), .B2(net_12001), .A(net_7138) );
AOI21_X2 inst_20968 ( .ZN(net_5271), .A(net_5270), .B2(net_5269), .B1(net_3710) );
OAI21_X2 inst_1962 ( .ZN(net_20342), .B1(net_12454), .A(net_4446), .B2(net_732) );
NOR2_X2 inst_4757 ( .A2(net_6426), .ZN(net_3822), .A1(net_2948) );
INV_X4 inst_13037 ( .A(net_16622), .ZN(net_16554) );
CLKBUF_X2 inst_21671 ( .A(net_21370), .Z(net_21543) );
INV_X4 inst_13582 ( .ZN(net_8979), .A(net_8978) );
NAND2_X2 inst_10492 ( .ZN(net_13943), .A2(net_6908), .A1(net_6611) );
NAND2_X2 inst_11551 ( .ZN(net_2863), .A1(net_2862), .A2(net_2797) );
INV_X4 inst_15334 ( .ZN(net_3405), .A(net_2601) );
NAND4_X2 inst_5283 ( .ZN(net_15954), .A4(net_15209), .A2(net_13777), .A1(net_10560), .A3(net_9899) );
INV_X4 inst_12925 ( .ZN(net_16810), .A(net_16513) );
INV_X4 inst_15635 ( .ZN(net_19008), .A(net_2140) );
CLKBUF_X2 inst_21570 ( .A(net_21334), .Z(net_21442) );
NAND3_X2 inst_6174 ( .ZN(net_13549), .A3(net_9213), .A2(net_4845), .A1(net_4281) );
NAND2_X2 inst_8168 ( .ZN(net_17959), .A2(net_17883), .A1(net_17837) );
XNOR2_X2 inst_194 ( .B(net_21137), .ZN(net_17677), .A(net_17673) );
CLKBUF_X2 inst_22856 ( .A(net_22727), .Z(net_22728) );
NAND2_X2 inst_8421 ( .ZN(net_17199), .A1(net_16924), .A2(net_16747) );
AND2_X4 inst_21205 ( .ZN(net_19046), .A1(net_13353), .A2(net_7818) );
NOR2_X2 inst_3453 ( .ZN(net_19717), .A2(net_14857), .A1(net_8808) );
NAND2_X4 inst_7686 ( .ZN(net_1301), .A2(net_776), .A1(net_185) );
INV_X4 inst_15594 ( .ZN(net_6407), .A(net_1603) );
INV_X2 inst_19721 ( .A(net_20785), .ZN(net_20784) );
INV_X4 inst_14181 ( .ZN(net_11278), .A(net_5987) );
NAND3_X2 inst_6136 ( .ZN(net_13723), .A3(net_12726), .A2(net_10546), .A1(net_7346) );
NAND2_X2 inst_8714 ( .A2(net_20968), .A1(net_20758), .ZN(net_16209) );
NAND2_X2 inst_11317 ( .ZN(net_6509), .A1(net_3766), .A2(net_1087) );
XNOR2_X2 inst_442 ( .ZN(net_15799), .A(net_15798), .B(net_14851) );
AOI21_X2 inst_20468 ( .ZN(net_14995), .B1(net_14994), .A(net_13552), .B2(net_11975) );
OAI211_X2 inst_2507 ( .ZN(net_12743), .B(net_12742), .C2(net_12741), .A(net_11784), .C1(net_7118) );
NAND2_X2 inst_8338 ( .A1(net_21149), .ZN(net_17496), .A2(net_17463) );
NAND2_X2 inst_9337 ( .A1(net_14458), .A2(net_13018), .ZN(net_12277) );
OAI21_X2 inst_2245 ( .ZN(net_7354), .A(net_4421), .B2(net_4420), .B1(net_1097) );
INV_X2 inst_19423 ( .ZN(net_1827), .A(net_1826) );
INV_X4 inst_14751 ( .ZN(net_6996), .A(net_3126) );
NAND4_X4 inst_5237 ( .ZN(net_18967), .A1(net_15078), .A3(net_14547), .A2(net_8668), .A4(net_7842) );
INV_X4 inst_12620 ( .ZN(net_17998), .A(net_17997) );
INV_X4 inst_15467 ( .ZN(net_20693), .A(net_2462) );
NAND3_X2 inst_6097 ( .ZN(net_13918), .A3(net_13161), .A2(net_10965), .A1(net_8615) );
CLKBUF_X2 inst_21434 ( .A(net_21287), .Z(net_21306) );
NOR2_X2 inst_4298 ( .A1(net_6637), .ZN(net_5961), .A2(net_4542) );
NAND2_X2 inst_11242 ( .ZN(net_4944), .A1(net_3929), .A2(net_2728) );
INV_X4 inst_14593 ( .ZN(net_15573), .A(net_14264) );
OAI22_X4 inst_1249 ( .ZN(net_9944), .B2(net_9943), .B1(net_9942), .A1(net_4963), .A2(net_3720) );
NAND2_X4 inst_7212 ( .ZN(net_11874), .A2(net_7890), .A1(net_7837) );
NOR2_X2 inst_4099 ( .ZN(net_8672), .A1(net_8533), .A2(net_5740) );
INV_X4 inst_15815 ( .A(net_5616), .ZN(net_1873) );
NOR2_X2 inst_4740 ( .A2(net_3073), .ZN(net_3050), .A1(net_3049) );
NAND4_X2 inst_5403 ( .ZN(net_14712), .A3(net_14711), .A2(net_12354), .A4(net_12033), .A1(net_11669) );
NAND3_X2 inst_5967 ( .ZN(net_20336), .A3(net_13415), .A1(net_11637), .A2(net_10857) );
OAI22_X2 inst_1318 ( .ZN(net_5242), .B1(net_5241), .B2(net_5240), .A1(net_5009), .A2(net_2640) );
NAND2_X4 inst_6894 ( .A2(net_20912), .ZN(net_18050), .A1(net_15933) );
NAND2_X4 inst_7219 ( .A2(net_20487), .ZN(net_20040), .A1(net_5833) );
AOI21_X2 inst_20740 ( .A(net_11482), .ZN(net_11429), .B2(net_7640), .B1(net_3577) );
CLKBUF_X2 inst_22149 ( .A(net_22020), .Z(net_22021) );
INV_X4 inst_16970 ( .ZN(net_3436), .A(net_1237) );
INV_X2 inst_18444 ( .ZN(net_19722), .A(net_12797) );
OR2_X4 inst_1070 ( .ZN(net_9769), .A1(net_9768), .A2(net_8917) );
NOR2_X2 inst_4584 ( .ZN(net_6555), .A2(net_3820), .A1(net_404) );
INV_X2 inst_19462 ( .ZN(net_2357), .A(net_1480) );
OAI211_X2 inst_2454 ( .ZN(net_19973), .C2(net_14430), .C1(net_13742), .A(net_10360), .B(net_10025) );
NAND2_X2 inst_12037 ( .ZN(net_1221), .A1(net_926), .A2(net_63) );
NOR2_X2 inst_3601 ( .ZN(net_12549), .A2(net_9600), .A1(net_6906) );
INV_X8 inst_12255 ( .ZN(net_3834), .A(net_1564) );
AOI21_X2 inst_20573 ( .ZN(net_14132), .A(net_12627), .B2(net_10471), .B1(net_9891) );
INV_X4 inst_14612 ( .A(net_5945), .ZN(net_4427) );
NAND2_X2 inst_9693 ( .ZN(net_15457), .A1(net_10231), .A2(net_8161) );
NOR2_X2 inst_4536 ( .ZN(net_5086), .A2(net_4210), .A1(net_154) );
INV_X2 inst_18840 ( .ZN(net_12825), .A(net_7221) );
NAND3_X4 inst_5601 ( .ZN(net_14450), .A3(net_14449), .A2(net_13515), .A1(net_3460) );
NAND2_X2 inst_11854 ( .A2(net_20859), .ZN(net_1685), .A1(net_1661) );
NAND3_X2 inst_6763 ( .ZN(net_20637), .A3(net_5385), .A2(net_3173), .A1(net_2394) );
OAI21_X2 inst_1673 ( .ZN(net_20305), .B2(net_14218), .A(net_10683), .B1(net_7718) );
NAND3_X2 inst_5745 ( .A3(net_20701), .A1(net_20700), .ZN(net_19561), .A2(net_9029) );
INV_X4 inst_15163 ( .ZN(net_19911), .A(net_4316) );
CLKBUF_X2 inst_22870 ( .A(net_22741), .Z(net_22742) );
INV_X2 inst_18832 ( .ZN(net_6773), .A(net_6772) );
CLKBUF_X2 inst_21614 ( .A(net_21485), .Z(net_21486) );
INV_X4 inst_14373 ( .ZN(net_8249), .A(net_5180) );
OR2_X2 inst_1153 ( .ZN(net_9659), .A2(net_9658), .A1(net_816) );
NOR2_X2 inst_3823 ( .ZN(net_19927), .A2(net_9776), .A1(net_3998) );
NAND2_X4 inst_7632 ( .A1(net_1990), .ZN(net_1578), .A2(net_913) );
NAND2_X2 inst_7959 ( .A2(net_18393), .ZN(net_18389), .A1(net_17910) );
CLKBUF_X2 inst_22096 ( .A(net_21967), .Z(net_21968) );
NAND2_X4 inst_7325 ( .ZN(net_8316), .A1(net_3984), .A2(net_2668) );
NAND2_X2 inst_10905 ( .ZN(net_8951), .A1(net_6945), .A2(net_5423) );
XNOR2_X2 inst_391 ( .ZN(net_16770), .A(net_16769), .B(net_13284) );
INV_X4 inst_18272 ( .ZN(net_19452), .A(net_16328) );
AOI21_X4 inst_20239 ( .ZN(net_11177), .B1(net_7528), .B2(net_6208), .A(net_6050) );
INV_X2 inst_19165 ( .ZN(net_3878), .A(net_3877) );
NOR2_X2 inst_4107 ( .ZN(net_7181), .A2(net_5310), .A1(net_861) );
INV_X4 inst_15020 ( .ZN(net_15297), .A(net_3398) );
INV_X4 inst_18014 ( .A(net_21197), .ZN(net_9255) );
AOI21_X2 inst_20729 ( .B1(net_11907), .ZN(net_11778), .B2(net_9441), .A(net_5036) );
INV_X4 inst_17939 ( .A(net_21222), .ZN(net_62) );
AOI21_X2 inst_20763 ( .ZN(net_10861), .A(net_7629), .B2(net_7378), .B1(net_1778) );
INV_X4 inst_14092 ( .ZN(net_6199), .A(net_6198) );
AOI21_X2 inst_20981 ( .B1(net_11460), .ZN(net_3204), .B2(net_3203), .A(net_3153) );
NAND2_X2 inst_8035 ( .ZN(net_18259), .A2(net_18258), .A1(net_17744) );
NAND2_X2 inst_10896 ( .A1(net_7661), .ZN(net_5396), .A2(net_4282) );
CLKBUF_X2 inst_22162 ( .A(net_21823), .Z(net_22034) );
CLKBUF_X2 inst_22765 ( .A(net_22636), .Z(net_22637) );
NAND3_X2 inst_6074 ( .ZN(net_14113), .A3(net_10458), .A2(net_7933), .A1(net_6783) );
CLKBUF_X2 inst_21577 ( .A(net_21448), .Z(net_21449) );
INV_X4 inst_17702 ( .ZN(net_1086), .A(net_242) );
INV_X4 inst_17045 ( .ZN(net_10417), .A(net_5951) );
NAND2_X2 inst_8403 ( .A2(net_17571), .ZN(net_17249), .A1(net_437) );
OAI21_X2 inst_1799 ( .ZN(net_14491), .A(net_14490), .B1(net_12187), .B2(net_11559) );
NOR2_X2 inst_4442 ( .ZN(net_4806), .A1(net_4805), .A2(net_4804) );
INV_X4 inst_15129 ( .A(net_14509), .ZN(net_3379) );
NAND2_X4 inst_7385 ( .A1(net_19286), .ZN(net_5177), .A2(net_3919) );
NAND2_X2 inst_9326 ( .ZN(net_13805), .A1(net_12307), .A2(net_9338) );
INV_X4 inst_17954 ( .A(net_21059), .ZN(net_626) );
NOR2_X2 inst_3458 ( .ZN(net_14767), .A2(net_14136), .A1(net_9328) );
INV_X2 inst_19584 ( .A(net_380), .ZN(net_369) );
CLKBUF_X2 inst_22728 ( .A(net_22599), .Z(net_22600) );
INV_X2 inst_19215 ( .ZN(net_7157), .A(net_3480) );
INV_X2 inst_19517 ( .A(net_1828), .ZN(net_1123) );
OAI22_X2 inst_1313 ( .A1(net_13940), .B2(net_8954), .ZN(net_8468), .A2(net_8467), .B1(net_7850) );
NOR2_X2 inst_4694 ( .ZN(net_5637), .A1(net_2225), .A2(net_193) );
DFF_X1 inst_19895 ( .D(net_16938), .CK(net_22077), .Q(x346) );
NAND2_X2 inst_8098 ( .A2(net_20444), .ZN(net_18122), .A1(net_17140) );
NAND2_X2 inst_11104 ( .ZN(net_13885), .A1(net_6647), .A2(net_4331) );
INV_X4 inst_14572 ( .ZN(net_7494), .A(net_4542) );
CLKBUF_X2 inst_21415 ( .A(net_21286), .Z(net_21287) );
NAND2_X2 inst_8632 ( .ZN(net_16591), .A1(net_16590), .A2(net_16476) );
INV_X4 inst_16192 ( .ZN(net_13093), .A(net_11088) );
NOR2_X4 inst_2886 ( .ZN(net_11039), .A2(net_9668), .A1(net_7577) );
NOR2_X2 inst_4116 ( .ZN(net_7056), .A2(net_6568), .A1(net_5637) );
INV_X4 inst_15146 ( .ZN(net_19202), .A(net_3028) );
INV_X4 inst_14851 ( .A(net_11221), .ZN(net_3826) );
AOI21_X2 inst_20352 ( .ZN(net_15707), .B1(net_15706), .B2(net_15019), .A(net_9543) );
NAND3_X2 inst_6523 ( .ZN(net_10624), .A1(net_10623), .A3(net_7857), .A2(net_5183) );
NOR2_X1 inst_5150 ( .ZN(net_8388), .A2(net_7149), .A1(net_3421) );
AND2_X4 inst_21235 ( .ZN(net_19382), .A2(net_12142), .A1(net_4113) );
NAND2_X2 inst_9613 ( .A1(net_15827), .ZN(net_10712), .A2(net_8547) );
INV_X4 inst_13747 ( .ZN(net_9226), .A(net_7623) );
NAND2_X2 inst_10978 ( .ZN(net_8141), .A1(net_6592), .A2(net_4247) );
OAI21_X2 inst_2081 ( .ZN(net_10517), .A(net_7914), .B1(net_7836), .B2(net_5325) );
NOR3_X2 inst_2773 ( .ZN(net_8498), .A3(net_6846), .A2(net_3421), .A1(net_2834) );
INV_X4 inst_13199 ( .ZN(net_19227), .A(net_13240) );
AOI22_X2 inst_19960 ( .A1(net_16359), .ZN(net_16194), .A2(net_15865), .B2(net_14155), .B1(net_12712) );
NOR2_X4 inst_3261 ( .ZN(net_20796), .A2(net_2170), .A1(net_1027) );
NAND2_X2 inst_8717 ( .ZN(net_16195), .A2(net_16020), .A1(net_15631) );
INV_X4 inst_16570 ( .A(net_1200), .ZN(net_1161) );
INV_X4 inst_13606 ( .ZN(net_19211), .A(net_8475) );
INV_X4 inst_15796 ( .A(net_10587), .ZN(net_1894) );
OR2_X2 inst_1211 ( .ZN(net_13955), .A1(net_9903), .A2(net_7743) );
OR2_X2 inst_1192 ( .ZN(net_4274), .A2(net_4273), .A1(net_3269) );
XNOR2_X1 inst_682 ( .ZN(net_17776), .A(net_17775), .B(net_17774) );
XNOR2_X2 inst_238 ( .B(net_18214), .ZN(net_17393), .A(net_16943) );
INV_X8 inst_12394 ( .ZN(net_244), .A(net_162) );
INV_X4 inst_16012 ( .ZN(net_13544), .A(net_10188) );
INV_X4 inst_16338 ( .ZN(net_6945), .A(net_4250) );
NOR2_X4 inst_3333 ( .ZN(net_20800), .A1(net_525), .A2(net_220) );
INV_X4 inst_15908 ( .A(net_12067), .ZN(net_8186) );
NAND2_X2 inst_10021 ( .ZN(net_10249), .A2(net_8811), .A1(net_8764) );
NOR2_X4 inst_3109 ( .ZN(net_6997), .A1(net_4073), .A2(net_2881) );
NAND2_X2 inst_10046 ( .ZN(net_13126), .A2(net_11151), .A1(net_8707) );
INV_X2 inst_18448 ( .ZN(net_20695), .A(net_12690) );
OAI21_X2 inst_2240 ( .B1(net_20575), .ZN(net_7384), .B2(net_3688), .A(net_1318) );
INV_X4 inst_14995 ( .ZN(net_14552), .A(net_2212) );
AOI21_X4 inst_20167 ( .B1(net_20621), .B2(net_15804), .ZN(net_15631), .A(net_11857) );
OR2_X2 inst_1210 ( .ZN(net_5362), .A1(net_4288), .A2(net_3160) );
NAND2_X2 inst_11680 ( .ZN(net_7026), .A2(net_4085), .A1(net_3737) );
NAND3_X2 inst_6090 ( .ZN(net_13944), .A2(net_13943), .A1(net_12557), .A3(net_11448) );
INV_X4 inst_12759 ( .ZN(net_17395), .A(net_17394) );
INV_X4 inst_14674 ( .ZN(net_5536), .A(net_4312) );
INV_X4 inst_17804 ( .A(net_312), .ZN(net_133) );
OAI211_X2 inst_2437 ( .C1(net_15340), .ZN(net_14985), .C2(net_11988), .B(net_11755), .A(net_10012) );
INV_X4 inst_15154 ( .ZN(net_14365), .A(net_1927) );
INV_X2 inst_18553 ( .A(net_11582), .ZN(net_10902) );
NOR2_X2 inst_4521 ( .A1(net_5565), .ZN(net_4133), .A2(net_4132) );
AND2_X4 inst_21218 ( .ZN(net_5960), .A1(net_5959), .A2(net_5958) );
NAND2_X2 inst_8324 ( .ZN(net_17555), .A1(net_17554), .A2(net_17302) );
OAI21_X2 inst_1981 ( .ZN(net_12114), .A(net_10188), .B1(net_10139), .B2(net_8349) );
CLKBUF_X2 inst_22264 ( .A(net_22135), .Z(net_22136) );
NAND3_X2 inst_6324 ( .ZN(net_12514), .A3(net_12513), .A2(net_6240), .A1(net_1506) );
NAND3_X2 inst_5960 ( .ZN(net_20664), .A3(net_14829), .A1(net_8418), .A2(net_5887) );
INV_X4 inst_18190 ( .A(net_20864), .ZN(net_16395) );
INV_X4 inst_15122 ( .ZN(net_3176), .A(net_2215) );
INV_X4 inst_17022 ( .ZN(net_1076), .A(net_955) );
CLKBUF_X2 inst_22375 ( .A(net_21473), .Z(net_22247) );
NAND2_X2 inst_8309 ( .ZN(net_19729), .A2(net_17333), .A1(net_2554) );
NOR2_X2 inst_3775 ( .ZN(net_10220), .A1(net_10219), .A2(net_10218) );
INV_X4 inst_16266 ( .ZN(net_7007), .A(net_4288) );
INV_X4 inst_13762 ( .ZN(net_10977), .A(net_9635) );
OAI211_X2 inst_2472 ( .C2(net_13878), .ZN(net_13845), .A(net_13778), .B(net_12229), .C1(net_6415) );
INV_X4 inst_14900 ( .ZN(net_14083), .A(net_13355) );
NAND2_X2 inst_11239 ( .ZN(net_6526), .A2(net_4092), .A1(net_226) );
NAND2_X2 inst_8293 ( .ZN(net_20665), .A2(net_17613), .A1(net_17521) );
SDFF_X2 inst_872 ( .Q(net_21227), .SI(net_17085), .SE(net_125), .CK(net_21456), .D(x7135) );
AOI221_X4 inst_20071 ( .C2(net_20656), .C1(net_20655), .ZN(net_20295), .A(net_13791), .B1(net_13310), .B2(net_12055) );
NAND3_X2 inst_6641 ( .ZN(net_8948), .A3(net_8947), .A1(net_6701), .A2(net_4564) );
INV_X4 inst_16795 ( .ZN(net_11407), .A(net_652) );
NAND2_X2 inst_11479 ( .ZN(net_3124), .A2(net_2744), .A1(net_2374) );
INV_X4 inst_14821 ( .ZN(net_6561), .A(net_3868) );
NAND2_X2 inst_9210 ( .A1(net_13483), .ZN(net_13047), .A2(net_13046) );
NAND4_X4 inst_5234 ( .A4(net_19820), .A1(net_19819), .ZN(net_18884), .A2(net_11233), .A3(net_10679) );
INV_X4 inst_12579 ( .ZN(net_18258), .A(net_18170) );
INV_X4 inst_14907 ( .ZN(net_6042), .A(net_3585) );
CLKBUF_X2 inst_21766 ( .A(net_21637), .Z(net_21638) );
OAI21_X2 inst_1667 ( .ZN(net_15665), .A(net_15452), .B2(net_14891), .B1(net_11056) );
INV_X4 inst_15375 ( .ZN(net_4619), .A(net_2566) );
INV_X4 inst_17985 ( .A(net_21188), .ZN(net_516) );
XNOR2_X2 inst_462 ( .ZN(net_13287), .B(net_13286), .A(net_9257) );
INV_X4 inst_15339 ( .ZN(net_3562), .A(net_2286) );
AOI22_X4 inst_19956 ( .A1(net_20458), .A2(net_15191), .B1(net_14793), .ZN(net_14577), .B2(net_9302) );
NAND2_X2 inst_10261 ( .ZN(net_7990), .A2(net_7989), .A1(net_2212) );
NAND3_X4 inst_5572 ( .ZN(net_15865), .A3(net_15335), .A1(net_14693), .A2(net_13671) );
NAND2_X2 inst_9398 ( .ZN(net_11700), .A2(net_11699), .A1(net_11164) );
AOI22_X2 inst_20002 ( .A1(net_14820), .ZN(net_13630), .A2(net_13629), .B1(net_10664), .B2(net_5822) );
NAND2_X2 inst_10579 ( .A1(net_8485), .ZN(net_6680), .A2(net_6679) );
NAND2_X4 inst_7223 ( .A2(net_19205), .ZN(net_10922), .A1(net_4396) );
INV_X2 inst_18975 ( .ZN(net_5207), .A(net_5206) );
INV_X2 inst_18641 ( .ZN(net_11484), .A(net_9376) );
INV_X4 inst_13381 ( .ZN(net_10786), .A(net_10785) );
NAND3_X2 inst_6661 ( .A3(net_19419), .ZN(net_8451), .A1(net_4880), .A2(net_2579) );
INV_X2 inst_18693 ( .ZN(net_10370), .A(net_8363) );
NAND2_X2 inst_10389 ( .A1(net_12496), .ZN(net_10732), .A2(net_7317) );
NOR2_X2 inst_4909 ( .ZN(net_2935), .A2(net_2187), .A1(net_1770) );
NAND2_X4 inst_7114 ( .ZN(net_13659), .A1(net_11086), .A2(net_11050) );
NAND2_X4 inst_6836 ( .A1(net_20472), .A2(net_19489), .ZN(net_18904) );
NAND2_X4 inst_7611 ( .A1(net_1803), .ZN(net_1374), .A2(net_606) );
OAI21_X2 inst_1914 ( .ZN(net_13066), .B1(net_13065), .A(net_11032), .B2(net_9715) );
OAI21_X2 inst_1975 ( .ZN(net_12192), .A(net_11236), .B2(net_8352), .B1(net_7587) );
NAND3_X2 inst_6219 ( .ZN(net_13244), .A1(net_10616), .A3(net_10053), .A2(net_5530) );
INV_X4 inst_14702 ( .ZN(net_8476), .A(net_4263) );
CLKBUF_X2 inst_22236 ( .A(net_21276), .Z(net_22108) );
AOI21_X2 inst_20615 ( .ZN(net_13656), .B1(net_13655), .B2(net_13654), .A(net_12426) );
INV_X4 inst_15855 ( .ZN(net_6854), .A(net_4952) );
NAND3_X2 inst_6647 ( .ZN(net_13919), .A3(net_7803), .A2(net_7597), .A1(net_3297) );
NOR2_X2 inst_4806 ( .ZN(net_8529), .A2(net_5859), .A1(net_2687) );
NAND2_X2 inst_9728 ( .ZN(net_10120), .A1(net_10119), .A2(net_10101) );
NAND2_X2 inst_9585 ( .A1(net_12658), .ZN(net_10916), .A2(net_10915) );
NAND2_X2 inst_8117 ( .A2(net_18147), .ZN(net_18091), .A1(net_17415) );
AOI22_X2 inst_20029 ( .ZN(net_9918), .A1(net_9917), .B1(net_9668), .A2(net_8171), .B2(net_4498) );
INV_X8 inst_12362 ( .ZN(net_954), .A(net_223) );
INV_X4 inst_17944 ( .A(net_21009), .ZN(net_533) );
INV_X4 inst_17155 ( .ZN(net_1207), .A(net_751) );
NAND2_X2 inst_11893 ( .ZN(net_2217), .A2(net_1593), .A1(net_539) );
NOR2_X4 inst_3017 ( .ZN(net_8221), .A1(net_5503), .A2(net_2828) );
NAND3_X2 inst_6389 ( .A3(net_13054), .ZN(net_12010), .A2(net_11970), .A1(net_5141) );
AOI21_X2 inst_20303 ( .A(net_16404), .ZN(net_16086), .B2(net_15558), .B1(net_15482) );
INV_X4 inst_17693 ( .A(net_1461), .ZN(net_1327) );
SDFF_X2 inst_845 ( .Q(net_21178), .SI(net_17315), .SE(net_125), .CK(net_22161), .D(x4603) );
AOI21_X4 inst_20122 ( .ZN(net_19602), .B2(net_15902), .A(net_15462), .B1(net_2573) );
NOR2_X2 inst_3554 ( .ZN(net_13035), .A2(net_10418), .A1(net_8733) );
OAI21_X4 inst_1367 ( .ZN(net_17596), .B2(net_17353), .A(net_17241), .B1(net_17189) );
INV_X4 inst_17613 ( .A(net_10514), .ZN(net_9581) );
INV_X4 inst_17289 ( .ZN(net_1813), .A(net_143) );
NAND2_X2 inst_10980 ( .ZN(net_4964), .A2(net_4804), .A1(net_2391) );
AOI21_X4 inst_20098 ( .ZN(net_18952), .B2(net_18067), .A(net_18056), .B1(net_16230) );
NAND2_X2 inst_9175 ( .ZN(net_13345), .A2(net_10538), .A1(net_3396) );
INV_X4 inst_16911 ( .A(net_15300), .ZN(net_15158) );
NAND2_X2 inst_10898 ( .A2(net_6684), .A1(net_6274), .ZN(net_5388) );
NOR2_X2 inst_3687 ( .A1(net_13702), .ZN(net_11414), .A2(net_9292) );
INV_X4 inst_15426 ( .A(net_16051), .ZN(net_2508) );
CLKBUF_X2 inst_21709 ( .A(net_21580), .Z(net_21581) );
NAND2_X2 inst_10837 ( .ZN(net_11661), .A1(net_9617), .A2(net_5480) );
INV_X2 inst_19477 ( .ZN(net_1407), .A(net_1406) );
NAND2_X2 inst_8434 ( .ZN(net_17158), .A1(net_16862), .A2(net_16861) );
CLKBUF_X2 inst_21820 ( .A(net_21691), .Z(net_21692) );
INV_X4 inst_17676 ( .ZN(net_4329), .A(net_242) );
NAND2_X2 inst_10103 ( .A1(net_13709), .ZN(net_8528), .A2(net_5470) );
NOR2_X4 inst_3053 ( .ZN(net_6148), .A2(net_3568), .A1(net_154) );
NAND2_X2 inst_7829 ( .ZN(net_19233), .A2(net_18649), .A1(net_16833) );
NAND2_X2 inst_10409 ( .ZN(net_19942), .A1(net_9626), .A2(net_7261) );
NOR2_X2 inst_4810 ( .A1(net_5712), .A2(net_3029), .ZN(net_2639) );
NAND2_X2 inst_9962 ( .ZN(net_8907), .A1(net_8906), .A2(net_5554) );
NAND2_X2 inst_10708 ( .ZN(net_8918), .A2(net_6000), .A1(net_5458) );
INV_X4 inst_17202 ( .ZN(net_1011), .A(net_167) );
NOR2_X4 inst_3103 ( .ZN(net_8541), .A1(net_4091), .A2(net_225) );
INV_X4 inst_16075 ( .ZN(net_7193), .A(net_6911) );
NAND2_X2 inst_11985 ( .ZN(net_1273), .A1(net_1272), .A2(net_1271) );
AOI22_X2 inst_20058 ( .A1(net_4783), .ZN(net_2943), .B1(net_2942), .A2(net_2402), .B2(net_1826) );
NOR2_X4 inst_3304 ( .A2(net_20876), .ZN(net_2325), .A1(net_839) );
NAND2_X4 inst_7520 ( .ZN(net_2794), .A1(net_2071), .A2(net_2070) );
CLKBUF_X2 inst_21797 ( .A(net_21384), .Z(net_21669) );
INV_X4 inst_16045 ( .ZN(net_1606), .A(net_1605) );
NAND2_X2 inst_7762 ( .ZN(net_18771), .A2(net_18728), .A1(net_18682) );
NAND4_X2 inst_5384 ( .ZN(net_15019), .A1(net_12625), .A4(net_11964), .A2(net_10549), .A3(net_5378) );
INV_X4 inst_17275 ( .A(net_4394), .ZN(net_4383) );
INV_X4 inst_16766 ( .ZN(net_1389), .A(net_1023) );
NOR2_X2 inst_4723 ( .A1(net_19424), .ZN(net_5487), .A2(net_1875) );
NOR2_X2 inst_3655 ( .ZN(net_14291), .A1(net_12542), .A2(net_11644) );
NAND2_X4 inst_7532 ( .ZN(net_2609), .A2(net_1955), .A1(net_1715) );
CLKBUF_X2 inst_21961 ( .A(net_21363), .Z(net_21833) );
NAND2_X1 inst_12145 ( .A2(net_17487), .ZN(net_16818), .A1(net_5792) );
NAND3_X2 inst_6692 ( .ZN(net_20617), .A3(net_7702), .A2(net_4229), .A1(net_2947) );
INV_X2 inst_19481 ( .A(net_6601), .ZN(net_1379) );
NAND3_X2 inst_6617 ( .ZN(net_9067), .A3(net_9066), .A2(net_9041), .A1(net_3522) );
OAI21_X2 inst_1888 ( .B2(net_19851), .B1(net_19850), .A(net_14160), .ZN(net_13502) );
NOR2_X4 inst_2843 ( .A2(net_19034), .A1(net_19033), .ZN(net_14591) );
OAI21_X2 inst_1763 ( .ZN(net_14705), .B1(net_14222), .B2(net_12161), .A(net_10504) );
NOR2_X2 inst_3379 ( .ZN(net_20689), .A2(net_16284), .A1(net_16282) );
INV_X4 inst_13071 ( .ZN(net_19318), .A(net_16217) );
INV_X4 inst_16061 ( .ZN(net_9183), .A(net_2660) );
AOI21_X4 inst_20134 ( .ZN(net_20309), .B1(net_19346), .B2(net_15087), .A(net_14030) );
INV_X2 inst_18473 ( .ZN(net_12656), .A(net_12655) );
NAND2_X4 inst_7190 ( .ZN(net_13764), .A1(net_7806), .A2(net_4155) );
INV_X4 inst_13685 ( .ZN(net_11847), .A(net_7972) );
OR2_X4 inst_1094 ( .A1(net_9668), .ZN(net_4015), .A2(net_4014) );
INV_X4 inst_14309 ( .A(net_10575), .ZN(net_5500) );
AOI21_X2 inst_20690 ( .ZN(net_12214), .A(net_10216), .B2(net_7991), .B1(net_2921) );
NOR2_X2 inst_4145 ( .ZN(net_6912), .A1(net_6911), .A2(net_4124) );
INV_X2 inst_19179 ( .ZN(net_6644), .A(net_5639) );
NOR2_X2 inst_4590 ( .A2(net_3847), .ZN(net_3796), .A1(net_117) );
NOR2_X2 inst_3680 ( .A2(net_19460), .ZN(net_11428), .A1(net_10386) );
NAND3_X2 inst_6376 ( .ZN(net_20108), .A1(net_12040), .A3(net_10435), .A2(net_2558) );
NAND2_X4 inst_7168 ( .A2(net_20528), .ZN(net_12995), .A1(net_9496) );
OAI21_X2 inst_1699 ( .A(net_15463), .ZN(net_15327), .B2(net_13643), .B1(net_9262) );
NOR2_X2 inst_4878 ( .ZN(net_5327), .A2(net_1397), .A1(net_1154) );
INV_X4 inst_12685 ( .ZN(net_17706), .A(net_17705) );
XOR2_X2 inst_50 ( .A(net_21191), .Z(net_403), .B(net_402) );
INV_X2 inst_18906 ( .ZN(net_7500), .A(net_6055) );
INV_X2 inst_19326 ( .A(net_8714), .ZN(net_2567) );
INV_X4 inst_16324 ( .ZN(net_8007), .A(net_4288) );
OAI211_X2 inst_2589 ( .ZN(net_5773), .A(net_5511), .C1(net_5510), .B(net_2465), .C2(net_2418) );
NAND2_X2 inst_11762 ( .ZN(net_2090), .A2(net_2089), .A1(net_168) );
NAND2_X2 inst_10626 ( .A2(net_14222), .ZN(net_11457), .A1(net_5479) );
INV_X4 inst_16849 ( .ZN(net_9309), .A(net_704) );
NAND2_X2 inst_8699 ( .A1(net_20952), .ZN(net_16317), .A2(net_16124) );
OAI21_X2 inst_1650 ( .A(net_16368), .ZN(net_15887), .B2(net_15320), .B1(net_10734) );
INV_X4 inst_18074 ( .A(net_21020), .ZN(net_714) );
INV_X2 inst_19098 ( .A(net_5972), .ZN(net_4540) );
NOR2_X2 inst_4439 ( .A2(net_20804), .ZN(net_5977), .A1(net_143) );
NAND2_X4 inst_7469 ( .ZN(net_8469), .A1(net_2610), .A2(net_661) );
NAND2_X2 inst_8250 ( .A1(net_20207), .ZN(net_17712), .A2(net_17711) );
NOR2_X4 inst_2872 ( .ZN(net_12334), .A2(net_10914), .A1(net_9156) );
NAND2_X2 inst_8683 ( .ZN(net_16448), .A2(net_16447), .A1(net_16424) );
INV_X2 inst_18702 ( .A(net_16009), .ZN(net_8298) );
NOR2_X2 inst_3380 ( .A2(net_19388), .A1(net_19387), .ZN(net_16376) );
INV_X4 inst_16887 ( .A(net_6525), .ZN(net_1895) );
AOI21_X2 inst_20868 ( .ZN(net_20348), .A(net_13343), .B2(net_8580), .B1(net_2907) );
SDFF_X2 inst_804 ( .Q(net_20914), .SE(net_18837), .SI(net_17960), .D(net_474), .CK(net_21265) );
INV_X4 inst_16147 ( .ZN(net_1463), .A(net_1462) );
INV_X2 inst_19285 ( .ZN(net_2898), .A(net_2897) );
INV_X4 inst_15965 ( .ZN(net_1691), .A(net_1690) );
NOR2_X4 inst_3290 ( .ZN(net_3292), .A2(net_2253), .A1(net_1556) );
NAND2_X2 inst_8824 ( .ZN(net_19160), .A2(net_14828), .A1(net_8230) );
XOR2_X2 inst_13 ( .B(net_21198), .Z(net_17030), .A(net_17029) );
OAI211_X2 inst_2584 ( .ZN(net_7664), .C2(net_7663), .B(net_6323), .C1(net_5358), .A(net_3721) );
CLKBUF_X2 inst_22298 ( .A(net_22169), .Z(net_22170) );
INV_X4 inst_14527 ( .ZN(net_19910), .A(net_4764) );
CLKBUF_X2 inst_21455 ( .A(net_21326), .Z(net_21327) );
NOR3_X2 inst_2755 ( .ZN(net_11355), .A3(net_11179), .A2(net_10030), .A1(net_9619) );
NAND2_X2 inst_9101 ( .ZN(net_13765), .A2(net_13764), .A1(net_12329) );
NAND2_X2 inst_9393 ( .ZN(net_11709), .A1(net_11708), .A2(net_11707) );
INV_X4 inst_17443 ( .ZN(net_3814), .A(net_761) );
OAI21_X2 inst_1819 ( .ZN(net_14161), .B2(net_10614), .A(net_10389), .B1(net_6985) );
INV_X4 inst_14718 ( .ZN(net_16054), .A(net_4189) );
INV_X4 inst_17080 ( .ZN(net_5459), .A(net_1345) );
XNOR2_X2 inst_453 ( .ZN(net_13952), .B(net_13951), .A(net_10495) );
XNOR2_X2 inst_493 ( .ZN(net_9237), .A(net_9236), .B(net_9235) );
XOR2_X2 inst_23 ( .A(net_21128), .Z(net_16678), .B(net_16677) );
OAI21_X2 inst_1822 ( .ZN(net_14154), .A(net_14153), .B2(net_10518), .B1(net_8760) );
NOR2_X2 inst_3790 ( .ZN(net_20058), .A1(net_8604), .A2(net_4153) );
INV_X2 inst_18765 ( .A(net_9274), .ZN(net_7607) );
INV_X4 inst_12551 ( .ZN(net_18332), .A(net_18280) );
AOI21_X2 inst_20751 ( .ZN(net_11350), .A(net_9591), .B2(net_7631), .B1(net_5010) );
INV_X4 inst_17282 ( .ZN(net_817), .A(net_217) );
NAND3_X2 inst_6701 ( .A3(net_10261), .A2(net_9695), .ZN(net_7360), .A1(net_1904) );
INV_X4 inst_15574 ( .ZN(net_9668), .A(net_4794) );
CLKBUF_X2 inst_22471 ( .A(net_21669), .Z(net_22343) );
NAND2_X2 inst_10340 ( .ZN(net_20267), .A1(net_5435), .A2(net_4396) );
INV_X4 inst_14798 ( .ZN(net_6716), .A(net_5386) );
DFFS_X1 inst_19929 ( .SN(x339831), .QN(net_21177), .D(net_18005), .CK(net_22478) );
SDFF_X2 inst_812 ( .Q(net_21153), .SI(net_17828), .SE(net_125), .CK(net_22251), .D(x5605) );
NAND2_X2 inst_10347 ( .ZN(net_7512), .A2(net_7511), .A1(net_809) );
INV_X4 inst_15535 ( .ZN(net_10976), .A(net_10829) );
XNOR2_X2 inst_179 ( .B(net_21161), .A(net_17771), .ZN(net_17770) );
AOI22_X2 inst_20020 ( .A1(net_12419), .ZN(net_11216), .A2(net_9806), .B1(net_6083), .B2(net_4666) );
INV_X4 inst_15603 ( .ZN(net_3256), .A(net_1736) );
OAI21_X2 inst_1730 ( .ZN(net_15083), .B2(net_12898), .B1(net_8905), .A(net_864) );
NAND3_X2 inst_5698 ( .A3(net_20819), .A1(net_20818), .ZN(net_16230), .A2(net_13859) );
NOR2_X2 inst_3799 ( .ZN(net_9881), .A1(net_6864), .A2(net_5389) );
XNOR2_X2 inst_76 ( .B(net_21159), .ZN(net_18708), .A(net_18652) );
NOR2_X2 inst_3734 ( .ZN(net_10807), .A2(net_7435), .A1(net_3967) );
AOI221_X4 inst_20074 ( .B1(net_19713), .ZN(net_15240), .C1(net_14490), .C2(net_13242), .A(net_12912), .B2(net_843) );
AND2_X2 inst_21311 ( .A1(net_12675), .A2(net_11906), .ZN(net_8610) );
XNOR2_X2 inst_172 ( .B(net_17876), .ZN(net_17817), .A(net_17334) );
NAND3_X2 inst_6769 ( .ZN(net_5298), .A2(net_5297), .A3(net_2513), .A1(net_2062) );
DFF_X1 inst_19920 ( .Q(net_21113), .D(net_14371), .CK(net_21693) );
NAND2_X2 inst_11228 ( .ZN(net_3953), .A1(net_3915), .A2(net_2761) );
INV_X4 inst_16870 ( .ZN(net_10592), .A(net_8502) );
XNOR2_X2 inst_277 ( .ZN(net_17174), .A(net_17170), .B(net_13286) );
NOR2_X2 inst_4366 ( .ZN(net_10219), .A1(net_6669), .A2(net_5491) );
XNOR2_X2 inst_83 ( .ZN(net_18575), .A(net_18536), .B(net_16841) );
NAND2_X2 inst_7787 ( .ZN(net_18722), .A2(net_18721), .A1(net_17083) );
CLKBUF_X2 inst_22877 ( .A(net_22056), .Z(net_22749) );
NOR2_X2 inst_4186 ( .ZN(net_8053), .A1(net_6750), .A2(net_6683) );
NAND3_X4 inst_5566 ( .ZN(net_15942), .A3(net_15219), .A1(net_14872), .A2(net_10712) );
CLKBUF_X2 inst_22177 ( .A(net_21803), .Z(net_22049) );
NAND2_X2 inst_7946 ( .ZN(net_18410), .A2(net_18286), .A1(net_17328) );
NOR2_X2 inst_3386 ( .ZN(net_16291), .A1(net_16115), .A2(net_15928) );
INV_X4 inst_13673 ( .ZN(net_9548), .A(net_8008) );
XNOR2_X2 inst_140 ( .B(net_21188), .ZN(net_18177), .A(net_18140) );
NAND2_X2 inst_7990 ( .A2(net_18332), .ZN(net_18324), .A1(net_17629) );
INV_X2 inst_19623 ( .A(net_21230), .ZN(net_36) );
INV_X4 inst_16880 ( .ZN(net_19038), .A(net_956) );
NOR2_X4 inst_2824 ( .A2(net_19275), .A1(net_19274), .ZN(net_16221) );
NAND3_X2 inst_5945 ( .ZN(net_14892), .A3(net_12693), .A2(net_10638), .A1(net_6584) );
NOR2_X2 inst_3594 ( .ZN(net_14913), .A2(net_12665), .A1(net_5486) );
NAND2_X2 inst_8155 ( .ZN(net_18001), .A2(net_17944), .A1(net_7385) );
CLKBUF_X2 inst_22570 ( .A(net_22441), .Z(net_22442) );
NOR2_X4 inst_3124 ( .A1(net_20578), .A2(net_19037), .ZN(net_4939) );
NAND2_X2 inst_7993 ( .ZN(net_18322), .A2(net_18266), .A1(net_18227) );
AND2_X4 inst_21158 ( .ZN(net_19405), .A2(net_13127), .A1(net_12652) );
NOR2_X4 inst_2952 ( .ZN(net_10695), .A2(net_5180), .A1(net_154) );
NAND2_X2 inst_11896 ( .A1(net_1848), .ZN(net_1585), .A2(net_913) );
INV_X4 inst_14990 ( .ZN(net_5282), .A(net_3399) );
INV_X4 inst_17621 ( .ZN(net_475), .A(net_300) );
XNOR2_X2 inst_174 ( .ZN(net_17781), .A(net_17754), .B(net_960) );
NAND2_X2 inst_11558 ( .A2(net_5884), .ZN(net_2832), .A1(net_2831) );
INV_X4 inst_17313 ( .ZN(net_4430), .A(net_601) );
INV_X4 inst_16462 ( .A(net_9972), .ZN(net_8874) );
CLKBUF_X2 inst_22408 ( .A(net_22279), .Z(net_22280) );
NAND2_X2 inst_8658 ( .A2(net_19432), .ZN(net_19130), .A1(net_9193) );
NAND2_X2 inst_8942 ( .ZN(net_14733), .A2(net_13502), .A1(net_10685) );
INV_X8 inst_12293 ( .ZN(net_4305), .A(net_3915) );
XOR2_X2 inst_5 ( .A(net_21190), .B(net_20444), .Z(net_18155) );
OAI21_X2 inst_2105 ( .A(net_10379), .ZN(net_10059), .B2(net_6151), .B1(net_2771) );
NAND2_X2 inst_11186 ( .A2(net_6446), .ZN(net_4106), .A1(net_2451) );
INV_X4 inst_17718 ( .ZN(net_10688), .A(net_10087) );
INV_X4 inst_17778 ( .A(net_20868), .ZN(net_3800) );
AOI21_X2 inst_20445 ( .ZN(net_15109), .A(net_15108), .B2(net_12918), .B1(net_6954) );
SDFF_X2 inst_729 ( .Q(net_20909), .SE(net_18859), .SI(net_18566), .D(net_4239), .CK(net_22711) );
NAND3_X2 inst_6567 ( .A2(net_10539), .ZN(net_10478), .A3(net_10477), .A1(net_2968) );
OAI21_X2 inst_2157 ( .A(net_12877), .ZN(net_9266), .B2(net_7503), .B1(net_4599) );
NAND3_X2 inst_6506 ( .ZN(net_10794), .A3(net_7233), .A2(net_6659), .A1(net_3272) );
NAND2_X2 inst_10891 ( .A1(net_6812), .ZN(net_6620), .A2(net_5351) );
NOR3_X2 inst_2783 ( .ZN(net_6458), .A3(net_6457), .A2(net_5127), .A1(net_2672) );
NOR2_X2 inst_4553 ( .ZN(net_6594), .A2(net_4010), .A1(net_3947) );
XNOR2_X2 inst_604 ( .A(net_17015), .B(net_16470), .ZN(net_16334) );
NAND3_X2 inst_5804 ( .ZN(net_15679), .A3(net_15093), .A1(net_12539), .A2(net_6653) );
NAND2_X2 inst_9004 ( .ZN(net_14282), .A2(net_13478), .A1(net_8820) );
NAND2_X4 inst_7085 ( .ZN(net_19368), .A2(net_15094), .A1(net_14964) );
NAND2_X4 inst_7539 ( .ZN(net_5385), .A2(net_2365), .A1(net_825) );
INV_X4 inst_13872 ( .ZN(net_7434), .A(net_7433) );
NOR2_X2 inst_4057 ( .A2(net_14314), .ZN(net_13788), .A1(net_8559) );
OR2_X2 inst_1179 ( .A1(net_13984), .ZN(net_5361), .A2(net_5360) );
INV_X2 inst_19367 ( .A(net_2908), .ZN(net_2227) );
AND3_X4 inst_21116 ( .ZN(net_13609), .A2(net_13608), .A3(net_13607), .A1(net_6687) );
XNOR2_X2 inst_292 ( .B(net_21136), .ZN(net_17133), .A(net_16973) );
NOR2_X2 inst_3650 ( .ZN(net_11672), .A1(net_11010), .A2(net_8281) );
NAND2_X2 inst_11661 ( .ZN(net_3231), .A2(net_1465), .A1(net_532) );
OAI21_X2 inst_2012 ( .ZN(net_11385), .A(net_11384), .B1(net_7581), .B2(net_7539) );
NAND2_X2 inst_11350 ( .A1(net_10993), .ZN(net_3649), .A2(net_3648) );
NAND2_X2 inst_10900 ( .ZN(net_6607), .A1(net_5799), .A2(net_5386) );
INV_X2 inst_19513 ( .ZN(net_1684), .A(net_851) );
AOI21_X2 inst_20370 ( .B1(net_19770), .ZN(net_15625), .B2(net_15044), .A(net_14002) );
INV_X4 inst_16768 ( .ZN(net_5438), .A(net_1604) );
NAND3_X2 inst_6605 ( .ZN(net_11695), .A3(net_9698), .A2(net_9542), .A1(net_904) );
SDFF_X2 inst_839 ( .Q(net_21142), .SI(net_17390), .SE(net_125), .CK(net_21403), .D(x3553) );
INV_X4 inst_16296 ( .ZN(net_15706), .A(net_15198) );
XNOR2_X2 inst_240 ( .B(net_21117), .ZN(net_17381), .A(net_17380) );
NAND4_X2 inst_5455 ( .ZN(net_13451), .A4(net_10016), .A3(net_9841), .A2(net_8832), .A1(net_4463) );
NOR2_X2 inst_3966 ( .ZN(net_8418), .A2(net_7818), .A1(net_7058) );
NAND2_X4 inst_7501 ( .ZN(net_3188), .A1(net_1781), .A2(net_1697) );
INV_X2 inst_19352 ( .ZN(net_2387), .A(net_2386) );
INV_X4 inst_13681 ( .ZN(net_12066), .A(net_7982) );
CLKBUF_X2 inst_21980 ( .A(net_21646), .Z(net_21852) );
AND2_X4 inst_21186 ( .ZN(net_20735), .A1(net_11041), .A2(net_11040) );
XNOR2_X2 inst_99 ( .ZN(net_18540), .A(net_18432), .B(net_18325) );
NAND3_X2 inst_6634 ( .ZN(net_8986), .A2(net_8985), .A1(net_5728), .A3(net_3004) );
NAND2_X2 inst_9997 ( .ZN(net_19755), .A1(net_8831), .A2(net_8114) );
INV_X4 inst_13210 ( .ZN(net_13666), .A(net_12889) );
INV_X4 inst_13152 ( .ZN(net_14888), .A(net_14374) );
NOR2_X2 inst_4384 ( .ZN(net_6132), .A2(net_3976), .A1(net_3890) );
NAND2_X2 inst_11050 ( .A1(net_11572), .ZN(net_4709), .A2(net_4708) );
OAI21_X2 inst_2059 ( .A(net_14759), .ZN(net_10700), .B1(net_8706), .B2(net_5577) );
INV_X4 inst_13851 ( .A(net_11175), .ZN(net_7467) );
NAND2_X4 inst_7023 ( .ZN(net_17236), .A1(net_16589), .A2(net_16460) );
NAND2_X2 inst_9445 ( .ZN(net_13814), .A1(net_11541), .A2(net_11540) );
NAND2_X2 inst_9473 ( .A2(net_12870), .ZN(net_11469), .A1(net_11468) );
XNOR2_X2 inst_311 ( .ZN(net_17087), .A(net_17086), .B(net_14421) );
NAND2_X2 inst_9656 ( .A1(net_13747), .ZN(net_10341), .A2(net_7944) );
AOI22_X2 inst_20022 ( .ZN(net_10516), .A1(net_10515), .B1(net_10514), .A2(net_6527), .B2(net_5969) );
INV_X4 inst_12461 ( .ZN(net_20007), .A(net_18851) );
INV_X4 inst_16390 ( .A(net_7975), .ZN(net_1274) );
CLKBUF_X2 inst_21486 ( .A(net_21357), .Z(net_21358) );
NAND2_X2 inst_9914 ( .A1(net_13620), .A2(net_9386), .ZN(net_9312) );
INV_X2 inst_18402 ( .A(net_16526), .ZN(net_16494) );
INV_X4 inst_13205 ( .ZN(net_13839), .A(net_13148) );
OAI21_X2 inst_2203 ( .A(net_9754), .ZN(net_8552), .B2(net_7000), .B1(net_4844) );
NAND2_X2 inst_8139 ( .ZN(net_18029), .A2(net_17990), .A1(net_17938) );
INV_X4 inst_13180 ( .ZN(net_14329), .A(net_13856) );
INV_X2 inst_18948 ( .A(net_16050), .ZN(net_5655) );
NAND2_X2 inst_10495 ( .ZN(net_13304), .A1(net_8644), .A2(net_4443) );
INV_X4 inst_14413 ( .A(net_6720), .ZN(net_6239) );
INV_X2 inst_19683 ( .A(net_20526), .ZN(net_20524) );
INV_X4 inst_17874 ( .ZN(net_20842), .A(net_874) );
OAI21_X2 inst_1930 ( .ZN(net_12942), .B1(net_12941), .B2(net_11775), .A(net_11511) );
INV_X4 inst_15002 ( .A(net_13350), .ZN(net_11541) );
INV_X2 inst_19534 ( .ZN(net_1258), .A(net_556) );
INV_X2 inst_19312 ( .ZN(net_2700), .A(net_2699) );
XNOR2_X2 inst_577 ( .B(net_17247), .ZN(net_614), .A(net_613) );
NAND3_X4 inst_5536 ( .A3(net_19983), .A1(net_19982), .ZN(net_17515), .A2(net_16121) );
INV_X8 inst_12305 ( .ZN(net_9254), .A(net_5875) );
INV_X4 inst_13497 ( .ZN(net_10933), .A(net_9446) );
NOR2_X2 inst_4975 ( .A1(net_20860), .ZN(net_1555), .A2(net_1141) );
INV_X4 inst_15269 ( .A(net_3819), .ZN(net_2765) );
NAND3_X2 inst_6760 ( .ZN(net_5617), .A3(net_5616), .A2(net_4348), .A1(net_3235) );
INV_X2 inst_19351 ( .A(net_3253), .ZN(net_2392) );
INV_X4 inst_17233 ( .ZN(net_667), .A(net_549) );
NOR2_X2 inst_3938 ( .ZN(net_10133), .A2(net_8670), .A1(net_81) );
NOR2_X4 inst_2865 ( .ZN(net_12402), .A1(net_11015), .A2(net_9943) );
NAND3_X2 inst_5986 ( .ZN(net_20397), .A2(net_14538), .A1(net_12296), .A3(net_11611) );
INV_X4 inst_14933 ( .ZN(net_6166), .A(net_3539) );
NOR2_X2 inst_4891 ( .ZN(net_3247), .A2(net_3027), .A1(net_168) );
AOI21_X2 inst_20731 ( .B1(net_14279), .ZN(net_11773), .B2(net_7894), .A(net_5014) );
INV_X4 inst_14520 ( .ZN(net_5814), .A(net_3496) );
NAND2_X4 inst_7460 ( .ZN(net_5131), .A1(net_2641), .A2(net_1797) );
NAND2_X2 inst_11016 ( .ZN(net_11167), .A1(net_4815), .A2(net_4814) );
NAND2_X2 inst_11092 ( .ZN(net_5125), .A2(net_4975), .A1(net_2859) );
NAND3_X2 inst_6264 ( .ZN(net_19468), .A1(net_12974), .A3(net_10437), .A2(net_7604) );
INV_X4 inst_17111 ( .A(net_786), .ZN(net_785) );
INV_X4 inst_17384 ( .A(net_3919), .ZN(net_3226) );
INV_X4 inst_14556 ( .A(net_4578), .ZN(net_4577) );
NAND2_X4 inst_7040 ( .ZN(net_16935), .A2(net_16401), .A1(net_16055) );
AND4_X4 inst_21089 ( .ZN(net_20254), .A4(net_14007), .A1(net_12737), .A3(net_11774), .A2(net_9765) );
NOR2_X2 inst_4905 ( .ZN(net_1971), .A2(net_1970), .A1(net_1969) );
INV_X4 inst_18350 ( .ZN(net_20794), .A(net_18107) );
INV_X4 inst_17855 ( .A(net_1790), .ZN(net_184) );
XNOR2_X2 inst_63 ( .ZN(net_18811), .A(net_18763), .B(net_17765) );
AOI21_X2 inst_20578 ( .ZN(net_14101), .B1(net_12419), .B2(net_10633), .A(net_7312) );
NAND2_X2 inst_7968 ( .A1(net_20762), .ZN(net_18364), .A2(net_18363) );
OR2_X2 inst_1233 ( .ZN(net_6784), .A2(net_6495), .A1(net_1543) );
NAND4_X2 inst_5469 ( .ZN(net_13219), .A1(net_12446), .A3(net_10986), .A4(net_10035), .A2(net_8879) );
NOR2_X4 inst_2924 ( .ZN(net_11735), .A1(net_7887), .A2(net_955) );
NAND2_X2 inst_10445 ( .A2(net_8947), .ZN(net_7180), .A1(net_4706) );
NAND2_X2 inst_11117 ( .ZN(net_11162), .A1(net_7489), .A2(net_4315) );
OAI21_X2 inst_2006 ( .A(net_14476), .ZN(net_11409), .B2(net_9234), .B1(net_2061) );
NAND2_X2 inst_10337 ( .ZN(net_12487), .A2(net_7511), .A1(net_6981) );
AOI21_X2 inst_20521 ( .B1(net_15345), .ZN(net_14562), .B2(net_11973), .A(net_10086) );
NOR3_X4 inst_2619 ( .ZN(net_20169), .A3(net_19873), .A1(net_19872), .A2(net_7768) );
INV_X4 inst_15625 ( .A(net_5300), .ZN(net_2150) );
NAND2_X4 inst_7057 ( .A1(net_19609), .ZN(net_18909), .A2(net_16394) );
OAI21_X2 inst_2033 ( .A(net_20484), .ZN(net_11309), .B1(net_10716), .B2(net_9777) );
NOR2_X2 inst_3465 ( .ZN(net_14602), .A2(net_13253), .A1(net_10253) );
INV_X4 inst_14131 ( .ZN(net_9625), .A(net_6109) );
NAND2_X2 inst_7850 ( .A2(net_20936), .ZN(net_18589), .A1(net_15932) );
NAND2_X4 inst_7675 ( .A1(net_1711), .ZN(net_1139), .A2(net_153) );
OAI211_X2 inst_2559 ( .C1(net_14554), .ZN(net_9922), .C2(net_9921), .B(net_4912), .A(net_3444) );
INV_X4 inst_13336 ( .ZN(net_12681), .A(net_11120) );
INV_X4 inst_13898 ( .ZN(net_20008), .A(net_7167) );
INV_X4 inst_16551 ( .ZN(net_2093), .A(net_778) );
NAND2_X2 inst_12039 ( .A2(net_20495), .ZN(net_1705), .A1(net_955) );
CLKBUF_X2 inst_21379 ( .A(net_21250), .Z(net_21251) );
NAND2_X2 inst_10201 ( .A2(net_20077), .ZN(net_10267), .A1(net_10037) );
NAND2_X4 inst_6997 ( .A2(net_20620), .A1(net_20619), .ZN(net_17200) );
NAND2_X2 inst_8386 ( .ZN(net_20410), .A1(net_17049), .A2(net_16903) );
NAND2_X2 inst_8837 ( .ZN(net_19116), .A2(net_14795), .A1(net_14278) );
NAND3_X2 inst_6125 ( .ZN(net_13748), .A1(net_13747), .A3(net_13746), .A2(net_8261) );
OAI22_X2 inst_1269 ( .B1(net_21167), .B2(net_20214), .A2(net_20213), .ZN(net_17038), .A1(net_16879) );
INV_X4 inst_12657 ( .ZN(net_17823), .A(net_17822) );
INV_X4 inst_13575 ( .A(net_12063), .ZN(net_9124) );
INV_X4 inst_14768 ( .A(net_5483), .ZN(net_5118) );
INV_X2 inst_18653 ( .A(net_11435), .ZN(net_9219) );
NAND2_X4 inst_7202 ( .A1(net_20618), .ZN(net_10235), .A2(net_6812) );
CLKBUF_X2 inst_22834 ( .A(net_22705), .Z(net_22706) );
INV_X4 inst_18301 ( .A(net_20480), .ZN(net_20479) );
NOR2_X4 inst_3241 ( .ZN(net_2889), .A2(net_2314), .A1(net_1796) );
INV_X4 inst_17253 ( .ZN(net_9350), .A(net_884) );
NAND2_X2 inst_11842 ( .ZN(net_1722), .A1(net_1018), .A2(net_957) );
OAI21_X2 inst_1620 ( .ZN(net_16073), .B2(net_15512), .A(net_14675), .B1(net_6866) );
NOR2_X2 inst_4958 ( .A1(net_3436), .ZN(net_2161), .A2(net_964) );
INV_X4 inst_16376 ( .A(net_10113), .ZN(net_8682) );
INV_X4 inst_13344 ( .ZN(net_13657), .A(net_11075) );
NAND2_X2 inst_10572 ( .ZN(net_6697), .A1(net_6696), .A2(net_6695) );
AND2_X4 inst_21199 ( .ZN(net_8821), .A1(net_8820), .A2(net_6473) );
XNOR2_X2 inst_347 ( .B(net_21131), .ZN(net_16941), .A(net_16438) );
AOI21_X2 inst_20417 ( .ZN(net_19608), .A(net_14238), .B2(net_5944), .B1(net_4892) );
NAND4_X2 inst_5438 ( .ZN(net_13915), .A3(net_13914), .A2(net_11206), .A4(net_8937), .A1(net_7187) );
NAND2_X2 inst_11600 ( .A2(net_2697), .ZN(net_2661), .A1(net_2300) );
SDFF_X2 inst_755 ( .Q(net_20864), .SE(net_18837), .SI(net_18526), .D(net_506), .CK(net_22456) );
AOI21_X2 inst_20820 ( .A(net_14319), .ZN(net_10005), .B1(net_6872), .B2(net_4518) );
OAI21_X2 inst_1724 ( .ZN(net_15093), .B2(net_13063), .B1(net_12808), .A(net_1774) );
NAND2_X2 inst_7918 ( .ZN(net_19693), .A2(net_18382), .A1(net_17888) );
NAND3_X2 inst_5855 ( .A1(net_19622), .ZN(net_15408), .A3(net_14897), .A2(net_8627) );
NOR2_X2 inst_4505 ( .A1(net_9984), .ZN(net_4220), .A2(net_2849) );
INV_X4 inst_13149 ( .ZN(net_19629), .A(net_14408) );
NOR3_X4 inst_2610 ( .A1(net_19019), .ZN(net_16060), .A2(net_15252), .A3(net_14936) );
NAND2_X2 inst_8819 ( .ZN(net_15574), .A1(net_15573), .A2(net_14845) );
SDFF_X2 inst_1043 ( .QN(net_21056), .D(net_394), .SE(net_263), .CK(net_22490), .SI(x2115) );
NOR2_X2 inst_4030 ( .ZN(net_7981), .A2(net_6222), .A1(net_2460) );
INV_X8 inst_12327 ( .ZN(net_8190), .A(net_165) );
NAND2_X4 inst_7230 ( .ZN(net_14092), .A1(net_9350), .A2(net_6843) );
NAND2_X2 inst_9234 ( .A1(net_14511), .ZN(net_14298), .A2(net_11130) );
CLKBUF_X2 inst_21872 ( .A(net_21743), .Z(net_21744) );
OAI21_X2 inst_1792 ( .ZN(net_14601), .A(net_14600), .B2(net_11791), .B1(net_9269) );
NAND2_X2 inst_9769 ( .ZN(net_9811), .A1(net_9810), .A2(net_6989) );
NOR2_X2 inst_4426 ( .ZN(net_6101), .A2(net_5054), .A1(net_409) );
INV_X2 inst_19439 ( .A(net_2089), .ZN(net_1704) );
CLKBUF_X2 inst_22303 ( .A(net_22174), .Z(net_22175) );
NAND3_X2 inst_6017 ( .ZN(net_14388), .A2(net_14387), .A3(net_14320), .A1(net_10019) );
NAND2_X2 inst_10231 ( .A1(net_9478), .ZN(net_8051), .A2(net_8050) );
NOR2_X2 inst_3353 ( .A2(net_19428), .ZN(net_17788), .A1(net_17429) );
NOR2_X2 inst_3634 ( .ZN(net_12190), .A2(net_12151), .A1(net_7616) );
INV_X4 inst_12877 ( .ZN(net_16930), .A(net_16929) );
INV_X2 inst_19719 ( .A(net_20782), .ZN(net_20781) );
NOR2_X2 inst_4598 ( .ZN(net_4744), .A1(net_3188), .A2(net_2569) );
INV_X2 inst_19450 ( .ZN(net_2167), .A(net_1265) );
NOR2_X2 inst_4681 ( .ZN(net_3220), .A2(net_3219), .A1(net_703) );
NAND2_X2 inst_9772 ( .ZN(net_19469), .A1(net_10454), .A2(net_9798) );
CLKBUF_X2 inst_21611 ( .A(net_21482), .Z(net_21483) );
NAND2_X2 inst_11204 ( .ZN(net_10593), .A1(net_5450), .A2(net_3864) );
INV_X4 inst_16157 ( .ZN(net_6482), .A(net_1455) );
AND2_X4 inst_21213 ( .ZN(net_6569), .A2(net_6568), .A1(net_2974) );
INV_X2 inst_18805 ( .ZN(net_7407), .A(net_7406) );
INV_X2 inst_18490 ( .ZN(net_12346), .A(net_12345) );
NOR2_X4 inst_3145 ( .A1(net_19508), .ZN(net_6076), .A2(net_170) );
NOR2_X2 inst_5144 ( .ZN(net_625), .A1(net_28), .A2(net_27) );
AND2_X4 inst_21251 ( .A2(net_2283), .A1(net_2264), .ZN(net_1594) );
XNOR2_X2 inst_648 ( .B(net_481), .ZN(net_385), .A(net_384) );
NAND2_X2 inst_10600 ( .ZN(net_7893), .A2(net_6740), .A1(net_6625) );
NAND2_X2 inst_7857 ( .ZN(net_18572), .A1(net_18557), .A2(net_18546) );
INV_X4 inst_13718 ( .ZN(net_11721), .A(net_7825) );
INV_X4 inst_16363 ( .ZN(net_7915), .A(net_1634) );
XNOR2_X2 inst_270 ( .B(net_21205), .A(net_20436), .ZN(net_17218) );
OAI21_X2 inst_1901 ( .B1(net_14572), .ZN(net_13333), .B2(net_9941), .A(net_7166) );
AND4_X2 inst_21103 ( .A4(net_12095), .ZN(net_11846), .A3(net_11845), .A2(net_7840), .A1(net_6287) );
AOI21_X4 inst_20223 ( .B2(net_20152), .B1(net_20151), .ZN(net_14054), .A(net_13076) );
AOI21_X2 inst_20845 ( .ZN(net_9261), .A(net_9260), .B2(net_4587), .B1(net_2309) );
NOR2_X2 inst_4104 ( .A1(net_13091), .ZN(net_7190), .A2(net_7189) );
CLKBUF_X2 inst_22749 ( .A(net_22620), .Z(net_22621) );
NAND2_X2 inst_11826 ( .ZN(net_5859), .A1(net_3830), .A2(net_1786) );
CLKBUF_X2 inst_21815 ( .A(net_21686), .Z(net_21687) );
NAND2_X2 inst_8608 ( .ZN(net_16645), .A1(net_16644), .A2(net_16643) );
OAI211_X2 inst_2552 ( .ZN(net_10809), .A(net_9282), .C1(net_7078), .C2(net_4613), .B(net_2177) );
INV_X2 inst_18914 ( .ZN(net_6012), .A(net_6011) );
XNOR2_X2 inst_631 ( .B(net_16644), .ZN(net_451), .A(net_450) );
NAND2_X2 inst_11809 ( .A2(net_2303), .ZN(net_1854), .A1(net_26) );
INV_X2 inst_18712 ( .ZN(net_8218), .A(net_8217) );
NAND3_X2 inst_6427 ( .ZN(net_11928), .A2(net_11927), .A3(net_9646), .A1(net_3676) );
INV_X4 inst_15070 ( .A(net_4151), .ZN(net_3400) );
NOR2_X2 inst_3674 ( .A1(net_12546), .A2(net_11603), .ZN(net_11475) );
AOI21_X2 inst_20975 ( .A(net_5239), .ZN(net_4454), .B2(net_4206), .B1(net_2196) );
INV_X4 inst_12835 ( .ZN(net_17120), .A(net_17119) );
NAND2_X2 inst_11346 ( .A1(net_7867), .ZN(net_3655), .A2(net_3654) );
INV_X4 inst_13505 ( .A(net_12284), .ZN(net_9417) );
INV_X4 inst_13789 ( .ZN(net_10958), .A(net_7566) );
CLKBUF_X2 inst_21531 ( .A(net_21372), .Z(net_21403) );
NOR2_X2 inst_3995 ( .ZN(net_8253), .A1(net_8252), .A2(net_8251) );
NOR2_X2 inst_5074 ( .ZN(net_11384), .A1(net_4329), .A2(net_910) );
INV_X2 inst_19198 ( .ZN(net_3597), .A(net_3596) );
XNOR2_X2 inst_102 ( .ZN(net_18533), .A(net_18424), .B(net_17259) );
INV_X4 inst_14749 ( .ZN(net_4549), .A(net_4076) );
OAI211_X2 inst_2527 ( .A(net_12647), .ZN(net_11780), .C1(net_11779), .B(net_10264), .C2(net_10238) );
CLKBUF_X2 inst_22251 ( .A(net_22122), .Z(net_22123) );
NOR2_X4 inst_3277 ( .ZN(net_2404), .A2(net_1697), .A1(net_1172) );
CLKBUF_X2 inst_22839 ( .A(net_22710), .Z(net_22711) );
NAND2_X2 inst_12042 ( .ZN(net_947), .A1(net_236), .A2(net_103) );
CLKBUF_X2 inst_21773 ( .A(net_21644), .Z(net_21645) );
AOI21_X2 inst_20388 ( .ZN(net_15469), .B1(net_15468), .B2(net_14587), .A(net_12112) );
NOR3_X2 inst_2786 ( .ZN(net_5583), .A2(net_4975), .A1(net_3776), .A3(net_3711) );
NAND4_X2 inst_5352 ( .ZN(net_15417), .A4(net_15416), .A1(net_14659), .A3(net_14092), .A2(net_7211) );
OR2_X2 inst_1224 ( .ZN(net_6782), .A1(net_2369), .A2(net_1325) );
NAND2_X2 inst_10043 ( .A1(net_9913), .ZN(net_8711), .A2(net_8710) );
NAND2_X2 inst_11045 ( .ZN(net_9958), .A1(net_4718), .A2(net_4717) );
INV_X4 inst_16040 ( .ZN(net_6580), .A(net_4838) );
NOR2_X2 inst_3905 ( .ZN(net_8884), .A2(net_8883), .A1(net_8064) );
NAND2_X4 inst_7666 ( .ZN(net_1178), .A1(net_1134), .A2(net_894) );
OR2_X2 inst_1170 ( .A2(net_10236), .ZN(net_6839), .A1(net_6838) );
NAND2_X2 inst_8929 ( .A1(net_15612), .ZN(net_14859), .A2(net_13603) );
NAND2_X2 inst_11797 ( .ZN(net_6004), .A1(net_5448), .A2(net_1940) );
INV_X4 inst_16886 ( .ZN(net_12609), .A(net_5735) );
CLKBUF_X2 inst_22397 ( .A(net_22268), .Z(net_22269) );
INV_X4 inst_14246 ( .ZN(net_7493), .A(net_5764) );
INV_X4 inst_15219 ( .ZN(net_4380), .A(net_2878) );
NAND2_X2 inst_11659 ( .A1(net_20556), .ZN(net_6971), .A2(net_1331) );
NAND2_X2 inst_8752 ( .ZN(net_15918), .A1(net_15917), .A2(net_15471) );
INV_X4 inst_17373 ( .A(net_949), .ZN(net_540) );
SDFF_X2 inst_785 ( .Q(net_20947), .SE(net_18858), .SI(net_18038), .D(net_569), .CK(net_21283) );
OAI21_X1 inst_2362 ( .ZN(net_10067), .A(net_10066), .B2(net_6169), .B1(net_2119) );
CLKBUF_X2 inst_21408 ( .A(net_21279), .Z(net_21280) );
INV_X2 inst_18389 ( .A(net_16789), .ZN(net_16635) );
NOR2_X4 inst_2856 ( .ZN(net_12290), .A2(net_9050), .A1(net_8847) );
NAND2_X2 inst_9280 ( .ZN(net_20139), .A1(net_9788), .A2(net_9508) );
NAND2_X2 inst_10417 ( .ZN(net_19926), .A1(net_10361), .A2(net_6755) );
NAND2_X2 inst_7945 ( .ZN(net_18416), .A2(net_18297), .A1(net_18257) );
XNOR2_X2 inst_527 ( .ZN(net_3435), .A(net_1948), .B(net_1942) );
XNOR2_X2 inst_226 ( .ZN(net_17501), .A(net_17184), .B(net_4450) );
OR2_X2 inst_1180 ( .ZN(net_13876), .A2(net_4987), .A1(net_4907) );
NAND4_X2 inst_5509 ( .A4(net_11359), .ZN(net_11235), .A3(net_11234), .A2(net_9041), .A1(net_1839) );
CLKBUF_X2 inst_22670 ( .A(net_22541), .Z(net_22542) );
INV_X2 inst_19066 ( .ZN(net_4639), .A(net_4638) );
NAND2_X2 inst_8223 ( .ZN(net_17872), .A2(net_17622), .A1(net_17559) );
INV_X4 inst_13861 ( .ZN(net_7460), .A(net_4823) );
NAND2_X2 inst_11232 ( .ZN(net_9076), .A1(net_4711), .A2(net_3946) );
XNOR2_X2 inst_212 ( .ZN(net_17546), .A(net_17149), .B(net_623) );
NAND2_X2 inst_11688 ( .ZN(net_2334), .A2(net_2332), .A1(net_193) );
CLKBUF_X2 inst_21878 ( .A(net_21555), .Z(net_21750) );
DFF_X1 inst_19792 ( .Q(net_20936), .D(net_18570), .CK(net_21699) );
NOR3_X2 inst_2732 ( .ZN(net_12848), .A3(net_12847), .A1(net_11127), .A2(net_11027) );
INV_X4 inst_16682 ( .A(net_10000), .ZN(net_8226) );
NAND3_X2 inst_6321 ( .ZN(net_12519), .A2(net_9212), .A3(net_5022), .A1(net_1578) );
NAND2_X2 inst_9323 ( .ZN(net_12325), .A1(net_11536), .A2(net_11422) );
INV_X4 inst_15293 ( .ZN(net_20152), .A(net_2715) );
INV_X2 inst_18627 ( .ZN(net_12538), .A(net_9547) );
DFF_X1 inst_19838 ( .D(net_17511), .CK(net_21355), .Q(x184) );
INV_X2 inst_18771 ( .ZN(net_12569), .A(net_7575) );
NAND2_X2 inst_10013 ( .ZN(net_8779), .A2(net_8159), .A1(net_7260) );
CLKBUF_X2 inst_21508 ( .A(net_21379), .Z(net_21380) );
NAND4_X2 inst_5431 ( .A2(net_19149), .A1(net_19148), .ZN(net_14109), .A4(net_11320), .A3(net_8022) );
AOI21_X2 inst_20485 ( .ZN(net_14835), .A(net_14600), .B2(net_13449), .B1(net_3778) );
NAND2_X2 inst_8330 ( .ZN(net_20236), .A2(net_17507), .A1(net_17392) );
INV_X4 inst_14638 ( .A(net_5485), .ZN(net_5113) );
NOR2_X4 inst_2966 ( .A2(net_11041), .ZN(net_7800), .A1(net_398) );
NOR2_X4 inst_3246 ( .ZN(net_4089), .A2(net_2294), .A1(net_1364) );
DFF_X1 inst_19805 ( .D(net_18177), .CK(net_22392), .Q(x833) );
NOR2_X2 inst_4904 ( .A2(net_2099), .ZN(net_1972), .A1(net_493) );
INV_X4 inst_16440 ( .ZN(net_1773), .A(net_809) );
INV_X2 inst_19059 ( .ZN(net_4699), .A(net_4698) );
INV_X4 inst_16803 ( .ZN(net_15666), .A(net_1006) );
NOR2_X2 inst_4887 ( .ZN(net_3406), .A2(net_1220), .A1(net_168) );
NAND2_X2 inst_11272 ( .ZN(net_3888), .A2(net_2083), .A1(net_674) );
OAI211_X4 inst_2381 ( .ZN(net_14744), .C1(net_14743), .B(net_13591), .C2(net_10602), .A(net_9637) );
NAND3_X2 inst_5823 ( .ZN(net_15570), .A2(net_15569), .A1(net_14812), .A3(net_14170) );
NAND2_X2 inst_11538 ( .A1(net_11443), .ZN(net_2921), .A2(net_1851) );
INV_X4 inst_16059 ( .ZN(net_3147), .A(net_1589) );
NAND2_X2 inst_11284 ( .A1(net_3924), .ZN(net_3851), .A2(net_3830) );
INV_X2 inst_19598 ( .A(net_20901), .ZN(net_19484) );
INV_X4 inst_16922 ( .ZN(net_1334), .A(net_1022) );
INV_X2 inst_18947 ( .A(net_8473), .ZN(net_7118) );
XNOR2_X2 inst_454 ( .ZN(net_13947), .B(net_13946), .A(net_10497) );
INV_X4 inst_13753 ( .ZN(net_10730), .A(net_7619) );
INV_X4 inst_13947 ( .ZN(net_9741), .A(net_6778) );
INV_X4 inst_14299 ( .ZN(net_8201), .A(net_5538) );
INV_X2 inst_18719 ( .ZN(net_8137), .A(net_8136) );
NAND2_X2 inst_8251 ( .A1(net_20462), .ZN(net_18888), .A2(net_17374) );
CLKBUF_X2 inst_22320 ( .A(net_21286), .Z(net_22192) );
INV_X4 inst_15475 ( .ZN(net_2859), .A(net_2457) );
INV_X2 inst_19379 ( .ZN(net_2157), .A(net_2156) );
INV_X4 inst_17035 ( .ZN(net_6221), .A(net_498) );
NAND2_X2 inst_7899 ( .ZN(net_18484), .A1(net_18381), .A2(net_18280) );
INV_X4 inst_16175 ( .ZN(net_5632), .A(net_1076) );
NAND2_X2 inst_11130 ( .A1(net_5330), .A2(net_4289), .ZN(net_4271) );
NAND2_X2 inst_11067 ( .ZN(net_10002), .A2(net_4580), .A1(net_4516) );
NAND2_X4 inst_6990 ( .A2(net_19840), .A1(net_19839), .ZN(net_17222) );
INV_X4 inst_13622 ( .A(net_8903), .ZN(net_8355) );
INV_X4 inst_12974 ( .A(net_16512), .ZN(net_16511) );
AOI211_X2 inst_21052 ( .ZN(net_11859), .C1(net_11858), .B(net_10300), .A(net_9558), .C2(net_2477) );
OAI211_X2 inst_2419 ( .ZN(net_15324), .A(net_14417), .B(net_11508), .C2(net_7779), .C1(net_4452) );
INV_X4 inst_14793 ( .ZN(net_4845), .A(net_4003) );
NAND2_X2 inst_9484 ( .A1(net_12888), .ZN(net_11452), .A2(net_10939) );
NAND2_X2 inst_11612 ( .ZN(net_2608), .A1(net_2607), .A2(net_2606) );
INV_X4 inst_17996 ( .A(net_21044), .ZN(net_467) );
NOR2_X2 inst_5041 ( .ZN(net_12053), .A2(net_8181), .A1(net_788) );
OAI21_X4 inst_1428 ( .B2(net_19685), .B1(net_19684), .ZN(net_18950), .A(net_16357) );
NAND2_X2 inst_11089 ( .A1(net_9183), .ZN(net_4365), .A2(net_2815) );
CLKBUF_X2 inst_22412 ( .A(net_22283), .Z(net_22284) );
INV_X4 inst_16467 ( .ZN(net_19488), .A(net_2948) );
NAND2_X2 inst_9456 ( .ZN(net_11506), .A1(net_11505), .A2(net_11504) );
NOR3_X2 inst_2739 ( .ZN(net_12758), .A2(net_12757), .A1(net_10205), .A3(net_6095) );
INV_X4 inst_12691 ( .ZN(net_17649), .A(net_17648) );
SDFF_X2 inst_1046 ( .QN(net_20993), .D(net_1862), .SE(net_263), .CK(net_21823), .SI(x3136) );
NAND3_X2 inst_5955 ( .ZN(net_19095), .A3(net_14829), .A1(net_12974), .A2(net_5090) );
NOR2_X2 inst_4355 ( .ZN(net_5608), .A2(net_5602), .A1(net_4736) );
NAND2_X2 inst_10152 ( .A1(net_18025), .ZN(net_8283), .A2(net_357) );
CLKBUF_X2 inst_22565 ( .A(net_22436), .Z(net_22437) );
NAND4_X2 inst_5426 ( .A2(net_20809), .A1(net_20808), .ZN(net_19663), .A4(net_9199), .A3(net_5116) );
NAND3_X2 inst_6206 ( .A2(net_13494), .ZN(net_13290), .A3(net_10288), .A1(net_5390) );
CLKBUF_X2 inst_22319 ( .A(net_22190), .Z(net_22191) );
NAND2_X2 inst_9515 ( .ZN(net_11146), .A2(net_9107), .A1(net_4140) );
CLKBUF_X2 inst_21510 ( .A(net_21330), .Z(net_21382) );
AOI21_X2 inst_20592 ( .ZN(net_13936), .B1(net_13080), .B2(net_11201), .A(net_5746) );
INV_X4 inst_16859 ( .ZN(net_1049), .A(net_964) );
INV_X4 inst_16454 ( .ZN(net_10470), .A(net_8629) );
SDFF_X2 inst_909 ( .Q(net_21155), .D(net_16770), .SE(net_263), .CK(net_22276), .SI(x5537) );
INV_X4 inst_17393 ( .ZN(net_9365), .A(net_4802) );
OAI211_X2 inst_2484 ( .C1(net_14315), .ZN(net_13480), .A(net_13479), .C2(net_12563), .B(net_6978) );
NAND3_X2 inst_5758 ( .ZN(net_15996), .A1(net_15707), .A3(net_14766), .A2(net_13073) );
NAND2_X2 inst_9927 ( .ZN(net_9192), .A1(net_9191), .A2(net_6454) );
AOI21_X4 inst_20211 ( .ZN(net_19092), .B2(net_11823), .A(net_11456), .B1(net_333) );
INV_X2 inst_19148 ( .A(net_5613), .ZN(net_4082) );
NAND3_X2 inst_6494 ( .A1(net_20510), .A2(net_14500), .A3(net_14395), .ZN(net_10859) );
NOR2_X4 inst_2919 ( .ZN(net_8082), .A1(net_8081), .A2(net_8080) );
OAI21_X2 inst_1872 ( .ZN(net_13708), .B2(net_13707), .B1(net_7164), .A(net_1831) );
NOR2_X2 inst_5039 ( .A1(net_5120), .ZN(net_2075), .A2(net_1101) );
NAND2_X2 inst_10795 ( .ZN(net_7261), .A1(net_5570), .A2(net_3213) );
NAND2_X2 inst_10827 ( .ZN(net_8971), .A1(net_7489), .A2(net_4058) );
NAND2_X2 inst_12003 ( .A1(net_3060), .ZN(net_2135), .A2(net_305) );
INV_X4 inst_15917 ( .ZN(net_2413), .A(net_1743) );
NOR2_X2 inst_4028 ( .A1(net_11494), .ZN(net_9543), .A2(net_8002) );
CLKBUF_X2 inst_22575 ( .A(net_22446), .Z(net_22447) );
NAND2_X2 inst_8478 ( .ZN(net_17009), .A1(net_17008), .A2(net_17007) );
INV_X4 inst_16658 ( .ZN(net_5265), .A(net_3792) );
INV_X4 inst_17640 ( .ZN(net_6377), .A(net_4850) );
INV_X4 inst_17608 ( .A(net_14029), .ZN(net_512) );
INV_X4 inst_17136 ( .ZN(net_1552), .A(net_764) );
INV_X4 inst_16083 ( .A(net_1548), .ZN(net_1537) );
INV_X4 inst_13556 ( .ZN(net_20313), .A(net_9161) );
INV_X4 inst_18200 ( .A(net_20915), .ZN(net_193) );
NOR2_X4 inst_3119 ( .ZN(net_6848), .A1(net_3199), .A2(net_2744) );
NOR2_X2 inst_3777 ( .ZN(net_13081), .A2(net_11983), .A1(net_10142) );
NOR2_X2 inst_5138 ( .A1(net_279), .A2(net_189), .ZN(net_180) );
INV_X4 inst_18109 ( .A(net_20872), .ZN(net_16357) );
XOR2_X2 inst_29 ( .A(net_21210), .B(net_21114), .Z(net_15587) );
INV_X4 inst_14515 ( .A(net_8515), .ZN(net_7852) );
NAND2_X2 inst_9900 ( .ZN(net_12168), .A2(net_9496), .A1(net_9364) );
DFF_X1 inst_19852 ( .D(net_17191), .CK(net_21759), .Q(x71) );
NAND2_X4 inst_6937 ( .A2(net_19269), .A1(net_19268), .ZN(net_17715) );
NAND2_X2 inst_8469 ( .ZN(net_17156), .A2(net_16695), .A1(net_16542) );
NAND2_X2 inst_7782 ( .ZN(net_20810), .A1(net_20208), .A2(net_18670) );
NAND2_X2 inst_9713 ( .ZN(net_10176), .A1(net_10175), .A2(net_7701) );
INV_X4 inst_16471 ( .ZN(net_4701), .A(net_1429) );
OAI21_X2 inst_2152 ( .ZN(net_9303), .A(net_7514), .B2(net_2964), .B1(net_933) );
NOR2_X2 inst_3947 ( .A1(net_9914), .A2(net_8710), .ZN(net_8620) );
NAND2_X2 inst_10540 ( .ZN(net_8112), .A2(net_5083), .A1(net_4228) );
INV_X4 inst_16232 ( .A(net_6635), .ZN(net_5330) );
NAND2_X2 inst_7740 ( .ZN(net_18800), .A2(net_18769), .A1(net_17810) );
INV_X4 inst_13270 ( .ZN(net_12550), .A(net_11337) );
INV_X4 inst_15712 ( .ZN(net_10664), .A(net_7610) );
NAND2_X2 inst_10590 ( .ZN(net_7932), .A2(net_6670), .A1(net_6655) );
NAND2_X2 inst_11152 ( .ZN(net_4204), .A2(net_4203), .A1(net_809) );
INV_X4 inst_12775 ( .ZN(net_17324), .A(net_17323) );
NAND3_X2 inst_6207 ( .ZN(net_13283), .A1(net_11729), .A3(net_10282), .A2(net_6204) );
AOI22_X2 inst_20040 ( .ZN(net_7117), .A1(net_7116), .B1(net_7115), .A2(net_5488), .B2(net_4236) );
NAND2_X2 inst_11396 ( .A2(net_7667), .ZN(net_6001), .A1(net_1911) );
XNOR2_X2 inst_538 ( .A(net_15798), .ZN(net_1510), .B(net_685) );
CLKBUF_X2 inst_22390 ( .A(net_21595), .Z(net_22262) );
NAND2_X2 inst_8344 ( .A2(net_20207), .A1(net_17485), .ZN(net_17484) );
INV_X4 inst_16277 ( .ZN(net_1808), .A(net_170) );
AOI21_X2 inst_20689 ( .ZN(net_12223), .B2(net_10715), .B1(net_8232), .A(net_4243) );
NOR2_X2 inst_4537 ( .ZN(net_4486), .A2(net_4026), .A1(net_940) );
NAND4_X2 inst_5280 ( .ZN(net_15997), .A2(net_15445), .A1(net_15264), .A4(net_14589), .A3(net_11503) );
CLKBUF_X2 inst_22814 ( .A(net_22685), .Z(net_22686) );
XOR2_X2 inst_35 ( .A(net_21182), .Z(net_687), .B(net_686) );
INV_X2 inst_19558 ( .ZN(net_1487), .A(net_839) );
CLKBUF_X2 inst_21650 ( .A(net_21262), .Z(net_21522) );
NOR2_X2 inst_4765 ( .ZN(net_7161), .A1(net_4301), .A2(net_2979) );
NAND2_X2 inst_8890 ( .ZN(net_15127), .A2(net_14161), .A1(net_14059) );
NAND2_X2 inst_10599 ( .A1(net_10898), .ZN(net_7895), .A2(net_6707) );
CLKBUF_X2 inst_22352 ( .A(net_22223), .Z(net_22224) );
NAND2_X2 inst_11146 ( .A1(net_6968), .ZN(net_6264), .A2(net_4221) );
NOR4_X2 inst_2600 ( .ZN(net_13724), .A1(net_12952), .A2(net_10851), .A3(net_10050), .A4(net_9338) );
INV_X4 inst_14158 ( .ZN(net_13702), .A(net_6020) );
CLKBUF_X2 inst_21633 ( .A(net_21504), .Z(net_21505) );
INV_X4 inst_16990 ( .ZN(net_1229), .A(net_877) );
OAI21_X2 inst_2274 ( .A(net_13734), .ZN(net_7135), .B1(net_5534), .B2(net_3465) );
NAND4_X4 inst_5178 ( .A3(net_19112), .A1(net_19111), .ZN(net_16689), .A4(net_16305), .A2(net_14884) );
NAND2_X2 inst_10055 ( .ZN(net_13161), .A2(net_8689), .A1(net_8138) );
INV_X4 inst_16671 ( .ZN(net_8276), .A(net_761) );
SDFF_X2 inst_695 ( .Q(net_20889), .SE(net_18862), .SI(net_18852), .D(net_545), .CK(net_22046) );
INV_X2 inst_19016 ( .ZN(net_4985), .A(net_4984) );
CLKBUF_X2 inst_22392 ( .A(net_22263), .Z(net_22264) );
AOI21_X2 inst_20465 ( .ZN(net_15001), .B2(net_12996), .B1(net_12339), .A(net_8902) );
NOR2_X2 inst_4038 ( .ZN(net_7910), .A1(net_5901), .A2(net_1634) );
NAND4_X2 inst_5492 ( .A3(net_20239), .A1(net_20238), .ZN(net_19925), .A2(net_12245), .A4(net_12217) );
NAND2_X2 inst_10606 ( .A1(net_10759), .ZN(net_10637), .A2(net_4822) );
NAND2_X2 inst_10663 ( .ZN(net_11854), .A2(net_5285), .A1(net_4292) );
INV_X4 inst_14001 ( .ZN(net_6375), .A(net_6374) );
NAND2_X4 inst_6877 ( .A2(net_20282), .A1(net_20281), .ZN(net_18239) );
NAND2_X2 inst_10782 ( .ZN(net_6966), .A2(net_5613), .A1(net_5594) );
INV_X4 inst_14376 ( .ZN(net_9999), .A(net_5176) );
NAND3_X2 inst_6154 ( .ZN(net_19565), .A2(net_13673), .A3(net_12390), .A1(net_3657) );
NOR2_X2 inst_3559 ( .ZN(net_12979), .A2(net_10184), .A1(net_8004) );
INV_X4 inst_17790 ( .ZN(net_673), .A(net_232) );
INV_X4 inst_17306 ( .ZN(net_5277), .A(net_4394) );
NAND3_X2 inst_5720 ( .ZN(net_20611), .A3(net_15704), .A2(net_15072), .A1(net_13809) );
INV_X8 inst_12277 ( .ZN(net_2315), .A(net_984) );
INV_X4 inst_17688 ( .A(net_20875), .ZN(net_1614) );
NAND2_X2 inst_9449 ( .A2(net_12528), .ZN(net_11525), .A1(net_7885) );
INV_X4 inst_17386 ( .ZN(net_5308), .A(net_1740) );
NAND2_X4 inst_7183 ( .A1(net_20008), .ZN(net_19492), .A2(net_4264) );
CLKBUF_X2 inst_22348 ( .A(net_22219), .Z(net_22220) );
NAND2_X2 inst_8328 ( .ZN(net_20596), .A2(net_18704), .A1(net_17216) );
NAND2_X2 inst_11772 ( .A2(net_3776), .ZN(net_3622), .A1(net_2646) );
INV_X4 inst_12790 ( .A(net_17852), .ZN(net_17286) );
INV_X4 inst_16315 ( .ZN(net_14694), .A(net_14171) );
NAND3_X2 inst_6001 ( .ZN(net_14431), .A3(net_12549), .A1(net_8888), .A2(net_8799) );
NAND2_X4 inst_7004 ( .ZN(net_17341), .A1(net_16737), .A2(net_16591) );
INV_X4 inst_12506 ( .ZN(net_18642), .A(net_18640) );
INV_X4 inst_18268 ( .A(net_19449), .ZN(net_19445) );
INV_X4 inst_16995 ( .ZN(net_1070), .A(net_816) );
NAND2_X2 inst_8193 ( .ZN(net_17895), .A2(net_17894), .A1(net_17832) );
INV_X2 inst_19102 ( .ZN(net_4532), .A(net_4531) );
INV_X4 inst_14086 ( .ZN(net_11179), .A(net_6210) );
NAND2_X2 inst_11646 ( .ZN(net_2482), .A2(net_2178), .A1(net_168) );
NAND2_X2 inst_10751 ( .ZN(net_5702), .A1(net_5701), .A2(net_5700) );
NAND2_X2 inst_11525 ( .ZN(net_20087), .A1(net_2974), .A2(net_2973) );
NAND2_X2 inst_10666 ( .A2(net_11220), .ZN(net_6272), .A1(net_4154) );
NAND3_X2 inst_6592 ( .ZN(net_9960), .A2(net_9959), .A3(net_9958), .A1(net_3204) );
NAND2_X4 inst_7209 ( .ZN(net_11983), .A2(net_7941), .A1(net_6074) );
INV_X4 inst_14865 ( .ZN(net_7258), .A(net_3323) );
NAND4_X4 inst_5217 ( .A4(net_20295), .A1(net_20294), .ZN(net_16622), .A3(net_16068), .A2(net_13997) );
NAND2_X2 inst_8069 ( .ZN(net_18178), .A2(net_18135), .A1(net_17097) );
INV_X4 inst_15307 ( .ZN(net_3396), .A(net_2212) );
NOR2_X2 inst_4600 ( .ZN(net_8575), .A1(net_6719), .A2(net_1578) );
NOR2_X2 inst_3872 ( .A1(net_11678), .ZN(net_11546), .A2(net_6612) );
NAND2_X4 inst_6923 ( .ZN(net_17784), .A1(net_17584), .A2(net_17518) );
NAND2_X2 inst_9273 ( .ZN(net_12601), .A2(net_10845), .A1(net_10386) );
NAND2_X2 inst_11574 ( .ZN(net_5490), .A2(net_2744), .A1(net_2409) );
CLKBUF_X2 inst_21617 ( .A(net_21397), .Z(net_21489) );
INV_X4 inst_17067 ( .A(net_1415), .ZN(net_1169) );
NAND2_X2 inst_10227 ( .A1(net_9466), .ZN(net_8059), .A2(net_6129) );
INV_X4 inst_17849 ( .ZN(net_96), .A(net_95) );
OAI21_X4 inst_1411 ( .B2(net_19007), .B1(net_19006), .A(net_16390), .ZN(net_16175) );
XNOR2_X2 inst_149 ( .ZN(net_18036), .A(net_17992), .B(net_17663) );
NAND2_X2 inst_11028 ( .A1(net_5458), .ZN(net_4776), .A2(net_3494) );
INV_X4 inst_12527 ( .ZN(net_18430), .A(net_18429) );
INV_X4 inst_18048 ( .A(net_20948), .ZN(net_268) );
NAND2_X2 inst_8854 ( .ZN(net_15364), .A1(net_15217), .A2(net_14368) );
AOI21_X2 inst_20623 ( .ZN(net_13474), .B2(net_12417), .B1(net_7988), .A(net_6035) );
NAND2_X4 inst_6924 ( .ZN(net_17782), .A1(net_17587), .A2(net_17519) );
INV_X4 inst_18134 ( .A(net_20918), .ZN(net_301) );
NAND2_X2 inst_9542 ( .ZN(net_13744), .A2(net_11054), .A1(net_6840) );
NAND2_X2 inst_7771 ( .ZN(net_18742), .A2(net_18741), .A1(net_17439) );
INV_X4 inst_15608 ( .A(net_7659), .ZN(net_7115) );
OAI21_X2 inst_2320 ( .A(net_13542), .ZN(net_5669), .B2(net_5288), .B1(net_1036) );
INV_X4 inst_15203 ( .ZN(net_3661), .A(net_2236) );
CLKBUF_X2 inst_21519 ( .A(net_21390), .Z(net_21391) );
INV_X4 inst_17582 ( .A(net_14022), .ZN(net_843) );
OAI211_X2 inst_2534 ( .C1(net_13576), .ZN(net_11259), .A(net_11258), .B(net_11257), .C2(net_10008) );
INV_X4 inst_17527 ( .A(net_2585), .ZN(net_1099) );
INV_X2 inst_19702 ( .A(net_20923), .ZN(net_20565) );
NAND4_X2 inst_5377 ( .ZN(net_19535), .A3(net_13888), .A4(net_13704), .A1(net_11409), .A2(net_11200) );
NAND2_X2 inst_10775 ( .A2(net_7149), .ZN(net_7016), .A1(net_1620) );
NOR2_X2 inst_3737 ( .ZN(net_10719), .A1(net_10718), .A2(net_7843) );
OAI21_X2 inst_1636 ( .ZN(net_15962), .B1(net_15369), .B2(net_15281), .A(net_12853) );
CLKBUF_X2 inst_22530 ( .A(net_22023), .Z(net_22402) );
CLKBUF_X2 inst_21421 ( .A(net_21292), .Z(net_21293) );
AOI21_X2 inst_20276 ( .B1(net_21236), .ZN(net_16327), .B2(net_16081), .A(net_15757) );
XNOR2_X2 inst_515 ( .ZN(net_5790), .A(net_5789), .B(net_5788) );
NAND2_X2 inst_8501 ( .ZN(net_17068), .A2(net_16604), .A1(net_16471) );
AOI21_X2 inst_20349 ( .ZN(net_15750), .A(net_15602), .B2(net_15042), .B1(net_4274) );
OAI21_X4 inst_1501 ( .B1(net_19379), .ZN(net_13851), .A(net_10113), .B2(net_10068) );
NAND2_X4 inst_7278 ( .ZN(net_9739), .A2(net_5845), .A1(net_2537) );
INV_X8 inst_12242 ( .ZN(net_5333), .A(net_1945) );
NOR2_X4 inst_3212 ( .A2(net_20495), .A1(net_4216), .ZN(net_3824) );
INV_X4 inst_14982 ( .ZN(net_3414), .A(net_3413) );
OAI21_X2 inst_1584 ( .A(net_21228), .ZN(net_16297), .B2(net_15994), .B1(net_15035) );
INV_X4 inst_14183 ( .A(net_7833), .ZN(net_5986) );
NAND2_X2 inst_9361 ( .ZN(net_12149), .A2(net_9889), .A1(net_7394) );
CLKBUF_X2 inst_21896 ( .A(net_21767), .Z(net_21768) );
AOI21_X2 inst_20636 ( .ZN(net_13339), .A(net_10797), .B2(net_9267), .B1(net_5536) );
NAND2_X2 inst_7933 ( .ZN(net_20153), .A2(net_18350), .A1(net_16998) );
NAND2_X2 inst_11023 ( .ZN(net_5954), .A1(net_4792), .A2(net_4791) );
CLKBUF_X2 inst_21882 ( .A(net_21753), .Z(net_21754) );
INV_X4 inst_15499 ( .A(net_13462), .ZN(net_7246) );
NAND2_X2 inst_8129 ( .A2(net_20880), .ZN(net_18045), .A1(net_16004) );
NOR2_X4 inst_2933 ( .ZN(net_9129), .A2(net_7459), .A1(net_1254) );
NAND3_X2 inst_6467 ( .ZN(net_11358), .A3(net_11357), .A2(net_6436), .A1(net_3691) );
NAND2_X2 inst_8706 ( .A2(net_20968), .A1(net_19992), .ZN(net_16298) );
INV_X4 inst_14641 ( .ZN(net_5670), .A(net_4377) );
NOR3_X2 inst_2713 ( .ZN(net_20148), .A1(net_12379), .A3(net_12259), .A2(net_8015) );
SDFF_X2 inst_1008 ( .QN(net_21083), .D(net_729), .SE(net_263), .CK(net_22578), .SI(x1674) );
XNOR2_X2 inst_559 ( .B(net_17262), .A(net_16644), .ZN(net_685) );
NAND2_X2 inst_7877 ( .ZN(net_18530), .A2(net_18479), .A1(net_18452) );
NAND2_X2 inst_8872 ( .ZN(net_15260), .A2(net_14668), .A1(net_10061) );
AOI21_X4 inst_20187 ( .B1(net_20715), .B2(net_15345), .ZN(net_15216), .A(net_14446) );
NAND3_X2 inst_6725 ( .ZN(net_6504), .A1(net_6487), .A3(net_5055), .A2(net_4828) );
NAND2_X2 inst_7706 ( .ZN(net_18869), .A2(net_18866), .A1(net_7388) );
NAND2_X2 inst_9476 ( .ZN(net_20636), .A2(net_12900), .A1(net_5779) );
NAND2_X2 inst_11596 ( .ZN(net_4801), .A2(net_3165), .A1(net_2671) );
INV_X2 inst_19012 ( .A(net_6672), .ZN(net_5004) );
NAND2_X2 inst_9250 ( .ZN(net_12667), .A2(net_12666), .A1(net_10398) );
INV_X4 inst_14940 ( .ZN(net_4610), .A(net_3532) );
AND2_X4 inst_21240 ( .A1(net_10714), .ZN(net_3072), .A2(net_3071) );
INV_X2 inst_18933 ( .ZN(net_8518), .A(net_5842) );
INV_X4 inst_16818 ( .ZN(net_997), .A(net_996) );
NOR2_X2 inst_3405 ( .A2(net_20249), .A1(net_20248), .ZN(net_19472) );
INV_X2 inst_19616 ( .A(net_21105), .ZN(net_42) );
NOR2_X2 inst_3888 ( .ZN(net_9244), .A2(net_5961), .A1(net_2310) );
NAND2_X2 inst_8979 ( .ZN(net_14506), .A2(net_12961), .A1(net_2484) );
INV_X4 inst_12831 ( .ZN(net_19974), .A(net_17138) );
CLKBUF_X2 inst_21500 ( .A(net_21368), .Z(net_21372) );
NAND2_X2 inst_9797 ( .A1(net_12968), .ZN(net_9706), .A2(net_9705) );
NAND2_X4 inst_7366 ( .ZN(net_5111), .A1(net_4272), .A2(net_3491) );
INV_X8 inst_12221 ( .ZN(net_9801), .A(net_5177) );
INV_X4 inst_15275 ( .ZN(net_14990), .A(net_6528) );
NOR2_X2 inst_4334 ( .ZN(net_7433), .A1(net_6812), .A2(net_5739) );
NAND2_X2 inst_8017 ( .A2(net_18283), .ZN(net_18281), .A1(net_17156) );
OR2_X4 inst_1075 ( .A1(net_13416), .A2(net_9955), .ZN(net_8314) );
INV_X2 inst_19038 ( .ZN(net_4830), .A(net_4829) );
CLKBUF_X2 inst_22655 ( .A(net_22526), .Z(net_22527) );
NAND2_X2 inst_9230 ( .ZN(net_20131), .A2(net_10411), .A1(net_7963) );
INV_X4 inst_12701 ( .ZN(net_17834), .A(net_17610) );
OAI21_X2 inst_2257 ( .A(net_12669), .ZN(net_7257), .B2(net_7256), .B1(net_2414) );
NAND2_X2 inst_11504 ( .ZN(net_3981), .A1(net_3426), .A2(net_3061) );
NAND2_X2 inst_11781 ( .ZN(net_6399), .A1(net_1790), .A2(net_1136) );
INV_X4 inst_16183 ( .ZN(net_1871), .A(net_1425) );
INV_X4 inst_15278 ( .ZN(net_5010), .A(net_2741) );
INV_X4 inst_13641 ( .ZN(net_10351), .A(net_8176) );
INV_X4 inst_14306 ( .ZN(net_6094), .A(net_5505) );
INV_X4 inst_15553 ( .A(net_12440), .ZN(net_8798) );
CLKBUF_X2 inst_22612 ( .A(net_22483), .Z(net_22484) );
CLKBUF_X2 inst_21626 ( .A(net_21349), .Z(net_21498) );
INV_X4 inst_15210 ( .ZN(net_2895), .A(net_2894) );
NAND3_X2 inst_6536 ( .A3(net_14544), .ZN(net_10581), .A2(net_10580), .A1(net_6782) );
NAND3_X2 inst_6110 ( .ZN(net_13890), .A3(net_13851), .A2(net_11929), .A1(net_9767) );
NAND3_X2 inst_6434 ( .ZN(net_11833), .A3(net_11832), .A2(net_10562), .A1(net_6943) );
XNOR2_X2 inst_494 ( .ZN(net_9195), .A(net_9194), .B(net_9193) );
XNOR2_X2 inst_329 ( .B(net_21114), .ZN(net_17308), .A(net_16983) );
CLKBUF_X2 inst_21934 ( .A(net_21805), .Z(net_21806) );
INV_X4 inst_17823 ( .ZN(net_271), .A(net_109) );
NAND3_X2 inst_5942 ( .ZN(net_14901), .A2(net_14900), .A3(net_14863), .A1(net_11331) );
OAI21_X2 inst_2347 ( .B2(net_4378), .ZN(net_4213), .A(net_3016), .B1(net_2720) );
INV_X4 inst_13845 ( .ZN(net_11023), .A(net_7476) );
INV_X4 inst_13085 ( .ZN(net_18970), .A(net_15938) );
INV_X4 inst_17117 ( .ZN(net_1353), .A(net_781) );
INV_X4 inst_14167 ( .A(net_12215), .ZN(net_6008) );
CLKBUF_X2 inst_22686 ( .A(net_22557), .Z(net_22558) );
NOR2_X4 inst_2894 ( .ZN(net_10912), .A1(net_9321), .A2(net_8341) );
CLKBUF_X2 inst_21452 ( .A(net_21321), .Z(net_21324) );
NAND3_X2 inst_5949 ( .A3(net_20427), .ZN(net_19785), .A2(net_14270), .A1(net_11414) );
NAND2_X4 inst_7045 ( .ZN(net_16491), .A1(net_16354), .A2(net_16221) );
NAND3_X2 inst_6085 ( .ZN(net_13958), .A3(net_11155), .A2(net_5671), .A1(net_4412) );
NAND2_X2 inst_10192 ( .A2(net_13876), .ZN(net_8153), .A1(net_8152) );
NOR2_X4 inst_2959 ( .ZN(net_8015), .A2(net_6733), .A1(net_6732) );
INV_X4 inst_15130 ( .ZN(net_4117), .A(net_3135) );
INV_X2 inst_18474 ( .ZN(net_12652), .A(net_12651) );
INV_X4 inst_13906 ( .A(net_10618), .ZN(net_8896) );
INV_X2 inst_19194 ( .ZN(net_6273), .A(net_4409) );
OAI21_X2 inst_1683 ( .ZN(net_20159), .A(net_14769), .B2(net_14422), .B1(net_11139) );
NAND2_X2 inst_10714 ( .ZN(net_19753), .A1(net_6028), .A2(net_3387) );
NOR2_X2 inst_3865 ( .ZN(net_9385), .A2(net_9384), .A1(net_7452) );
INV_X4 inst_18003 ( .A(net_21089), .ZN(net_707) );
AOI21_X2 inst_20915 ( .B2(net_10630), .A(net_10022), .ZN(net_7332), .B1(net_3066) );
INV_X4 inst_16983 ( .ZN(net_2137), .A(net_445) );
NAND2_X2 inst_10459 ( .ZN(net_7019), .A1(net_7018), .A2(net_4101) );
INV_X4 inst_13109 ( .ZN(net_15673), .A(net_15473) );
NAND2_X2 inst_9896 ( .ZN(net_12171), .A1(net_9367), .A2(net_4823) );
INV_X4 inst_15099 ( .ZN(net_3229), .A(net_3228) );
NOR2_X2 inst_3543 ( .ZN(net_13317), .A2(net_10346), .A1(net_9030) );
INV_X4 inst_15486 ( .ZN(net_14472), .A(net_11550) );
NAND3_X2 inst_6712 ( .ZN(net_7102), .A2(net_4216), .A3(net_4060), .A1(net_3892) );
NAND2_X2 inst_10737 ( .A1(net_5785), .ZN(net_5762), .A2(net_4732) );
NAND2_X2 inst_11361 ( .ZN(net_3611), .A2(net_3472), .A1(net_2953) );
INV_X4 inst_13867 ( .ZN(net_12501), .A(net_7452) );
NAND2_X2 inst_8158 ( .ZN(net_17987), .A2(net_17931), .A1(net_17885) );
INV_X4 inst_15080 ( .A(net_14279), .ZN(net_13348) );
INV_X8 inst_12423 ( .A(net_20910), .ZN(net_234) );
AND2_X4 inst_21173 ( .ZN(net_19526), .A2(net_12665), .A1(net_9738) );
NOR2_X2 inst_3461 ( .ZN(net_14683), .A2(net_13163), .A1(net_1052) );
NAND2_X2 inst_10974 ( .ZN(net_4968), .A2(net_2668), .A1(net_86) );
NAND2_X2 inst_9754 ( .ZN(net_10027), .A2(net_10026), .A1(net_5578) );
NOR2_X2 inst_4969 ( .A1(net_6712), .ZN(net_3153), .A2(net_1588) );
NAND2_X2 inst_8546 ( .A2(net_19452), .ZN(net_16809), .A1(net_16808) );
CLKBUF_X2 inst_22275 ( .A(net_22146), .Z(net_22147) );
INV_X2 inst_18409 ( .ZN(net_16350), .A(net_16289) );
NOR2_X2 inst_4692 ( .ZN(net_8581), .A1(net_3929), .A2(net_3178) );
NAND2_X2 inst_8244 ( .ZN(net_17801), .A1(net_17553), .A2(net_17465) );
NOR2_X2 inst_4883 ( .ZN(net_2172), .A1(net_1216), .A2(net_1035) );
CLKBUF_X2 inst_22628 ( .A(net_21851), .Z(net_22500) );
AOI21_X2 inst_20933 ( .B1(net_6867), .ZN(net_6547), .A(net_4177), .B2(net_2939) );
NAND2_X2 inst_10487 ( .ZN(net_6935), .A1(net_6934), .A2(net_6468) );
NAND2_X2 inst_8580 ( .ZN(net_16723), .A1(net_16689), .A2(net_16576) );
NAND2_X4 inst_7538 ( .A1(net_19418), .ZN(net_1924), .A2(net_786) );
CLKBUF_X2 inst_22674 ( .A(net_22545), .Z(net_22546) );
CLKBUF_X2 inst_22432 ( .A(net_21393), .Z(net_22304) );
OAI21_X2 inst_2178 ( .ZN(net_8869), .A(net_8868), .B2(net_8867), .B1(net_1706) );
XNOR2_X2 inst_185 ( .ZN(net_17822), .A(net_17762), .B(net_17517) );
NAND2_X2 inst_9498 ( .A2(net_12847), .A1(net_11617), .ZN(net_11427) );
AND2_X2 inst_21320 ( .ZN(net_7003), .A1(net_7002), .A2(net_5158) );
INV_X4 inst_17474 ( .ZN(net_3033), .A(net_252) );
XNOR2_X2 inst_166 ( .B(net_21129), .ZN(net_17835), .A(net_17834) );
NOR2_X2 inst_3815 ( .ZN(net_9820), .A2(net_9819), .A1(net_9368) );
NOR2_X2 inst_4786 ( .ZN(net_4011), .A2(net_2836), .A1(net_573) );
INV_X4 inst_12617 ( .A(net_20912), .ZN(net_18067) );
INV_X4 inst_13822 ( .A(net_9388), .ZN(net_7509) );
OAI21_X2 inst_1757 ( .ZN(net_14787), .A(net_14563), .B2(net_13271), .B1(net_6831) );
CLKBUF_X2 inst_21548 ( .A(net_21300), .Z(net_21420) );
NOR2_X2 inst_3851 ( .ZN(net_9530), .A1(net_9529), .A2(net_7574) );
NAND3_X2 inst_6370 ( .A1(net_12737), .ZN(net_12064), .A2(net_12063), .A3(net_10655) );
NAND3_X2 inst_6772 ( .ZN(net_5150), .A2(net_5149), .A3(net_2798), .A1(net_1742) );
INV_X8 inst_12358 ( .A(net_20901), .ZN(net_987) );
INV_X4 inst_15683 ( .ZN(net_3695), .A(net_2038) );
INV_X4 inst_16143 ( .ZN(net_4655), .A(net_1523) );
CLKBUF_X2 inst_22699 ( .A(net_22570), .Z(net_22571) );
NAND3_X2 inst_6359 ( .ZN(net_12089), .A2(net_12088), .A3(net_11824), .A1(net_11077) );
NAND2_X2 inst_12026 ( .ZN(net_5511), .A2(net_1065), .A1(x7654) );
OAI21_X2 inst_1605 ( .A(net_20872), .B2(net_20203), .B1(net_20202), .ZN(net_19603) );
INV_X4 inst_18280 ( .ZN(net_20072), .A(net_20068) );
NAND2_X2 inst_10206 ( .ZN(net_8116), .A1(net_8115), .A2(net_4650) );
NAND2_X2 inst_11635 ( .ZN(net_4249), .A2(net_2519), .A1(net_2179) );
INV_X4 inst_13593 ( .ZN(net_11178), .A(net_8791) );
INV_X2 inst_18518 ( .A(net_14535), .ZN(net_11545) );
NOR2_X2 inst_4649 ( .ZN(net_4470), .A1(net_3356), .A2(net_3355) );
INV_X4 inst_14508 ( .ZN(net_7847), .A(net_6591) );
INV_X2 inst_18462 ( .ZN(net_18948), .A(net_11803) );
INV_X4 inst_12904 ( .ZN(net_19151), .A(net_16549) );
NAND2_X2 inst_10558 ( .ZN(net_10472), .A2(net_5070), .A1(net_4430) );
INV_X4 inst_17975 ( .A(net_21152), .ZN(net_17404) );
INV_X4 inst_12922 ( .ZN(net_16859), .A(net_16688) );
INV_X4 inst_17774 ( .A(net_161), .ZN(net_150) );
NAND4_X2 inst_5308 ( .ZN(net_15795), .A4(net_14787), .A1(net_13066), .A3(net_12115), .A2(net_9927) );
INV_X4 inst_15770 ( .A(net_15699), .ZN(net_15612) );
INV_X4 inst_14634 ( .ZN(net_9502), .A(net_4385) );
AOI22_X2 inst_20017 ( .ZN(net_11233), .A2(net_9680), .B1(net_9537), .B2(net_5856), .A1(net_308) );
NOR2_X2 inst_4475 ( .ZN(net_8429), .A1(net_3820), .A2(net_703) );
INV_X4 inst_17059 ( .ZN(net_1213), .A(net_821) );
CLKBUF_X2 inst_22801 ( .A(net_22672), .Z(net_22673) );
NAND2_X2 inst_7757 ( .ZN(net_18766), .A2(net_18742), .A1(net_18714) );
NAND2_X2 inst_11077 ( .ZN(net_4472), .A1(net_2744), .A2(net_2605) );
INV_X4 inst_16837 ( .ZN(net_1535), .A(net_1343) );
INV_X4 inst_15925 ( .ZN(net_2208), .A(net_1737) );
INV_X4 inst_17514 ( .ZN(net_6982), .A(net_4394) );
NAND4_X4 inst_5201 ( .A4(net_19970), .A1(net_19969), .ZN(net_16577), .A3(net_15884), .A2(net_7684) );
INV_X4 inst_14831 ( .A(net_5527), .ZN(net_4756) );
INV_X4 inst_16121 ( .ZN(net_1489), .A(net_1488) );
INV_X4 inst_16705 ( .A(net_7976), .ZN(net_6702) );
OAI211_X4 inst_2373 ( .C2(net_20920), .C1(net_19094), .ZN(net_16552), .B(net_16171), .A(net_8065) );
NAND2_X2 inst_11436 ( .ZN(net_3508), .A1(net_2007), .A2(net_1064) );
INV_X4 inst_15321 ( .ZN(net_3533), .A(net_2631) );
OAI221_X2 inst_1331 ( .ZN(net_19835), .C1(net_15688), .B1(net_14990), .C2(net_14438), .A(net_12791), .B2(net_12175) );
NAND2_X2 inst_9215 ( .ZN(net_18999), .A2(net_11390), .A1(net_5528) );
NAND2_X4 inst_7604 ( .A1(net_19340), .ZN(net_3101), .A2(net_1347) );
INV_X8 inst_12322 ( .ZN(net_1264), .A(net_131) );
INV_X4 inst_15779 ( .ZN(net_8179), .A(net_6963) );
NAND2_X4 inst_7404 ( .A2(net_20536), .ZN(net_5781), .A1(net_4016) );
NOR2_X4 inst_3223 ( .ZN(net_3395), .A1(net_3068), .A2(net_2597) );
NOR2_X2 inst_3560 ( .ZN(net_12978), .A1(net_12681), .A2(net_10391) );
NOR3_X2 inst_2683 ( .ZN(net_19367), .A2(net_12333), .A1(net_10424), .A3(net_9204) );
INV_X4 inst_13736 ( .ZN(net_7655), .A(net_5777) );
AOI21_X2 inst_20539 ( .A(net_15048), .ZN(net_14482), .B2(net_11680), .B1(net_10079) );
INV_X4 inst_17442 ( .ZN(net_3862), .A(net_3800) );
NOR2_X2 inst_4223 ( .ZN(net_13005), .A2(net_7204), .A1(net_1378) );
AND2_X2 inst_21318 ( .ZN(net_7039), .A1(net_5275), .A2(net_5155) );
INV_X4 inst_18235 ( .A(net_21154), .ZN(net_16833) );
INV_X4 inst_16910 ( .ZN(net_20457), .A(net_940) );
INV_X4 inst_14152 ( .A(net_8189), .ZN(net_6027) );
INV_X4 inst_14277 ( .A(net_12238), .ZN(net_9374) );
INV_X4 inst_17182 ( .ZN(net_951), .A(net_143) );
INV_X2 inst_19255 ( .ZN(net_4241), .A(net_2226) );
INV_X4 inst_13283 ( .ZN(net_12434), .A(net_11160) );
NAND3_X2 inst_6677 ( .ZN(net_7749), .A2(net_7748), .A3(net_3878), .A1(net_2978) );
CLKBUF_X2 inst_21383 ( .A(net_21254), .Z(net_21255) );
CLKBUF_X2 inst_21784 ( .A(net_21655), .Z(net_21656) );
INV_X4 inst_15931 ( .ZN(net_1729), .A(net_1728) );
OAI21_X2 inst_1910 ( .A(net_14038), .ZN(net_13087), .B1(net_9412), .B2(net_6977) );
INV_X4 inst_13420 ( .ZN(net_10250), .A(net_10249) );
INV_X4 inst_14461 ( .ZN(net_6086), .A(net_4940) );
INV_X4 inst_16091 ( .A(net_2321), .ZN(net_1525) );
AND2_X4 inst_21225 ( .A1(net_13554), .A2(net_9931), .ZN(net_5192) );
NAND2_X2 inst_10272 ( .ZN(net_7971), .A2(net_6215), .A1(net_4931) );
NAND2_X2 inst_9265 ( .ZN(net_14270), .A2(net_12303), .A1(net_9109) );
NOR2_X4 inst_3115 ( .ZN(net_5083), .A2(net_4022), .A1(net_3056) );
NAND3_X2 inst_5814 ( .ZN(net_15643), .A1(net_15033), .A2(net_13234), .A3(net_10746) );
INV_X4 inst_15887 ( .A(net_14759), .ZN(net_14572) );
NOR2_X4 inst_3219 ( .ZN(net_2703), .A2(net_2702), .A1(net_809) );
NAND2_X2 inst_10867 ( .A2(net_20541), .ZN(net_9045), .A1(net_5400) );
NAND3_X2 inst_5673 ( .ZN(net_16370), .A3(net_16159), .A1(net_14973), .A2(net_12754) );
NAND2_X2 inst_10025 ( .ZN(net_8760), .A1(net_8759), .A2(net_8758) );
INV_X2 inst_18659 ( .ZN(net_9202), .A(net_9201) );
OAI21_X2 inst_1991 ( .ZN(net_12008), .A(net_12007), .B1(net_12006), .B2(net_11841) );
INV_X4 inst_14872 ( .ZN(net_6317), .A(net_3692) );
INV_X4 inst_13054 ( .A(net_16479), .ZN(net_16378) );
NOR2_X4 inst_3066 ( .ZN(net_5993), .A1(net_4833), .A2(net_896) );
NAND2_X2 inst_7861 ( .ZN(net_18561), .A2(net_18528), .A1(net_18509) );
AOI21_X2 inst_20312 ( .ZN(net_16012), .B1(net_16011), .B2(net_15426), .A(net_14901) );
INV_X4 inst_14129 ( .ZN(net_7524), .A(net_6111) );
INV_X4 inst_15441 ( .ZN(net_3295), .A(net_2014) );
CLKBUF_X2 inst_21901 ( .A(net_21554), .Z(net_21773) );
NAND2_X2 inst_11630 ( .ZN(net_3838), .A2(net_2232), .A1(net_1080) );
NAND2_X4 inst_7419 ( .A2(net_20492), .ZN(net_5598), .A1(net_2285) );
NAND3_X2 inst_6771 ( .ZN(net_5258), .A3(net_4677), .A2(net_4306), .A1(net_2999) );
NOR2_X2 inst_4703 ( .A1(net_9254), .ZN(net_4128), .A2(net_3169) );
NAND3_X2 inst_6640 ( .ZN(net_8950), .A3(net_8949), .A1(net_6694), .A2(net_3316) );
NAND2_X2 inst_8173 ( .ZN(net_17948), .A1(net_17857), .A2(net_17796) );
NOR3_X2 inst_2672 ( .ZN(net_14816), .A2(net_14274), .A3(net_12389), .A1(net_10923) );
NOR2_X2 inst_3527 ( .ZN(net_13597), .A2(net_13596), .A1(net_13571) );
INV_X4 inst_13924 ( .ZN(net_8192), .A(net_5546) );
INV_X4 inst_13637 ( .ZN(net_11792), .A(net_8192) );
AOI21_X4 inst_20245 ( .ZN(net_11302), .B2(net_9981), .B1(net_8580), .A(net_495) );
NAND2_X2 inst_9558 ( .ZN(net_14276), .A1(net_11236), .A2(net_11023) );
NAND3_X2 inst_6045 ( .ZN(net_14258), .A3(net_12365), .A2(net_8947), .A1(net_7445) );
NOR2_X2 inst_3764 ( .ZN(net_20151), .A2(net_6771), .A1(net_6213) );
NAND3_X2 inst_6408 ( .ZN(net_11965), .A2(net_11964), .A1(net_9961), .A3(net_9375) );
NAND2_X2 inst_9042 ( .ZN(net_20015), .A2(net_12020), .A1(net_1663) );
NAND2_X2 inst_8764 ( .A1(net_16242), .ZN(net_15882), .A2(net_15645) );
NAND2_X2 inst_11912 ( .A2(net_9090), .ZN(net_1553), .A1(net_1552) );
NAND2_X4 inst_7330 ( .ZN(net_6155), .A2(net_4826), .A1(net_885) );
INV_X4 inst_13101 ( .ZN(net_15826), .A(net_15648) );
NAND2_X4 inst_7581 ( .ZN(net_3023), .A2(net_1581), .A1(net_247) );
OAI21_X2 inst_2340 ( .B1(net_5402), .ZN(net_4674), .A(net_4673), .B2(net_2103) );
AND2_X2 inst_21368 ( .ZN(net_344), .A2(net_123), .A1(net_46) );
INV_X4 inst_17589 ( .ZN(net_343), .A(net_108) );
INV_X4 inst_18324 ( .A(net_20923), .ZN(net_20539) );
INV_X4 inst_15492 ( .ZN(net_19491), .A(net_2433) );
INV_X4 inst_17496 ( .ZN(net_3120), .A(net_167) );
CLKBUF_X2 inst_22062 ( .A(net_21933), .Z(net_21934) );
INV_X4 inst_18027 ( .A(net_21230), .ZN(net_60) );
XOR2_X2 inst_16 ( .B(net_21138), .A(net_20513), .Z(net_17021) );
INV_X2 inst_18562 ( .A(net_11532), .ZN(net_10795) );
INV_X4 inst_15362 ( .ZN(net_3478), .A(net_2579) );
INV_X4 inst_14173 ( .ZN(net_11281), .A(net_5353) );
CLKBUF_X2 inst_22462 ( .A(net_21955), .Z(net_22334) );
XNOR2_X2 inst_156 ( .ZN(net_17984), .B(net_17958), .A(net_17861) );
NOR2_X4 inst_2808 ( .ZN(net_17811), .A1(net_17560), .A2(net_17486) );
AOI211_X2 inst_21025 ( .ZN(net_14609), .C2(net_12460), .C1(net_10536), .A(net_9870), .B(net_8800) );
INV_X4 inst_17530 ( .ZN(net_6571), .A(net_117) );
CLKBUF_X2 inst_22805 ( .A(net_21373), .Z(net_22677) );
NAND3_X2 inst_6239 ( .ZN(net_19246), .A3(net_12172), .A1(net_8626), .A2(net_7994) );
AOI21_X4 inst_20149 ( .B2(net_19612), .B1(net_19611), .ZN(net_19517), .A(net_789) );
NOR2_X2 inst_3442 ( .ZN(net_20325), .A2(net_13905), .A1(net_10554) );
NOR3_X2 inst_2693 ( .ZN(net_14223), .A2(net_14222), .A1(net_12645), .A3(net_10996) );
INV_X4 inst_14920 ( .ZN(net_19483), .A(net_3562) );
INV_X4 inst_17228 ( .ZN(net_683), .A(net_279) );
NAND2_X2 inst_10307 ( .ZN(net_7863), .A1(net_7862), .A2(net_5919) );
INV_X4 inst_18133 ( .A(net_21072), .ZN(net_563) );
NAND4_X2 inst_5380 ( .ZN(net_15060), .A4(net_13852), .A2(net_13545), .A1(net_13330), .A3(net_12833) );
INV_X4 inst_14838 ( .ZN(net_4841), .A(net_3132) );
NAND2_X2 inst_10936 ( .A1(net_9785), .ZN(net_7338), .A2(net_3006) );
NAND3_X2 inst_6473 ( .ZN(net_11288), .A1(net_8519), .A2(net_7586), .A3(net_6195) );
OAI21_X2 inst_1549 ( .ZN(net_17732), .A(net_17471), .B1(net_17470), .B2(net_17469) );
NOR2_X4 inst_3020 ( .A2(net_20548), .A1(net_19911), .ZN(net_7235) );
NAND3_X2 inst_6186 ( .A3(net_20625), .A1(net_20624), .ZN(net_13468), .A2(net_9526) );
NAND2_X2 inst_9239 ( .ZN(net_12693), .A2(net_10850), .A1(net_8252) );
INV_X4 inst_12894 ( .ZN(net_17658), .A(net_16864) );
NAND2_X2 inst_10576 ( .A2(net_14222), .A1(net_12864), .ZN(net_6687) );
INV_X4 inst_13477 ( .ZN(net_11638), .A(net_10190) );
SDFF_X2 inst_821 ( .Q(net_21209), .SI(net_17671), .SE(net_125), .CK(net_22448), .D(x5853) );
NOR2_X4 inst_2881 ( .ZN(net_20641), .A2(net_19821), .A1(net_8891) );
NAND2_X2 inst_9113 ( .A1(net_14242), .ZN(net_13579), .A2(net_12335) );
NAND2_X2 inst_8879 ( .A1(net_15214), .ZN(net_15194), .A2(net_14527) );
INV_X4 inst_16225 ( .A(net_1826), .ZN(net_1381) );
SDFF_X2 inst_980 ( .QN(net_21103), .D(net_346), .SE(net_263), .CK(net_21768), .SI(x1354) );
INV_X4 inst_15750 ( .ZN(net_1943), .A(net_1942) );
CLKBUF_X2 inst_22942 ( .A(net_22813), .Z(net_22814) );
CLKBUF_X2 inst_21861 ( .A(net_21732), .Z(net_21733) );
AOI22_X2 inst_19994 ( .ZN(net_14553), .A1(net_14552), .B1(net_14551), .A2(net_11931), .B2(net_9506) );
INV_X4 inst_16021 ( .ZN(net_2307), .A(net_933) );
NAND2_X2 inst_8486 ( .ZN(net_20188), .A1(net_16808), .A2(net_16638) );
AOI21_X4 inst_20142 ( .ZN(net_20607), .B1(net_18881), .B2(net_15178), .A(net_10489) );
INV_X4 inst_16714 ( .ZN(net_2365), .A(net_1057) );
OAI21_X2 inst_1785 ( .ZN(net_14651), .B1(net_12490), .B2(net_11810), .A(net_1052) );
NAND2_X2 inst_10104 ( .A1(net_12928), .ZN(net_8497), .A2(net_7283) );
INV_X4 inst_12939 ( .ZN(net_16784), .A(net_16637) );
NOR2_X2 inst_4213 ( .A1(net_9438), .ZN(net_7923), .A2(net_6643) );
NAND2_X2 inst_9341 ( .ZN(net_12211), .A2(net_8914), .A1(net_2267) );
INV_X4 inst_15180 ( .ZN(net_19375), .A(net_3882) );
NAND2_X2 inst_9575 ( .ZN(net_10948), .A1(net_10947), .A2(net_7657) );
AOI22_X2 inst_20045 ( .A1(net_9014), .ZN(net_6378), .B1(net_6377), .B2(net_6376), .A2(net_4928) );
OAI21_X2 inst_2286 ( .A(net_10593), .ZN(net_6539), .B1(net_6538), .B2(net_6537) );
NAND3_X2 inst_6022 ( .A3(net_20822), .A1(net_20821), .ZN(net_20009), .A2(net_12994) );
NAND2_X2 inst_10694 ( .ZN(net_6073), .A2(net_4584), .A1(net_2585) );
NAND2_X2 inst_12118 ( .ZN(net_213), .A1(net_212), .A2(net_211) );
INV_X2 inst_19158 ( .ZN(net_5001), .A(net_3976) );
NAND2_X4 inst_7142 ( .ZN(net_12061), .A2(net_10914), .A1(net_9806) );
NAND2_X4 inst_7512 ( .ZN(net_2637), .A2(net_2137), .A1(net_1278) );
OAI21_X2 inst_2137 ( .ZN(net_9982), .B2(net_8830), .A(net_5974), .B1(net_2744) );
NAND2_X2 inst_9406 ( .ZN(net_20833), .A2(net_12582), .A1(net_11681) );
CLKBUF_X2 inst_21741 ( .A(net_21311), .Z(net_21613) );
NAND2_X4 inst_7107 ( .ZN(net_14448), .A1(net_11108), .A2(net_7298) );
OAI21_X2 inst_1613 ( .A(net_16260), .ZN(net_16110), .B1(net_15657), .B2(net_15410) );
NAND3_X2 inst_6624 ( .A3(net_19056), .ZN(net_9049), .A1(net_6762), .A2(net_2995) );
INV_X4 inst_16503 ( .ZN(net_2193), .A(net_1501) );
NAND3_X2 inst_5659 ( .ZN(net_16846), .A1(net_16319), .A3(net_16288), .A2(net_15965) );
INV_X4 inst_15508 ( .ZN(net_4750), .A(net_4018) );
NAND3_X2 inst_5965 ( .ZN(net_14779), .A3(net_13357), .A2(net_12071), .A1(net_11922) );
INV_X4 inst_15098 ( .A(net_4032), .ZN(net_3230) );
INV_X4 inst_17002 ( .ZN(net_19340), .A(net_867) );
OR2_X2 inst_1141 ( .ZN(net_20137), .A2(net_11478), .A1(net_4957) );
INV_X4 inst_15982 ( .ZN(net_2374), .A(net_1324) );
OAI211_X2 inst_2488 ( .A(net_14226), .ZN(net_13200), .B(net_13199), .C1(net_13198), .C2(net_6142) );
NOR2_X2 inst_3589 ( .ZN(net_20275), .A2(net_12350), .A1(net_10869) );
INV_X2 inst_18379 ( .ZN(net_16894), .A(net_16704) );
SDFF_X2 inst_932 ( .QN(net_21019), .D(net_402), .SE(net_253), .CK(net_21907), .SI(x2688) );
XNOR2_X2 inst_180 ( .A(net_17771), .ZN(net_17769), .B(net_9241) );
INV_X4 inst_12891 ( .A(net_17244), .ZN(net_16807) );
INV_X4 inst_13472 ( .A(net_9646), .ZN(net_9645) );
NAND2_X2 inst_9057 ( .ZN(net_14000), .A1(net_13999), .A2(net_12024) );
INV_X2 inst_18762 ( .A(net_12976), .ZN(net_7626) );
INV_X4 inst_16584 ( .ZN(net_7414), .A(net_2994) );
NAND2_X2 inst_8003 ( .A2(net_18310), .ZN(net_18306), .A1(net_17387) );
INV_X4 inst_15474 ( .ZN(net_13534), .A(net_11562) );
AOI21_X2 inst_20422 ( .ZN(net_19901), .B1(net_15864), .B2(net_14088), .A(net_11543) );
NAND2_X2 inst_8475 ( .A1(net_20767), .ZN(net_17013), .A2(net_16807) );
NAND2_X2 inst_11995 ( .ZN(net_1452), .A1(net_417), .A2(net_56) );
NAND3_X2 inst_6455 ( .ZN(net_20667), .A3(net_11717), .A1(net_9513), .A2(net_3544) );
INV_X4 inst_12635 ( .ZN(net_17918), .A(net_17917) );
INV_X4 inst_12654 ( .ZN(net_17842), .A(net_17841) );
INV_X4 inst_17870 ( .A(net_888), .ZN(net_320) );
CLKBUF_X2 inst_22846 ( .A(net_22717), .Z(net_22718) );
NAND2_X2 inst_10318 ( .ZN(net_9346), .A1(net_7836), .A2(net_4834) );
INV_X4 inst_13527 ( .ZN(net_12802), .A(net_9316) );
INV_X4 inst_15214 ( .ZN(net_4332), .A(net_2888) );
AOI21_X2 inst_20817 ( .ZN(net_10017), .B2(net_6571), .B1(net_6270), .A(net_3796) );
INV_X16 inst_19744 ( .ZN(net_20557), .A(net_20548) );
NOR2_X4 inst_3287 ( .A2(net_20567), .ZN(net_2685), .A1(net_61) );
XNOR2_X2 inst_211 ( .ZN(net_17547), .A(net_17151), .B(net_723) );
NAND3_X2 inst_5892 ( .ZN(net_20639), .A3(net_14039), .A2(net_8719), .A1(net_8586) );
NAND2_X2 inst_11628 ( .ZN(net_3329), .A1(net_2114), .A2(net_1692) );
NOR2_X2 inst_4659 ( .ZN(net_3291), .A2(net_3290), .A1(net_3054) );
NOR2_X4 inst_3120 ( .ZN(net_6919), .A1(net_4027), .A2(net_2431) );
NAND3_X2 inst_5735 ( .ZN(net_16053), .A1(net_15778), .A3(net_13691), .A2(net_12696) );
NAND3_X2 inst_5917 ( .ZN(net_19696), .A1(net_14000), .A3(net_12065), .A2(net_11097) );
INV_X2 inst_18579 ( .ZN(net_10382), .A(net_8892) );
INV_X2 inst_18934 ( .A(net_6030), .ZN(net_5838) );
NAND2_X2 inst_11565 ( .A2(net_2952), .ZN(net_2801), .A1(net_2349) );
CLKBUF_X2 inst_21602 ( .A(net_21473), .Z(net_21474) );
AOI21_X2 inst_20280 ( .ZN(net_19848), .B1(net_16125), .B2(net_16006), .A(net_15460) );
INV_X4 inst_15243 ( .ZN(net_3574), .A(net_2813) );
INV_X4 inst_17004 ( .A(net_4810), .ZN(net_4286) );
NAND2_X4 inst_6945 ( .A2(net_20098), .A1(net_20097), .ZN(net_17618) );
INV_X4 inst_12806 ( .A(net_17214), .ZN(net_17213) );
NOR3_X2 inst_2736 ( .ZN(net_12796), .A2(net_12795), .A3(net_12794), .A1(net_10244) );
NAND2_X4 inst_7178 ( .ZN(net_10883), .A2(net_9356), .A1(net_8115) );
INV_X4 inst_18138 ( .A(net_20988), .ZN(net_2473) );
NAND2_X4 inst_7636 ( .ZN(net_2422), .A1(net_1442), .A2(net_841) );
NOR2_X2 inst_4489 ( .ZN(net_6583), .A2(net_3829), .A1(net_1187) );
INV_X4 inst_17015 ( .ZN(net_19278), .A(net_857) );
NAND3_X4 inst_5523 ( .A3(net_19193), .A1(net_19192), .ZN(net_18183), .A2(net_16034) );
NAND2_X2 inst_10637 ( .A1(net_14226), .ZN(net_6423), .A2(net_3461) );
OAI21_X4 inst_1403 ( .ZN(net_16211), .A(net_16210), .B1(net_15879), .B2(net_15239) );
NAND2_X4 inst_7155 ( .ZN(net_11705), .A1(net_10914), .A2(net_9574) );
INV_X4 inst_14811 ( .ZN(net_6917), .A(net_3962) );
CLKBUF_X2 inst_22090 ( .A(net_21961), .Z(net_21962) );
INV_X4 inst_15100 ( .ZN(net_14460), .A(net_10229) );
INV_X4 inst_14684 ( .ZN(net_18847), .A(net_18025) );
DFF_X1 inst_19882 ( .D(net_17131), .CK(net_21978), .Q(x957) );
INV_X2 inst_18745 ( .ZN(net_7894), .A(net_7893) );
XOR2_X2 inst_42 ( .A(net_21183), .Z(net_579), .B(net_578) );
NAND2_X2 inst_10521 ( .ZN(net_11763), .A1(net_6856), .A2(net_6855) );
INV_X4 inst_13535 ( .A(net_9212), .ZN(net_9211) );
INV_X4 inst_15880 ( .ZN(net_13538), .A(net_6905) );
INV_X4 inst_16009 ( .ZN(net_14009), .A(net_7170) );
INV_X1 inst_19748 ( .A(net_12694), .ZN(net_12410) );
INV_X4 inst_17732 ( .ZN(net_693), .A(net_182) );
NOR2_X2 inst_4084 ( .A1(net_14166), .A2(net_12035), .ZN(net_10718) );
INV_X4 inst_16154 ( .ZN(net_12306), .A(net_8222) );
OAI21_X4 inst_1479 ( .B2(net_19501), .B1(net_19500), .ZN(net_14661), .A(net_12398) );
INV_X4 inst_18346 ( .ZN(net_20778), .A(net_4031) );
INV_X2 inst_19641 ( .A(net_19438), .ZN(net_19433) );
XNOR2_X2 inst_437 ( .ZN(net_16096), .A(net_16095), .B(net_15586) );
NAND2_X2 inst_11606 ( .A1(net_3780), .ZN(net_2626), .A2(net_2037) );
INV_X4 inst_16664 ( .ZN(net_3311), .A(net_61) );
INV_X4 inst_13307 ( .ZN(net_11815), .A(net_10486) );
NAND2_X2 inst_8316 ( .ZN(net_17574), .A2(net_17351), .A1(net_17228) );
INV_X4 inst_14489 ( .ZN(net_13855), .A(net_4848) );
INV_X4 inst_14391 ( .ZN(net_5133), .A(net_5132) );
INV_X4 inst_16034 ( .A(net_2332), .ZN(net_2210) );
CLKBUF_X2 inst_21523 ( .A(net_21272), .Z(net_21395) );
AOI21_X4 inst_20252 ( .B1(net_14334), .ZN(net_7127), .A(net_6078), .B2(net_3144) );
INV_X4 inst_17513 ( .A(net_14308), .ZN(net_410) );
INV_X4 inst_12782 ( .ZN(net_17304), .A(net_17303) );
NAND2_X2 inst_9425 ( .ZN(net_20733), .A1(net_9325), .A2(net_9284) );
NAND2_X2 inst_10451 ( .ZN(net_7045), .A1(net_7044), .A2(net_7043) );
OAI21_X2 inst_1706 ( .A(net_15876), .ZN(net_15255), .B2(net_14129), .B1(net_12599) );
INV_X2 inst_19400 ( .A(net_2642), .ZN(net_2028) );
NAND3_X2 inst_6733 ( .ZN(net_6479), .A2(net_6478), .A1(net_3183), .A3(net_1694) );
NAND3_X2 inst_6778 ( .A2(net_9342), .A3(net_5260), .ZN(net_4506), .A1(net_2733) );
INV_X4 inst_17638 ( .ZN(net_2636), .A(net_310) );
OAI21_X2 inst_2220 ( .B2(net_11090), .B1(net_9768), .ZN(net_8513), .A(net_5355) );
AOI21_X2 inst_20653 ( .ZN(net_13042), .B2(net_9486), .A(net_8563), .B1(net_2902) );
INV_X2 inst_18769 ( .ZN(net_7585), .A(net_7584) );
INV_X4 inst_17075 ( .ZN(net_3852), .A(net_1269) );
NAND2_X2 inst_9958 ( .ZN(net_20022), .A1(net_8917), .A2(net_8916) );
OAI21_X2 inst_2247 ( .A(net_10319), .ZN(net_7327), .B2(net_6919), .B1(net_1149) );
INV_X4 inst_13517 ( .ZN(net_13001), .A(net_9394) );
NAND2_X2 inst_9706 ( .A1(net_14051), .ZN(net_13121), .A2(net_10200) );
NAND2_X2 inst_11852 ( .A1(net_20493), .ZN(net_3217), .A2(net_2710) );
INV_X4 inst_17302 ( .A(net_3309), .ZN(net_607) );
NAND3_X2 inst_5786 ( .A3(net_18892), .A1(net_18891), .ZN(net_15779), .A2(net_13230) );
NOR2_X2 inst_3418 ( .A1(net_15969), .ZN(net_15577), .A2(net_14807) );
INV_X4 inst_17784 ( .A(net_20875), .ZN(net_140) );
NOR2_X4 inst_3334 ( .A2(net_766), .ZN(net_200), .A1(net_199) );
XNOR2_X2 inst_407 ( .A(net_16650), .ZN(net_16647), .B(net_16646) );
NOR2_X2 inst_3558 ( .ZN(net_12982), .A1(net_10738), .A2(net_10321) );
AOI21_X4 inst_20201 ( .B2(net_20393), .ZN(net_19806), .A(net_14612), .B1(net_13814) );
OR2_X2 inst_1208 ( .ZN(net_3316), .A1(net_3315), .A2(net_3314) );
NAND3_X2 inst_5843 ( .ZN(net_20047), .A3(net_14494), .A1(net_11411), .A2(net_10501) );
AOI211_X2 inst_21013 ( .ZN(net_15682), .C1(net_15681), .C2(net_14928), .A(net_11475), .B(net_7907) );
CLKBUF_X2 inst_21642 ( .A(net_21513), .Z(net_21514) );
XNOR2_X2 inst_652 ( .B(net_500), .ZN(net_371), .A(net_370) );
AOI21_X2 inst_20346 ( .ZN(net_15759), .A(net_15345), .B2(net_15054), .B1(net_11427) );
NAND2_X4 inst_7642 ( .ZN(net_1413), .A2(net_1009), .A1(net_515) );
INV_X4 inst_15643 ( .A(net_7044), .ZN(net_2119) );
CLKBUF_X2 inst_22047 ( .A(net_21918), .Z(net_21919) );
NAND2_X2 inst_9935 ( .ZN(net_20757), .A1(net_9148), .A2(net_7103) );
XNOR2_X2 inst_677 ( .B(net_20768), .ZN(net_18872), .A(net_11891) );
XNOR2_X2 inst_130 ( .B(net_21195), .ZN(net_18249), .A(net_18136) );
NAND2_X1 inst_12155 ( .A2(net_10950), .A1(net_9387), .ZN(net_6609) );
OAI21_X2 inst_1566 ( .A(net_16644), .ZN(net_16525), .B2(net_16366), .B1(net_14965) );
AOI21_X2 inst_20530 ( .ZN(net_14525), .B1(net_12546), .B2(net_11706), .A(net_11100) );
INV_X4 inst_12468 ( .ZN(net_18786), .A(net_18785) );
NAND2_X2 inst_7711 ( .ZN(net_18854), .A2(net_18845), .A1(net_18829) );
NAND2_X2 inst_10829 ( .A1(net_7976), .ZN(net_6774), .A2(net_4049) );
INV_X4 inst_14892 ( .A(net_5189), .ZN(net_3650) );
NAND2_X2 inst_10489 ( .ZN(net_6932), .A2(net_5086), .A1(net_70) );
INV_X4 inst_18247 ( .A(net_20959), .ZN(net_211) );
SDFF_X2 inst_1054 ( .QN(net_20977), .D(net_1843), .SE(net_263), .CK(net_22640), .SI(x3346) );
INV_X2 inst_18650 ( .A(net_10208), .ZN(net_9225) );
NAND2_X2 inst_11420 ( .A1(net_20536), .ZN(net_9073), .A2(net_4339) );
SDFF_X2 inst_972 ( .QN(net_21012), .D(net_422), .SE(net_263), .CK(net_22730), .SI(x2835) );
AOI21_X2 inst_20864 ( .ZN(net_8749), .B1(net_5100), .B2(net_4734), .A(net_948) );
INV_X4 inst_15227 ( .ZN(net_4741), .A(net_2857) );
INV_X4 inst_13992 ( .ZN(net_10619), .A(net_6507) );
CLKBUF_X2 inst_22705 ( .A(net_22576), .Z(net_22577) );
OAI21_X2 inst_1843 ( .ZN(net_19240), .B2(net_11610), .B1(net_3285), .A(net_1070) );
INV_X4 inst_16897 ( .ZN(net_4250), .A(net_2985) );
INV_X4 inst_16639 ( .ZN(net_9542), .A(net_154) );
CLKBUF_X2 inst_21887 ( .A(net_21758), .Z(net_21759) );
INV_X16 inst_19738 ( .ZN(net_1730), .A(net_981) );
INV_X2 inst_19631 ( .A(net_21226), .ZN(net_291) );
NAND2_X2 inst_11113 ( .ZN(net_4318), .A2(net_2741), .A1(net_143) );
AOI21_X2 inst_20287 ( .A(net_16743), .ZN(net_16237), .B2(net_15899), .B1(net_8715) );
INV_X2 inst_18853 ( .ZN(net_6517), .A(net_5318) );
NAND2_X2 inst_10224 ( .ZN(net_10368), .A2(net_5117), .A1(net_1670) );
NAND2_X2 inst_11951 ( .ZN(net_1416), .A1(net_1415), .A2(net_954) );
NAND2_X2 inst_11480 ( .ZN(net_7111), .A1(net_2585), .A2(net_2133) );
INV_X4 inst_14679 ( .ZN(net_12532), .A(net_4307) );
INV_X4 inst_15392 ( .ZN(net_10709), .A(net_8667) );
INV_X4 inst_12717 ( .ZN(net_17548), .A(net_17334) );
XNOR2_X2 inst_204 ( .ZN(net_17608), .A(net_17544), .B(net_16267) );
OAI21_X2 inst_1550 ( .ZN(net_17726), .B2(net_17578), .A(net_17461), .B1(net_17460) );
SDFF_X2 inst_910 ( .Q(net_21160), .D(net_16533), .SE(net_263), .CK(net_21528), .SI(x5328) );
INV_X4 inst_14816 ( .ZN(net_8511), .A(net_3935) );
NAND2_X4 inst_7586 ( .ZN(net_3136), .A2(net_1787), .A1(net_782) );
NAND2_X2 inst_10134 ( .ZN(net_8339), .A1(net_8338), .A2(net_5167) );
NAND2_X2 inst_8772 ( .A1(net_15880), .ZN(net_15835), .A2(net_15584) );
INV_X4 inst_13080 ( .ZN(net_19187), .A(net_16049) );
INV_X4 inst_16207 ( .ZN(net_8485), .A(net_5776) );
AOI21_X2 inst_20859 ( .B2(net_10174), .ZN(net_8900), .A(net_6867), .B1(net_4620) );
INV_X4 inst_12494 ( .A(net_18670), .ZN(net_18652) );
NAND2_X4 inst_7562 ( .ZN(net_3025), .A1(net_1687), .A2(net_1533) );
AOI21_X2 inst_20409 ( .B2(net_20177), .B1(net_20176), .ZN(net_15328), .A(net_15113) );
INV_X8 inst_12344 ( .A(net_1192), .ZN(net_387) );
NAND2_X2 inst_11515 ( .ZN(net_2997), .A1(net_2996), .A2(net_1064) );
SDFF_X2 inst_937 ( .QN(net_21070), .D(net_644), .SE(net_263), .CK(net_21741), .SI(x1912) );
NAND2_X4 inst_7401 ( .ZN(net_5908), .A1(net_3766), .A2(net_3115) );
CLKBUF_X2 inst_22362 ( .A(net_22233), .Z(net_22234) );
INV_X4 inst_15315 ( .A(net_3409), .ZN(net_2644) );
AOI222_X2 inst_20060 ( .A1(net_20612), .A2(net_16644), .ZN(net_16288), .B1(net_16287), .B2(net_13823), .C2(net_13480), .C1(net_7284) );
XNOR2_X2 inst_355 ( .ZN(net_16892), .A(net_16887), .B(net_14910) );
NAND2_X2 inst_9259 ( .ZN(net_19127), .A1(net_12640), .A2(net_12614) );
INV_X2 inst_19275 ( .ZN(net_5378), .A(net_2480) );
NAND3_X2 inst_6584 ( .A3(net_19862), .ZN(net_10434), .A1(net_10433), .A2(net_6825) );
NOR2_X2 inst_3498 ( .ZN(net_14079), .A1(net_14078), .A2(net_11932) );
NAND3_X2 inst_6753 ( .A1(net_7822), .ZN(net_5715), .A2(net_5714), .A3(net_5483) );
INV_X4 inst_16139 ( .ZN(net_3703), .A(net_3381) );
NOR2_X2 inst_3693 ( .ZN(net_11268), .A2(net_7813), .A1(net_5581) );
NAND3_X2 inst_6806 ( .A1(net_3276), .ZN(net_3059), .A2(net_2585), .A3(net_2445) );
NAND2_X4 inst_7655 ( .ZN(net_1672), .A1(net_322), .A2(net_108) );
NAND2_X2 inst_11309 ( .ZN(net_4760), .A1(net_4155), .A2(net_3010) );
INV_X4 inst_14619 ( .ZN(net_8101), .A(net_7985) );
INV_X4 inst_15655 ( .ZN(net_4201), .A(net_2101) );
DFF_X1 inst_19868 ( .D(net_17070), .CK(net_22099), .Q(x323) );
INV_X2 inst_18614 ( .ZN(net_11635), .A(net_9615) );
NOR2_X2 inst_3769 ( .ZN(net_11625), .A1(net_10292), .A2(net_10291) );
INV_X4 inst_16466 ( .ZN(net_1523), .A(net_85) );
NOR2_X2 inst_4053 ( .A2(net_13320), .ZN(net_11753), .A1(net_9014) );
OAI21_X2 inst_1747 ( .ZN(net_14943), .B2(net_13527), .A(net_9611), .B1(net_3799) );
NOR2_X2 inst_5109 ( .A2(net_1271), .ZN(net_941), .A1(net_550) );
NAND2_X2 inst_9066 ( .ZN(net_13985), .A1(net_13984), .A2(net_12012) );
NAND2_X2 inst_10477 ( .A1(net_13673), .ZN(net_6979), .A2(net_4262) );
NAND2_X2 inst_11834 ( .ZN(net_11845), .A2(net_1753), .A1(net_168) );
NAND2_X2 inst_11978 ( .ZN(net_1324), .A2(net_931), .A1(net_817) );
CLKBUF_X2 inst_21587 ( .A(net_21458), .Z(net_21459) );
INV_X4 inst_13026 ( .A(net_16465), .ZN(net_16415) );
INV_X4 inst_13352 ( .ZN(net_12673), .A(net_10987) );
NOR2_X2 inst_3917 ( .ZN(net_10295), .A1(net_8803), .A2(net_8219) );
NAND2_X2 inst_9419 ( .A1(net_12528), .ZN(net_11641), .A2(net_11640) );
INV_X4 inst_13243 ( .ZN(net_13299), .A(net_13298) );
NAND2_X4 inst_7601 ( .ZN(net_2153), .A2(net_1456), .A1(net_1442) );
CLKBUF_X2 inst_22025 ( .A(net_21858), .Z(net_21897) );
OAI211_X2 inst_2574 ( .C1(net_9966), .ZN(net_8964), .A(net_8963), .B(net_8962), .C2(net_8446) );
OAI21_X2 inst_2229 ( .A(net_13538), .ZN(net_8266), .B1(net_3877), .B2(net_3593) );
NAND2_X2 inst_11456 ( .ZN(net_5139), .A1(net_3060), .A2(net_2600) );
INV_X4 inst_16613 ( .ZN(net_6797), .A(net_154) );
INV_X4 inst_16966 ( .ZN(net_1308), .A(net_1272) );
NAND3_X2 inst_6252 ( .ZN(net_13009), .A3(net_12944), .A1(net_12566), .A2(net_7628) );
INV_X4 inst_14587 ( .ZN(net_7992), .A(net_4479) );
OR2_X2 inst_1245 ( .ZN(net_10345), .A1(net_824), .A2(net_43) );
DFF_X1 inst_19887 ( .D(net_17122), .CK(net_21819), .Q(x1247) );
INV_X2 inst_19131 ( .ZN(net_4831), .A(net_4224) );
INV_X4 inst_12560 ( .ZN(net_18245), .A(net_18244) );
INV_X4 inst_16941 ( .ZN(net_12363), .A(net_7801) );
NOR2_X2 inst_3788 ( .ZN(net_10086), .A2(net_7766), .A1(net_652) );
NAND4_X2 inst_5409 ( .ZN(net_14615), .A4(net_12511), .A2(net_12043), .A3(net_10998), .A1(net_9686) );
NOR2_X2 inst_3663 ( .A2(net_12835), .ZN(net_11563), .A1(net_11562) );
NAND2_X2 inst_11977 ( .ZN(net_1458), .A1(net_692), .A2(net_70) );
INV_X4 inst_15526 ( .ZN(net_2394), .A(net_2243) );
NOR2_X4 inst_3008 ( .ZN(net_6058), .A1(net_5658), .A2(net_5042) );
CLKBUF_X2 inst_21848 ( .A(net_21719), .Z(net_21720) );
NAND4_X2 inst_5515 ( .A3(net_20784), .ZN(net_10500), .A4(net_10499), .A2(net_6552), .A1(net_6329) );
NAND3_X2 inst_5900 ( .ZN(net_15149), .A3(net_13403), .A2(net_10390), .A1(net_5747) );
NAND2_X2 inst_8234 ( .A1(net_20711), .ZN(net_17755), .A2(net_17754) );
CLKBUF_X2 inst_22827 ( .A(net_22698), .Z(net_22699) );
NAND2_X2 inst_10640 ( .ZN(net_6419), .A2(net_6418), .A1(net_2466) );
AOI211_X2 inst_21047 ( .ZN(net_12860), .B(net_12859), .C1(net_11860), .A(net_9226), .C2(net_3208) );
NOR2_X2 inst_4071 ( .ZN(net_7640), .A1(net_4605), .A2(net_2937) );
NAND2_X2 inst_8738 ( .A1(net_16242), .ZN(net_16024), .A2(net_15720) );
INV_X4 inst_13614 ( .A(net_10613), .ZN(net_10393) );
CLKBUF_X2 inst_21790 ( .A(net_21661), .Z(net_21662) );
NAND2_X2 inst_11363 ( .ZN(net_6100), .A2(net_3607), .A1(net_2163) );
NAND2_X2 inst_8249 ( .ZN(net_17713), .A2(net_17533), .A1(net_811) );
CLKBUF_X2 inst_22061 ( .A(net_21932), .Z(net_21933) );
OAI211_X2 inst_2469 ( .ZN(net_13875), .B(net_13842), .C1(net_12620), .C2(net_7543), .A(net_5138) );
NAND2_X2 inst_7868 ( .ZN(net_18552), .A2(net_18510), .A1(net_18481) );
NAND2_X2 inst_9287 ( .ZN(net_12536), .A2(net_9562), .A1(net_1409) );
CLKBUF_X2 inst_21568 ( .A(net_21439), .Z(net_21440) );
INV_X4 inst_13230 ( .ZN(net_13511), .A(net_12498) );
NOR2_X2 inst_4736 ( .A1(net_20802), .ZN(net_3936), .A2(net_3284) );
INV_X4 inst_16509 ( .ZN(net_13619), .A(net_8293) );
CLKBUF_X2 inst_22428 ( .A(net_21946), .Z(net_22300) );
NAND2_X2 inst_8437 ( .ZN(net_19352), .A2(net_17125), .A1(net_17031) );
INV_X4 inst_14442 ( .ZN(net_4993), .A(net_4992) );
INV_X4 inst_14761 ( .ZN(net_6956), .A(net_4060) );
NAND3_X2 inst_6259 ( .ZN(net_12996), .A3(net_12995), .A2(net_8546), .A1(net_6545) );
AOI211_X2 inst_20999 ( .C1(net_16035), .ZN(net_15966), .C2(net_15568), .B(net_11679), .A(net_11477) );
INV_X4 inst_17417 ( .ZN(net_1607), .A(net_970) );
NAND2_X2 inst_10330 ( .ZN(net_7722), .A1(net_4515), .A2(net_3114) );
NOR2_X2 inst_3715 ( .A2(net_11435), .ZN(net_10979), .A1(net_7688) );
NAND2_X4 inst_6983 ( .ZN(net_17576), .A2(net_16918), .A1(net_16736) );
NAND2_X2 inst_10929 ( .ZN(net_6338), .A1(net_5217), .A2(net_3661) );
CLKBUF_X2 inst_21868 ( .A(net_21287), .Z(net_21740) );
INV_X4 inst_16733 ( .ZN(net_9537), .A(net_5572) );
NOR2_X4 inst_3042 ( .ZN(net_6222), .A2(net_5043), .A1(net_3578) );
INV_X4 inst_17328 ( .A(net_1545), .ZN(net_925) );
CLKBUF_X2 inst_22574 ( .A(net_22445), .Z(net_22446) );
SDFF_X2 inst_981 ( .QN(net_21072), .D(net_563), .SE(net_253), .CK(net_21728), .SI(x1878) );
NAND2_X2 inst_7735 ( .ZN(net_18813), .A2(net_18765), .A1(net_17720) );
NAND2_X2 inst_11940 ( .ZN(net_6480), .A1(net_991), .A2(net_667) );
AOI222_X2 inst_20065 ( .ZN(net_11923), .A2(net_8684), .B1(net_8488), .B2(net_5654), .C1(net_5438), .C2(net_4072), .A1(net_60) );
NAND2_X2 inst_8815 ( .ZN(net_15581), .A2(net_14824), .A1(net_5758) );
AOI21_X2 inst_20832 ( .ZN(net_9734), .A(net_9733), .B1(net_9294), .B2(net_2892) );
INV_X4 inst_17746 ( .ZN(net_3493), .A(net_965) );
CLKBUF_X2 inst_21789 ( .A(net_21634), .Z(net_21661) );
NAND3_X2 inst_6189 ( .ZN(net_13424), .A2(net_12226), .A1(net_10897), .A3(net_10270) );
INV_X8 inst_12260 ( .ZN(net_3882), .A(net_2143) );
NAND2_X2 inst_12064 ( .ZN(net_1211), .A1(net_856), .A2(net_153) );
INV_X4 inst_15056 ( .ZN(net_11866), .A(net_8311) );
CLKBUF_X2 inst_22583 ( .A(net_22454), .Z(net_22455) );
OAI21_X2 inst_2094 ( .ZN(net_10123), .A(net_10122), .B1(net_7422), .B2(net_5569) );
NOR2_X2 inst_3417 ( .ZN(net_15592), .A2(net_14903), .A1(net_14297) );
NAND3_X2 inst_6279 ( .ZN(net_20609), .A2(net_12903), .A3(net_12902), .A1(net_11203) );
AOI21_X2 inst_20950 ( .B2(net_13002), .A(net_11087), .ZN(net_5771), .B1(net_2930) );
NAND3_X2 inst_6794 ( .ZN(net_3460), .A2(net_3459), .A3(net_3458), .A1(net_1321) );
INV_X4 inst_13347 ( .A(net_12851), .ZN(net_11061) );
NAND4_X2 inst_5406 ( .ZN(net_19698), .A2(net_18899), .A1(net_18898), .A4(net_7565), .A3(net_3304) );
INV_X4 inst_14337 ( .ZN(net_10207), .A(net_5383) );
NAND3_X2 inst_6292 ( .ZN(net_20133), .A2(net_12830), .A3(net_12829), .A1(net_11035) );
INV_X4 inst_14947 ( .ZN(net_11786), .A(net_9263) );
INV_X4 inst_13959 ( .ZN(net_6748), .A(net_6747) );
NAND4_X2 inst_5324 ( .ZN(net_15725), .A4(net_14975), .A1(net_14519), .A3(net_14296), .A2(net_13481) );
NOR2_X2 inst_3491 ( .ZN(net_14249), .A1(net_12611), .A2(net_9946) );
OAI211_X2 inst_2393 ( .C2(net_20401), .C1(net_20400), .ZN(net_19209), .B(net_15547), .A(net_15029) );
XNOR2_X2 inst_71 ( .ZN(net_18754), .B(net_18732), .A(net_17635) );
INV_X4 inst_14787 ( .ZN(net_4528), .A(net_4013) );
INV_X2 inst_19455 ( .A(net_9656), .ZN(net_1528) );
NOR2_X2 inst_4079 ( .ZN(net_7382), .A1(net_6267), .A2(net_4646) );
NAND2_X2 inst_10114 ( .ZN(net_8424), .A2(net_5012), .A1(net_4127) );
NOR2_X4 inst_3231 ( .ZN(net_4075), .A1(net_1734), .A2(net_107) );
NAND2_X2 inst_9084 ( .ZN(net_19321), .A1(net_13813), .A2(net_13812) );
CLKBUF_X2 inst_22544 ( .A(net_22415), .Z(net_22416) );
CLKBUF_X2 inst_22045 ( .A(net_21448), .Z(net_21917) );
INV_X4 inst_16902 ( .ZN(net_5836), .A(net_946) );
INV_X4 inst_12884 ( .A(net_17029), .ZN(net_16820) );
INV_X4 inst_14407 ( .ZN(net_7777), .A(net_6927) );
INV_X4 inst_16833 ( .ZN(net_7121), .A(net_986) );
XNOR2_X2 inst_336 ( .B(net_21208), .A(net_17370), .ZN(net_16987) );
NAND2_X1 inst_12129 ( .A2(net_18649), .ZN(net_18637), .A1(net_16866) );
INV_X4 inst_16923 ( .ZN(net_1220), .A(net_221) );
CLKBUF_X2 inst_22775 ( .A(net_22646), .Z(net_22647) );
NAND3_X2 inst_6479 ( .ZN(net_11274), .A2(net_11273), .A3(net_11272), .A1(net_2664) );
INV_X2 inst_19565 ( .A(net_15178), .ZN(net_789) );
OAI21_X2 inst_1939 ( .ZN(net_12862), .B1(net_12861), .B2(net_11189), .A(net_5601) );
NOR2_X1 inst_5157 ( .A1(net_10093), .ZN(net_5349), .A2(net_5348) );
INV_X2 inst_18872 ( .ZN(net_7592), .A(net_6242) );
NOR2_X4 inst_2902 ( .ZN(net_12428), .A2(net_9106), .A1(net_5107) );
INV_X4 inst_14503 ( .A(net_6624), .ZN(net_4834) );
CLKBUF_X2 inst_22850 ( .A(net_22721), .Z(net_22722) );
NAND2_X2 inst_7844 ( .A1(net_21161), .A2(net_18626), .ZN(net_18613) );
INV_X4 inst_17424 ( .A(net_3309), .ZN(net_909) );
NAND2_X2 inst_8726 ( .A1(net_20928), .ZN(net_20116), .A2(net_15768) );
DFF_X1 inst_19825 ( .D(net_17684), .CK(net_21364), .Q(x304) );
AOI211_X2 inst_21001 ( .ZN(net_20261), .C1(net_15889), .B(net_15251), .A(net_14908), .C2(net_14247) );
NAND4_X4 inst_5174 ( .A4(net_18975), .A1(net_18974), .ZN(net_17099), .A3(net_14956), .A2(net_13104) );
NAND2_X2 inst_8508 ( .ZN(net_16923), .A2(net_16922), .A1(net_5274) );
NAND2_X2 inst_9553 ( .ZN(net_12689), .A1(net_11018), .A2(net_11017) );
INV_X4 inst_13450 ( .ZN(net_12872), .A(net_9747) );
NAND2_X2 inst_11736 ( .ZN(net_6391), .A2(net_2477), .A1(net_168) );
NAND2_X2 inst_8263 ( .ZN(net_19120), .A2(net_17775), .A1(net_792) );
NAND3_X2 inst_5870 ( .A2(net_19293), .A1(net_19292), .ZN(net_19141), .A3(net_12831) );
INV_X4 inst_17218 ( .ZN(net_692), .A(net_154) );
NAND3_X2 inst_5998 ( .ZN(net_14435), .A1(net_12760), .A3(net_11219), .A2(net_9544) );
INV_X2 inst_18432 ( .ZN(net_20241), .A(net_14128) );
AOI21_X2 inst_20649 ( .ZN(net_13059), .A(net_13058), .B2(net_9836), .B1(net_6547) );
INV_X4 inst_17352 ( .ZN(net_1343), .A(net_213) );
INV_X2 inst_18593 ( .ZN(net_10129), .A(net_10128) );
NOR2_X2 inst_3752 ( .ZN(net_10410), .A1(net_10409), .A2(net_7317) );
XNOR2_X2 inst_284 ( .B(net_21207), .ZN(net_17161), .A(net_16970) );
INV_X4 inst_13809 ( .ZN(net_12561), .A(net_7541) );
INV_X4 inst_16756 ( .ZN(net_12067), .A(net_8533) );
OAI211_X2 inst_2579 ( .ZN(net_7684), .B(net_7399), .C1(net_4361), .A(net_3960), .C2(net_3317) );
OAI21_X2 inst_1713 ( .ZN(net_15193), .A(net_14720), .B2(net_13918), .B1(net_8728) );
INV_X4 inst_12668 ( .ZN(net_20006), .A(net_17793) );
NAND3_X2 inst_5650 ( .A2(net_20274), .A1(net_20273), .ZN(net_16706), .A3(net_16434) );
NAND2_X4 inst_6970 ( .A2(net_19959), .A1(net_19958), .ZN(net_17408) );
NOR2_X2 inst_4527 ( .A2(net_6404), .ZN(net_5132), .A1(net_111) );
NAND2_X2 inst_9532 ( .ZN(net_11092), .A1(net_11091), .A2(net_11090) );
NOR2_X4 inst_3137 ( .ZN(net_7065), .A2(net_3915), .A1(net_3791) );
INV_X4 inst_16632 ( .ZN(net_1847), .A(net_1109) );
NAND2_X2 inst_11668 ( .ZN(net_2382), .A1(net_1645), .A2(net_1319) );
CLKBUF_X2 inst_21975 ( .A(net_21287), .Z(net_21847) );
INV_X4 inst_18337 ( .A(net_20584), .ZN(net_20583) );
NAND4_X2 inst_5437 ( .ZN(net_13916), .A1(net_10097), .A4(net_8931), .A2(net_8456), .A3(net_6620) );
NAND2_X4 inst_7544 ( .ZN(net_3963), .A2(net_1836), .A1(net_834) );
AOI21_X2 inst_20737 ( .ZN(net_11551), .A(net_11550), .B2(net_7408), .B1(net_3598) );
NOR2_X2 inst_4496 ( .ZN(net_4954), .A2(net_3986), .A1(net_168) );
NAND2_X4 inst_7357 ( .A2(net_19583), .ZN(net_7183), .A1(net_3606) );
NAND3_X2 inst_6344 ( .ZN(net_19322), .A2(net_12248), .A1(net_9362), .A3(net_5730) );
SDFF_X2 inst_951 ( .QN(net_21097), .D(net_727), .SE(net_263), .CK(net_21790), .SI(x1446) );
INV_X4 inst_12565 ( .ZN(net_18278), .A(net_18222) );
NAND2_X2 inst_7727 ( .ZN(net_18829), .A2(net_18802), .A1(net_17566) );
NAND2_X2 inst_9836 ( .ZN(net_11597), .A2(net_9572), .A1(net_7465) );
NAND3_X2 inst_5831 ( .ZN(net_15516), .A1(net_14773), .A3(net_14672), .A2(net_13185) );
INV_X4 inst_15414 ( .ZN(net_15991), .A(net_15666) );
NAND2_X2 inst_10268 ( .ZN(net_9522), .A1(net_7976), .A2(net_6080) );
NAND2_X2 inst_11253 ( .A1(net_20851), .ZN(net_20333), .A2(net_2270) );
NAND2_X2 inst_8938 ( .ZN(net_14840), .A2(net_14096), .A1(net_11665) );
NOR2_X4 inst_3188 ( .ZN(net_5465), .A2(net_3109), .A1(net_3047) );
NAND2_X4 inst_7358 ( .ZN(net_6198), .A2(net_4641), .A1(net_1524) );
NAND2_X4 inst_7351 ( .ZN(net_4812), .A1(net_3446), .A2(net_2621) );
NAND2_X4 inst_7435 ( .ZN(net_4445), .A1(net_3127), .A2(net_2274) );
NAND2_X2 inst_11545 ( .ZN(net_2904), .A1(net_2903), .A2(net_2607) );
NOR2_X4 inst_3129 ( .ZN(net_6878), .A2(net_6221), .A1(net_3883) );
INV_X2 inst_19577 ( .ZN(net_886), .A(net_266) );
NOR2_X2 inst_4674 ( .ZN(net_3731), .A2(net_3241), .A1(net_146) );
INV_X4 inst_12590 ( .ZN(net_18138), .A(net_18086) );
CLKBUF_X2 inst_22192 ( .A(net_22063), .Z(net_22064) );
INV_X4 inst_16048 ( .ZN(net_14634), .A(net_8842) );
AOI21_X2 inst_20699 ( .ZN(net_12139), .A(net_11678), .B2(net_8026), .B1(net_6280) );
NAND3_X4 inst_5581 ( .A1(net_20185), .ZN(net_19373), .A3(net_13659), .A2(net_4173) );
SDFF_X2 inst_921 ( .Q(net_21171), .D(net_16483), .SE(net_263), .CK(net_21376), .SI(x4848) );
INV_X4 inst_14202 ( .ZN(net_5944), .A(net_5943) );
INV_X2 inst_19617 ( .A(net_20914), .ZN(net_41) );
INV_X4 inst_17914 ( .A(net_229), .ZN(net_192) );
NAND2_X4 inst_7618 ( .A1(net_19718), .ZN(net_1332), .A2(net_981) );
NAND2_X2 inst_10772 ( .A1(net_8376), .ZN(net_5628), .A2(net_3972) );
NOR2_X2 inst_3970 ( .ZN(net_8409), .A1(net_8408), .A2(net_4094) );
NAND2_X4 inst_7425 ( .ZN(net_5940), .A2(net_3509), .A1(net_548) );
INV_X4 inst_16633 ( .ZN(net_20755), .A(net_4526) );
NAND2_X2 inst_11499 ( .ZN(net_3074), .A2(net_3073), .A1(net_1982) );
NAND3_X2 inst_6395 ( .ZN(net_11996), .A3(net_11995), .A1(net_9064), .A2(net_7407) );
NAND2_X2 inst_8825 ( .ZN(net_19316), .A1(net_15542), .A2(net_15127) );
INV_X4 inst_16273 ( .A(net_1895), .ZN(net_1814) );
AOI211_X2 inst_21066 ( .B(net_12805), .ZN(net_8992), .C1(net_8991), .A(net_5135), .C2(net_3281) );
SDFF_X2 inst_790 ( .Q(net_20881), .SE(net_18581), .SI(net_18035), .D(net_708), .CK(net_22623) );
INV_X2 inst_18686 ( .A(net_12932), .ZN(net_8669) );
SDFF_X2 inst_1009 ( .QN(net_21004), .SE(net_17277), .D(net_2041), .CK(net_21889), .SI(x2985) );
NAND2_X2 inst_10515 ( .ZN(net_8209), .A2(net_6940), .A1(net_6877) );
NAND2_X2 inst_8931 ( .ZN(net_20147), .A1(net_14858), .A2(net_11523) );
NAND2_X2 inst_8024 ( .ZN(net_18272), .A2(net_18271), .A1(net_17420) );
INV_X4 inst_13217 ( .ZN(net_13636), .A(net_12801) );
INV_X2 inst_19610 ( .A(net_20959), .ZN(net_51) );
SDFF_X2 inst_733 ( .Q(net_20931), .SE(net_18585), .SI(net_18561), .D(net_403), .CK(net_21497) );
NAND3_X2 inst_5885 ( .A3(net_20675), .A1(net_20674), .ZN(net_15241), .A2(net_13529) );
OAI21_X2 inst_1959 ( .ZN(net_12524), .A(net_12523), .B1(net_12522), .B2(net_12475) );
INV_X4 inst_16106 ( .ZN(net_12658), .A(net_7087) );
INV_X4 inst_14294 ( .ZN(net_8965), .A(net_5562) );
INV_X4 inst_16753 ( .ZN(net_1041), .A(net_1040) );
AOI21_X2 inst_20935 ( .B1(net_7071), .ZN(net_6502), .A(net_6451), .B2(net_6445) );
NAND2_X2 inst_8020 ( .ZN(net_18277), .A2(net_18219), .A1(net_17805) );
NAND2_X2 inst_7892 ( .ZN(net_18499), .A2(net_18442), .A1(net_18388) );
INV_X4 inst_18162 ( .A(net_20974), .ZN(net_153) );
NAND3_X2 inst_6416 ( .ZN(net_11947), .A3(net_10221), .A1(net_5774), .A2(net_5041) );
CLKBUF_X2 inst_22144 ( .A(net_22015), .Z(net_22016) );
INV_X4 inst_16690 ( .A(net_10286), .ZN(net_6889) );
NOR2_X2 inst_4471 ( .A1(net_11062), .ZN(net_4425), .A2(net_4424) );
XNOR2_X2 inst_615 ( .B(net_17253), .A(net_17113), .ZN(net_15798) );
INV_X8 inst_12182 ( .ZN(net_17239), .A(net_16911) );
INV_X2 inst_19297 ( .A(net_4066), .ZN(net_2803) );
INV_X4 inst_12597 ( .A(net_18118), .ZN(net_18096) );
NAND2_X2 inst_9157 ( .ZN(net_13385), .A1(net_11440), .A2(net_10605) );
INV_X4 inst_16877 ( .ZN(net_2050), .A(net_282) );
NAND2_X2 inst_8456 ( .A1(net_19459), .ZN(net_17057), .A2(net_16485) );
NAND2_X2 inst_7906 ( .ZN(net_18472), .A2(net_18396), .A1(net_18331) );
CLKBUF_X2 inst_21724 ( .A(net_21595), .Z(net_21596) );
NOR2_X2 inst_3843 ( .ZN(net_9595), .A2(net_9594), .A1(net_8616) );
NAND2_X2 inst_11583 ( .ZN(net_4798), .A1(net_4020), .A2(net_2745) );
NAND2_X2 inst_10621 ( .ZN(net_7830), .A2(net_6573), .A1(net_81) );
INV_X4 inst_17360 ( .A(net_2744), .ZN(net_548) );
INV_X4 inst_13632 ( .A(net_8659), .ZN(net_8238) );
CLKBUF_X2 inst_21918 ( .A(net_21789), .Z(net_21790) );
CLKBUF_X2 inst_22780 ( .A(net_21906), .Z(net_22652) );
NAND3_X4 inst_5593 ( .A3(net_20430), .A1(net_20429), .ZN(net_15016), .A2(net_11609) );
CLKBUF_X2 inst_22951 ( .A(net_22528), .Z(net_22823) );
NAND2_X2 inst_10255 ( .ZN(net_7998), .A1(net_5023), .A2(net_4932) );
CLKBUF_X2 inst_21696 ( .A(net_21541), .Z(net_21568) );
CLKBUF_X2 inst_22465 ( .A(net_22336), .Z(net_22337) );
NOR2_X2 inst_4941 ( .ZN(net_3089), .A1(net_1719), .A2(net_1503) );
INV_X2 inst_18631 ( .ZN(net_9444), .A(net_9443) );
NAND2_X2 inst_7835 ( .ZN(net_19766), .A2(net_18632), .A1(net_16774) );
NOR2_X2 inst_5133 ( .ZN(net_204), .A1(net_203), .A2(net_202) );
NAND2_X4 inst_7095 ( .A1(net_20233), .ZN(net_14487), .A2(net_333) );
AOI22_X2 inst_19984 ( .ZN(net_15209), .A2(net_14111), .B1(net_13940), .B2(net_8551), .A1(net_855) );
NAND2_X2 inst_9986 ( .A1(net_10052), .ZN(net_8849), .A2(net_6504) );
OAI211_X2 inst_2412 ( .ZN(net_15521), .B(net_14654), .A(net_14545), .C1(net_14348), .C2(net_12858) );
NOR2_X2 inst_4928 ( .A1(net_14308), .ZN(net_8717), .A2(net_5432) );
NAND2_X2 inst_10384 ( .A2(net_10523), .ZN(net_7334), .A1(net_7333) );
AOI21_X2 inst_20660 ( .ZN(net_12984), .B1(net_12714), .B2(net_9296), .A(net_5815) );
INV_X2 inst_19357 ( .ZN(net_3302), .A(net_3095) );
OAI21_X2 inst_2214 ( .A(net_15375), .ZN(net_8525), .B2(net_8524), .B1(net_5545) );
AND2_X4 inst_21267 ( .ZN(net_4687), .A2(net_703), .A1(net_152) );
AOI21_X4 inst_20179 ( .ZN(net_19028), .B2(net_14586), .A(net_13269), .B1(net_1244) );
INV_X2 inst_18956 ( .A(net_5713), .ZN(net_5524) );
CLKBUF_X2 inst_22664 ( .A(net_22535), .Z(net_22536) );
NAND2_X2 inst_10018 ( .ZN(net_8773), .A1(net_8772), .A2(net_8771) );
INV_X4 inst_14051 ( .ZN(net_6251), .A(net_6250) );
DFF_X1 inst_19793 ( .D(net_18870), .CK(net_22834), .Q(x1032) );
OAI211_X2 inst_2495 ( .ZN(net_13061), .C2(net_11300), .B(net_8380), .A(net_8056), .C1(net_1864) );
NOR2_X2 inst_4019 ( .A2(net_20077), .ZN(net_8026), .A1(net_8025) );
AND2_X4 inst_21168 ( .A1(net_15413), .ZN(net_13141), .A2(net_13140) );
AOI21_X2 inst_20677 ( .ZN(net_12453), .B1(net_11770), .B2(net_9206), .A(net_2639) );
NAND2_X4 inst_6902 ( .ZN(net_17962), .A1(net_17812), .A2(net_17643) );
NAND2_X2 inst_11265 ( .ZN(net_9626), .A1(net_6613), .A2(net_4192) );
CLKBUF_X2 inst_21706 ( .A(net_21577), .Z(net_21578) );
INV_X4 inst_18147 ( .A(net_21193), .ZN(net_18141) );
NAND2_X2 inst_11697 ( .A2(net_3045), .ZN(net_2316), .A1(net_954) );
NOR2_X4 inst_3236 ( .ZN(net_4304), .A2(net_1700), .A1(net_310) );
NAND2_X2 inst_11219 ( .A1(net_8611), .A2(net_5209), .ZN(net_3968) );
NAND2_X2 inst_10474 ( .A2(net_8469), .ZN(net_6984), .A1(net_6983) );
NAND2_X2 inst_11096 ( .ZN(net_7282), .A1(net_4301), .A2(net_3324) );
INV_X4 inst_15759 ( .A(net_2436), .ZN(net_1928) );
NOR2_X2 inst_3408 ( .ZN(net_19913), .A2(net_15378), .A1(net_15148) );
CLKBUF_X2 inst_22036 ( .A(net_21755), .Z(net_21908) );
XNOR2_X2 inst_88 ( .ZN(net_18565), .A(net_18499), .B(net_17766) );
DFF_X1 inst_19815 ( .D(net_17835), .CK(net_21371), .Q(x222) );
INV_X4 inst_17369 ( .ZN(net_3342), .A(net_640) );
NAND3_X2 inst_6054 ( .ZN(net_14231), .A2(net_14216), .A1(net_12343), .A3(net_8771) );
NAND2_X2 inst_10397 ( .ZN(net_7287), .A2(net_5286), .A1(net_4071) );
NAND2_X2 inst_10356 ( .ZN(net_10998), .A2(net_7443), .A1(net_4915) );
NAND2_X2 inst_11190 ( .ZN(net_6683), .A1(net_4093), .A2(net_4092) );
XNOR2_X2 inst_360 ( .ZN(net_16886), .A(net_16885), .B(net_14916) );
INV_X4 inst_14646 ( .ZN(net_18582), .A(net_18025) );
NAND3_X2 inst_6604 ( .ZN(net_9876), .A3(net_9875), .A2(net_5996), .A1(net_3046) );
NAND2_X2 inst_10876 ( .A1(net_11311), .ZN(net_5424), .A2(net_5423) );
INV_X2 inst_18786 ( .ZN(net_20642), .A(net_9696) );
NOR2_X2 inst_3908 ( .A1(net_12067), .A2(net_10597), .ZN(net_8861) );
INV_X4 inst_12574 ( .ZN(net_18265), .A(net_18226) );
NAND3_X2 inst_6797 ( .A3(net_9903), .A2(net_4931), .ZN(net_3450), .A1(net_3449) );
OR2_X4 inst_1129 ( .ZN(net_4802), .A2(net_703), .A1(net_152) );
NAND2_X2 inst_8922 ( .ZN(net_14954), .A2(net_13737), .A1(net_8717) );
SDFF_X2 inst_744 ( .Q(net_20879), .SE(net_18585), .SI(net_18549), .D(net_8993), .CK(net_22697) );
INV_X4 inst_13116 ( .ZN(net_19876), .A(net_15305) );
INV_X4 inst_17104 ( .ZN(net_2129), .A(net_1101) );
INV_X4 inst_13375 ( .ZN(net_10879), .A(net_10878) );
NOR2_X2 inst_3827 ( .ZN(net_9749), .A1(net_9748), .A2(net_7572) );
INV_X2 inst_18720 ( .A(net_8721), .ZN(net_8130) );
INV_X8 inst_12385 ( .ZN(net_336), .A(net_202) );
INV_X4 inst_17362 ( .ZN(net_4090), .A(net_3780) );
NOR2_X2 inst_4112 ( .ZN(net_7067), .A2(net_6662), .A1(net_4159) );
INV_X4 inst_13492 ( .A(net_11834), .ZN(net_9483) );
INV_X4 inst_16357 ( .ZN(net_12203), .A(net_1292) );
AOI21_X2 inst_20903 ( .ZN(net_7697), .B2(net_4626), .B1(net_2004), .A(net_1140) );
AOI21_X2 inst_20620 ( .ZN(net_20362), .A(net_14743), .B2(net_9153), .B1(net_7457) );
INV_X4 inst_17898 ( .ZN(net_14029), .A(net_78) );
NAND2_X2 inst_11002 ( .ZN(net_4888), .A2(net_3629), .A1(net_874) );
INV_X4 inst_15487 ( .ZN(net_2587), .A(net_2436) );
XNOR2_X2 inst_536 ( .ZN(net_1517), .B(net_1516), .A(net_553) );
INV_X4 inst_12711 ( .ZN(net_17827), .A(net_17459) );
CLKBUF_X2 inst_21829 ( .A(net_21700), .Z(net_21701) );
AOI21_X2 inst_20557 ( .A(net_15289), .ZN(net_14273), .B2(net_12430), .B1(net_5340) );
INV_X4 inst_16243 ( .A(net_2735), .ZN(net_1840) );
NAND2_X2 inst_11032 ( .ZN(net_7264), .A2(net_4419), .A1(net_1072) );
OAI21_X2 inst_2027 ( .ZN(net_11316), .B1(net_11315), .A(net_9894), .B2(net_9640) );
NAND2_X2 inst_8146 ( .ZN(net_18019), .A2(net_17984), .A1(net_17725) );
NAND3_X2 inst_5882 ( .ZN(net_15257), .A2(net_14187), .A3(net_14176), .A1(net_12628) );
NAND2_X4 inst_7487 ( .ZN(net_3898), .A2(net_2445), .A1(net_66) );
XNOR2_X2 inst_416 ( .B(net_21191), .ZN(net_17448), .A(net_16571) );
INV_X4 inst_15773 ( .A(net_16051), .ZN(net_1919) );
NAND2_X2 inst_9169 ( .A1(net_13517), .ZN(net_13357), .A2(net_10533) );
NAND2_X2 inst_10871 ( .A2(net_5525), .ZN(net_5430), .A1(net_809) );
OAI21_X4 inst_1406 ( .A(net_20856), .B2(net_18883), .B1(net_18882), .ZN(net_16183) );
NAND2_X2 inst_8396 ( .ZN(net_17400), .A2(net_16976), .A1(net_16818) );
NAND4_X2 inst_5500 ( .ZN(net_11838), .A1(net_11837), .A4(net_11836), .A3(net_10355), .A2(net_5000) );
NAND4_X2 inst_5330 ( .A4(net_19040), .A1(net_19039), .ZN(net_15571), .A2(net_10700), .A3(net_9918) );
NOR2_X2 inst_4319 ( .A1(net_7357), .A2(net_5914), .ZN(net_5871) );
NAND2_X2 inst_9520 ( .ZN(net_11141), .A2(net_10838), .A1(net_3973) );
NAND2_X2 inst_10943 ( .ZN(net_5154), .A1(net_5153), .A2(net_4398) );
INV_X2 inst_19395 ( .ZN(net_4664), .A(net_3194) );
INV_X2 inst_18392 ( .ZN(net_17082), .A(net_16732) );
NAND2_X2 inst_8046 ( .ZN(net_18230), .A2(net_18226), .A1(net_17186) );
INV_X4 inst_18257 ( .A(net_20958), .ZN(net_212) );
NOR2_X2 inst_4432 ( .A2(net_7096), .ZN(net_4891), .A1(net_4890) );
NAND2_X2 inst_11039 ( .ZN(net_9969), .A1(net_6358), .A2(net_4368) );
INV_X4 inst_13014 ( .ZN(net_16724), .A(net_16569) );
SDFF_X2 inst_973 ( .QN(net_21081), .D(net_739), .SE(net_263), .CK(net_22594), .SI(x1701) );
NOR2_X4 inst_3058 ( .ZN(net_8109), .A2(net_4963), .A1(net_4962) );
INV_X4 inst_13374 ( .ZN(net_20253), .A(net_10883) );
NAND2_X2 inst_11258 ( .ZN(net_4923), .A1(net_3990), .A2(net_3380) );
NAND2_X2 inst_11884 ( .ZN(net_1610), .A2(net_1282), .A1(net_268) );
NAND2_X2 inst_11771 ( .ZN(net_2062), .A2(net_1105), .A1(net_994) );
NOR2_X4 inst_3089 ( .ZN(net_5700), .A1(net_4295), .A2(net_4288) );
INV_X4 inst_18309 ( .A(net_20501), .ZN(net_20500) );
OR2_X4 inst_1122 ( .ZN(net_4805), .A2(net_193), .A1(net_41) );
INV_X4 inst_15009 ( .ZN(net_15582), .A(net_14465) );
INV_X8 inst_12170 ( .ZN(net_20320), .A(net_18377) );
NOR2_X4 inst_3324 ( .A1(net_2001), .ZN(net_1107), .A2(net_826) );
DFF_X1 inst_19848 ( .D(net_17217), .CK(net_22107), .Q(x445) );
NAND2_X4 inst_7478 ( .ZN(net_5006), .A1(net_3331), .A2(net_225) );
NAND2_X2 inst_7987 ( .ZN(net_18329), .A2(net_18328), .A1(net_17223) );
CLKBUF_X2 inst_21757 ( .A(net_21628), .Z(net_21629) );
AOI22_X2 inst_20033 ( .ZN(net_8489), .B1(net_8488), .B2(net_6053), .A2(net_3718), .A1(net_60) );
INV_X4 inst_14351 ( .ZN(net_6121), .A(net_3952) );
NOR2_X4 inst_2981 ( .ZN(net_9746), .A2(net_6172), .A1(net_703) );
INV_X4 inst_15677 ( .ZN(net_2655), .A(net_2049) );
NOR2_X2 inst_4998 ( .A2(net_3276), .ZN(net_1366), .A1(net_718) );
INV_X4 inst_15403 ( .ZN(net_11050), .A(net_10898) );
NAND4_X2 inst_5390 ( .ZN(net_14923), .A1(net_12688), .A2(net_8701), .A4(net_8274), .A3(net_6820) );
NAND2_X2 inst_9240 ( .ZN(net_12692), .A2(net_12402), .A1(net_6513) );
CLKBUF_X2 inst_22213 ( .A(net_21438), .Z(net_22085) );
NOR2_X2 inst_4406 ( .A1(net_5435), .ZN(net_5096), .A2(net_5013) );
AOI21_X2 inst_20267 ( .B2(net_20880), .ZN(net_18062), .B1(net_16141), .A(net_13050) );
NAND3_X2 inst_6169 ( .A2(net_20763), .ZN(net_13615), .A3(net_12830), .A1(net_12392) );
NAND3_X2 inst_6696 ( .ZN(net_7673), .A3(net_7672), .A2(net_6098), .A1(net_3349) );
INV_X2 inst_19125 ( .ZN(net_7313), .A(net_5478) );
INV_X16 inst_19735 ( .ZN(net_868), .A(net_504) );
XNOR2_X2 inst_90 ( .ZN(net_18559), .A(net_18476), .B(net_17650) );
AOI21_X2 inst_20498 ( .A(net_15174), .ZN(net_14674), .B2(net_11917), .B1(net_9311) );
NAND2_X2 inst_11166 ( .ZN(net_20045), .A1(net_8330), .A2(net_4174) );
INV_X4 inst_14950 ( .A(net_4735), .ZN(net_3511) );
INV_X4 inst_16348 ( .A(net_13514), .ZN(net_7170) );
INV_X4 inst_17875 ( .A(net_2744), .ZN(net_758) );
NAND2_X4 inst_6858 ( .ZN(net_18418), .A1(net_18405), .A2(net_18344) );
NAND2_X2 inst_10850 ( .A1(net_6201), .ZN(net_5466), .A2(net_5465) );
INV_X2 inst_18910 ( .ZN(net_9665), .A(net_8085) );
NOR2_X2 inst_4650 ( .A1(net_19439), .ZN(net_4531), .A2(net_3391) );
NAND2_X2 inst_8860 ( .ZN(net_15346), .A1(net_15345), .A2(net_14426) );
NAND2_X4 inst_7197 ( .ZN(net_10372), .A2(net_9148), .A1(net_8284) );
NOR2_X2 inst_5093 ( .ZN(net_10061), .A1(net_522), .A2(net_78) );
NAND2_X4 inst_7625 ( .A2(net_2071), .ZN(net_1727), .A1(net_751) );
NOR2_X2 inst_3833 ( .ZN(net_9715), .A2(net_9714), .A1(net_6905) );
CLKBUF_X2 inst_22874 ( .A(net_21551), .Z(net_22746) );
OAI211_X2 inst_2460 ( .ZN(net_14155), .C2(net_9210), .A(net_6057), .B(net_3840), .C1(net_3364) );
NAND2_X2 inst_8457 ( .A2(net_19459), .ZN(net_17056), .A1(net_16526) );
INV_X2 inst_18893 ( .A(net_7958), .ZN(net_6104) );
OR2_X2 inst_1217 ( .ZN(net_2760), .A2(net_2759), .A1(net_2218) );
INV_X4 inst_15936 ( .A(net_1911), .ZN(net_1724) );
NAND2_X2 inst_10832 ( .ZN(net_7239), .A2(net_5485), .A1(net_703) );
CLKBUF_X2 inst_21928 ( .A(net_21799), .Z(net_21800) );
INV_X2 inst_18706 ( .ZN(net_8248), .A(net_8247) );
NAND2_X2 inst_10788 ( .ZN(net_5586), .A1(net_5585), .A2(net_5584) );
INV_X4 inst_16372 ( .A(net_7298), .ZN(net_6886) );
NAND2_X2 inst_10285 ( .A1(net_10515), .ZN(net_10243), .A2(net_5030) );
NAND2_X4 inst_6938 ( .A2(net_19159), .A1(net_19158), .ZN(net_18252) );
NAND2_X4 inst_7126 ( .A1(net_19211), .ZN(net_12319), .A2(net_10898) );
NAND2_X2 inst_10187 ( .A1(net_9909), .ZN(net_8172), .A2(net_8171) );
INV_X4 inst_15545 ( .A(net_9510), .ZN(net_2363) );
INV_X2 inst_19698 ( .A(net_20554), .ZN(net_20553) );
NOR2_X4 inst_3027 ( .A2(net_6604), .ZN(net_6367), .A1(net_5232) );
NAND3_X2 inst_5907 ( .ZN(net_19792), .A3(net_12922), .A1(net_8869), .A2(net_8619) );
INV_X4 inst_17762 ( .ZN(net_1299), .A(net_295) );
NAND2_X2 inst_8614 ( .ZN(net_20620), .A2(net_16614), .A1(net_500) );
INV_X4 inst_14016 ( .ZN(net_11927), .A(net_6302) );
INV_X4 inst_14059 ( .A(net_8050), .ZN(net_7606) );
AND2_X4 inst_21201 ( .ZN(net_19689), .A1(net_8394), .A2(net_8393) );
INV_X4 inst_18283 ( .ZN(net_20077), .A(net_3427) );
NAND2_X2 inst_10235 ( .ZN(net_8043), .A2(net_6125), .A1(net_5517) );
INV_X4 inst_15843 ( .ZN(net_1841), .A(net_1840) );
NAND2_X4 inst_7480 ( .ZN(net_2879), .A1(net_2285), .A2(net_1785) );
XNOR2_X2 inst_68 ( .ZN(net_18796), .A(net_18740), .B(net_17488) );
NAND2_X2 inst_8029 ( .ZN(net_18266), .A2(net_18265), .A1(net_17430) );
INV_X2 inst_18725 ( .ZN(net_20380), .A(net_12838) );
INV_X4 inst_18289 ( .A(net_20214), .ZN(net_20213) );
OAI22_X2 inst_1253 ( .B2(net_18211), .A1(net_18182), .ZN(net_17877), .A2(net_17876), .B1(net_17875) );
NAND2_X2 inst_10913 ( .ZN(net_5352), .A2(net_5351), .A1(net_4329) );
NAND2_X2 inst_10689 ( .ZN(net_11247), .A1(net_6091), .A2(net_6044) );
NAND2_X2 inst_11943 ( .A2(net_20581), .ZN(net_1443), .A1(net_110) );
NOR3_X2 inst_2793 ( .A2(net_14033), .A3(net_9681), .A1(net_8394), .ZN(net_4235) );
INV_X4 inst_15647 ( .A(net_4655), .ZN(net_3264) );
OAI21_X2 inst_2018 ( .ZN(net_11346), .A(net_11345), .B1(net_9748), .B2(net_6279) );
OAI21_X2 inst_1884 ( .A(net_15119), .ZN(net_13524), .B1(net_9811), .B2(net_9042) );
NAND3_X2 inst_6488 ( .ZN(net_11173), .A2(net_11172), .A3(net_8918), .A1(net_3048) );
CLKBUF_X2 inst_22600 ( .A(net_22471), .Z(net_22472) );
AND2_X2 inst_21346 ( .A2(net_2685), .ZN(net_2666), .A1(net_1184) );
INV_X4 inst_13172 ( .A(net_21109), .ZN(net_16445) );
NAND2_X2 inst_8540 ( .A1(net_21153), .A2(net_17126), .ZN(net_16826) );
INV_X2 inst_19387 ( .ZN(net_2103), .A(net_2102) );
OAI21_X2 inst_1690 ( .ZN(net_15378), .B1(net_14949), .B2(net_13892), .A(net_10689) );
NAND3_X2 inst_6413 ( .ZN(net_11953), .A2(net_9380), .A1(net_8434), .A3(net_5084) );
NAND2_X2 inst_9815 ( .ZN(net_9662), .A1(net_9661), .A2(net_9660) );
NAND4_X2 inst_5312 ( .ZN(net_19383), .A4(net_15089), .A3(net_15018), .A1(net_14645), .A2(net_13797) );
NAND2_X2 inst_9540 ( .ZN(net_11063), .A1(net_11062), .A2(net_11006) );
INV_X4 inst_13015 ( .ZN(net_16431), .A(net_16399) );
OAI22_X2 inst_1287 ( .A1(net_19460), .B1(net_13512), .ZN(net_12889), .A2(net_12888), .B2(net_12887) );
NOR2_X2 inst_4231 ( .ZN(net_8735), .A2(net_8448), .A1(net_948) );
INV_X4 inst_16840 ( .A(net_13058), .ZN(net_977) );
AOI21_X2 inst_20782 ( .B1(net_14038), .ZN(net_10558), .A(net_10557), .B2(net_6417) );
INV_X4 inst_17333 ( .ZN(net_4111), .A(net_1682) );
OR2_X2 inst_1169 ( .A2(net_10593), .ZN(net_6929), .A1(net_81) );
NOR2_X2 inst_4266 ( .ZN(net_9774), .A2(net_6177), .A1(net_6176) );
NAND3_X2 inst_5826 ( .ZN(net_19708), .A1(net_14814), .A2(net_13220), .A3(net_12118) );
DFF_X1 inst_19784 ( .D(net_18708), .CK(net_21631), .Q(x556) );
NOR2_X2 inst_3483 ( .A1(net_14678), .ZN(net_14307), .A2(net_13521) );
INV_X4 inst_17921 ( .A(net_20937), .ZN(net_67) );
NAND3_X2 inst_5704 ( .ZN(net_16205), .A3(net_15863), .A2(net_15101), .A1(net_14598) );
NAND2_X2 inst_8634 ( .A1(net_19445), .A2(net_16602), .ZN(net_16586) );
NAND2_X2 inst_9440 ( .ZN(net_19995), .A2(net_11555), .A1(net_11090) );
AOI21_X2 inst_20661 ( .B1(net_13565), .ZN(net_12966), .A(net_12965), .B2(net_6953) );
CLKBUF_X2 inst_22172 ( .A(net_22043), .Z(net_22044) );
INV_X4 inst_17522 ( .ZN(net_6318), .A(net_112) );
INV_X8 inst_12251 ( .ZN(net_4826), .A(net_2441) );
INV_X4 inst_17788 ( .ZN(net_14557), .A(net_171) );
NOR2_X4 inst_2877 ( .A1(net_13265), .ZN(net_11610), .A2(net_10119) );
AOI211_X2 inst_21039 ( .ZN(net_13874), .C1(net_13873), .B(net_13105), .C2(net_13005), .A(net_9549) );
DFF_X1 inst_19891 ( .D(net_16873), .CK(net_21321), .Q(x215) );
AND3_X2 inst_21137 ( .ZN(net_19415), .A2(net_13170), .A3(net_13169), .A1(net_6711) );
INV_X4 inst_12908 ( .ZN(net_17187), .A(net_16698) );
INV_X4 inst_15150 ( .ZN(net_4902), .A(net_3566) );
INV_X4 inst_16331 ( .ZN(net_1554), .A(net_1303) );
NAND3_X2 inst_6514 ( .ZN(net_10656), .A1(net_10655), .A2(net_10654), .A3(net_10499) );
NAND2_X2 inst_11221 ( .A2(net_9748), .ZN(net_5178), .A1(net_732) );
INV_X4 inst_16561 ( .ZN(net_2627), .A(net_2431) );
NAND2_X4 inst_7502 ( .A1(net_2402), .ZN(net_2284), .A2(net_1662) );
CLKBUF_X2 inst_22491 ( .A(net_22362), .Z(net_22363) );
NAND2_X2 inst_11709 ( .ZN(net_8446), .A2(net_1490), .A1(net_222) );
NAND2_X2 inst_12062 ( .A2(net_1165), .ZN(net_1084), .A1(net_166) );
INV_X2 inst_18983 ( .A(net_9913), .ZN(net_5130) );
OAI21_X4 inst_1418 ( .B2(net_19311), .B1(net_19310), .A(net_16187), .ZN(net_16142) );
NAND2_X2 inst_9095 ( .ZN(net_13784), .A2(net_12470), .A1(net_761) );
INV_X4 inst_14124 ( .ZN(net_6124), .A(net_6123) );
OAI21_X2 inst_1740 ( .ZN(net_15034), .A(net_14764), .B2(net_12789), .B1(net_6412) );
NAND2_X2 inst_10171 ( .ZN(net_8223), .A1(net_8222), .A2(net_8221) );
INV_X4 inst_14499 ( .ZN(net_13479), .A(net_6597) );
NAND3_X2 inst_5663 ( .ZN(net_19208), .A3(net_16262), .A2(net_15882), .A1(net_9248) );
INV_X2 inst_19638 ( .A(net_19428), .ZN(net_19427) );
INV_X4 inst_16433 ( .ZN(net_4872), .A(net_2744) );
INV_X4 inst_16126 ( .ZN(net_4038), .A(net_1322) );
NAND2_X2 inst_7822 ( .ZN(net_19163), .A1(net_18648), .A2(net_17763) );
NAND2_X2 inst_11176 ( .ZN(net_7050), .A1(net_4155), .A2(net_2228) );
OAI21_X2 inst_2001 ( .ZN(net_11650), .A(net_11482), .B2(net_7632), .B1(net_2496) );
NOR2_X2 inst_4836 ( .A1(net_4945), .ZN(net_2565), .A2(net_1710) );
INV_X2 inst_18602 ( .ZN(net_20245), .A(net_10314) );
OAI21_X2 inst_1657 ( .ZN(net_15789), .B2(net_14785), .A(net_14643), .B1(net_14079) );
NAND2_X2 inst_10321 ( .ZN(net_9335), .A1(net_7487), .A2(net_6006) );
INV_X4 inst_12982 ( .A(net_17763), .ZN(net_17372) );
INV_X4 inst_14385 ( .ZN(net_5161), .A(net_5160) );
DFF_X2 inst_19778 ( .Q(net_21106), .D(net_6688), .CK(net_22191) );
INV_X4 inst_15570 ( .ZN(net_4184), .A(net_1421) );
AOI21_X2 inst_20587 ( .ZN(net_14015), .A(net_14014), .B2(net_10384), .B1(net_10078) );
OAI21_X2 inst_2077 ( .ZN(net_10572), .A(net_9940), .B1(net_9573), .B2(net_7891) );
NAND2_X2 inst_10085 ( .A1(net_11466), .ZN(net_8630), .A2(net_8060) );
INV_X4 inst_17057 ( .ZN(net_9396), .A(net_5472) );
INV_X4 inst_14473 ( .ZN(net_8168), .A(net_4896) );
NAND2_X2 inst_8078 ( .A1(net_20442), .ZN(net_19137), .A2(net_18153) );
INV_X4 inst_12729 ( .ZN(net_17771), .A(net_17340) );
AOI21_X2 inst_20571 ( .ZN(net_14142), .B1(net_14141), .B2(net_10656), .A(net_8814) );
INV_X4 inst_13704 ( .ZN(net_12246), .A(net_7876) );
AOI211_X2 inst_21006 ( .ZN(net_15848), .C2(net_15317), .B(net_14503), .A(net_6534), .C1(net_3164) );
INV_X4 inst_13930 ( .A(net_8191), .ZN(net_7623) );
NAND3_X2 inst_6656 ( .ZN(net_8493), .A3(net_8492), .A2(net_8395), .A1(net_5332) );
INV_X8 inst_12179 ( .ZN(net_16969), .A(net_16810) );
OAI21_X4 inst_1495 ( .B1(net_19617), .ZN(net_14327), .A(net_12100), .B2(net_7161) );
SDFF_X2 inst_797 ( .Q(net_20882), .SE(net_18858), .SI(net_17987), .D(net_677), .CK(net_21797) );
NOR2_X2 inst_5051 ( .ZN(net_2412), .A2(net_1397), .A1(net_222) );
NAND3_X4 inst_5546 ( .A3(net_20369), .A1(net_20368), .A2(net_20250), .ZN(net_16808) );
CLKBUF_X2 inst_22789 ( .A(net_22660), .Z(net_22661) );
NAND2_X2 inst_9310 ( .ZN(net_12362), .A2(net_12361), .A1(net_4460) );
INV_X4 inst_17318 ( .ZN(net_6358), .A(net_703) );
NOR2_X4 inst_3032 ( .A1(net_18976), .ZN(net_8397), .A2(net_7941) );
AOI21_X2 inst_20339 ( .ZN(net_20303), .B1(net_20011), .B2(net_15790), .A(net_9009) );
NAND2_X2 inst_8882 ( .ZN(net_15177), .A2(net_14681), .A1(net_13021) );
CLKBUF_X2 inst_21841 ( .A(net_21620), .Z(net_21713) );
INV_X4 inst_17489 ( .ZN(net_428), .A(net_146) );
NAND2_X2 inst_12069 ( .ZN(net_822), .A1(net_808), .A2(net_129) );
CLKBUF_X2 inst_22371 ( .A(net_22242), .Z(net_22243) );
NAND2_X4 inst_6856 ( .ZN(net_18445), .A2(net_18324), .A1(net_18275) );
NAND3_X2 inst_6787 ( .ZN(net_4223), .A2(net_4222), .A1(net_1929), .A3(net_1520) );
INV_X4 inst_13195 ( .ZN(net_14081), .A(net_13410) );
INV_X4 inst_14699 ( .ZN(net_8504), .A(net_4265) );
NOR2_X2 inst_3583 ( .A1(net_14350), .ZN(net_12672), .A2(net_10991) );
INV_X2 inst_19665 ( .A(net_20476), .ZN(net_20475) );
INV_X4 inst_13242 ( .ZN(net_14274), .A(net_13364) );
NAND2_X2 inst_8446 ( .ZN(net_18478), .A2(net_16779), .A1(net_16626) );
INV_X2 inst_19399 ( .ZN(net_19647), .A(net_2033) );
OR2_X4 inst_1115 ( .ZN(net_5565), .A1(net_824), .A2(net_809) );
NOR2_X2 inst_4933 ( .A1(net_2942), .ZN(net_1760), .A2(net_1144) );
AOI21_X2 inst_20703 ( .A(net_20889), .ZN(net_12128), .B1(net_7785), .B2(net_7034) );
INV_X4 inst_17793 ( .ZN(net_3107), .A(net_896) );
NAND3_X2 inst_6234 ( .ZN(net_13215), .A3(net_13167), .A2(net_12409), .A1(net_8309) );
SDFF_X2 inst_1021 ( .QN(net_21061), .D(net_483), .SE(net_263), .CK(net_21712), .SI(x2035) );
NOR2_X4 inst_2976 ( .ZN(net_9536), .A2(net_3588), .A1(net_1848) );
INV_X4 inst_17662 ( .ZN(net_19372), .A(net_255) );
NAND2_X2 inst_9140 ( .ZN(net_19098), .A1(net_14086), .A2(net_10786) );
NOR2_X2 inst_4204 ( .ZN(net_15950), .A2(net_6794), .A1(net_6682) );
INV_X4 inst_18116 ( .A(net_20975), .ZN(net_265) );
NAND2_X2 inst_12095 ( .A2(net_2274), .ZN(net_567), .A1(net_97) );
NOR2_X2 inst_4827 ( .ZN(net_2825), .A2(net_1749), .A1(net_874) );
AOI21_X2 inst_20459 ( .A(net_15312), .ZN(net_15035), .B2(net_12796), .B1(net_6416) );
XNOR2_X2 inst_572 ( .B(net_16879), .ZN(net_627), .A(net_626) );
INV_X4 inst_12699 ( .ZN(net_17628), .A(net_17627) );
INV_X8 inst_12392 ( .A(net_318), .ZN(net_255) );
XNOR2_X2 inst_257 ( .A(net_19436), .ZN(net_17285), .B(net_16546) );
NOR2_X2 inst_5036 ( .A1(net_1697), .ZN(net_1120), .A2(net_919) );
INV_X4 inst_15062 ( .ZN(net_3634), .A(net_3299) );
INV_X4 inst_17449 ( .ZN(net_1261), .A(net_332) );
XNOR2_X2 inst_485 ( .B(net_21183), .ZN(net_10497), .A(net_10496) );
INV_X4 inst_12971 ( .ZN(net_16887), .A(net_16515) );
AOI21_X2 inst_20775 ( .B2(net_19757), .B1(net_19756), .ZN(net_10616), .A(net_5393) );
NAND2_X2 inst_10684 ( .ZN(net_11820), .A2(net_3722), .A1(net_2694) );
INV_X4 inst_14655 ( .ZN(net_18858), .A(net_18025) );
OR2_X2 inst_1205 ( .A2(net_19440), .ZN(net_3534), .A1(net_2221) );
INV_X2 inst_19659 ( .A(net_20437), .ZN(net_20436) );
INV_X4 inst_17609 ( .ZN(net_2712), .A(net_310) );
INV_X4 inst_18043 ( .A(net_20980), .ZN(net_1860) );
NOR2_X2 inst_5085 ( .A2(net_20923), .ZN(net_1359), .A1(net_146) );
INV_X4 inst_16286 ( .ZN(net_6601), .A(net_732) );
NAND2_X2 inst_11048 ( .A1(net_11614), .A2(net_4736), .ZN(net_4714) );
CLKBUF_X2 inst_22317 ( .A(net_22188), .Z(net_22189) );
INV_X2 inst_18558 ( .ZN(net_10870), .A(net_10869) );
AOI21_X2 inst_20325 ( .ZN(net_20344), .B1(net_20289), .A(net_13834), .B2(net_8734) );
INV_X4 inst_17064 ( .ZN(net_8644), .A(net_6648) );
NAND2_X2 inst_8310 ( .A2(net_17662), .ZN(net_17585), .A1(net_17402) );
INV_X4 inst_15012 ( .ZN(net_13569), .A(net_10141) );
NAND2_X2 inst_8641 ( .A1(net_16799), .ZN(net_16575), .A2(net_16574) );
INV_X2 inst_19593 ( .A(net_889), .ZN(net_259) );
INV_X4 inst_14409 ( .ZN(net_6161), .A(net_4043) );
NAND2_X4 inst_6929 ( .A2(net_19097), .A1(net_19096), .ZN(net_17730) );
NOR2_X2 inst_3716 ( .ZN(net_19191), .A2(net_7607), .A1(net_7262) );
INV_X4 inst_15903 ( .A(net_2178), .ZN(net_1767) );
XNOR2_X2 inst_253 ( .ZN(net_17437), .A(net_17287), .B(net_17066) );
INV_X4 inst_16239 ( .ZN(net_16700), .A(net_2554) );
INV_X4 inst_16219 ( .A(net_2321), .ZN(net_2160) );
CLKBUF_X2 inst_21623 ( .A(net_21494), .Z(net_21495) );
INV_X4 inst_14080 ( .A(net_7900), .ZN(net_6219) );
INV_X4 inst_16052 ( .ZN(net_2225), .A(net_1120) );
XNOR2_X2 inst_589 ( .B(net_16607), .ZN(net_566), .A(net_565) );
NAND4_X4 inst_5229 ( .A2(net_20653), .A1(net_20652), .ZN(net_19618), .A4(net_19011), .A3(net_12541) );
INV_X2 inst_18671 ( .ZN(net_13509), .A(net_11393) );
NOR2_X2 inst_4868 ( .ZN(net_3905), .A2(net_2240), .A1(net_1163) );
NAND2_X2 inst_10176 ( .ZN(net_8200), .A1(net_8199), .A2(net_6309) );
NAND2_X2 inst_11969 ( .ZN(net_1825), .A1(net_448), .A2(net_252) );
NOR2_X2 inst_4273 ( .ZN(net_7537), .A2(net_4555), .A1(net_3284) );
INV_X2 inst_18461 ( .ZN(net_12827), .A(net_11817) );
INV_X4 inst_17347 ( .ZN(net_13089), .A(net_1471) );
NAND2_X2 inst_9829 ( .ZN(net_11606), .A2(net_9618), .A1(net_5479) );
NAND2_X2 inst_9822 ( .ZN(net_9641), .A2(net_9640), .A1(net_6993) );
OAI21_X2 inst_1877 ( .A(net_15649), .ZN(net_13687), .B2(net_13641), .B1(net_11109) );
XNOR2_X2 inst_59 ( .ZN(net_18834), .A(net_18781), .B(net_18687) );
INV_X2 inst_19463 ( .ZN(net_1476), .A(net_1475) );
OAI211_X4 inst_2367 ( .C2(net_20912), .ZN(net_18073), .B(net_18049), .C1(net_16372), .A(net_10373) );
CLKBUF_X2 inst_21473 ( .A(net_21344), .Z(net_21345) );
NAND2_X2 inst_9182 ( .ZN(net_13258), .A2(net_10615), .A1(net_6582) );
NAND2_X2 inst_10533 ( .A1(net_10238), .A2(net_8476), .ZN(net_6814) );
NOR2_X4 inst_3256 ( .A1(net_8490), .ZN(net_2263), .A2(net_252) );
CLKBUF_X2 inst_21419 ( .A(net_21290), .Z(net_21291) );
NAND2_X2 inst_9050 ( .ZN(net_14019), .A2(net_11949), .A1(net_816) );
INV_X4 inst_12867 ( .A(net_17014), .ZN(net_16977) );
OAI21_X2 inst_1865 ( .ZN(net_13757), .B2(net_11111), .A(net_10098), .B1(net_6292) );
INV_X4 inst_15715 ( .ZN(net_2573), .A(net_333) );
XOR2_X2 inst_37 ( .A(net_21168), .Z(net_654), .B(net_653) );
NAND3_X2 inst_6390 ( .ZN(net_12009), .A3(net_9520), .A2(net_7939), .A1(net_6466) );
NAND2_X2 inst_11960 ( .ZN(net_3219), .A1(net_1848), .A2(net_1583) );
OAI21_X2 inst_1664 ( .ZN(net_19890), .A(net_15612), .B2(net_15095), .B1(net_14510) );
OAI21_X4 inst_1447 ( .ZN(net_19361), .B1(net_15692), .B2(net_15037), .A(net_13838) );
INV_X4 inst_14881 ( .A(net_5208), .ZN(net_3680) );
NAND2_X2 inst_9601 ( .ZN(net_13431), .A1(net_10756), .A2(net_7369) );
AOI21_X2 inst_20391 ( .ZN(net_15464), .A(net_15463), .B1(net_14466), .B2(net_14455) );
NOR2_X2 inst_4730 ( .ZN(net_3982), .A2(net_3082), .A1(net_3014) );
NOR2_X4 inst_3075 ( .A2(net_20572), .ZN(net_5904), .A1(net_4735) );
NOR3_X1 inst_2800 ( .A3(net_11088), .A2(net_10891), .ZN(net_6534), .A1(net_6533) );
NAND2_X2 inst_9487 ( .ZN(net_14336), .A1(net_13462), .A2(net_9393) );
SDFF_X2 inst_766 ( .Q(net_20964), .SE(net_18847), .SI(net_18508), .D(net_423), .CK(net_22176) );
OAI21_X2 inst_1908 ( .ZN(net_13109), .A(net_12440), .B1(net_9740), .B2(net_6678) );
NOR2_X4 inst_3270 ( .ZN(net_4322), .A1(net_3054), .A2(net_2294) );
INV_X4 inst_14879 ( .ZN(net_12474), .A(net_4670) );
INV_X4 inst_15957 ( .ZN(net_11451), .A(net_7087) );
DFF_X1 inst_19870 ( .D(net_17037), .CK(net_22098), .Q(x392) );
NOR2_X4 inst_3273 ( .ZN(net_2143), .A1(net_1314), .A2(net_129) );
CLKBUF_X2 inst_22568 ( .A(net_22439), .Z(net_22440) );
NAND3_X2 inst_6139 ( .ZN(net_20135), .A2(net_19998), .A1(net_13716), .A3(net_8069) );
NAND2_X2 inst_9943 ( .ZN(net_9065), .A1(net_9064), .A2(net_5705) );
CLKBUF_X2 inst_22105 ( .A(net_21976), .Z(net_21977) );
INV_X2 inst_19527 ( .A(net_1503), .ZN(net_1045) );
INV_X4 inst_14282 ( .ZN(net_6075), .A(net_5643) );
NAND3_X2 inst_6552 ( .A3(net_14384), .ZN(net_10529), .A2(net_9690), .A1(net_6378) );
OAI21_X2 inst_1619 ( .ZN(net_20353), .A(net_16187), .B1(net_15606), .B2(net_15484) );
INV_X4 inst_15344 ( .ZN(net_10690), .A(net_6990) );
XNOR2_X2 inst_441 ( .ZN(net_15960), .A(net_15959), .B(net_15295) );
NOR2_X4 inst_3110 ( .ZN(net_6851), .A2(net_4066), .A1(net_874) );
INV_X2 inst_19001 ( .A(net_6443), .ZN(net_6195) );
NAND3_X2 inst_6201 ( .A3(net_20600), .ZN(net_13305), .A2(net_13304), .A1(net_13170) );
NAND2_X2 inst_8425 ( .A2(net_19458), .ZN(net_17181), .A1(net_16727) );
NAND2_X2 inst_11414 ( .A2(net_7077), .ZN(net_3407), .A1(net_3406) );
NAND4_X4 inst_5228 ( .A4(net_18935), .A1(net_18934), .ZN(net_18908), .A2(net_15268), .A3(net_12953) );
INV_X4 inst_16256 ( .ZN(net_4762), .A(net_874) );
CLKBUF_X2 inst_22863 ( .A(net_22734), .Z(net_22735) );
SDFF_X2 inst_808 ( .Q(net_20944), .SE(net_18025), .D(net_17935), .SI(net_564), .CK(net_21255) );
INV_X2 inst_18622 ( .ZN(net_9568), .A(net_9567) );
NOR2_X2 inst_3859 ( .A1(net_11536), .ZN(net_11454), .A2(net_10610) );
INV_X4 inst_18159 ( .A(net_21060), .ZN(net_653) );
NAND2_X2 inst_9683 ( .A1(net_11918), .ZN(net_10258), .A2(net_6703) );
INV_X4 inst_16068 ( .ZN(net_3246), .A(net_1287) );
OAI21_X4 inst_1383 ( .A(net_16357), .ZN(net_16346), .B1(net_16101), .B2(net_15232) );
NOR2_X4 inst_2838 ( .A2(net_20366), .A1(net_20365), .ZN(net_19591) );
NAND3_X2 inst_6153 ( .ZN(net_13674), .A3(net_12413), .A1(net_9245), .A2(net_6179) );
CLKBUF_X2 inst_22962 ( .A(net_22833), .Z(net_22834) );
AOI21_X2 inst_20861 ( .B1(net_19252), .ZN(net_8840), .B2(net_5899), .A(net_1061) );
NOR2_X4 inst_2833 ( .A2(net_20127), .A1(net_20126), .ZN(net_19266) );
NOR2_X2 inst_3423 ( .ZN(net_19794), .A2(net_15144), .A1(net_15080) );
INV_X4 inst_15349 ( .A(net_3819), .ZN(net_2592) );
INV_X4 inst_16212 ( .ZN(net_14186), .A(net_3156) );
OAI21_X2 inst_2042 ( .ZN(net_11200), .B1(net_5925), .B2(net_4800), .A(net_178) );
CLKBUF_X2 inst_22604 ( .A(net_22475), .Z(net_22476) );
INV_X2 inst_19201 ( .A(net_4991), .ZN(net_4416) );
NAND2_X2 inst_8383 ( .ZN(net_17443), .A1(net_17050), .A2(net_16908) );
INV_X4 inst_16070 ( .ZN(net_1569), .A(net_1453) );
NAND2_X2 inst_8248 ( .A2(net_20463), .ZN(net_17714), .A1(net_17320) );
AND2_X2 inst_21352 ( .ZN(net_2191), .A2(net_2190), .A1(net_1791) );
INV_X2 inst_19186 ( .ZN(net_3732), .A(net_3731) );
AOI21_X4 inst_20107 ( .B1(net_19302), .ZN(net_18956), .B2(net_16187), .A(net_16070) );
INV_X4 inst_15503 ( .ZN(net_4252), .A(net_2420) );
CLKBUF_X2 inst_22853 ( .A(net_22724), .Z(net_22725) );
NOR2_X1 inst_5156 ( .ZN(net_20734), .A2(net_6585), .A1(net_4696) );
INV_X4 inst_13361 ( .ZN(net_10942), .A(net_10941) );
INV_X4 inst_15383 ( .A(net_15183), .ZN(net_2553) );
NAND3_X2 inst_6107 ( .ZN(net_13894), .A3(net_12117), .A1(net_11415), .A2(net_9675) );
NAND2_X2 inst_10758 ( .A2(net_12915), .ZN(net_7214), .A1(net_6712) );
NOR3_X2 inst_2796 ( .A2(net_6905), .A3(net_5265), .ZN(net_3215), .A1(net_3214) );
NOR3_X2 inst_2729 ( .ZN(net_13243), .A2(net_12770), .A1(net_10594), .A3(net_4692) );
NAND2_X2 inst_10587 ( .A1(net_9968), .A2(net_8429), .ZN(net_6660) );
NAND2_X2 inst_8364 ( .ZN(net_17375), .A2(net_17344), .A1(net_17294) );
NAND2_X2 inst_8842 ( .A1(net_15501), .ZN(net_15440), .A2(net_15023) );
OAI21_X2 inst_1815 ( .ZN(net_14169), .B2(net_10729), .B1(net_5353), .A(net_3396) );
NAND4_X2 inst_5267 ( .ZN(net_16168), .A4(net_15695), .A2(net_13860), .A1(net_13722), .A3(net_12936) );
INV_X4 inst_13187 ( .ZN(net_14220), .A(net_13618) );
NAND2_X2 inst_10422 ( .A1(net_14055), .ZN(net_7225), .A2(net_5501) );
INV_X4 inst_16826 ( .A(net_995), .ZN(net_991) );
INV_X4 inst_16788 ( .ZN(net_19229), .A(net_1014) );
AND2_X2 inst_21285 ( .A1(net_14301), .ZN(net_12967), .A2(net_10201) );
NAND2_X4 inst_7010 ( .A2(net_19263), .A1(net_19262), .ZN(net_17178) );
INV_X4 inst_17850 ( .ZN(net_791), .A(net_703) );
INV_X8 inst_12379 ( .ZN(net_684), .A(net_212) );
NAND3_X2 inst_6708 ( .ZN(net_7112), .A3(net_7111), .A1(net_3917), .A2(net_3898) );
INV_X2 inst_19710 ( .A(net_20708), .ZN(net_20707) );
NAND2_X2 inst_10840 ( .ZN(net_7203), .A1(net_6089), .A2(net_5560) );
NAND2_X2 inst_10319 ( .A1(net_11617), .A2(net_11057), .ZN(net_10172) );
NAND4_X2 inst_5442 ( .ZN(net_13886), .A2(net_13885), .A3(net_13697), .A4(net_11330), .A1(net_4882) );
INV_X4 inst_17555 ( .ZN(net_5754), .A(net_809) );
AOI21_X2 inst_20794 ( .B1(net_11654), .ZN(net_10469), .B2(net_7904), .A(net_5038) );
NOR2_X2 inst_4758 ( .ZN(net_5492), .A1(net_3063), .A2(net_2082) );
NAND2_X2 inst_9857 ( .A1(net_10108), .ZN(net_9508), .A2(net_5858) );
NOR2_X2 inst_3875 ( .ZN(net_20821), .A2(net_9359), .A1(net_3005) );
INV_X4 inst_15187 ( .A(net_4162), .ZN(net_2937) );
NOR3_X4 inst_2629 ( .A3(net_20338), .A1(net_20337), .ZN(net_14832), .A2(net_9352) );
NAND2_X2 inst_8989 ( .ZN(net_14468), .A2(net_12747), .A1(net_1864) );
INV_X4 inst_16421 ( .ZN(net_12620), .A(net_11311) );
INV_X4 inst_13658 ( .ZN(net_9628), .A(net_8134) );
CLKBUF_X2 inst_22911 ( .A(net_22782), .Z(net_22783) );
INV_X2 inst_19542 ( .ZN(net_1818), .A(net_1785) );
NAND2_X2 inst_9732 ( .ZN(net_10112), .A2(net_10111), .A1(net_8236) );
INV_X4 inst_14342 ( .ZN(net_20412), .A(net_5357) );
AOI211_X2 inst_21059 ( .ZN(net_10811), .B(net_10810), .C2(net_7681), .A(net_4453), .C1(net_2240) );
NAND2_X2 inst_9595 ( .ZN(net_10846), .A2(net_9220), .A1(net_3942) );
INV_X2 inst_19585 ( .ZN(net_345), .A(net_344) );
NAND2_X4 inst_7235 ( .A2(net_10034), .ZN(net_8371), .A1(net_3682) );
OAI221_X2 inst_1341 ( .C1(net_15340), .ZN(net_13928), .B1(net_13565), .A(net_11544), .B2(net_11338), .C2(net_6460) );
XNOR2_X2 inst_587 ( .B(net_11888), .ZN(net_575), .A(net_574) );
CLKBUF_X2 inst_21851 ( .A(net_21722), .Z(net_21723) );
XNOR2_X2 inst_666 ( .B(net_21149), .A(net_21117), .ZN(net_12268) );
NAND2_X2 inst_10798 ( .ZN(net_10477), .A2(net_5563), .A1(net_2996) );
INV_X2 inst_18673 ( .ZN(net_9119), .A(net_9118) );
NAND3_X2 inst_5937 ( .ZN(net_14920), .A1(net_13624), .A2(net_12233), .A3(net_12126) );
NAND2_X4 inst_7182 ( .ZN(net_10867), .A2(net_10139), .A1(net_7230) );
INV_X2 inst_19432 ( .ZN(net_1769), .A(net_1768) );
OAI21_X2 inst_1829 ( .ZN(net_14137), .B2(net_10466), .B1(net_9910), .A(net_8734) );
NAND3_X2 inst_6446 ( .ZN(net_11796), .A2(net_11795), .A3(net_11794), .A1(net_8139) );
NAND2_X2 inst_9868 ( .ZN(net_9482), .A1(net_7903), .A2(net_6164) );
NAND2_X4 inst_7368 ( .A1(net_20693), .ZN(net_5180), .A2(net_4090) );
AOI21_X2 inst_20824 ( .ZN(net_9877), .B1(net_7661), .B2(net_5075), .A(net_3050) );
INV_X8 inst_12376 ( .A(net_1697), .ZN(net_310) );
NAND4_X2 inst_5252 ( .A4(net_19021), .A1(net_19020), .ZN(net_18608), .A2(net_16122), .A3(net_10365) );
NAND2_X4 inst_7594 ( .A1(net_19038), .ZN(net_3287), .A2(net_321) );
NAND2_X2 inst_11217 ( .ZN(net_8444), .A2(net_3944), .A1(net_2375) );
NAND2_X2 inst_11939 ( .ZN(net_3178), .A2(net_1451), .A1(net_225) );
INV_X8 inst_12210 ( .ZN(net_7466), .A(net_4827) );
INV_X4 inst_13547 ( .ZN(net_9186), .A(net_9185) );
INV_X2 inst_19052 ( .A(net_6700), .ZN(net_4734) );
INV_X4 inst_17507 ( .ZN(net_1018), .A(net_916) );
NOR2_X4 inst_3315 ( .ZN(net_2590), .A2(net_987), .A1(net_894) );
NAND2_X4 inst_7347 ( .A1(net_5291), .ZN(net_4827), .A2(net_4099) );
AOI211_X2 inst_21032 ( .ZN(net_14376), .C1(net_13996), .B(net_12795), .A(net_12059), .C2(net_6456) );
NAND2_X2 inst_7753 ( .ZN(net_18773), .A2(net_18747), .A1(net_18725) );
INV_X4 inst_15783 ( .ZN(net_10298), .A(net_8186) );
INV_X2 inst_18426 ( .ZN(net_15080), .A(net_14679) );
NAND2_X2 inst_11652 ( .ZN(net_2446), .A1(net_2077), .A2(net_1763) );
INV_X4 inst_13094 ( .ZN(net_15875), .A(net_15743) );
INV_X4 inst_14809 ( .ZN(net_4998), .A(net_3969) );
CLKBUF_X2 inst_21803 ( .A(net_21674), .Z(net_21675) );
XNOR2_X2 inst_343 ( .ZN(net_16962), .A(net_16952), .B(net_16095) );
NAND2_X2 inst_10431 ( .ZN(net_7211), .A1(net_7210), .A2(net_5441) );
NOR2_X2 inst_4739 ( .ZN(net_5488), .A2(net_3057), .A1(net_1962) );
OR2_X4 inst_1106 ( .ZN(net_8563), .A1(net_1740), .A2(net_573) );
XNOR2_X2 inst_543 ( .ZN(net_747), .A(net_746), .B(net_745) );
AND4_X2 inst_21104 ( .A4(net_12093), .ZN(net_11844), .A2(net_11843), .A1(net_4345), .A3(net_2622) );
INV_X2 inst_19498 ( .A(net_15649), .ZN(net_1275) );
NAND2_X1 inst_12131 ( .ZN(net_18274), .A2(net_18273), .A1(net_17752) );
INV_X2 inst_19270 ( .A(net_4295), .ZN(net_3058) );
INV_X4 inst_14194 ( .ZN(net_10449), .A(net_7921) );
NAND2_X4 inst_6882 ( .ZN(net_18256), .A1(net_18117), .A2(net_18100) );
INV_X4 inst_13122 ( .ZN(net_15405), .A(net_15149) );
AND2_X2 inst_21367 ( .A2(net_1339), .ZN(net_711), .A1(net_170) );
INV_X4 inst_16915 ( .ZN(net_8521), .A(net_4111) );
OAI21_X2 inst_2070 ( .A(net_13984), .ZN(net_10626), .B2(net_10625), .B1(net_8583) );
NAND2_X4 inst_7697 ( .A2(net_20702), .ZN(net_760), .A1(net_513) );
NOR2_X4 inst_2890 ( .ZN(net_9607), .A1(net_7507), .A2(net_6585) );
NAND3_X2 inst_5765 ( .ZN(net_20136), .A1(net_15487), .A3(net_14753), .A2(net_7137) );
INV_X4 inst_13858 ( .ZN(net_13910), .A(net_7834) );
AOI21_X4 inst_20115 ( .B1(net_20043), .ZN(net_16285), .B2(net_15731), .A(net_14944) );
NAND3_X2 inst_6337 ( .ZN(net_12432), .A3(net_12431), .A2(net_11826), .A1(net_4875) );
INV_X4 inst_12538 ( .ZN(net_18358), .A(net_18357) );
INV_X4 inst_18292 ( .A(net_20219), .ZN(net_20218) );
INV_X4 inst_16109 ( .ZN(net_15917), .A(net_15831) );
AOI22_X2 inst_19976 ( .ZN(net_15486), .B1(net_14617), .A2(net_14615), .B2(net_11392), .A1(net_1340) );
NAND2_X4 inst_7555 ( .A1(net_20601), .ZN(net_2031), .A2(net_1741) );
CLKBUF_X2 inst_22937 ( .A(net_22808), .Z(net_22809) );
NAND2_X2 inst_8347 ( .ZN(net_19313), .A1(net_17474), .A2(net_17233) );
CLKBUF_X2 inst_22791 ( .A(net_22662), .Z(net_22663) );
NOR2_X2 inst_4304 ( .ZN(net_5936), .A2(net_5935), .A1(net_138) );
NAND2_X4 inst_6848 ( .ZN(net_18640), .A2(net_18602), .A1(net_18588) );
AOI21_X2 inst_20550 ( .B2(net_20815), .B1(net_20814), .ZN(net_14309), .A(net_14308) );
NOR3_X2 inst_2745 ( .ZN(net_12579), .A1(net_11368), .A2(net_11135), .A3(net_4451) );
INV_X4 inst_13810 ( .ZN(net_10636), .A(net_7540) );
AOI21_X2 inst_20413 ( .ZN(net_15292), .B1(net_14190), .B2(net_12722), .A(net_9656) );
INV_X4 inst_16719 ( .ZN(net_6586), .A(net_5565) );
NAND2_X4 inst_7253 ( .ZN(net_10762), .A1(net_4323), .A2(net_3774) );
NAND2_X2 inst_11802 ( .ZN(net_2579), .A1(net_2315), .A2(net_992) );
NAND2_X2 inst_11297 ( .ZN(net_4780), .A2(net_4201), .A1(net_732) );
INV_X4 inst_13125 ( .ZN(net_15387), .A(net_15135) );
INV_X8 inst_12452 ( .A(net_20923), .ZN(net_20558) );
INV_X4 inst_15959 ( .ZN(net_14687), .A(net_14663) );
OR2_X2 inst_1244 ( .ZN(net_647), .A2(net_225), .A1(net_94) );
NOR2_X2 inst_4410 ( .A1(net_9478), .ZN(net_6202), .A2(net_4961) );
NAND2_X2 inst_8134 ( .ZN(net_18037), .A2(net_18026), .A1(net_18018) );
CLKBUF_X2 inst_22327 ( .A(net_22198), .Z(net_22199) );
AND2_X4 inst_21180 ( .A1(net_11898), .ZN(net_11586), .A2(net_9781) );
AND4_X2 inst_21096 ( .ZN(net_14121), .A4(net_13843), .A3(net_11790), .A2(net_11344), .A1(net_7525) );
CLKBUF_X2 inst_22383 ( .A(net_22254), .Z(net_22255) );
XNOR2_X2 inst_582 ( .A(net_21139), .ZN(net_13296), .B(net_595) );
NOR2_X2 inst_4515 ( .ZN(net_13025), .A1(net_8462), .A2(net_4162) );
OAI21_X2 inst_1850 ( .A(net_14203), .ZN(net_14008), .B1(net_11183), .B2(net_8646) );
NOR2_X2 inst_3477 ( .ZN(net_14419), .A1(net_14418), .A2(net_13038) );
OAI21_X2 inst_1950 ( .ZN(net_12571), .B2(net_11114), .A(net_10292), .B1(net_3993) );
NAND2_X2 inst_12057 ( .A2(net_2585), .ZN(net_891), .A1(net_890) );
NAND4_X2 inst_5287 ( .ZN(net_15943), .A4(net_15194), .A1(net_15034), .A2(net_14708), .A3(net_12571) );
NAND2_X4 inst_7690 ( .ZN(net_1023), .A2(net_766), .A1(net_177) );
NAND2_X2 inst_9402 ( .ZN(net_11686), .A2(net_11070), .A1(net_6194) );
INV_X4 inst_16606 ( .ZN(net_15524), .A(net_60) );
NAND2_X4 inst_7292 ( .ZN(net_9066), .A2(net_7149), .A1(net_1033) );
INV_X4 inst_12673 ( .ZN(net_17743), .A(net_17742) );
INV_X4 inst_14727 ( .A(net_5547), .ZN(net_4124) );
INV_X4 inst_17907 ( .ZN(net_1711), .A(net_856) );
INV_X4 inst_17094 ( .A(net_15454), .ZN(net_14046) );
OAI21_X2 inst_1779 ( .ZN(net_14667), .B2(net_11938), .B1(net_10214), .A(net_652) );
INV_X2 inst_19025 ( .ZN(net_8086), .A(net_6825) );
NAND2_X4 inst_7299 ( .ZN(net_10475), .A2(net_9785), .A1(net_5559) );
OAI21_X2 inst_2115 ( .ZN(net_10033), .B2(net_9832), .B1(net_5820), .A(net_308) );
INV_X2 inst_18638 ( .ZN(net_11480), .A(net_9383) );
INV_X4 inst_15910 ( .ZN(net_1757), .A(net_1756) );
OAI21_X2 inst_1728 ( .ZN(net_15086), .B2(net_12855), .B1(net_6731), .A(net_333) );
XNOR2_X2 inst_112 ( .ZN(net_18513), .A(net_18372), .B(net_17497) );
NOR2_X4 inst_3251 ( .ZN(net_2540), .A2(net_1493), .A1(net_63) );
NAND2_X2 inst_11161 ( .ZN(net_5229), .A1(net_4301), .A2(net_4184) );
INV_X2 inst_19538 ( .A(net_4211), .ZN(net_966) );
AOI21_X2 inst_20563 ( .ZN(net_19510), .A(net_14572), .B2(net_12421), .B1(net_4354) );
NAND2_X2 inst_9824 ( .ZN(net_20452), .A1(net_9634), .A2(net_9633) );
NAND2_X2 inst_9523 ( .ZN(net_11127), .A1(net_11126), .A2(net_7554) );
NAND2_X4 inst_7441 ( .ZN(net_4291), .A1(net_2934), .A2(net_2289) );
NAND2_X2 inst_8376 ( .ZN(net_19009), .A1(net_17355), .A2(net_17215) );
CLKBUF_X2 inst_22093 ( .A(net_21964), .Z(net_21965) );
NOR3_X2 inst_2724 ( .ZN(net_13251), .A2(net_13246), .A1(net_10586), .A3(net_4362) );
AOI21_X2 inst_20893 ( .ZN(net_20627), .B1(net_9617), .B2(net_6357), .A(net_6348) );
AOI21_X4 inst_20192 ( .B1(net_19657), .ZN(net_15165), .B2(net_12133), .A(net_9757) );
NAND2_X2 inst_9353 ( .ZN(net_12170), .A1(net_12169), .A2(net_12168) );
NAND2_X4 inst_7067 ( .A2(net_20848), .A1(net_19087), .ZN(net_16239) );
NAND2_X2 inst_11334 ( .ZN(net_8094), .A2(net_3658), .A1(net_2104) );
NAND2_X2 inst_12010 ( .A1(net_3862), .ZN(net_1140), .A2(net_341) );
NAND3_X2 inst_5751 ( .ZN(net_16005), .A3(net_15623), .A2(net_13989), .A1(net_8794) );
NAND2_X2 inst_8062 ( .ZN(net_18196), .A2(net_18131), .A1(net_18114) );
AND2_X4 inst_21257 ( .ZN(net_1754), .A2(net_1630), .A1(net_1002) );
NAND2_X2 inst_10213 ( .ZN(net_8092), .A1(net_8091), .A2(net_6048) );
XNOR2_X2 inst_382 ( .ZN(net_16803), .A(net_16802), .B(net_15799) );
NAND2_X2 inst_9387 ( .ZN(net_11934), .A1(net_9452), .A2(net_7327) );
OAI21_X2 inst_2329 ( .ZN(net_5286), .B1(net_5285), .B2(net_5284), .A(net_3867) );
AOI221_X2 inst_20086 ( .ZN(net_15841), .C1(net_15840), .B1(net_15522), .C2(net_14926), .B2(net_14881), .A(net_9481) );
CLKBUF_X2 inst_22072 ( .A(net_21943), .Z(net_21944) );
INV_X4 inst_18294 ( .ZN(net_20438), .A(net_20434) );
NAND3_X2 inst_6101 ( .ZN(net_20347), .A2(net_12992), .A3(net_10353), .A1(net_9471) );
NAND2_X4 inst_7161 ( .A1(net_9754), .ZN(net_9524), .A2(net_6223) );
NAND2_X2 inst_10361 ( .ZN(net_7429), .A1(net_7428), .A2(net_4533) );
INV_X4 inst_17548 ( .A(net_442), .ZN(net_368) );
NAND3_X2 inst_6067 ( .ZN(net_14129), .A3(net_10559), .A2(net_7194), .A1(net_5753) );
NAND2_X2 inst_10560 ( .ZN(net_8710), .A2(net_6855), .A1(net_6719) );
INV_X4 inst_15040 ( .ZN(net_4407), .A(net_3341) );
SDFF_X2 inst_1049 ( .QN(net_20994), .SE(net_2426), .D(net_1856), .CK(net_22645), .SI(x3117) );
NAND2_X2 inst_8418 ( .ZN(net_17469), .A1(net_16915), .A2(net_16726) );
NOR2_X2 inst_5116 ( .A1(net_972), .ZN(net_326), .A2(net_325) );
INV_X4 inst_17421 ( .ZN(net_3886), .A(net_146) );
NAND2_X2 inst_8085 ( .A1(net_21204), .ZN(net_20279), .A2(net_18140) );
NOR2_X2 inst_4575 ( .ZN(net_6855), .A1(net_1848), .A2(net_1578) );
INV_X4 inst_17085 ( .ZN(net_812), .A(net_811) );
NAND3_X2 inst_6037 ( .ZN(net_14328), .A3(net_14327), .A2(net_11474), .A1(net_7990) );
INV_X4 inst_13819 ( .A(net_9741), .ZN(net_7516) );
NAND2_X2 inst_10547 ( .A1(net_7489), .ZN(net_6753), .A2(net_5268) );
NAND3_X4 inst_5613 ( .ZN(net_20082), .A3(net_8922), .A2(net_8072), .A1(net_8043) );
INV_X8 inst_12258 ( .ZN(net_3501), .A(net_2430) );
INV_X2 inst_18749 ( .ZN(net_7843), .A(net_7842) );
CLKBUF_X2 inst_22199 ( .A(net_21566), .Z(net_22071) );
NAND2_X2 inst_9643 ( .ZN(net_19868), .A1(net_10383), .A2(net_9814) );
INV_X4 inst_15113 ( .ZN(net_3494), .A(net_3188) );
XNOR2_X2 inst_580 ( .B(net_11888), .ZN(net_605), .A(net_604) );
NAND2_X2 inst_9249 ( .A1(net_12784), .ZN(net_12668), .A2(net_10984) );
INV_X4 inst_13533 ( .ZN(net_10779), .A(net_9215) );
INV_X4 inst_16519 ( .ZN(net_1424), .A(net_1403) );
INV_X4 inst_16384 ( .ZN(net_1278), .A(net_807) );
INV_X4 inst_18217 ( .A(net_20978), .ZN(net_2277) );
NAND2_X4 inst_7336 ( .ZN(net_7902), .A2(net_4910), .A1(net_4324) );
INV_X4 inst_12647 ( .ZN(net_17973), .A(net_17874) );
NAND2_X2 inst_11304 ( .ZN(net_4547), .A2(net_3530), .A1(net_809) );
INV_X2 inst_19646 ( .A(net_19447), .ZN(net_19446) );
INV_X4 inst_18128 ( .A(net_21125), .ZN(net_738) );
NOR2_X2 inst_3616 ( .ZN(net_20814), .A1(net_12372), .A2(net_6574) );
NAND2_X2 inst_8746 ( .ZN(net_19071), .A1(net_15826), .A2(net_14737) );
NAND2_X2 inst_9103 ( .ZN(net_13736), .A1(net_12394), .A2(net_11383) );
INV_X4 inst_13842 ( .A(net_9574), .ZN(net_9156) );
NOR3_X2 inst_2692 ( .ZN(net_20379), .A1(net_12648), .A2(net_12148), .A3(net_8070) );
INV_X4 inst_17101 ( .ZN(net_1934), .A(net_825) );
INV_X4 inst_13580 ( .ZN(net_11422), .A(net_8084) );
OAI21_X2 inst_1599 ( .A(net_21228), .ZN(net_16180), .B2(net_15794), .B1(net_10043) );
NOR2_X2 inst_3565 ( .ZN(net_12831), .A1(net_10147), .A2(net_7290) );
NOR2_X2 inst_5026 ( .ZN(net_3776), .A2(net_1164), .A1(net_133) );
NAND2_X4 inst_7348 ( .ZN(net_5991), .A1(net_4826), .A2(net_498) );
NAND2_X2 inst_8055 ( .ZN(net_20615), .A1(net_19902), .A2(net_18211) );
INV_X4 inst_14141 ( .ZN(net_9410), .A(net_6075) );
NAND3_X2 inst_5687 ( .ZN(net_16296), .A3(net_16018), .A1(net_15915), .A2(net_15640) );
NAND2_X2 inst_7922 ( .ZN(net_18452), .A1(net_18451), .A2(net_18373) );
INV_X2 inst_18744 ( .ZN(net_7896), .A(net_7895) );
NAND2_X4 inst_6960 ( .ZN(net_17552), .A1(net_17051), .A2(net_16914) );
NOR2_X2 inst_3977 ( .ZN(net_8396), .A1(net_6303), .A2(net_4765) );
NAND2_X2 inst_8629 ( .ZN(net_16595), .A2(net_16594), .A1(net_16517) );
OAI211_X2 inst_2593 ( .B(net_5511), .C2(net_5510), .ZN(net_5267), .A(net_1854), .C1(net_455) );
NAND2_X2 inst_11717 ( .A1(net_4108), .ZN(net_3717), .A2(net_1921) );
NOR2_X2 inst_5021 ( .A2(net_20868), .ZN(net_1198), .A1(net_779) );
NAND2_X2 inst_9850 ( .A1(net_11468), .A2(net_11418), .ZN(net_9531) );
INV_X4 inst_13550 ( .ZN(net_10742), .A(net_9171) );
CLKBUF_X2 inst_21666 ( .A(net_21537), .Z(net_21538) );
XNOR2_X2 inst_318 ( .ZN(net_17043), .A(net_17040), .B(net_13946) );
INV_X2 inst_19494 ( .A(net_10381), .ZN(net_1286) );
INV_X4 inst_18055 ( .A(net_21189), .ZN(net_9235) );
AOI22_X2 inst_19996 ( .ZN(net_14366), .A1(net_14365), .A2(net_12479), .B2(net_5650), .B1(net_2682) );
NOR2_X2 inst_4065 ( .A1(net_10947), .ZN(net_7792), .A2(net_7791) );
OAI21_X4 inst_1486 ( .ZN(net_19283), .A(net_13703), .B1(net_13657), .B2(net_11739) );
INV_X4 inst_13790 ( .ZN(net_9200), .A(net_7565) );
OAI21_X2 inst_2281 ( .ZN(net_6865), .A(net_6097), .B2(net_2643), .B1(net_2216) );
INV_X4 inst_13449 ( .ZN(net_14902), .A(net_9755) );
OR2_X2 inst_1175 ( .ZN(net_8969), .A1(net_5734), .A2(net_5733) );
INV_X4 inst_12666 ( .ZN(net_17802), .A(net_17801) );
INV_X4 inst_13929 ( .A(net_8982), .ZN(net_6866) );
INV_X4 inst_16778 ( .ZN(net_19347), .A(net_1022) );
NAND3_X2 inst_5877 ( .ZN(net_19836), .A1(net_14506), .A3(net_12280), .A2(net_2536) );
NAND4_X2 inst_5256 ( .ZN(net_19438), .A3(net_16311), .A4(net_16235), .A1(net_15973), .A2(net_14353) );
MUX2_X2 inst_12164 ( .Z(net_11911), .B(net_11910), .S(net_11909), .A(net_11836) );
INV_X8 inst_12208 ( .ZN(net_10647), .A(net_7337) );
NAND2_X2 inst_8305 ( .A2(net_20509), .ZN(net_17587), .A1(net_16839) );
NOR2_X2 inst_4509 ( .ZN(net_6633), .A1(net_3791), .A2(net_381) );
NAND2_X2 inst_8962 ( .ZN(net_14688), .A1(net_14687), .A2(net_13313) );
XNOR2_X2 inst_395 ( .A(net_16769), .ZN(net_16763), .B(net_13285) );
INV_X4 inst_17634 ( .A(net_20851), .ZN(net_732) );
SDFF_X2 inst_841 ( .Q(net_21144), .SI(net_17319), .SE(net_125), .CK(net_21665), .D(x3491) );
INV_X4 inst_14106 ( .ZN(net_12566), .A(net_6168) );
NOR2_X2 inst_3963 ( .ZN(net_8578), .A1(net_5417), .A2(net_3871) );
NAND2_X4 inst_7328 ( .ZN(net_5059), .A1(net_5057), .A2(net_4108) );
INV_X4 inst_13682 ( .ZN(net_10197), .A(net_7978) );
INV_X4 inst_13412 ( .ZN(net_10329), .A(net_10328) );
NOR2_X2 inst_4895 ( .ZN(net_4177), .A1(net_2585), .A2(net_1183) );
NAND3_X2 inst_6361 ( .ZN(net_12084), .A1(net_10502), .A2(net_8240), .A3(net_7924) );
INV_X4 inst_13538 ( .ZN(net_9205), .A(net_9204) );
AOI22_X2 inst_20011 ( .ZN(net_12441), .B1(net_12440), .A2(net_11104), .A1(net_8485), .B2(net_6019) );
INV_X4 inst_17457 ( .A(net_2001), .ZN(net_819) );
NOR2_X2 inst_3896 ( .ZN(net_9144), .A2(net_6441), .A1(net_4453) );
NOR2_X2 inst_3679 ( .A1(net_14363), .A2(net_12842), .ZN(net_11431) );
OAI21_X2 inst_1558 ( .ZN(net_17563), .B1(net_17404), .A(net_17246), .B2(net_17245) );
INV_X4 inst_14212 ( .ZN(net_9504), .A(net_7906) );
NOR2_X4 inst_2906 ( .ZN(net_8921), .A2(net_6500), .A1(net_5225) );
NAND3_X2 inst_5848 ( .A3(net_19226), .A1(net_19225), .ZN(net_18968), .A2(net_8663) );
INV_X4 inst_14622 ( .ZN(net_8306), .A(net_4407) );
INV_X4 inst_13398 ( .ZN(net_20039), .A(net_9049) );
INV_X4 inst_14206 ( .A(net_7264), .ZN(net_5929) );
NOR2_X2 inst_3886 ( .ZN(net_9246), .A2(net_6306), .A1(net_3330) );
INV_X4 inst_12836 ( .A(net_17275), .ZN(net_17112) );
NAND2_X2 inst_8797 ( .ZN(net_15674), .A2(net_15274), .A1(net_12153) );
NAND2_X2 inst_9072 ( .ZN(net_13974), .A2(net_12199), .A1(net_7162) );
AOI21_X2 inst_20768 ( .ZN(net_10687), .A(net_10686), .B2(net_7036), .B1(net_5341) );
INV_X4 inst_13201 ( .ZN(net_13860), .A(net_13180) );
NAND2_X2 inst_9505 ( .ZN(net_11333), .A2(net_10484), .A1(net_8255) );
NAND2_X2 inst_11692 ( .A1(net_3707), .ZN(net_3103), .A2(net_2325) );
NAND2_X2 inst_10643 ( .A2(net_7787), .ZN(net_7647), .A1(net_4211) );
NAND2_X2 inst_11510 ( .A1(net_6982), .ZN(net_5355), .A2(net_2120) );
NAND2_X2 inst_9890 ( .ZN(net_10909), .A2(net_5986), .A1(net_1790) );
INV_X2 inst_19552 ( .A(net_2788), .ZN(net_893) );
CLKBUF_X2 inst_21834 ( .A(net_21400), .Z(net_21706) );
NAND2_X2 inst_12127 ( .A2(net_2585), .ZN(net_2371), .A1(net_156) );
SDFF_X2 inst_920 ( .Q(net_21235), .SI(net_16478), .SE(net_125), .CK(net_22137), .D(x6832) );
NOR2_X2 inst_3454 ( .ZN(net_14855), .A2(net_14144), .A1(net_1297) );
NAND3_X2 inst_6298 ( .ZN(net_12815), .A2(net_10876), .A3(net_10524), .A1(net_8121) );
INV_X4 inst_18010 ( .A(net_21001), .ZN(net_2511) );
NAND3_X2 inst_5741 ( .ZN(net_20262), .A3(net_19746), .A1(net_19745), .A2(net_15466) );
CLKBUF_X2 inst_22166 ( .A(net_22037), .Z(net_22038) );
NAND3_X2 inst_6571 ( .ZN(net_10466), .A3(net_10465), .A2(net_9041), .A1(net_5890) );
INV_X4 inst_16903 ( .ZN(net_14593), .A(net_14175) );
NAND3_X2 inst_6116 ( .A2(net_14301), .ZN(net_13868), .A3(net_12177), .A1(net_8683) );
NAND2_X2 inst_11629 ( .ZN(net_4295), .A1(net_3332), .A2(net_2296) );
INV_X4 inst_13797 ( .ZN(net_20277), .A(net_9540) );
AOI21_X2 inst_20273 ( .B2(net_20960), .ZN(net_19739), .B1(net_19572), .A(net_13055) );
NOR2_X4 inst_2889 ( .A1(net_14642), .ZN(net_11009), .A2(net_10937) );
INV_X4 inst_14203 ( .ZN(net_9472), .A(net_5942) );
INV_X2 inst_18839 ( .A(net_7280), .ZN(net_6726) );
CLKBUF_X2 inst_22456 ( .A(net_21669), .Z(net_22328) );
INV_X4 inst_16935 ( .ZN(net_7325), .A(net_4900) );
NAND2_X2 inst_10109 ( .ZN(net_8430), .A2(net_5924), .A1(net_1995) );
NAND2_X2 inst_11380 ( .ZN(net_5926), .A2(net_3609), .A1(net_2618) );
INV_X4 inst_15265 ( .A(net_3823), .ZN(net_3541) );
NAND2_X2 inst_8034 ( .ZN(net_19863), .A2(net_18258), .A1(net_89) );
INV_X4 inst_13743 ( .A(net_10348), .ZN(net_7634) );
OAI21_X2 inst_2189 ( .B1(net_20381), .ZN(net_8740), .A(net_8739), .B2(net_6126) );
NAND4_X2 inst_5448 ( .ZN(net_13592), .A1(net_13591), .A3(net_13192), .A2(net_10855), .A4(net_10317) );
XNOR2_X2 inst_315 ( .B(net_21182), .A(net_20500), .ZN(net_17074) );
NOR2_X2 inst_4198 ( .ZN(net_7972), .A2(net_6837), .A1(net_6702) );
CLKBUF_X2 inst_22557 ( .A(net_22428), .Z(net_22429) );
INV_X4 inst_13176 ( .ZN(net_14356), .A(net_13870) );
INV_X4 inst_14989 ( .ZN(net_13023), .A(net_12419) );
XNOR2_X2 inst_216 ( .B(net_20086), .A(net_20085), .ZN(net_17536) );
NAND2_X2 inst_8992 ( .ZN(net_14461), .A1(net_14460), .A2(net_12943) );
CLKBUF_X2 inst_22708 ( .A(net_22579), .Z(net_22580) );
INV_X4 inst_16708 ( .ZN(net_15742), .A(net_1062) );
INV_X4 inst_15126 ( .ZN(net_5752), .A(net_3212) );
INV_X4 inst_14858 ( .ZN(net_4535), .A(net_3788) );
INV_X4 inst_13099 ( .ZN(net_15839), .A(net_15674) );
OAI21_X2 inst_2060 ( .ZN(net_19675), .A(net_10699), .B1(net_8708), .B2(net_6901) );
INV_X4 inst_12987 ( .A(net_17483), .ZN(net_17370) );
NOR3_X2 inst_2680 ( .A3(net_20603), .A1(net_20602), .ZN(net_14579), .A2(net_10281) );
NAND2_X2 inst_8771 ( .ZN(net_19084), .A2(net_15430), .A1(net_12224) );
NAND2_X4 inst_7321 ( .ZN(net_6156), .A1(net_5291), .A2(net_3491) );
NAND2_X2 inst_9225 ( .ZN(net_19364), .A2(net_10165), .A1(net_7355) );
OAI21_X2 inst_1795 ( .ZN(net_14521), .A(net_14083), .B1(net_12427), .B2(net_10356) );
SDFF_X2 inst_828 ( .Q(net_21130), .SI(net_17535), .SE(net_125), .CK(net_21411), .D(x3989) );
INV_X2 inst_19589 ( .A(net_3745), .ZN(net_297) );
NOR2_X2 inst_4697 ( .ZN(net_5646), .A1(net_5516), .A2(net_3175) );
INV_X4 inst_18173 ( .A(net_21000), .ZN(net_450) );
INV_X4 inst_13522 ( .ZN(net_12764), .A(net_9344) );
NAND2_X4 inst_7218 ( .A2(net_19844), .ZN(net_11918), .A1(net_5826) );
INV_X4 inst_17072 ( .ZN(net_7941), .A(net_1099) );
CLKBUF_X2 inst_22500 ( .A(net_22371), .Z(net_22372) );
NOR2_X2 inst_4164 ( .ZN(net_8795), .A2(net_6872), .A1(net_4212) );
INV_X4 inst_15852 ( .ZN(net_3347), .A(net_1016) );
INV_X2 inst_19427 ( .A(net_2328), .ZN(net_1807) );
INV_X4 inst_16446 ( .A(net_9191), .ZN(net_1449) );
INV_X4 inst_17540 ( .ZN(net_19037), .A(net_2744) );
AOI211_X2 inst_21064 ( .C1(net_20845), .ZN(net_9013), .C2(net_4750), .A(net_4551), .B(net_3040) );
NAND2_X2 inst_8899 ( .ZN(net_15101), .A2(net_13945), .A1(net_3943) );
AOI21_X2 inst_20969 ( .B1(net_20573), .ZN(net_19858), .B2(net_3856), .A(net_3125) );
INV_X4 inst_13919 ( .A(net_11587), .ZN(net_8657) );
NAND2_X2 inst_8052 ( .ZN(net_18216), .A2(net_18213), .A1(net_16996) );
NAND2_X2 inst_10854 ( .ZN(net_6738), .A1(net_5458), .A2(net_4266) );
INV_X4 inst_17766 ( .A(net_20875), .ZN(net_547) );
NAND3_X2 inst_6182 ( .ZN(net_13498), .A3(net_13497), .A2(net_12378), .A1(net_6134) );
NAND2_X4 inst_7382 ( .ZN(net_4542), .A1(net_2168), .A2(net_225) );
NAND2_X2 inst_8749 ( .A2(net_19986), .A1(net_19985), .ZN(net_19255) );
CLKBUF_X2 inst_22959 ( .A(net_22830), .Z(net_22831) );
NAND3_X2 inst_6240 ( .ZN(net_19271), .A3(net_12166), .A2(net_11603), .A1(net_8624) );
NAND2_X2 inst_9629 ( .ZN(net_10545), .A2(net_7205), .A1(net_652) );
NAND2_X2 inst_11426 ( .A2(net_3658), .ZN(net_3349), .A1(net_1933) );
NAND2_X2 inst_10127 ( .ZN(net_8353), .A2(net_5156), .A1(net_761) );
NAND2_X2 inst_9137 ( .ZN(net_13443), .A1(net_13442), .A2(net_13371) );
NAND2_X2 inst_10794 ( .A1(net_9754), .ZN(net_5578), .A2(net_4120) );
NAND2_X2 inst_10951 ( .ZN(net_5100), .A1(net_4616), .A2(net_3630) );
NOR2_X4 inst_3050 ( .ZN(net_6169), .A2(net_4394), .A1(net_3524) );
NAND2_X2 inst_11349 ( .ZN(net_3651), .A2(net_3614), .A1(net_1792) );
INV_X4 inst_13916 ( .A(net_14402), .ZN(net_6916) );
NAND2_X2 inst_8491 ( .A1(net_17123), .ZN(net_16956), .A2(net_16801) );
INV_X4 inst_18276 ( .A(net_19458), .ZN(net_19457) );
NOR2_X2 inst_3913 ( .A1(net_13348), .A2(net_10604), .ZN(net_8848) );
INV_X2 inst_19137 ( .ZN(net_4142), .A(net_4141) );
NAND3_X2 inst_5807 ( .ZN(net_15657), .A3(net_14869), .A2(net_13453), .A1(net_11408) );
INV_X4 inst_12625 ( .ZN(net_20234), .A(net_17983) );
NAND2_X4 inst_7484 ( .ZN(net_3308), .A2(net_2117), .A1(net_1990) );
AOI21_X2 inst_20715 ( .ZN(net_12027), .B1(net_11376), .A(net_9761), .B2(net_7733) );
OAI21_X2 inst_1941 ( .A(net_13514), .ZN(net_12769), .B1(net_9108), .B2(net_3223) );
NAND3_X2 inst_6247 ( .ZN(net_13143), .A3(net_12899), .A2(net_10798), .A1(net_4691) );
XOR2_X2 inst_9 ( .B(net_21133), .Z(net_17106), .A(net_17099) );
NOR2_X2 inst_3358 ( .ZN(net_20316), .A2(net_17541), .A1(net_17466) );
NAND3_X2 inst_6719 ( .A3(net_14962), .A1(net_7035), .ZN(net_6535), .A2(net_1447) );
CLKBUF_X2 inst_22308 ( .A(net_22179), .Z(net_22180) );
CLKBUF_X2 inst_21788 ( .A(net_21659), .Z(net_21660) );
INV_X2 inst_18751 ( .ZN(net_10195), .A(net_7810) );
OAI21_X2 inst_1594 ( .A(net_20848), .B2(net_19140), .B1(net_19139), .ZN(net_16234) );
AOI21_X2 inst_20302 ( .B1(net_20944), .ZN(net_19889), .B2(net_15572), .A(net_15531) );
SDFF_X2 inst_902 ( .Q(net_21136), .SE(net_17277), .D(net_16837), .CK(net_21643), .SI(x3771) );
INV_X4 inst_15810 ( .ZN(net_2543), .A(net_1551) );
INV_X2 inst_19266 ( .ZN(net_3104), .A(net_3103) );
NOR2_X2 inst_3489 ( .ZN(net_14266), .A1(net_14201), .A2(net_7340) );
INV_X8 inst_12224 ( .ZN(net_8014), .A(net_5111) );
SDFF_X2 inst_778 ( .Q(net_20904), .SE(net_18863), .SI(net_18406), .D(net_362), .CK(net_22689) );
NAND2_X2 inst_10118 ( .A2(net_10627), .ZN(net_8383), .A1(net_4506) );
INV_X4 inst_16581 ( .ZN(net_1502), .A(net_1152) );
INV_X4 inst_17405 ( .ZN(net_3069), .A(net_732) );
NAND2_X2 inst_7912 ( .ZN(net_18490), .A2(net_18347), .A1(net_18296) );
INV_X4 inst_14842 ( .ZN(net_3853), .A(net_3764) );
NAND2_X2 inst_11486 ( .ZN(net_3117), .A2(net_2891), .A1(net_2102) );
CLKBUF_X2 inst_22949 ( .A(net_22820), .Z(net_22821) );
NAND2_X2 inst_7810 ( .ZN(net_18677), .A2(net_18647), .A1(net_18637) );
NAND2_X2 inst_8845 ( .ZN(net_15421), .A1(net_15100), .A2(net_14601) );
INV_X4 inst_17945 ( .A(net_20887), .ZN(net_202) );
NAND2_X2 inst_8353 ( .A1(net_20774), .ZN(net_17465), .A2(net_17357) );
INV_X4 inst_12855 ( .ZN(net_17061), .A(net_17060) );
INV_X4 inst_13895 ( .ZN(net_7278), .A(net_7277) );
SDFF_X2 inst_781 ( .Q(net_20917), .SE(net_18576), .SI(net_18043), .D(net_592), .CK(net_21289) );
INV_X4 inst_18034 ( .A(net_20935), .ZN(net_121) );
NAND2_X2 inst_12033 ( .ZN(net_1110), .A1(net_949), .A2(net_221) );
NOR2_X2 inst_4042 ( .ZN(net_11150), .A1(net_8068), .A2(net_7899) );
INV_X8 inst_12368 ( .ZN(net_1333), .A(net_255) );
NAND2_X4 inst_7629 ( .ZN(net_1372), .A2(net_1195), .A1(net_879) );
INV_X4 inst_13409 ( .ZN(net_10340), .A(net_10339) );
AOI21_X2 inst_20501 ( .B1(net_15481), .ZN(net_14652), .B2(net_12094), .A(net_11625) );
NOR2_X2 inst_3696 ( .A2(net_20748), .A1(net_20747), .ZN(net_11185) );
NAND2_X2 inst_9450 ( .A2(net_11642), .ZN(net_11524), .A1(net_5403) );
INV_X4 inst_17593 ( .ZN(net_331), .A(net_330) );
CLKBUF_X2 inst_22675 ( .A(net_22094), .Z(net_22547) );
INV_X2 inst_18731 ( .ZN(net_8028), .A(net_8027) );
NAND2_X2 inst_9971 ( .ZN(net_20460), .A1(net_10056), .A2(net_6506) );
INV_X4 inst_16883 ( .ZN(net_1144), .A(net_446) );
NAND2_X4 inst_7053 ( .ZN(net_16422), .A1(net_16312), .A2(net_16292) );
OAI21_X2 inst_1928 ( .A(net_15087), .ZN(net_12953), .B1(net_12952), .B2(net_11593) );
OAI21_X2 inst_1967 ( .B1(net_19144), .ZN(net_12257), .A(net_10981), .B2(net_6334) );
NOR2_X2 inst_4485 ( .A2(net_20467), .A1(net_4707), .ZN(net_4692) );
INV_X4 inst_13733 ( .ZN(net_7730), .A(net_6431) );
NAND2_X4 inst_7659 ( .ZN(net_1503), .A1(net_931), .A2(net_930) );
INV_X4 inst_12944 ( .ZN(net_16632), .A(net_16631) );
OAI21_X2 inst_1947 ( .A(net_12737), .ZN(net_12584), .B1(net_12050), .B2(net_5857) );
NAND2_X2 inst_10967 ( .ZN(net_12908), .A2(net_5032), .A1(net_165) );
NAND2_X4 inst_7318 ( .A2(net_20492), .ZN(net_5137), .A1(net_5109) );
NAND2_X2 inst_8030 ( .ZN(net_18264), .A2(net_18263), .A1(net_17628) );
AOI211_X2 inst_21072 ( .ZN(net_7689), .A(net_7688), .B(net_4802), .C2(net_3308), .C1(net_2593) );
NAND3_X2 inst_6285 ( .A3(net_19927), .A1(net_19460), .ZN(net_12846), .A2(net_12782) );
INV_X4 inst_18186 ( .A(net_21043), .ZN(net_613) );
NOR2_X2 inst_4585 ( .A2(net_4273), .ZN(net_3817), .A1(net_3816) );
NAND2_X2 inst_8105 ( .ZN(net_18114), .A2(net_18093), .A1(net_16882) );
CLKBUF_X2 inst_22668 ( .A(net_22539), .Z(net_22540) );
INV_X4 inst_15143 ( .ZN(net_5437), .A(net_4290) );
INV_X4 inst_18102 ( .A(net_20853), .ZN(net_129) );
NAND2_X2 inst_9126 ( .ZN(net_19812), .A2(net_10788), .A1(net_10082) );
NAND2_X2 inst_9539 ( .A1(net_11505), .ZN(net_11064), .A2(net_11004) );
INV_X2 inst_19141 ( .ZN(net_4127), .A(net_4126) );
INV_X4 inst_15304 ( .ZN(net_4023), .A(net_2335) );
NAND2_X2 inst_11294 ( .A2(net_20801), .ZN(net_11811), .A1(net_3818) );
NAND2_X4 inst_7573 ( .ZN(net_2979), .A2(net_1513), .A1(net_276) );
INV_X4 inst_16830 ( .ZN(net_2524), .A(net_253) );
XNOR2_X2 inst_659 ( .B(net_1896), .A(net_745), .ZN(net_342) );
INV_X4 inst_17194 ( .ZN(net_19661), .A(net_938) );
NAND2_X4 inst_6890 ( .ZN(net_18118), .A2(net_18076), .A1(net_18044) );
INV_X2 inst_19725 ( .A(net_20794), .ZN(net_20793) );
NAND2_X2 inst_11747 ( .ZN(net_3940), .A1(net_2123), .A2(net_2053) );
INV_X4 inst_12868 ( .ZN(net_16971), .A(net_16970) );
INV_X4 inst_12883 ( .ZN(net_17014), .A(net_16821) );
CLKBUF_X2 inst_22243 ( .A(net_22114), .Z(net_22115) );
NAND4_X2 inst_5273 ( .ZN(net_19548), .A1(net_15809), .A4(net_15564), .A3(net_10378), .A2(net_9027) );
NAND2_X2 inst_8094 ( .A2(net_18128), .ZN(net_18127), .A1(net_16576) );
NAND4_X2 inst_5505 ( .A1(net_11379), .ZN(net_11283), .A2(net_11282), .A4(net_11281), .A3(net_3961) );
NAND2_X2 inst_10289 ( .ZN(net_9468), .A1(net_8376), .A2(net_6075) );
NOR2_X4 inst_3199 ( .ZN(net_5559), .A2(net_3034), .A1(net_85) );
NAND3_X2 inst_6178 ( .ZN(net_13540), .A3(net_12962), .A1(net_12478), .A2(net_5821) );
NOR2_X2 inst_3612 ( .ZN(net_12395), .A2(net_9654), .A1(net_7475) );
CLKBUF_X2 inst_22758 ( .A(net_22629), .Z(net_22630) );
OAI21_X2 inst_1581 ( .B2(net_19070), .B1(net_19069), .A(net_16357), .ZN(net_16311) );
INV_X4 inst_17952 ( .A(net_21097), .ZN(net_727) );
OAI21_X2 inst_2312 ( .A(net_8169), .ZN(net_5742), .B2(net_4302), .B1(net_2666) );
NAND4_X2 inst_5336 ( .ZN(net_15518), .A1(net_14518), .A4(net_14517), .A2(net_14334), .A3(net_13122) );
NOR2_X2 inst_3500 ( .ZN(net_14065), .A2(net_11846), .A1(net_4350) );
INV_X4 inst_17248 ( .A(net_2493), .ZN(net_912) );
NAND3_X2 inst_6381 ( .ZN(net_18943), .A1(net_12031), .A2(net_11767), .A3(net_8094) );
NAND2_X2 inst_10526 ( .ZN(net_11915), .A1(net_7528), .A2(net_6841) );
NAND2_X4 inst_7103 ( .ZN(net_13369), .A1(net_7475), .A2(net_2124) );
INV_X2 inst_19232 ( .A(net_7133), .ZN(net_5835) );
AND2_X4 inst_21230 ( .ZN(net_20338), .A2(net_4171), .A1(net_1037) );
OAI21_X2 inst_2241 ( .ZN(net_7383), .A(net_5034), .B1(net_3423), .B2(net_1164) );
INV_X4 inst_13419 ( .ZN(net_20197), .A(net_8770) );
NAND2_X2 inst_8165 ( .ZN(net_17966), .A2(net_17920), .A1(net_17272) );
OAI21_X2 inst_2182 ( .ZN(net_8843), .A(net_8842), .B1(net_4617), .B2(net_4303) );
NAND2_X2 inst_8334 ( .A2(net_20508), .ZN(net_17518), .A1(net_17517) );
INV_X2 inst_19601 ( .A(net_329), .ZN(net_148) );
NOR3_X2 inst_2667 ( .ZN(net_14932), .A2(net_14931), .A1(net_13633), .A3(net_9934) );
INV_X4 inst_17049 ( .ZN(net_12307), .A(net_832) );
SDFF_X2 inst_987 ( .QN(net_21057), .D(net_544), .SE(net_263), .CK(net_22506), .SI(x2103) );
NOR2_X2 inst_4194 ( .ZN(net_6717), .A2(net_6716), .A1(net_3248) );
NAND2_X2 inst_9376 ( .ZN(net_11981), .A1(net_11466), .A2(net_8695) );
NOR2_X4 inst_3006 ( .A2(net_19882), .A1(net_19881), .ZN(net_5763) );
CLKBUF_X2 inst_22200 ( .A(net_22071), .Z(net_22072) );
INV_X4 inst_17026 ( .ZN(net_10810), .A(net_849) );
AOI21_X2 inst_20652 ( .ZN(net_13051), .B2(net_9835), .A(net_8128), .B1(net_5335) );
AND4_X2 inst_21110 ( .A2(net_11629), .ZN(net_11226), .A1(net_11225), .A4(net_11224), .A3(net_8039) );
NAND2_X2 inst_9703 ( .ZN(net_10209), .A1(net_10208), .A2(net_10207) );
INV_X4 inst_18044 ( .A(net_20897), .ZN(net_68) );
INV_X4 inst_15350 ( .A(net_7688), .ZN(net_4200) );
XNOR2_X2 inst_371 ( .A(net_16996), .ZN(net_16844), .B(net_4453) );
AOI21_X2 inst_20309 ( .ZN(net_16036), .B1(net_16035), .B2(net_15518), .A(net_14952) );
NOR2_X2 inst_4962 ( .ZN(net_2657), .A2(net_1615), .A1(net_115) );
NAND3_X2 inst_6498 ( .ZN(net_10850), .A1(net_10844), .A2(net_7370), .A3(net_4798) );
AOI21_X4 inst_20106 ( .B2(net_20888), .B1(net_19218), .ZN(net_16386), .A(net_14271) );
NAND2_X2 inst_10768 ( .ZN(net_5633), .A1(net_5632), .A2(net_4139) );
AOI21_X2 inst_20810 ( .ZN(net_19000), .A(net_15077), .B1(net_11181), .B2(net_4519) );
NOR2_X2 inst_4619 ( .A1(net_4711), .ZN(net_3623), .A2(net_3622) );
CLKBUF_X2 inst_22934 ( .A(net_21631), .Z(net_22806) );
AOI21_X2 inst_20745 ( .A(net_14175), .ZN(net_11402), .B2(net_9082), .B1(net_5704) );
INV_X2 inst_18511 ( .ZN(net_11605), .A(net_10266) );
INV_X4 inst_17301 ( .ZN(net_936), .A(net_801) );
NOR2_X2 inst_3684 ( .ZN(net_11419), .A1(net_11418), .A2(net_9290) );
XNOR2_X2 inst_628 ( .B(net_16680), .ZN(net_14420), .A(net_604) );
NAND2_X4 inst_7470 ( .ZN(net_3583), .A1(net_2641), .A2(net_1014) );
INV_X2 inst_19447 ( .A(net_4457), .ZN(net_1620) );
NOR2_X2 inst_3642 ( .ZN(net_12049), .A1(net_9696), .A2(net_8840) );
NAND2_X2 inst_11873 ( .A2(net_20580), .ZN(net_1631), .A1(net_1630) );
INV_X4 inst_17883 ( .ZN(net_3789), .A(net_77) );
CLKBUF_X2 inst_22188 ( .A(net_22059), .Z(net_22060) );
AOI22_X2 inst_20018 ( .B1(net_20570), .ZN(net_11231), .B2(net_11230), .A1(net_10093), .A2(net_8168) );
NOR2_X4 inst_3092 ( .ZN(net_5421), .A2(net_2541), .A1(net_912) );
NAND3_X2 inst_6587 ( .ZN(net_11564), .A3(net_10225), .A2(net_9571), .A1(net_7568) );
INV_X4 inst_14162 ( .ZN(net_9363), .A(net_4919) );
AOI21_X1 inst_20986 ( .B2(net_10773), .ZN(net_9084), .A(net_9083), .B1(net_9082) );
INV_X4 inst_17911 ( .A(net_1469), .ZN(net_57) );
NOR2_X2 inst_3395 ( .ZN(net_18918), .A1(net_15803), .A2(net_15182) );
OR2_X4 inst_1130 ( .ZN(net_7450), .A2(net_896), .A1(net_117) );
NAND2_X2 inst_9300 ( .A1(net_13538), .ZN(net_12385), .A2(net_11493) );
INV_X4 inst_18239 ( .A(net_21227), .ZN(net_312) );
INV_X2 inst_18617 ( .ZN(net_9604), .A(net_9603) );
INV_X2 inst_18405 ( .A(net_16562), .ZN(net_16409) );
NAND3_X2 inst_6304 ( .ZN(net_12797), .A3(net_10943), .A2(net_9323), .A1(net_8132) );
INV_X4 inst_12706 ( .ZN(net_17589), .A(net_17588) );
INV_X4 inst_17341 ( .ZN(net_6750), .A(net_3842) );
NAND2_X2 inst_7851 ( .A2(net_20936), .ZN(net_18588), .A1(net_16200) );
NAND2_X2 inst_8996 ( .ZN(net_14401), .A2(net_13045), .A1(net_7289) );
INV_X4 inst_15748 ( .A(net_8618), .ZN(net_6990) );
NAND2_X2 inst_11823 ( .ZN(net_2272), .A2(net_1519), .A1(net_167) );
INV_X2 inst_18506 ( .ZN(net_12730), .A(net_11690) );
NAND4_X2 inst_5425 ( .A4(net_19703), .A1(net_19702), .ZN(net_14191), .A2(net_11172), .A3(net_8764) );
NAND2_X2 inst_9304 ( .A1(net_20485), .ZN(net_20376), .A2(net_9221) );
OAI21_X4 inst_1363 ( .A(net_20880), .ZN(net_19883), .B2(net_18902), .B1(net_18901) );
NOR2_X2 inst_4851 ( .ZN(net_13019), .A1(net_8961), .A2(net_6387) );
CLKBUF_X2 inst_22743 ( .A(net_22221), .Z(net_22615) );
INV_X4 inst_18097 ( .A(net_21007), .ZN(net_2403) );
INV_X4 inst_17038 ( .ZN(net_1681), .A(net_956) );
INV_X4 inst_17357 ( .ZN(net_4862), .A(net_3904) );
NAND2_X2 inst_8059 ( .ZN(net_18200), .A1(net_18150), .A2(net_18126) );
INV_X8 inst_12388 ( .ZN(net_880), .A(net_513) );
AOI221_X2 inst_20077 ( .ZN(net_19412), .C1(net_15561), .C2(net_15435), .B2(net_13927), .A(net_13079), .B1(net_4370) );
NAND2_X2 inst_11372 ( .ZN(net_3573), .A1(net_3355), .A2(net_1628) );
NAND2_X2 inst_11806 ( .A2(net_20797), .A1(net_2099), .ZN(net_1891) );
NAND2_X2 inst_11992 ( .ZN(net_7357), .A1(net_1215), .A2(net_1214) );
INV_X4 inst_15736 ( .ZN(net_2762), .A(net_1639) );
OAI21_X2 inst_2127 ( .ZN(net_10001), .B1(net_8250), .A(net_5766), .B2(net_3210) );
NAND3_X2 inst_6688 ( .ZN(net_7708), .A2(net_4232), .A3(net_3245), .A1(net_2538) );
INV_X4 inst_13626 ( .A(net_10440), .ZN(net_9787) );
INV_X4 inst_13689 ( .ZN(net_11717), .A(net_7949) );
NAND2_X2 inst_10611 ( .ZN(net_7857), .A1(net_6599), .A2(net_6572) );
INV_X4 inst_16974 ( .ZN(net_7436), .A(net_3297) );
OAI21_X2 inst_2268 ( .A(net_11018), .ZN(net_7145), .B1(net_7144), .B2(net_5611) );
OAI21_X4 inst_1373 ( .ZN(net_16802), .B1(net_16402), .A(net_16350), .B2(net_16198) );
OAI211_X2 inst_2458 ( .ZN(net_14213), .C2(net_14164), .B(net_13260), .A(net_12647), .C1(net_12457) );
NAND2_X4 inst_7285 ( .A1(net_20497), .ZN(net_7233), .A2(net_6571) );
NAND2_X2 inst_8474 ( .ZN(net_20051), .A2(net_17014), .A1(net_604) );
INV_X4 inst_14303 ( .A(net_11995), .ZN(net_5522) );
NOR2_X4 inst_3155 ( .ZN(net_4057), .A2(net_3225), .A1(net_1011) );
NAND2_X2 inst_9923 ( .ZN(net_9270), .A2(net_6249), .A1(net_3896) );
AOI21_X4 inst_20160 ( .B1(net_19536), .ZN(net_15698), .B2(net_15697), .A(net_13837) );
NOR2_X4 inst_3134 ( .ZN(net_4813), .A1(net_3205), .A2(net_2782) );
NAND4_X2 inst_5481 ( .ZN(net_12749), .A3(net_10204), .A4(net_9568), .A1(net_6612), .A2(net_6096) );
NOR2_X2 inst_4043 ( .ZN(net_9431), .A2(net_5992), .A1(net_703) );
NAND3_X2 inst_6710 ( .ZN(net_7105), .A3(net_7104), .A1(net_3891), .A2(net_3073) );
NAND2_X2 inst_11787 ( .ZN(net_2640), .A2(net_2445), .A1(net_1991) );
AOI22_X2 inst_19965 ( .ZN(net_16038), .B1(net_16037), .A2(net_15520), .B2(net_13153), .A1(net_4467) );
NAND2_X2 inst_8407 ( .ZN(net_17240), .A1(net_17239), .A2(net_17237) );
INV_X2 inst_18647 ( .ZN(net_10798), .A(net_9234) );
NAND2_X2 inst_11999 ( .ZN(net_3027), .A1(net_363), .A2(net_221) );
CLKBUF_X2 inst_22909 ( .A(net_22780), .Z(net_22781) );
NAND3_X2 inst_5755 ( .ZN(net_16002), .A3(net_15626), .A1(net_15489), .A2(net_8525) );
NAND2_X2 inst_11933 ( .A1(net_2636), .ZN(net_2175), .A2(net_836) );
INV_X4 inst_16163 ( .ZN(net_12366), .A(net_8222) );
INV_X4 inst_17432 ( .ZN(net_4795), .A(net_662) );
NAND2_X2 inst_8122 ( .A2(net_18067), .ZN(net_18059), .A1(net_15781) );
AOI21_X2 inst_20340 ( .ZN(net_15782), .B2(net_15142), .A(net_13944), .B1(net_828) );
INV_X4 inst_17620 ( .ZN(net_6669), .A(net_3789) );
CLKBUF_X2 inst_22524 ( .A(net_21602), .Z(net_22396) );
INV_X4 inst_15077 ( .ZN(net_3270), .A(net_3269) );
INV_X4 inst_13435 ( .ZN(net_11136), .A(net_9821) );
INV_X4 inst_15728 ( .ZN(net_10815), .A(net_1960) );
AOI21_X4 inst_20236 ( .ZN(net_12116), .A(net_10714), .B1(net_9140), .B2(net_6959) );
INV_X8 inst_12349 ( .ZN(net_3861), .A(net_315) );
INV_X4 inst_12490 ( .ZN(net_18666), .A(net_18665) );
AND2_X4 inst_21209 ( .A2(net_19324), .ZN(net_8903), .A1(net_6995) );
NOR2_X2 inst_4588 ( .ZN(net_6575), .A2(net_2699), .A1(net_405) );
INV_X4 inst_12755 ( .ZN(net_17690), .A(net_17421) );
INV_X4 inst_13746 ( .A(net_7628), .ZN(net_7627) );
NAND2_X2 inst_9099 ( .ZN(net_13769), .A2(net_13768), .A1(net_12995) );
NOR2_X2 inst_4049 ( .ZN(net_20747), .A2(net_7183), .A1(net_4305) );
NOR3_X2 inst_2702 ( .A3(net_15831), .A2(net_14751), .ZN(net_13924), .A1(net_12019) );
NOR2_X2 inst_5067 ( .ZN(net_12001), .A1(net_475), .A2(net_117) );
INV_X4 inst_15063 ( .ZN(net_5197), .A(net_3298) );
INV_X4 inst_12820 ( .ZN(net_17492), .A(net_17374) );
NOR2_X4 inst_2910 ( .ZN(net_20205), .A2(net_8369), .A1(net_8351) );
NOR2_X2 inst_4670 ( .ZN(net_4297), .A2(net_3162), .A1(net_154) );
NAND3_X2 inst_5701 ( .ZN(net_16218), .A3(net_15906), .A2(net_15259), .A1(net_13833) );
INV_X4 inst_15178 ( .ZN(net_3001), .A(net_3000) );
INV_X4 inst_16586 ( .ZN(net_7087), .A(net_1147) );
XNOR2_X2 inst_145 ( .ZN(net_18168), .A(net_18142), .B(net_18141) );
INV_X4 inst_13703 ( .ZN(net_12903), .A(net_7879) );
NOR2_X2 inst_4594 ( .A1(net_7862), .ZN(net_4764), .A2(net_3784) );
NAND4_X2 inst_5355 ( .ZN(net_15414), .A3(net_15413), .A1(net_14662), .A4(net_13107), .A2(net_8686) );
NAND2_X2 inst_9689 ( .ZN(net_10244), .A1(net_10243), .A2(net_10242) );
INV_X4 inst_15223 ( .A(net_3864), .ZN(net_2866) );
AOI21_X4 inst_20241 ( .B1(net_18964), .ZN(net_11154), .B2(net_10233), .A(net_3485) );
NAND3_X2 inst_6214 ( .A2(net_19769), .ZN(net_19033), .A1(net_13265), .A3(net_13176) );
CLKBUF_X2 inst_22181 ( .A(net_22052), .Z(net_22053) );
NAND2_X2 inst_10199 ( .A1(net_8222), .ZN(net_8132), .A2(net_8131) );
INV_X4 inst_17338 ( .ZN(net_5107), .A(net_4205) );
CLKBUF_X2 inst_21824 ( .A(net_21695), .Z(net_21696) );
OAI21_X4 inst_1437 ( .A(net_16395), .ZN(net_15919), .B1(net_15179), .B2(net_15164) );
NAND4_X2 inst_5345 ( .ZN(net_15436), .A1(net_15413), .A2(net_14362), .A4(net_13090), .A3(net_7160) );
INV_X8 inst_12240 ( .ZN(net_4989), .A(net_2814) );
INV_X4 inst_18006 ( .A(net_21129), .ZN(net_678) );
INV_X4 inst_17483 ( .A(net_731), .ZN(net_433) );
NAND2_X2 inst_9119 ( .ZN(net_13563), .A1(net_13562), .A2(net_13561) );
NAND2_X2 inst_9292 ( .ZN(net_19081), .A2(net_9166), .A1(net_5069) );
NAND2_X2 inst_10557 ( .ZN(net_8942), .A1(net_6706), .A2(net_4953) );
INV_X4 inst_13661 ( .ZN(net_9614), .A(net_8112) );
OAI211_X2 inst_2533 ( .C1(net_11430), .ZN(net_11261), .A(net_11260), .C2(net_9969), .B(net_5194) );
XOR2_X2 inst_27 ( .A(net_21156), .B(net_16501), .Z(net_16499) );
NAND2_X2 inst_8790 ( .ZN(net_18955), .A1(net_15747), .A2(net_15381) );
NAND2_X2 inst_10741 ( .A1(net_10676), .ZN(net_5726), .A2(net_4231) );
NOR2_X2 inst_4446 ( .ZN(net_10285), .A1(net_6599), .A2(net_6466) );
INV_X4 inst_14849 ( .A(net_5629), .ZN(net_3837) );
INV_X2 inst_19600 ( .A(net_304), .ZN(net_151) );
INV_X4 inst_16721 ( .A(net_8724), .ZN(net_8278) );
NAND2_X2 inst_11761 ( .ZN(net_3841), .A2(net_1716), .A1(net_1376) );
NAND2_X2 inst_10063 ( .A1(net_15270), .ZN(net_8677), .A2(net_6804) );
INV_X4 inst_16060 ( .ZN(net_2349), .A(net_1586) );
INV_X4 inst_15397 ( .ZN(net_5468), .A(net_2541) );
INV_X4 inst_15807 ( .ZN(net_2552), .A(net_1374) );
NAND3_X2 inst_6420 ( .ZN(net_20021), .A3(net_11943), .A2(net_9956), .A1(net_9244) );
INV_X4 inst_15879 ( .ZN(net_6135), .A(net_1962) );
NAND4_X4 inst_5230 ( .A2(net_19335), .A1(net_19334), .ZN(net_19218), .A4(net_15836), .A3(net_14237) );
INV_X2 inst_19349 ( .ZN(net_2411), .A(net_2410) );
XNOR2_X2 inst_639 ( .B(net_16842), .ZN(net_416), .A(net_415) );
NAND2_X2 inst_9045 ( .ZN(net_14045), .A2(net_12074), .A1(net_10170) );
INV_X4 inst_14687 ( .ZN(net_4591), .A(net_3583) );
CLKBUF_X2 inst_22506 ( .A(net_22377), .Z(net_22378) );
NOR2_X2 inst_3939 ( .A1(net_8706), .ZN(net_8650), .A2(net_8649) );
INV_X2 inst_19095 ( .ZN(net_4546), .A(net_4545) );
INV_X4 inst_17819 ( .ZN(net_113), .A(net_112) );
OAI21_X2 inst_2167 ( .ZN(net_8953), .B1(net_8952), .B2(net_8951), .A(net_4884) );
NAND2_X4 inst_7008 ( .ZN(net_17154), .A1(net_16692), .A2(net_16691) );
INV_X8 inst_12193 ( .ZN(net_16594), .A(net_16340) );
NAND2_X4 inst_7412 ( .ZN(net_11245), .A2(net_6982), .A1(net_3989) );
NAND3_X2 inst_6328 ( .ZN(net_12491), .A3(net_11138), .A2(net_8831), .A1(net_5837) );
OAI21_X2 inst_1651 ( .A(net_16395), .ZN(net_15886), .B2(net_15318), .B1(net_13130) );
NOR2_X2 inst_4248 ( .A1(net_9558), .ZN(net_6425), .A2(net_1882) );
INV_X4 inst_12561 ( .ZN(net_18243), .A(net_18242) );
INV_X8 inst_12176 ( .ZN(net_18313), .A(net_17215) );
NAND2_X2 inst_8281 ( .ZN(net_19687), .A2(net_17618), .A1(net_17485) );
NAND2_X2 inst_9758 ( .ZN(net_13211), .A1(net_10091), .A2(net_6590) );
INV_X4 inst_15695 ( .ZN(net_3233), .A(net_2020) );
AND2_X2 inst_21306 ( .ZN(net_9554), .A1(net_9553), .A2(net_9552) );
NAND3_X2 inst_6451 ( .ZN(net_11758), .A2(net_11757), .A3(net_10247), .A1(net_3743) );
NAND2_X2 inst_11159 ( .A1(net_7976), .ZN(net_4193), .A2(net_4192) );
OR2_X2 inst_1137 ( .ZN(net_11575), .A1(net_11574), .A2(net_10150) );
INV_X4 inst_15254 ( .ZN(net_3559), .A(net_2138) );
OAI21_X4 inst_1389 ( .A(net_20856), .ZN(net_19899), .B2(net_18931), .B1(net_18930) );
INV_X2 inst_18361 ( .A(net_18183), .ZN(net_18144) );
NAND2_X2 inst_9032 ( .ZN(net_14071), .A1(net_14070), .A2(net_11875) );
INV_X4 inst_14043 ( .ZN(net_7616), .A(net_6260) );
AOI21_X2 inst_20789 ( .A(net_14171), .ZN(net_10544), .B2(net_6718), .B1(net_6251) );
NOR2_X4 inst_3065 ( .ZN(net_8175), .A2(net_3493), .A1(net_2514) );
SDFF_X2 inst_715 ( .Q(net_20890), .SE(net_18837), .SI(net_18780), .D(net_478), .CK(net_22014) );
NAND4_X4 inst_5206 ( .ZN(net_20215), .A3(net_16243), .A4(net_16236), .A1(net_15848), .A2(net_13874) );
INV_X4 inst_14936 ( .A(net_4910), .ZN(net_4569) );
INV_X2 inst_18890 ( .ZN(net_11352), .A(net_6128) );
NAND3_X2 inst_6354 ( .ZN(net_12097), .A2(net_12096), .A3(net_12095), .A1(net_10597) );
NAND2_X4 inst_7333 ( .ZN(net_5901), .A1(net_4208), .A2(net_2809) );
NAND2_X2 inst_8941 ( .ZN(net_14750), .A2(net_13503), .A1(net_12340) );
NAND4_X4 inst_5213 ( .ZN(net_16469), .A4(net_16263), .A1(net_16135), .A3(net_15883), .A2(net_9249) );
INV_X4 inst_14113 ( .ZN(net_6152), .A(net_6151) );
OAI21_X2 inst_1682 ( .B2(net_20831), .B1(net_20830), .ZN(net_15455), .A(net_15454) );
NOR2_X2 inst_5077 ( .ZN(net_10066), .A2(net_888), .A1(net_602) );
CLKBUF_X2 inst_22680 ( .A(net_22325), .Z(net_22552) );
INV_X2 inst_18810 ( .ZN(net_7366), .A(net_7365) );
NAND2_X2 inst_10630 ( .A2(net_8486), .ZN(net_6511), .A1(net_1530) );
INV_X4 inst_13778 ( .A(net_9341), .ZN(net_9150) );
CLKBUF_X2 inst_22582 ( .A(net_22453), .Z(net_22454) );
INV_X4 inst_18191 ( .A(net_20873), .ZN(net_76) );
NOR2_X2 inst_3505 ( .ZN(net_13982), .A2(net_11756), .A1(net_8765) );
XOR2_X2 inst_31 ( .A(net_21160), .Z(net_737), .B(net_736) );
INV_X4 inst_15136 ( .ZN(net_3517), .A(net_2301) );
CLKBUF_X2 inst_21376 ( .A(net_21247), .Z(net_21248) );
INV_X4 inst_15751 ( .A(net_9401), .ZN(net_1941) );
CLKBUF_X2 inst_22920 ( .A(net_22791), .Z(net_22792) );
NAND2_X2 inst_10937 ( .A2(net_10819), .ZN(net_9291), .A1(net_3229) );
INV_X4 inst_12730 ( .ZN(net_17762), .A(net_17458) );
NOR2_X2 inst_3537 ( .ZN(net_13426), .A2(net_10860), .A1(net_8953) );
NAND2_X2 inst_9787 ( .ZN(net_11099), .A2(net_9746), .A1(net_4931) );
INV_X4 inst_12606 ( .ZN(net_18086), .A(net_18083) );
NOR2_X2 inst_4556 ( .A1(net_20547), .ZN(net_4948), .A2(net_3992) );
INV_X2 inst_19157 ( .ZN(net_3978), .A(net_3934) );
INV_X4 inst_14449 ( .A(net_6594), .ZN(net_6111) );
OAI21_X2 inst_1833 ( .B1(net_19749), .ZN(net_14053), .A(net_11614), .B2(net_8090) );
OAI21_X2 inst_2122 ( .ZN(net_10020), .A(net_9146), .B2(net_7957), .B1(net_5927) );
NAND4_X2 inst_5301 ( .ZN(net_19413), .A4(net_15330), .A2(net_13995), .A1(net_13590), .A3(net_8315) );
NAND2_X2 inst_8160 ( .ZN(net_17980), .A1(net_17979), .A2(net_17978) );
NOR2_X2 inst_3520 ( .ZN(net_13754), .A1(net_13584), .A2(net_7336) );
NAND2_X2 inst_9809 ( .ZN(net_9682), .A1(net_9681), .A2(net_9680) );
NAND2_X2 inst_11601 ( .ZN(net_5364), .A1(net_2660), .A2(net_2116) );
INV_X4 inst_13041 ( .A(net_16562), .ZN(net_16408) );
NOR2_X2 inst_3573 ( .A1(net_20205), .ZN(net_12722), .A2(net_12348) );
INV_X4 inst_17739 ( .A(net_20860), .ZN(net_391) );
XNOR2_X2 inst_623 ( .B(net_17404), .ZN(net_468), .A(net_467) );
NAND2_X2 inst_11306 ( .A1(net_10737), .ZN(net_9717), .A2(net_3787) );
INV_X4 inst_13453 ( .A(net_12099), .ZN(net_11493) );
INV_X4 inst_15612 ( .ZN(net_2864), .A(net_1653) );
AND3_X4 inst_21120 ( .ZN(net_12869), .A2(net_12488), .A3(net_11580), .A1(net_6370) );
NAND2_X2 inst_8557 ( .A1(net_21197), .A2(net_20501), .ZN(net_16752) );
OAI21_X2 inst_1621 ( .A(net_16385), .ZN(net_16072), .B1(net_15494), .B2(net_15436) );
NAND2_X2 inst_10373 ( .ZN(net_12511), .A1(net_7394), .A2(net_7393) );
INV_X2 inst_18881 ( .ZN(net_6188), .A(net_6187) );
INV_X4 inst_14877 ( .ZN(net_6366), .A(net_2653) );
NOR2_X4 inst_3226 ( .ZN(net_5563), .A2(net_2979), .A1(net_252) );
NAND2_X2 inst_8435 ( .A1(net_21142), .ZN(net_17148), .A2(net_16977) );
NAND2_X2 inst_10674 ( .ZN(net_9053), .A1(net_6221), .A2(net_3408) );
NAND2_X2 inst_9609 ( .ZN(net_19182), .A1(net_9617), .A2(net_8453) );
INV_X4 inst_13224 ( .A(net_14302), .ZN(net_13603) );
INV_X2 inst_19338 ( .ZN(net_2464), .A(net_2463) );
INV_X4 inst_15523 ( .A(net_3219), .ZN(net_2398) );
NOR2_X4 inst_3125 ( .ZN(net_6670), .A2(net_3963), .A1(net_3035) );
NAND2_X2 inst_10571 ( .A2(net_7256), .ZN(net_6699), .A1(net_6698) );
INV_X4 inst_14130 ( .ZN(net_7522), .A(net_6110) );
INV_X4 inst_16494 ( .ZN(net_2089), .A(net_1196) );
INV_X2 inst_18998 ( .ZN(net_5065), .A(net_5064) );
INV_X4 inst_16546 ( .A(net_9254), .ZN(net_4694) );
SDFF_X2 inst_760 ( .Q(net_20960), .SE(net_18577), .SI(net_18523), .D(net_566), .CK(net_22452) );
NAND2_X2 inst_10562 ( .ZN(net_6715), .A2(net_4935), .A1(net_3079) );
NAND2_X2 inst_10750 ( .A2(net_11530), .A1(net_6643), .ZN(net_5703) );
AOI21_X2 inst_20432 ( .ZN(net_15172), .B1(net_14678), .B2(net_13896), .A(net_10140) );
AOI21_X2 inst_20582 ( .ZN(net_14056), .A(net_14055), .B2(net_10302), .B1(net_1877) );
NAND2_X2 inst_10814 ( .A2(net_5573), .ZN(net_5518), .A1(net_5517) );
INV_X4 inst_12842 ( .ZN(net_17357), .A(net_17231) );
NAND2_X2 inst_8867 ( .ZN(net_15321), .A2(net_14380), .A1(net_12276) );
INV_X2 inst_18799 ( .ZN(net_7421), .A(net_7420) );
CLKBUF_X2 inst_21793 ( .A(net_21664), .Z(net_21665) );
AND2_X2 inst_21315 ( .A1(net_13996), .ZN(net_7200), .A2(net_5253) );
OAI21_X2 inst_1696 ( .ZN(net_15354), .A(net_15353), .B2(net_13681), .B1(net_11531) );
INV_X4 inst_15863 ( .ZN(net_1806), .A(net_1805) );
INV_X4 inst_16591 ( .ZN(net_1472), .A(net_1144) );
INV_X4 inst_14519 ( .ZN(net_4788), .A(net_4787) );
NAND2_X2 inst_9347 ( .ZN(net_12200), .A1(net_10702), .A2(net_9939) );
INV_X4 inst_17171 ( .ZN(net_735), .A(net_112) );
INV_X4 inst_17203 ( .ZN(net_3151), .A(net_955) );
NOR2_X2 inst_3727 ( .ZN(net_12662), .A2(net_7498), .A1(net_761) );
NAND2_X2 inst_9831 ( .ZN(net_9612), .A1(net_9611), .A2(net_5860) );
NAND2_X2 inst_10812 ( .ZN(net_7227), .A1(net_5754), .A2(net_5525) );
INV_X8 inst_12237 ( .ZN(net_10141), .A(net_7219) );
INV_X4 inst_17189 ( .ZN(net_1821), .A(net_193) );
NAND2_X4 inst_7258 ( .ZN(net_11948), .A2(net_7917), .A1(net_7258) );
CLKBUF_X2 inst_21605 ( .A(net_21320), .Z(net_21477) );
NOR2_X2 inst_3989 ( .ZN(net_9755), .A2(net_6394), .A1(net_6156) );
NAND2_X2 inst_10000 ( .A1(net_13274), .ZN(net_12028), .A2(net_6916) );
INV_X4 inst_14973 ( .ZN(net_4450), .A(net_3422) );
INV_X4 inst_12934 ( .ZN(net_17820), .A(net_16641) );
NOR2_X2 inst_3569 ( .ZN(net_12735), .A1(net_12734), .A2(net_11044) );
NAND2_X4 inst_7268 ( .ZN(net_9751), .A1(net_4918), .A2(net_3572) );
NOR2_X2 inst_3411 ( .ZN(net_15654), .A2(net_15328), .A1(net_14713) );
NAND2_X2 inst_10436 ( .ZN(net_7199), .A1(net_7198), .A2(net_5251) );
OAI211_X2 inst_2524 ( .A(net_12958), .C1(net_12006), .ZN(net_11793), .B(net_11792), .C2(net_4219) );
INV_X2 inst_19486 ( .ZN(net_19259), .A(net_1301) );
OAI21_X4 inst_1446 ( .B2(net_20106), .B1(net_20105), .ZN(net_15745), .A(net_15366) );
NAND2_X2 inst_9486 ( .ZN(net_13761), .A1(net_12551), .A2(net_10899) );
OAI211_X2 inst_2421 ( .ZN(net_15317), .C1(net_14458), .A(net_14419), .C2(net_10861), .B(net_10172) );
XNOR2_X2 inst_390 ( .ZN(net_16771), .A(net_16764), .B(net_14917) );
INV_X4 inst_16866 ( .ZN(net_19616), .A(net_1030) );
INV_X4 inst_17754 ( .ZN(net_5516), .A(net_271) );
OR3_X2 inst_1062 ( .ZN(net_3167), .A1(net_2047), .A2(net_824), .A3(net_85) );
NAND2_X2 inst_8181 ( .A2(net_20705), .A1(net_20704), .ZN(net_17931) );
INV_X4 inst_14455 ( .ZN(net_6105), .A(net_4953) );
INV_X4 inst_16669 ( .A(net_15463), .ZN(net_1077) );
NAND2_X2 inst_7996 ( .ZN(net_18317), .A2(net_18271), .A1(net_17433) );
INV_X4 inst_13757 ( .ZN(net_11535), .A(net_10610) );
AOI21_X2 inst_20920 ( .A(net_10550), .ZN(net_7245), .B2(net_5413), .B1(net_3716) );
CLKBUF_X2 inst_21402 ( .A(net_21250), .Z(net_21274) );
INV_X4 inst_12814 ( .ZN(net_17463), .A(net_17344) );
CLKBUF_X2 inst_21528 ( .A(net_21399), .Z(net_21400) );
INV_X4 inst_14361 ( .ZN(net_5227), .A(net_5226) );
INV_X4 inst_16745 ( .ZN(net_15039), .A(net_1052) );
NAND2_X2 inst_10277 ( .ZN(net_7956), .A1(net_7439), .A2(net_6101) );
AOI21_X2 inst_20511 ( .ZN(net_14618), .B1(net_14617), .A(net_12653), .B2(net_12032) );
INV_X4 inst_15944 ( .ZN(net_2753), .A(net_1715) );
CLKBUF_X2 inst_22111 ( .A(net_21982), .Z(net_21983) );
CLKBUF_X2 inst_21651 ( .A(net_21434), .Z(net_21523) );
INV_X8 inst_12440 ( .A(net_20488), .ZN(net_20487) );
NAND2_X4 inst_7063 ( .A2(net_20310), .A1(net_20309), .ZN(net_20003) );
NOR3_X2 inst_2642 ( .ZN(net_15901), .A3(net_15407), .A1(net_14132), .A2(net_10698) );
INV_X4 inst_12539 ( .ZN(net_18356), .A(net_18355) );
INV_X4 inst_15974 ( .ZN(net_9387), .A(net_1233) );
INV_X2 inst_18817 ( .ZN(net_7119), .A(net_7118) );
INV_X4 inst_18317 ( .A(net_20523), .ZN(net_20521) );
INV_X2 inst_18995 ( .ZN(net_5075), .A(net_5074) );
INV_X4 inst_14394 ( .ZN(net_5126), .A(net_5125) );
XNOR2_X2 inst_123 ( .ZN(net_18341), .B(net_18278), .A(net_17862) );
NAND4_X4 inst_5250 ( .ZN(net_19247), .A3(net_11285), .A1(net_10922), .A2(net_8511), .A4(net_7506) );
OAI21_X2 inst_2160 ( .ZN(net_9248), .B1(net_9247), .A(net_6965), .B2(net_4628) );
NAND4_X4 inst_5181 ( .A2(net_19603), .A1(net_19602), .A4(net_19073), .ZN(net_17487), .A3(net_16346) );
AOI221_X2 inst_20094 ( .ZN(net_9032), .C2(net_9031), .B1(net_8664), .C1(net_7667), .B2(net_5932), .A(net_2756) );
NAND2_X2 inst_10981 ( .ZN(net_9981), .A2(net_3480), .A1(net_3356) );
OAI21_X2 inst_2298 ( .B1(net_7679), .ZN(net_6431), .A(net_6430), .B2(net_6429) );
INV_X4 inst_14355 ( .ZN(net_8235), .A(net_5268) );
INV_X4 inst_14546 ( .A(net_5899), .ZN(net_4614) );
XNOR2_X2 inst_167 ( .B(net_21121), .ZN(net_17830), .A(net_17827) );
NAND2_X2 inst_11660 ( .ZN(net_10635), .A1(net_2627), .A2(net_2260) );
NAND2_X2 inst_11354 ( .ZN(net_3631), .A2(net_3630), .A1(net_3449) );
INV_X4 inst_13138 ( .ZN(net_15129), .A(net_14744) );
CLKBUF_X2 inst_22031 ( .A(net_21507), .Z(net_21903) );
NOR2_X2 inst_4913 ( .ZN(net_3538), .A1(net_1922), .A2(net_1780) );
NAND2_X2 inst_8524 ( .ZN(net_16904), .A2(net_16535), .A1(net_16510) );
OAI211_X2 inst_2475 ( .ZN(net_20080), .C1(net_19968), .B(net_11457), .A(net_11073), .C2(net_2355) );
NOR2_X2 inst_4874 ( .A1(net_20859), .ZN(net_4164), .A2(net_1227) );
INV_X2 inst_19574 ( .ZN(net_878), .A(net_699) );
CLKBUF_X2 inst_21810 ( .A(net_21461), .Z(net_21682) );
INV_X2 inst_19607 ( .A(net_21235), .ZN(net_54) );
NAND3_X1 inst_6824 ( .A2(net_13855), .A3(net_10247), .ZN(net_9052), .A1(net_8244) );
INV_X4 inst_13033 ( .A(net_16721), .ZN(net_16413) );
CLKBUF_X2 inst_22696 ( .A(net_22567), .Z(net_22568) );
INV_X4 inst_17848 ( .A(net_896), .ZN(net_321) );
NAND2_X2 inst_9195 ( .ZN(net_13096), .A1(net_13095), .A2(net_11246) );
INV_X4 inst_13131 ( .ZN(net_15268), .A(net_14879) );
XNOR2_X2 inst_331 ( .ZN(net_17001), .A(net_17000), .B(net_12265) );
NAND2_X2 inst_10691 ( .ZN(net_6087), .A1(net_5714), .A2(net_4596) );
INV_X4 inst_13312 ( .ZN(net_19744), .A(net_10327) );
NAND2_X2 inst_8948 ( .ZN(net_14727), .A2(net_13239), .A1(net_10683) );
INV_X4 inst_14317 ( .ZN(net_9020), .A(net_7351) );
NAND2_X2 inst_11227 ( .A1(net_20923), .ZN(net_8546), .A2(net_7147) );
OAI21_X2 inst_2353 ( .ZN(net_3283), .A(net_3282), .B2(net_3281), .B1(net_1567) );
DFF_X1 inst_19796 ( .D(net_18246), .CK(net_22826), .Q(x1146) );
NAND2_X2 inst_11921 ( .ZN(net_1520), .A1(net_1519), .A2(net_1518) );
AOI21_X4 inst_20226 ( .B1(net_20654), .ZN(net_13721), .B2(net_9768), .A(net_4080) );
INV_X4 inst_17552 ( .ZN(net_4810), .A(net_547) );
INV_X2 inst_19340 ( .ZN(net_12925), .A(net_2452) );
INV_X4 inst_13483 ( .ZN(net_9546), .A(net_9545) );
CLKBUF_X2 inst_22399 ( .A(net_22270), .Z(net_22271) );
NOR3_X2 inst_2762 ( .A3(net_13654), .ZN(net_10474), .A1(net_8257), .A2(net_6751) );
CLKBUF_X2 inst_21985 ( .A(net_21856), .Z(net_21857) );
CLKBUF_X2 inst_22757 ( .A(net_22628), .Z(net_22629) );
SDFF_X2 inst_997 ( .QN(net_21066), .D(net_424), .SE(net_263), .CK(net_21723), .SI(x1975) );
SDFF_X2 inst_857 ( .Q(net_21125), .D(net_17150), .SE(net_263), .CK(net_21252), .SI(x4215) );
INV_X4 inst_16235 ( .A(net_2070), .ZN(net_2047) );
NOR2_X2 inst_4824 ( .A1(net_5217), .ZN(net_2989), .A2(net_2422) );
NAND3_X2 inst_6403 ( .ZN(net_11976), .A1(net_8494), .A2(net_7964), .A3(net_6654) );
CLKBUF_X2 inst_21990 ( .A(net_21798), .Z(net_21862) );
NOR2_X2 inst_4179 ( .A1(net_8226), .ZN(net_8105), .A2(net_6799) );
INV_X4 inst_12721 ( .ZN(net_17533), .A(net_17532) );
AOI21_X4 inst_20154 ( .B2(net_19132), .B1(net_19131), .ZN(net_15756), .A(net_14195) );
NAND3_X2 inst_5951 ( .ZN(net_14883), .A2(net_14541), .A1(net_13573), .A3(net_13369) );
NOR2_X2 inst_4006 ( .ZN(net_9603), .A1(net_8097), .A2(net_8096) );
NAND2_X2 inst_7988 ( .A2(net_18328), .ZN(net_18327), .A1(net_17911) );
INV_X4 inst_15918 ( .ZN(net_2727), .A(net_1249) );
CLKBUF_X2 inst_21552 ( .A(net_21423), .Z(net_21424) );
INV_X2 inst_18532 ( .A(net_11501), .ZN(net_11080) );
NOR2_X4 inst_3203 ( .ZN(net_5353), .A2(net_3182), .A1(net_3047) );
INV_X4 inst_15368 ( .ZN(net_10816), .A(net_2574) );
AOI21_X2 inst_20942 ( .A(net_9926), .ZN(net_6409), .B1(net_5775), .B2(net_2816) );
INV_X2 inst_19651 ( .ZN(net_20069), .A(net_20068) );
NOR2_X2 inst_5073 ( .ZN(net_10052), .A1(net_115), .A2(net_67) );
CLKBUF_X2 inst_22830 ( .A(net_22701), .Z(net_22702) );
INV_X4 inst_13951 ( .ZN(net_8635), .A(net_7203) );
OAI22_X2 inst_1310 ( .B1(net_10490), .A1(net_9581), .ZN(net_8955), .B2(net_8954), .A2(net_6595) );
INV_X2 inst_19246 ( .A(net_14279), .ZN(net_3266) );
NOR2_X4 inst_3280 ( .ZN(net_2243), .A1(net_1645), .A2(net_1178) );
NOR2_X2 inst_4491 ( .A1(net_9064), .ZN(net_5496), .A2(net_4694) );
INV_X2 inst_19281 ( .ZN(net_5198), .A(net_2935) );
NAND2_X4 inst_7397 ( .A2(net_19026), .ZN(net_6807), .A1(net_3255) );
NOR2_X4 inst_2823 ( .ZN(net_20368), .A2(net_16065), .A1(net_16033) );
NAND2_X2 inst_11594 ( .ZN(net_2679), .A1(net_1629), .A2(net_1331) );
INV_X4 inst_13981 ( .ZN(net_10506), .A(net_5388) );
INV_X4 inst_13413 ( .ZN(net_17144), .A(net_12872) );
INV_X4 inst_15171 ( .ZN(net_5343), .A(net_4249) );
INV_X4 inst_16711 ( .ZN(net_4025), .A(net_1262) );
INV_X4 inst_14464 ( .ZN(net_4927), .A(net_4926) );
XNOR2_X2 inst_136 ( .B(net_21194), .ZN(net_18223), .A(net_18162) );
NAND3_X2 inst_5839 ( .ZN(net_19592), .A3(net_14604), .A2(net_8650), .A1(net_8172) );
NAND2_X2 inst_11733 ( .ZN(net_2196), .A2(net_1833), .A1(net_819) );
CLKBUF_X2 inst_22207 ( .A(net_22078), .Z(net_22079) );
INV_X4 inst_13837 ( .ZN(net_9161), .A(net_7486) );
OAI21_X2 inst_1526 ( .A(net_18582), .ZN(net_18032), .B2(net_17981), .B1(net_17957) );
OAI211_X2 inst_2547 ( .ZN(net_10822), .B(net_9309), .C2(net_4636), .A(net_4456), .C1(net_3165) );
NOR2_X2 inst_4637 ( .ZN(net_3485), .A2(net_3484), .A1(net_3481) );
CLKBUF_X2 inst_22332 ( .A(net_22203), .Z(net_22204) );
INV_X4 inst_16800 ( .ZN(net_10415), .A(net_7230) );
SDFF_X2 inst_1047 ( .QN(net_20980), .D(net_1860), .SE(net_263), .CK(net_22648), .SI(x3322) );
INV_X4 inst_15790 ( .A(net_15659), .ZN(net_1902) );
NAND2_X4 inst_6860 ( .A2(net_20719), .A1(net_20718), .ZN(net_18384) );
NAND2_X2 inst_8507 ( .A2(net_20500), .ZN(net_16924), .A1(net_9235) );
AND2_X4 inst_21163 ( .ZN(net_19936), .A1(net_15602), .A2(net_13586) );
NAND2_X2 inst_11768 ( .ZN(net_7094), .A2(net_2073), .A1(net_184) );
NOR2_X2 inst_3700 ( .ZN(net_11115), .A1(net_11114), .A2(net_11113) );
NAND3_X2 inst_6744 ( .ZN(net_6393), .A2(net_6392), .A3(net_6391), .A1(net_3746) );
INV_X8 inst_12432 ( .ZN(net_19459), .A(net_16541) );
INV_X4 inst_15519 ( .A(net_9018), .ZN(net_6083) );
INV_X4 inst_16955 ( .ZN(net_1187), .A(net_120) );
OAI21_X2 inst_1858 ( .ZN(net_13816), .A(net_11404), .B2(net_11110), .B1(net_9124) );
INV_X4 inst_17120 ( .A(net_2179), .ZN(net_1200) );
NOR2_X2 inst_3846 ( .ZN(net_9582), .A1(net_9581), .A2(net_7623) );
INV_X4 inst_13668 ( .ZN(net_9125), .A(net_8061) );
OAI221_X2 inst_1334 ( .ZN(net_15376), .B1(net_15375), .C1(net_15374), .A(net_13839), .C2(net_13339), .B2(net_11855) );
AOI21_X2 inst_20426 ( .ZN(net_15208), .B1(net_14600), .B2(net_14113), .A(net_10673) );
AOI21_X2 inst_20547 ( .ZN(net_14390), .B2(net_12519), .B1(net_9365), .A(net_8028) );
INV_X4 inst_17491 ( .ZN(net_6648), .A(net_522) );
CLKBUF_X2 inst_22536 ( .A(net_22407), .Z(net_22408) );
NAND3_X2 inst_5944 ( .ZN(net_20156), .A1(net_13712), .A2(net_5722), .A3(net_588) );
NAND4_X2 inst_5383 ( .ZN(net_20386), .A2(net_12984), .A4(net_10060), .A3(net_9657), .A1(net_9519) );
NAND3_X2 inst_6129 ( .ZN(net_13741), .A3(net_10942), .A2(net_8238), .A1(net_4351) );
INV_X4 inst_14735 ( .ZN(net_5186), .A(net_4154) );
CLKBUF_X2 inst_21533 ( .A(net_21404), .Z(net_21405) );
AOI21_X2 inst_20541 ( .ZN(net_14423), .B2(net_11462), .A(net_8821), .B1(net_909) );
NAND2_X4 inst_7273 ( .ZN(net_9658), .A1(net_6041), .A2(net_6040) );
NAND2_X1 inst_12130 ( .ZN(net_18284), .A2(net_18283), .A1(net_18138) );
CLKBUF_X2 inst_21716 ( .A(net_21587), .Z(net_21588) );
INV_X4 inst_15567 ( .ZN(net_2804), .A(net_2289) );
NAND2_X2 inst_11453 ( .ZN(net_4424), .A1(net_3915), .A2(net_3292) );
XNOR2_X2 inst_265 ( .ZN(net_17255), .A(net_17254), .B(net_17253) );
OAI21_X2 inst_2055 ( .ZN(net_10839), .A(net_10838), .B2(net_10837), .B1(net_2311) );
NAND2_X2 inst_11702 ( .ZN(net_2774), .A1(net_1472), .A2(net_1216) );
NAND2_X2 inst_7783 ( .ZN(net_18726), .A2(net_18673), .A1(net_16653) );
NAND3_X4 inst_5554 ( .ZN(net_16219), .A3(net_15920), .A2(net_14852), .A1(net_12210) );
CLKBUF_X2 inst_21375 ( .A(x7698), .Z(net_21247) );
AOI21_X2 inst_20642 ( .ZN(net_13229), .B1(net_12105), .B2(net_8970), .A(net_253) );
INV_X2 inst_18667 ( .A(net_11826), .ZN(net_9172) );
NOR2_X4 inst_3262 ( .A1(net_2585), .ZN(net_2151), .A2(net_1499) );
AOI21_X2 inst_20283 ( .B1(net_20904), .ZN(net_20027), .B2(net_15944), .A(net_12123) );
INV_X4 inst_17932 ( .A(net_20983), .ZN(net_1855) );
NOR2_X2 inst_4566 ( .ZN(net_4881), .A2(net_3884), .A1(net_60) );
INV_X4 inst_12993 ( .ZN(net_16789), .A(net_16489) );
NAND2_X2 inst_10653 ( .ZN(net_11910), .A2(net_6317), .A1(net_5149) );
NAND3_X2 inst_6301 ( .ZN(net_12808), .A2(net_12807), .A1(net_10918), .A3(net_10280) );
CLKBUF_X2 inst_22159 ( .A(net_21537), .Z(net_22031) );
INV_X2 inst_19510 ( .A(net_13206), .ZN(net_2454) );
NAND2_X4 inst_7249 ( .ZN(net_12286), .A1(net_6797), .A2(net_5066) );
NAND2_X2 inst_7975 ( .ZN(net_18349), .A2(net_18285), .A1(net_17329) );
NOR2_X2 inst_3954 ( .ZN(net_8601), .A2(net_7098), .A1(net_5916) );
INV_X4 inst_12956 ( .A(net_16727), .ZN(net_16538) );
NAND2_X2 inst_9367 ( .ZN(net_12121), .A2(net_12120), .A1(net_9423) );
XNOR2_X2 inst_222 ( .ZN(net_17508), .A(net_17502), .B(net_16334) );
INV_X2 inst_18857 ( .ZN(net_9188), .A(net_7459) );
NAND3_X2 inst_6372 ( .ZN(net_12060), .A1(net_10452), .A2(net_8833), .A3(net_8371) );
NAND3_X2 inst_6073 ( .ZN(net_14115), .A3(net_10487), .A2(net_8792), .A1(net_8331) );
CLKBUF_X2 inst_21999 ( .A(net_21870), .Z(net_21871) );
INV_X4 inst_13166 ( .ZN(net_14805), .A(net_14212) );
INV_X8 inst_12218 ( .A(net_10144), .ZN(net_8588) );
NAND3_X2 inst_6728 ( .ZN(net_6490), .A2(net_6489), .A3(net_6488), .A1(net_2970) );
CLKBUF_X2 inst_22382 ( .A(net_22253), .Z(net_22254) );
OAI22_X2 inst_1302 ( .ZN(net_10522), .B1(net_10521), .B2(net_10520), .A1(net_8682), .A2(net_6540) );
INV_X4 inst_18220 ( .A(net_20991), .ZN(net_2458) );
NAND2_X2 inst_10609 ( .ZN(net_7868), .A1(net_6611), .A2(net_4852) );
OAI21_X2 inst_1648 ( .B2(net_19977), .B1(net_19976), .A(net_16385), .ZN(net_15906) );
OR2_X4 inst_1079 ( .ZN(net_12088), .A2(net_7665), .A1(net_6325) );
NAND3_X2 inst_5847 ( .ZN(net_15435), .A1(net_14997), .A2(net_14544), .A3(net_12109) );
INV_X4 inst_13958 ( .ZN(net_10625), .A(net_6749) );
INV_X4 inst_13833 ( .A(net_9321), .ZN(net_9165) );
INV_X2 inst_19144 ( .ZN(net_4101), .A(net_4100) );
INV_X4 inst_16857 ( .ZN(net_1501), .A(net_967) );
NOR2_X2 inst_3925 ( .ZN(net_10232), .A1(net_9917), .A2(net_8937) );
INV_X2 inst_18918 ( .ZN(net_5949), .A(net_5948) );
NOR3_X4 inst_2606 ( .ZN(net_19930), .A1(net_15999), .A3(net_14456), .A2(net_7516) );
NOR2_X2 inst_4314 ( .A1(net_8341), .ZN(net_7418), .A2(net_5894) );
NAND2_X2 inst_9837 ( .ZN(net_10981), .A1(net_9350), .A2(net_7521) );
OAI211_X2 inst_2523 ( .C1(net_13070), .ZN(net_11809), .A(net_11808), .B(net_11807), .C2(net_5926) );
XNOR2_X2 inst_506 ( .B(net_21184), .ZN(net_7741), .A(net_7740) );
NAND2_X2 inst_10662 ( .ZN(net_11853), .A1(net_6295), .A2(net_3147) );
INV_X4 inst_13569 ( .A(net_9134), .ZN(net_9133) );
INV_X4 inst_17834 ( .ZN(net_14022), .A(net_126) );
NAND2_X2 inst_11782 ( .A2(net_7676), .ZN(net_5297), .A1(net_1599) );
NAND2_X2 inst_8572 ( .ZN(net_16735), .A2(net_16734), .A1(net_16444) );
NAND2_X2 inst_10835 ( .ZN(net_10373), .A1(net_9148), .A2(net_4055) );
OAI22_X1 inst_1323 ( .A2(net_17815), .B2(net_17752), .ZN(net_16981), .A1(net_5786), .B1(net_3520) );
OR2_X4 inst_1085 ( .ZN(net_11224), .A2(net_3341), .A1(net_90) );
INV_X4 inst_14048 ( .A(net_11315), .ZN(net_6254) );
CLKBUF_X2 inst_21969 ( .A(net_21272), .Z(net_21841) );
INV_X2 inst_19656 ( .A(net_20220), .ZN(net_20219) );
INV_X4 inst_18177 ( .A(net_21220), .ZN(net_16404) );
NAND2_X2 inst_8791 ( .ZN(net_20843), .A2(net_15399), .A1(net_10683) );
NAND2_X2 inst_10464 ( .ZN(net_8363), .A1(net_7007), .A2(net_7006) );
CLKBUF_X2 inst_22393 ( .A(net_22264), .Z(net_22265) );
NOR3_X2 inst_2655 ( .ZN(net_15431), .A3(net_14313), .A1(net_11401), .A2(net_8666) );
CLKBUF_X2 inst_21698 ( .A(net_21569), .Z(net_21570) );
OAI21_X2 inst_1720 ( .ZN(net_15150), .B1(net_15064), .B2(net_13262), .A(net_13182) );
XNOR2_X2 inst_160 ( .ZN(net_17942), .A(net_17824), .B(net_17570) );
INV_X2 inst_19522 ( .A(net_1543), .ZN(net_1106) );
NAND2_X2 inst_8889 ( .ZN(net_15133), .A2(net_14163), .A1(net_14063) );
INV_X4 inst_14420 ( .ZN(net_5053), .A(net_5052) );
NAND2_X2 inst_9243 ( .A2(net_12694), .ZN(net_12683), .A1(net_4716) );
INV_X2 inst_18494 ( .ZN(net_13564), .A(net_12314) );
XNOR2_X2 inst_370 ( .B(net_21200), .A(net_20075), .ZN(net_16845) );
NAND2_X4 inst_7450 ( .ZN(net_14334), .A1(net_3224), .A2(net_2274) );
NAND2_X2 inst_7825 ( .ZN(net_18644), .A1(net_18624), .A2(net_18618) );
NAND2_X2 inst_10414 ( .A2(net_7337), .ZN(net_7249), .A1(net_7248) );
OAI22_X2 inst_1265 ( .A2(net_17487), .B2(net_17371), .ZN(net_17131), .A1(net_6459), .B1(net_5761) );
INV_X4 inst_14480 ( .ZN(net_11057), .A(net_11041) );
NAND2_X2 inst_10669 ( .ZN(net_6238), .A1(net_6237), .A2(net_5894) );
NAND2_X2 inst_8371 ( .ZN(net_17368), .A1(net_17366), .A2(net_17365) );
AOI22_X2 inst_19999 ( .ZN(net_14140), .A2(net_10770), .A1(net_9438), .B2(net_9188), .B1(net_5479) );
NAND2_X2 inst_8176 ( .ZN(net_17939), .A1(net_17938), .A2(net_17854) );
NAND2_X2 inst_11288 ( .A2(net_3933), .ZN(net_3835), .A1(net_573) );
OAI22_X2 inst_1321 ( .A1(net_6201), .B2(net_5265), .ZN(net_2944), .B1(net_2862), .A2(net_1294) );
SDFF_X2 inst_1012 ( .QN(net_20985), .SE(net_17277), .D(net_2030), .CK(net_22654), .SI(x3242) );
NAND4_X2 inst_5255 ( .ZN(net_16496), .A1(net_16367), .A2(net_16298), .A4(net_13898), .A3(net_9408) );
INV_X4 inst_12768 ( .ZN(net_17675), .A(net_17337) );
INV_X4 inst_16082 ( .ZN(net_3804), .A(net_1538) );
NAND2_X2 inst_8341 ( .A1(net_20071), .ZN(net_17491), .A2(net_17490) );
NOR2_X2 inst_3492 ( .ZN(net_14229), .A1(net_12637), .A2(net_7273) );
INV_X2 inst_18542 ( .ZN(net_10992), .A(net_10991) );
INV_X4 inst_14032 ( .ZN(net_10414), .A(net_8325) );
INV_X4 inst_14724 ( .ZN(net_19575), .A(net_4145) );
INV_X2 inst_19594 ( .A(net_314), .ZN(net_210) );
NAND2_X2 inst_9015 ( .ZN(net_14256), .A2(net_12670), .A1(net_8730) );
NOR2_X4 inst_3149 ( .A2(net_20578), .ZN(net_6841), .A1(net_2744) );
INV_X4 inst_17644 ( .A(net_955), .ZN(net_628) );
NOR2_X2 inst_4034 ( .A2(net_13320), .ZN(net_10150), .A1(net_1233) );
AOI21_X2 inst_20894 ( .ZN(net_7784), .B2(net_4652), .A(net_4166), .B1(net_308) );
XNOR2_X2 inst_377 ( .B(net_21168), .A(net_16848), .ZN(net_16835) );
INV_X4 inst_13570 ( .ZN(net_12497), .A(net_9129) );
NAND2_X4 inst_6993 ( .ZN(net_20585), .A1(net_16740), .A2(net_16595) );
NAND2_X2 inst_10157 ( .A1(net_10000), .ZN(net_8263), .A2(net_6305) );
NOR2_X2 inst_3946 ( .ZN(net_14412), .A1(net_12620), .A2(net_8713) );
NOR2_X2 inst_4760 ( .ZN(net_5625), .A1(net_2994), .A2(net_2993) );
INV_X4 inst_15703 ( .ZN(net_4326), .A(net_2650) );
NOR2_X2 inst_3920 ( .ZN(net_10282), .A1(net_8796), .A2(net_8795) );
NAND2_X4 inst_6953 ( .ZN(net_18994), .A1(net_18493), .A2(net_16967) );
NAND2_X4 inst_6920 ( .ZN(net_19686), .A1(net_17711), .A2(net_16985) );
NOR2_X4 inst_3018 ( .ZN(net_6276), .A2(net_5459), .A1(net_3636) );
NOR2_X4 inst_3078 ( .ZN(net_6220), .A2(net_5131), .A1(net_1713) );
INV_X4 inst_13750 ( .A(net_9594), .ZN(net_9222) );
NAND3_X2 inst_5792 ( .ZN(net_20202), .A3(net_15008), .A1(net_14177), .A2(net_8899) );
INV_X4 inst_12779 ( .ZN(net_17557), .A(net_17474) );
DFF_X1 inst_19919 ( .D(net_16529), .CK(net_22779), .Q(x1204) );
CLKBUF_X2 inst_21504 ( .A(net_21375), .Z(net_21376) );
NAND2_X2 inst_9731 ( .ZN(net_13852), .A1(net_10113), .A2(net_9404) );
INV_X4 inst_13579 ( .ZN(net_9103), .A(net_9102) );
INV_X2 inst_19442 ( .ZN(net_2470), .A(net_1969) );
INV_X2 inst_18481 ( .ZN(net_12558), .A(net_11354) );
NOR2_X2 inst_5054 ( .ZN(net_2523), .A2(net_1562), .A1(net_1376) );
NAND3_X2 inst_5926 ( .ZN(net_19918), .A1(net_14049), .A3(net_10413), .A2(net_3723) );
INV_X4 inst_16113 ( .A(net_2258), .ZN(net_1494) );
NOR2_X2 inst_4627 ( .ZN(net_3602), .A2(net_3326), .A1(net_2406) );
INV_X4 inst_17018 ( .A(net_3342), .ZN(net_1182) );
INV_X8 inst_12414 ( .A(net_20867), .ZN(net_2585) );
INV_X4 inst_13559 ( .A(net_9158), .ZN(net_9157) );
INV_X4 inst_14429 ( .A(net_13147), .ZN(net_5031) );
INV_X4 inst_16110 ( .ZN(net_1496), .A(net_1216) );
XNOR2_X2 inst_107 ( .ZN(net_18523), .A(net_18458), .B(net_17363) );
INV_X4 inst_14191 ( .ZN(net_11159), .A(net_5504) );
INV_X4 inst_16166 ( .ZN(net_3278), .A(net_1911) );
SDFF_X2 inst_990 ( .QN(net_21023), .D(net_485), .SE(net_263), .CK(net_21892), .SI(x2639) );
INV_X8 inst_12381 ( .A(net_199), .ZN(net_177) );
AOI21_X2 inst_20798 ( .ZN(net_10416), .A(net_10415), .B2(net_10414), .B1(net_3674) );
INV_X4 inst_16807 ( .ZN(net_1753), .A(net_397) );
NAND2_X4 inst_7225 ( .A1(net_19961), .ZN(net_9128), .A2(net_4020) );
NAND2_X2 inst_10412 ( .ZN(net_14537), .A1(net_6911), .A2(net_6844) );
NOR2_X2 inst_4710 ( .ZN(net_6530), .A1(net_4464), .A2(net_3150) );
NOR2_X2 inst_3628 ( .ZN(net_12278), .A1(net_9144), .A2(net_5979) );
AOI22_X2 inst_19981 ( .ZN(net_15391), .B1(net_14634), .A2(net_13967), .A1(net_13023), .B2(net_7381) );
INV_X4 inst_15632 ( .A(net_2491), .ZN(net_2142) );
OAI21_X1 inst_2366 ( .ZN(net_19833), .A(net_8338), .B2(net_4942), .B1(net_3071) );
NAND2_X2 inst_10093 ( .A2(net_8651), .ZN(net_8619), .A1(net_8618) );
INV_X4 inst_14886 ( .ZN(net_3668), .A(net_3667) );
NOR2_X2 inst_5049 ( .ZN(net_2343), .A1(net_1376), .A2(net_1155) );
NAND2_X2 inst_11343 ( .ZN(net_3674), .A2(net_3673), .A1(net_2917) );
INV_X4 inst_14155 ( .ZN(net_7482), .A(net_6024) );
CLKBUF_X2 inst_22745 ( .A(net_22616), .Z(net_22617) );
INV_X4 inst_13998 ( .ZN(net_6383), .A(net_5247) );
NOR2_X2 inst_4605 ( .A2(net_20468), .ZN(net_6410), .A1(net_3748) );
NAND2_X2 inst_10351 ( .ZN(net_7491), .A2(net_7443), .A1(net_6884) );
NAND2_X2 inst_11207 ( .ZN(net_4727), .A2(net_4035), .A1(net_154) );
OR2_X2 inst_1237 ( .ZN(net_8568), .A1(net_235), .A2(net_130) );
AOI21_X2 inst_20564 ( .B1(net_14515), .ZN(net_14248), .A(net_13516), .B2(net_6630) );
INV_X4 inst_12873 ( .ZN(net_17146), .A(net_17007) );
INV_X4 inst_15196 ( .ZN(net_11893), .A(net_10664) );
NAND2_X4 inst_7175 ( .ZN(net_11552), .A1(net_9392), .A2(net_732) );
INV_X2 inst_19413 ( .A(net_2827), .ZN(net_1939) );
NOR2_X4 inst_3310 ( .ZN(net_1748), .A1(net_1101), .A2(net_1080) );
NOR2_X4 inst_3062 ( .ZN(net_6778), .A1(net_5042), .A2(net_4945) );
NAND3_X2 inst_6267 ( .ZN(net_12963), .A2(net_12962), .A3(net_6772), .A1(net_5385) );
AOI21_X4 inst_20188 ( .ZN(net_15213), .A(net_14300), .B2(net_13455), .B1(net_1030) );
INV_X4 inst_14249 ( .A(net_10709), .ZN(net_5760) );
INV_X4 inst_13459 ( .ZN(net_11499), .A(net_9721) );
NOR2_X2 inst_5100 ( .ZN(net_1518), .A2(net_167), .A1(net_86) );
NAND2_X2 inst_8536 ( .A1(net_19434), .ZN(net_16856), .A2(net_16724) );
AND4_X4 inst_21085 ( .ZN(net_16769), .A4(net_16324), .A2(net_16106), .A1(net_15741), .A3(net_15236) );
INV_X4 inst_15239 ( .ZN(net_6265), .A(net_2825) );
AND2_X2 inst_21357 ( .ZN(net_4413), .A2(net_1623), .A1(net_703) );
INV_X4 inst_13967 ( .ZN(net_6704), .A(net_6703) );
INV_X4 inst_14745 ( .ZN(net_6545), .A(net_5593) );
NAND3_X2 inst_6013 ( .ZN(net_14409), .A1(net_14209), .A3(net_11592), .A2(net_7620) );
XNOR2_X2 inst_383 ( .B(net_21164), .ZN(net_17470), .A(net_16801) );
INV_X4 inst_15017 ( .ZN(net_14085), .A(net_13651) );
AOI21_X2 inst_20890 ( .B1(net_10091), .ZN(net_7788), .B2(net_7787), .A(net_6351) );
NAND2_X2 inst_11793 ( .ZN(net_20697), .A1(net_5009), .A2(net_2489) );
INV_X4 inst_13561 ( .A(net_11251), .ZN(net_9154) );
NOR2_X2 inst_4132 ( .ZN(net_6957), .A2(net_5123), .A1(net_4100) );
NAND2_X4 inst_7031 ( .ZN(net_16860), .A2(net_16859), .A1(net_16813) );
NAND2_X4 inst_7670 ( .A1(net_20901), .ZN(net_1122), .A2(net_210) );
NAND2_X4 inst_7679 ( .ZN(net_1314), .A2(net_808), .A1(net_807) );
NAND2_X2 inst_9765 ( .ZN(net_9825), .A1(net_9824), .A2(net_4103) );
INV_X2 inst_19588 ( .A(net_792), .ZN(net_324) );
CLKBUF_X2 inst_22356 ( .A(net_22227), .Z(net_22228) );
INV_X4 inst_17908 ( .ZN(net_1861), .A(net_834) );
INV_X2 inst_19115 ( .A(net_15897), .ZN(net_4449) );
INV_X4 inst_16651 ( .A(net_1144), .ZN(net_1093) );
NAND2_X2 inst_11801 ( .ZN(net_20470), .A2(net_2053), .A1(net_286) );
INV_X4 inst_15972 ( .ZN(net_2409), .A(net_1238) );
NAND4_X2 inst_5372 ( .ZN(net_15232), .A4(net_14021), .A3(net_11772), .A2(net_8653), .A1(net_6950) );
CLKBUF_X2 inst_21615 ( .A(net_21486), .Z(net_21487) );
NOR2_X2 inst_3375 ( .ZN(net_16495), .A2(net_16389), .A1(net_16058) );
XNOR2_X2 inst_234 ( .B(net_21117), .A(net_17480), .ZN(net_17407) );
CLKBUF_X2 inst_22593 ( .A(net_22464), .Z(net_22465) );
INV_X4 inst_16428 ( .A(net_9656), .ZN(net_1402) );
AOI21_X2 inst_20461 ( .ZN(net_15021), .B1(net_15020), .A(net_13911), .B2(net_6423) );
NAND4_X2 inst_5293 ( .ZN(net_15930), .A4(net_15185), .A1(net_13359), .A3(net_12111), .A2(net_11600) );
INV_X4 inst_16893 ( .ZN(net_10037), .A(net_3049) );
INV_X8 inst_12398 ( .ZN(net_304), .A(net_94) );
INV_X2 inst_18604 ( .ZN(net_11584), .A(net_9784) );
INV_X4 inst_13975 ( .A(net_6652), .ZN(net_6651) );
NOR2_X2 inst_3429 ( .ZN(net_19900), .A1(net_15102), .A2(net_14603) );
OAI221_X2 inst_1328 ( .B1(net_21220), .ZN(net_16220), .A(net_15819), .B2(net_15721), .C2(net_15675), .C1(net_1947) );
INV_X4 inst_18204 ( .A(net_20960), .ZN(net_16242) );
NAND2_X2 inst_8429 ( .A1(net_20789), .A2(net_20071), .ZN(net_19655) );
INV_X4 inst_15434 ( .ZN(net_12885), .A(net_12884) );
OAI21_X2 inst_1776 ( .A(net_14684), .ZN(net_14680), .B2(net_11940), .B1(net_11685) );
OAI21_X2 inst_2335 ( .ZN(net_4684), .B2(net_4029), .B1(net_3736), .A(net_1612) );
NAND2_X2 inst_7715 ( .ZN(net_18848), .A2(net_18830), .A1(net_18816) );
INV_X4 inst_13157 ( .ZN(net_14870), .A(net_14326) );
CLKBUF_X2 inst_22001 ( .A(net_21872), .Z(net_21873) );
CLKBUF_X2 inst_21811 ( .A(net_21682), .Z(net_21683) );
INV_X2 inst_18699 ( .A(net_8876), .ZN(net_8321) );
XNOR2_X2 inst_598 ( .B(net_16759), .ZN(net_13291), .A(net_675) );
OAI21_X2 inst_1624 ( .ZN(net_16047), .B1(net_16046), .A(net_15630), .B2(net_15477) );
INV_X4 inst_14868 ( .A(net_5386), .ZN(net_3728) );
NAND2_X2 inst_10595 ( .ZN(net_7920), .A1(net_6635), .A2(net_6634) );
CLKBUF_X2 inst_22625 ( .A(net_22496), .Z(net_22497) );
NAND2_X2 inst_10728 ( .ZN(net_5837), .A1(net_5836), .A2(net_5835) );
AOI21_X4 inst_20170 ( .ZN(net_20222), .A(net_15454), .B2(net_14627), .B1(net_14106) );
NOR2_X4 inst_3167 ( .ZN(net_5575), .A1(net_3110), .A2(net_85) );
INV_X4 inst_13501 ( .A(net_11869), .ZN(net_9432) );
INV_X4 inst_14029 ( .ZN(net_6282), .A(net_6281) );
NAND2_X4 inst_7205 ( .A1(net_9801), .ZN(net_9630), .A2(net_5595) );
AOI21_X2 inst_20311 ( .B1(net_19592), .ZN(net_16032), .B2(net_13827), .A(net_9011) );
CLKBUF_X2 inst_22239 ( .A(net_22105), .Z(net_22111) );
XNOR2_X2 inst_325 ( .B(net_21135), .ZN(net_17699), .A(net_17025) );
INV_X4 inst_14861 ( .ZN(net_3774), .A(net_3773) );
NAND3_X2 inst_6502 ( .ZN(net_10833), .A2(net_5322), .A1(net_4657), .A3(net_4562) );
INV_X4 inst_16579 ( .A(net_2948), .ZN(net_1725) );
NAND2_X2 inst_8858 ( .ZN(net_20701), .A1(net_15356), .A2(net_14424) );
NOR2_X2 inst_4769 ( .ZN(net_4282), .A2(net_2970), .A1(net_117) );
CLKBUF_X2 inst_21562 ( .A(net_21433), .Z(net_21434) );
OR2_X2 inst_1197 ( .A1(net_7950), .ZN(net_6823), .A2(net_4010) );
INV_X2 inst_18371 ( .ZN(net_17482), .A(net_17368) );
NAND2_X4 inst_6958 ( .ZN(net_20520), .A2(net_19221), .A1(net_19220) );
NAND2_X2 inst_10544 ( .ZN(net_10480), .A2(net_6781), .A1(net_6648) );
SDFF_X2 inst_955 ( .QN(net_21002), .D(net_2437), .SE(net_253), .CK(net_21848), .SI(x3007) );
INV_X4 inst_15793 ( .ZN(net_2566), .A(net_1899) );
NAND2_X2 inst_11041 ( .ZN(net_10008), .A1(net_9943), .A2(net_4366) );
NAND2_X2 inst_9519 ( .ZN(net_11142), .A1(net_9842), .A2(net_9104) );
INV_X4 inst_18264 ( .A(net_19436), .ZN(net_19435) );
INV_X4 inst_15157 ( .ZN(net_3052), .A(net_3051) );
NAND3_X2 inst_5851 ( .ZN(net_15423), .A3(net_14396), .A2(net_11159), .A1(net_7398) );
INV_X2 inst_18418 ( .ZN(net_15670), .A(net_15470) );
INV_X4 inst_16364 ( .ZN(net_2053), .A(net_1010) );
INV_X2 inst_19627 ( .A(net_21239), .ZN(net_90) );
NAND3_X2 inst_6665 ( .ZN(net_8441), .A3(net_8440), .A2(net_4831), .A1(net_3888) );
INV_X4 inst_12502 ( .A(net_18649), .ZN(net_18648) );
CLKBUF_X2 inst_21622 ( .A(net_21493), .Z(net_21494) );
NAND2_X4 inst_7117 ( .ZN(net_12390), .A1(net_11023), .A2(net_6274) );
NOR2_X4 inst_2842 ( .ZN(net_14592), .A2(net_13267), .A1(net_12139) );
NAND2_X2 inst_11142 ( .A1(net_8700), .ZN(net_4234), .A2(net_3875) );
INV_X4 inst_13663 ( .ZN(net_10190), .A(net_8103) );
CLKBUF_X2 inst_21930 ( .A(net_21613), .Z(net_21802) );
INV_X2 inst_19715 ( .ZN(net_20769), .A(net_20766) );
NOR2_X2 inst_3792 ( .ZN(net_10078), .A2(net_6333), .A1(net_5418) );
OAI21_X2 inst_2084 ( .ZN(net_10457), .B1(net_7822), .B2(net_6623), .A(net_4237) );
NAND3_X2 inst_5711 ( .A3(net_19559), .A1(net_19558), .ZN(net_16185), .A2(net_15913) );
INV_X4 inst_16179 ( .A(net_7865), .ZN(net_5387) );
NAND2_X2 inst_11534 ( .A1(net_10875), .ZN(net_2928), .A2(net_2034) );
INV_X8 inst_12310 ( .ZN(net_1583), .A(net_460) );
INV_X2 inst_18715 ( .ZN(net_10291), .A(net_8795) );
INV_X4 inst_17143 ( .ZN(net_9146), .A(net_5877) );
NAND2_X2 inst_8203 ( .ZN(net_17978), .A2(net_17793), .A1(net_17610) );
INV_X4 inst_16686 ( .ZN(net_11016), .A(net_3760) );
INV_X2 inst_19489 ( .ZN(net_2340), .A(net_1556) );
AOI211_X2 inst_21056 ( .C1(net_14653), .ZN(net_11219), .A(net_11218), .B(net_11217), .C2(net_7122) );
SDFF_X2 inst_803 ( .Q(net_20950), .SE(net_18856), .SI(net_17974), .D(net_379), .CK(net_22614) );
NAND2_X2 inst_12011 ( .ZN(net_1548), .A2(net_1136), .A1(net_639) );
INV_X2 inst_18943 ( .A(net_7283), .ZN(net_5685) );
AOI21_X2 inst_20802 ( .ZN(net_10349), .B2(net_10348), .A(net_10286), .B1(net_2425) );
AOI21_X2 inst_20454 ( .ZN(net_15059), .B1(net_15058), .B2(net_12988), .A(net_7683) );
INV_X4 inst_15167 ( .ZN(net_3665), .A(net_3017) );
INV_X2 inst_19549 ( .ZN(net_2710), .A(net_882) );
NAND2_X2 inst_10312 ( .A1(net_10490), .ZN(net_9380), .A2(net_5392) );
AOI21_X2 inst_20974 ( .ZN(net_4658), .A(net_1888), .B2(net_1640), .B1(net_1076) );
NAND2_X2 inst_11936 ( .A1(net_20860), .A2(net_1661), .ZN(net_1460) );
XNOR2_X2 inst_662 ( .A(net_21183), .B(net_21119), .ZN(net_306) );
INV_X4 inst_15590 ( .ZN(net_4065), .A(net_2250) );
CLKBUF_X2 inst_22579 ( .A(net_21710), .Z(net_22451) );
AOI21_X2 inst_20979 ( .B1(net_20553), .ZN(net_3709), .A(net_2015), .B2(net_1669) );
NOR2_X2 inst_3495 ( .ZN(net_19843), .A2(net_13468), .A1(net_9336) );
OAI21_X2 inst_1533 ( .B1(net_18003), .ZN(net_17976), .B2(net_17848), .A(net_2029) );
NAND2_X4 inst_7156 ( .ZN(net_11710), .A1(net_9573), .A2(net_4794) );
NAND2_X2 inst_7741 ( .ZN(net_18799), .A1(net_18756), .A2(net_18736) );
CLKBUF_X2 inst_22722 ( .A(net_22593), .Z(net_22594) );
CLKBUF_X2 inst_21778 ( .A(net_21649), .Z(net_21650) );
NAND2_X2 inst_11046 ( .A1(net_6601), .A2(net_5165), .ZN(net_4716) );
INV_X4 inst_12491 ( .ZN(net_18656), .A(net_18655) );
INV_X4 inst_17720 ( .ZN(net_3682), .A(net_194) );
INV_X2 inst_18574 ( .ZN(net_10682), .A(net_10681) );
INV_X4 inst_18243 ( .A(net_20994), .ZN(net_1856) );
INV_X2 inst_19050 ( .A(net_6695), .ZN(net_4739) );
XOR2_X1 inst_53 ( .B(net_21162), .Z(net_18651), .A(net_18649) );
NOR2_X2 inst_5030 ( .ZN(net_1587), .A1(net_956), .A2(net_764) );
INV_X4 inst_12653 ( .ZN(net_17854), .A(net_17853) );
AND2_X4 inst_21170 ( .ZN(net_13100), .A1(net_13099), .A2(net_13098) );
AOI21_X2 inst_20849 ( .B1(net_11943), .A(net_9972), .ZN(net_9095), .B2(net_9094) );
NOR2_X4 inst_3337 ( .ZN(net_699), .A2(net_164), .A1(net_163) );
NOR3_X4 inst_2614 ( .ZN(net_19939), .A1(net_15084), .A3(net_15007), .A2(net_10544) );
NOR2_X2 inst_4090 ( .A1(net_9917), .ZN(net_7255), .A2(net_6745) );
NAND2_X2 inst_10513 ( .ZN(net_8213), .A2(net_6939), .A1(net_6911) );
AOI21_X2 inst_20770 ( .B2(net_20647), .B1(net_20646), .ZN(net_10678), .A(net_146) );
OAI21_X2 inst_2111 ( .ZN(net_10040), .B2(net_6115), .B1(net_3994), .A(net_60) );
INV_X4 inst_14512 ( .ZN(net_5981), .A(net_4817) );
NAND2_X2 inst_8419 ( .ZN(net_17305), .A1(net_16926), .A2(net_16752) );
INV_X4 inst_13943 ( .A(net_12782), .ZN(net_8678) );
OAI21_X4 inst_1463 ( .B2(net_20348), .B1(net_20347), .ZN(net_15192), .A(net_1171) );
INV_X4 inst_14242 ( .ZN(net_7262), .A(net_5783) );
NAND2_X2 inst_9665 ( .ZN(net_12970), .A2(net_9755), .A1(net_8724) );
INV_X4 inst_16311 ( .ZN(net_2058), .A(net_892) );
INV_X4 inst_13463 ( .ZN(net_9704), .A(net_9703) );
SDFF_X2 inst_759 ( .Q(net_20940), .SE(net_18859), .SI(net_18524), .D(net_11877), .CK(net_22746) );
NAND2_X2 inst_11655 ( .ZN(net_2839), .A2(net_2439), .A1(net_868) );
INV_X4 inst_13192 ( .ZN(net_20044), .A(net_13467) );
DFF_X1 inst_19855 ( .D(net_17165), .CK(net_22105), .Q(x492) );
AND2_X2 inst_21272 ( .ZN(net_18942), .A2(net_14272), .A1(net_12999) );
INV_X2 inst_18776 ( .ZN(net_7546), .A(net_7545) );
NAND3_X2 inst_6596 ( .ZN(net_9907), .A1(net_6925), .A2(net_6165), .A3(net_6067) );
NAND2_X2 inst_9274 ( .ZN(net_12600), .A1(net_10930), .A2(net_10843) );
AOI21_X2 inst_20725 ( .A(net_14552), .ZN(net_11961), .B1(net_11849), .B2(net_7905) );
INV_X4 inst_18330 ( .A(net_20923), .ZN(net_20559) );
NOR2_X2 inst_3586 ( .ZN(net_20130), .A1(net_10971), .A2(net_9784) );
INV_X4 inst_13652 ( .ZN(net_11837), .A(net_8150) );
NAND2_X2 inst_7744 ( .ZN(net_18794), .A2(net_18759), .A1(net_18675) );
INV_X4 inst_14625 ( .A(net_15027), .ZN(net_12208) );
NAND2_X4 inst_7203 ( .ZN(net_10237), .A1(net_8867), .A2(net_4794) );
NAND2_X2 inst_9974 ( .A2(net_10637), .ZN(net_8880), .A1(net_8879) );
OAI21_X2 inst_2282 ( .A(net_8839), .ZN(net_6802), .B2(net_6801), .B1(net_1926) );
CLKBUF_X2 inst_21431 ( .A(net_21247), .Z(net_21303) );
INV_X4 inst_14594 ( .ZN(net_9258), .A(net_7740) );
NAND3_X2 inst_5718 ( .ZN(net_16138), .A3(net_15687), .A2(net_14861), .A1(net_12005) );
XNOR2_X2 inst_169 ( .B(net_21153), .A(net_17827), .ZN(net_17826) );
NAND3_X2 inst_6158 ( .A3(net_20025), .ZN(net_13647), .A1(net_12319), .A2(net_11995) );
AOI21_X2 inst_20873 ( .ZN(net_8540), .B1(net_8539), .A(net_8181), .B2(net_5391) );
INV_X4 inst_12880 ( .ZN(net_16854), .A(net_16853) );
NAND2_X2 inst_11748 ( .ZN(net_20786), .A2(net_2070), .A1(net_85) );
XNOR2_X2 inst_555 ( .A(net_17522), .B(net_17404), .ZN(net_12264) );
NAND2_X2 inst_8014 ( .ZN(net_18292), .A1(net_18291), .A2(net_18290) );
NAND2_X2 inst_10293 ( .A1(net_8868), .ZN(net_7914), .A2(net_5906) );
INV_X4 inst_12978 ( .A(net_17010), .ZN(net_16866) );
OR2_X2 inst_1184 ( .A1(net_6482), .A2(net_5564), .ZN(net_4710) );
INV_X4 inst_17148 ( .ZN(net_20601), .A(net_962) );
NAND2_X2 inst_9352 ( .ZN(net_12176), .A1(net_12175), .A2(net_12174) );
NOR2_X2 inst_4685 ( .ZN(net_5596), .A1(net_3368), .A2(net_3196) );
INV_X4 inst_14325 ( .A(net_11530), .ZN(net_5441) );
NAND3_X2 inst_6157 ( .A3(net_13744), .ZN(net_13664), .A2(net_9024), .A1(net_5624) );
CLKBUF_X2 inst_22810 ( .A(net_22681), .Z(net_22682) );
CLKBUF_X2 inst_22154 ( .A(net_22025), .Z(net_22026) );
CLKBUF_X2 inst_21661 ( .A(net_21405), .Z(net_21533) );
NAND2_X2 inst_7796 ( .ZN(net_18706), .A2(net_18693), .A1(net_17868) );
NAND2_X2 inst_8197 ( .A1(net_20519), .ZN(net_17886), .A2(net_17808) );
INV_X4 inst_12523 ( .ZN(net_18474), .A(net_18473) );
INV_X4 inst_14999 ( .A(net_5333), .ZN(net_4575) );
AOI21_X2 inst_20260 ( .B2(net_20936), .ZN(net_18592), .B1(net_15571), .A(net_15533) );
NAND3_X2 inst_6580 ( .ZN(net_10441), .A3(net_10440), .A2(net_6090), .A1(net_6069) );
INV_X2 inst_18754 ( .ZN(net_7738), .A(net_6465) );
NOR2_X2 inst_5140 ( .A1(net_1339), .A2(net_1009), .ZN(net_157) );
NAND2_X2 inst_9480 ( .A1(net_11642), .ZN(net_11458), .A2(net_11457) );
NAND2_X2 inst_11863 ( .ZN(net_3168), .A2(net_1778), .A1(net_1655) );
AND2_X4 inst_21255 ( .ZN(net_2278), .A2(net_783), .A1(net_279) );
NAND2_X2 inst_11578 ( .A1(net_4038), .ZN(net_3528), .A2(net_2735) );
NAND2_X2 inst_8756 ( .A1(net_16359), .ZN(net_15911), .A2(net_15514) );
INV_X8 inst_12273 ( .ZN(net_4820), .A(net_1622) );
NAND2_X4 inst_7521 ( .A2(net_20851), .ZN(net_20465), .A1(net_2066) );
NAND2_X2 inst_8952 ( .ZN(net_20371), .A2(net_13301), .A1(net_12203) );
AOI21_X4 inst_20215 ( .B1(net_19810), .ZN(net_14394), .A(net_12337), .B2(net_10142) );
INV_X4 inst_12931 ( .A(net_16876), .ZN(net_16653) );
NOR2_X2 inst_3991 ( .ZN(net_8277), .A1(net_8276), .A2(net_5662) );
NAND2_X2 inst_9546 ( .A1(net_12133), .ZN(net_11037), .A2(net_10929) );
INV_X4 inst_13620 ( .ZN(net_9808), .A(net_8359) );
INV_X4 inst_14812 ( .ZN(net_4544), .A(net_3951) );
NAND3_X2 inst_6203 ( .ZN(net_13301), .A3(net_9866), .A2(net_7702), .A1(net_5608) );
INV_X4 inst_15661 ( .A(net_2676), .ZN(net_2085) );
NOR2_X2 inst_3343 ( .ZN(net_18174), .A1(net_18102), .A2(net_18087) );
NAND2_X2 inst_8617 ( .ZN(net_20454), .A1(net_16648), .A2(net_16614) );
NOR2_X2 inst_4140 ( .ZN(net_8308), .A1(net_6930), .A2(net_5051) );
INV_X4 inst_13340 ( .ZN(net_11095), .A(net_11094) );
INV_X2 inst_19676 ( .A(net_20504), .ZN(net_20503) );
INV_X4 inst_16654 ( .ZN(net_6127), .A(net_3707) );
NOR3_X1 inst_2801 ( .A2(net_14628), .A3(net_6415), .ZN(net_5316), .A1(net_5315) );
NOR2_X2 inst_4219 ( .A1(net_9183), .ZN(net_7904), .A2(net_4911) );
OAI21_X2 inst_2303 ( .A(net_8472), .ZN(net_5860), .B2(net_5859), .B1(net_2861) );
NAND2_X2 inst_9153 ( .ZN(net_13392), .A1(net_11380), .A2(net_10583) );
INV_X4 inst_13714 ( .ZN(net_7835), .A(net_7834) );
NAND2_X2 inst_8090 ( .ZN(net_18132), .A2(net_18129), .A1(net_17760) );
INV_X4 inst_14765 ( .ZN(net_5657), .A(net_4055) );
INV_X4 inst_16991 ( .ZN(net_6812), .A(net_2630) );
INV_X4 inst_16369 ( .ZN(net_1775), .A(net_1282) );
INV_X2 inst_19375 ( .ZN(net_2176), .A(net_2175) );
NOR2_X2 inst_3771 ( .ZN(net_10287), .A1(net_10286), .A2(net_7738) );
INV_X4 inst_17895 ( .ZN(net_7489), .A(net_70) );
OAI21_X2 inst_1695 ( .B2(net_19777), .B1(net_19776), .ZN(net_15355), .A(net_14160) );
NAND3_X4 inst_5557 ( .ZN(net_19109), .A3(net_15745), .A1(net_15213), .A2(net_14907) );
AND2_X2 inst_21297 ( .ZN(net_10187), .A1(net_10186), .A2(net_10185) );
INV_X4 inst_17957 ( .A(net_21211), .ZN(net_15585) );
NAND2_X2 inst_8954 ( .A1(net_15044), .ZN(net_14719), .A2(net_13215) );
CLKBUF_X2 inst_21514 ( .A(net_21385), .Z(net_21386) );
INV_X2 inst_19322 ( .ZN(net_2603), .A(net_2602) );
NAND2_X2 inst_9724 ( .A2(net_11878), .ZN(net_10143), .A1(net_6021) );
INV_X4 inst_15851 ( .ZN(net_3171), .A(net_1115) );
AOI21_X4 inst_20138 ( .B1(net_16260), .ZN(net_16043), .B2(net_15508), .A(net_14286) );
OAI221_X2 inst_1339 ( .ZN(net_14247), .C2(net_13542), .A(net_13461), .B1(net_10292), .C1(net_8574), .B2(net_7352) );
NOR2_X2 inst_4284 ( .ZN(net_6054), .A1(net_6053), .A2(net_6052) );
NAND2_X2 inst_11235 ( .ZN(net_12096), .A1(net_11858), .A2(net_3944) );
NOR2_X2 inst_4971 ( .ZN(net_3094), .A1(net_1645), .A2(net_1122) );
NOR2_X2 inst_4724 ( .ZN(net_20779), .A1(net_20662), .A2(net_3101) );
INV_X4 inst_17672 ( .A(net_7489), .ZN(net_690) );
NOR2_X2 inst_4467 ( .A1(net_9478), .ZN(net_4489), .A2(net_3441) );
INV_X4 inst_13512 ( .ZN(net_11580), .A(net_9404) );
AOI21_X2 inst_20322 ( .B1(net_20591), .ZN(net_20263), .B2(net_15692), .A(net_11074) );
NOR2_X2 inst_3654 ( .ZN(net_11665), .A2(net_11664), .A1(net_5496) );
INV_X2 inst_18971 ( .ZN(net_11269), .A(net_5225) );
SDFF_X2 inst_977 ( .QN(net_21036), .D(net_356), .SE(net_263), .CK(net_21966), .SI(x2382) );
DFF_X1 inst_19925 ( .QN(net_21112), .D(net_13229), .CK(net_21685) );
NAND2_X4 inst_6901 ( .A1(net_20006), .ZN(net_17979), .A2(net_17834) );
AND2_X2 inst_21332 ( .A2(net_11217), .A1(net_8981), .ZN(net_5152) );
AOI21_X4 inst_20126 ( .B2(net_20889), .ZN(net_19166), .B1(net_18988), .A(net_14011) );
NOR2_X2 inst_4802 ( .ZN(net_5129), .A1(net_2499), .A2(net_107) );
XNOR2_X2 inst_297 ( .ZN(net_17122), .A(net_16633), .B(net_16404) );
INV_X4 inst_15402 ( .A(net_15183), .ZN(net_8734) );
NAND2_X2 inst_11728 ( .ZN(net_7669), .A1(net_3226), .A2(net_2229) );
INV_X4 inst_13145 ( .ZN(net_15055), .A(net_14624) );
INV_X4 inst_13933 ( .ZN(net_12282), .A(net_6845) );
INV_X4 inst_16334 ( .A(net_1625), .ZN(net_1302) );
DFF_X1 inst_19845 ( .D(net_17396), .CK(net_21348), .Q(x277) );
NOR2_X2 inst_3436 ( .ZN(net_15261), .A2(net_14665), .A1(net_1257) );
OAI21_X2 inst_2188 ( .ZN(net_8742), .A(net_8741), .B2(net_4856), .B1(net_4396) );
NOR2_X2 inst_3351 ( .A1(net_19427), .ZN(net_17839), .A2(net_17428) );
NAND2_X2 inst_10466 ( .ZN(net_7001), .A2(net_6992), .A1(net_5255) );
INV_X4 inst_13057 ( .ZN(net_19094), .A(net_16330) );
INV_X4 inst_17692 ( .ZN(net_11395), .A(net_333) );
XNOR2_X2 inst_162 ( .ZN(net_17899), .A(net_17843), .B(net_16265) );
INV_X4 inst_17645 ( .A(net_20889), .ZN(net_14476) );
NOR2_X4 inst_3308 ( .A2(net_20495), .ZN(net_1115), .A1(net_1114) );
CLKBUF_X2 inst_21769 ( .A(net_21288), .Z(net_21641) );
NAND2_X4 inst_7373 ( .ZN(net_10562), .A2(net_4304), .A1(net_3844) );
INV_X4 inst_14903 ( .ZN(net_4612), .A(net_3601) );
NAND2_X4 inst_7302 ( .ZN(net_11165), .A1(net_4914), .A2(net_4478) );
INV_X4 inst_17697 ( .A(net_992), .ZN(net_572) );
INV_X4 inst_13387 ( .ZN(net_13371), .A(net_10740) );
NOR2_X2 inst_3819 ( .ZN(net_19560), .A2(net_6174), .A1(net_5089) );
NOR2_X4 inst_2829 ( .A2(net_19880), .A1(net_19879), .ZN(net_19054) );
INV_X4 inst_15939 ( .ZN(net_12006), .A(net_8685) );
INV_X2 inst_18902 ( .ZN(net_6065), .A(net_6064) );
NOR2_X2 inst_3668 ( .ZN(net_11544), .A1(net_11543), .A2(net_7831) );
NAND2_X2 inst_11383 ( .ZN(net_9663), .A2(net_3949), .A1(net_1604) );
INV_X4 inst_16790 ( .ZN(net_5162), .A(net_4228) );
NAND2_X2 inst_12086 ( .ZN(net_5673), .A2(net_1376), .A1(net_93) );
AOI21_X2 inst_20720 ( .ZN(net_11986), .B1(net_8822), .B2(net_7716), .A(net_4517) );
NAND2_X2 inst_8143 ( .ZN(net_18022), .A2(net_17989), .A1(net_17967) );
INV_X4 inst_17681 ( .ZN(net_935), .A(net_248) );
OR2_X4 inst_1098 ( .ZN(net_8481), .A2(net_3294), .A1(net_573) );
INV_X2 inst_19473 ( .ZN(net_1428), .A(net_1427) );
NOR2_X2 inst_4149 ( .ZN(net_6906), .A1(net_6905), .A2(net_4115) );
NAND2_X4 inst_7077 ( .A1(net_19368), .ZN(net_18878), .A2(net_15880) );
OAI211_X2 inst_2443 ( .ZN(net_20384), .C1(net_20284), .C2(net_14820), .B(net_13558), .A(net_9724) );
NAND2_X2 inst_10051 ( .A1(net_12658), .ZN(net_8693), .A2(net_8150) );
SDFF_X2 inst_723 ( .Q(net_20873), .SE(net_18863), .SI(net_18573), .D(net_9003), .CK(net_21865) );
NAND2_X2 inst_8921 ( .ZN(net_14955), .A2(net_13739), .A1(net_10162) );
NAND2_X2 inst_10990 ( .ZN(net_9915), .A1(net_4931), .A2(net_4930) );
CLKBUF_X2 inst_21892 ( .A(net_21763), .Z(net_21764) );
NOR2_X2 inst_3893 ( .ZN(net_9189), .A2(net_9188), .A1(net_3548) );
NAND2_X2 inst_11055 ( .ZN(net_8594), .A1(net_2652), .A2(net_1804) );
NAND2_X2 inst_11616 ( .ZN(net_2583), .A2(net_2008), .A1(net_1769) );
NAND3_X2 inst_5777 ( .ZN(net_15867), .A1(net_15431), .A3(net_15342), .A2(net_14345) );
INV_X4 inst_13274 ( .ZN(net_12493), .A(net_11259) );
INV_X2 inst_18836 ( .A(net_9020), .ZN(net_6751) );
CLKBUF_X2 inst_22015 ( .A(net_21496), .Z(net_21887) );
AOI22_X2 inst_20006 ( .A1(net_15012), .B1(net_13198), .ZN(net_12895), .A2(net_9303), .B2(net_7207) );
OAI21_X2 inst_2067 ( .A(net_10945), .ZN(net_10663), .B2(net_8659), .B1(net_6339) );
NAND2_X2 inst_7894 ( .ZN(net_18492), .A2(net_18410), .A1(net_18349) );
DFF_X1 inst_19923 ( .QN(net_21114), .D(net_13224), .CK(net_21688) );
INV_X4 inst_14651 ( .ZN(net_12238), .A(net_6592) );
INV_X4 inst_18018 ( .A(net_21010), .ZN(net_686) );
INV_X4 inst_17851 ( .A(net_396), .ZN(net_215) );
NAND2_X2 inst_8268 ( .A1(net_17775), .ZN(net_17656), .A2(net_17590) );
INV_X4 inst_13075 ( .ZN(net_16226), .A(net_16169) );
AND2_X2 inst_21290 ( .ZN(net_12167), .A1(net_12166), .A2(net_12165) );
NOR3_X2 inst_2777 ( .ZN(net_7747), .A3(net_4545), .A1(net_3757), .A2(net_2145) );
INV_X8 inst_12283 ( .A(net_5043), .ZN(net_3184) );
NAND3_X2 inst_6784 ( .ZN(net_20671), .A1(net_4232), .A2(net_3175), .A3(net_3057) );
NAND2_X4 inst_6830 ( .ZN(net_18819), .A2(net_18789), .A1(net_17573) );
INV_X4 inst_17031 ( .A(net_4917), .ZN(net_4270) );
INV_X2 inst_19692 ( .A(net_20545), .ZN(net_20544) );
INV_X2 inst_18360 ( .A(net_18295), .ZN(net_18241) );
OAI211_X2 inst_2446 ( .ZN(net_14668), .C2(net_13713), .B(net_5998), .A(net_4904), .C1(net_4325) );
NOR2_X2 inst_5046 ( .A2(net_4099), .A1(net_1214), .ZN(net_1073) );
INV_X4 inst_13602 ( .ZN(net_8608), .A(net_7184) );
NAND2_X2 inst_7840 ( .ZN(net_18622), .A2(net_18608), .A1(net_17426) );
NAND2_X2 inst_8452 ( .ZN(net_17198), .A1(net_16731), .A2(net_16578) );
AND2_X2 inst_21343 ( .ZN(net_2845), .A1(net_2676), .A2(net_2424) );
INV_X2 inst_19094 ( .ZN(net_4548), .A(net_4547) );
INV_X4 inst_14128 ( .A(net_7948), .ZN(net_7527) );
INV_X4 inst_13070 ( .ZN(net_18936), .A(net_16219) );
AOI21_X2 inst_20698 ( .ZN(net_19673), .B1(net_9628), .B2(net_5819), .A(net_145) );
INV_X4 inst_15549 ( .ZN(net_4206), .A(net_1557) );
INV_X4 inst_14260 ( .ZN(net_5738), .A(net_5737) );
NAND4_X4 inst_5210 ( .ZN(net_19432), .A1(net_16240), .A4(net_16059), .A2(net_15886), .A3(net_10827) );
NAND3_X2 inst_6613 ( .A1(net_9759), .ZN(net_9077), .A2(net_9076), .A3(net_9075) );
INV_X4 inst_12767 ( .ZN(net_17458), .A(net_17339) );
INV_X4 inst_17820 ( .ZN(net_303), .A(net_189) );
INV_X4 inst_16611 ( .A(net_14684), .ZN(net_1125) );
NAND4_X2 inst_5464 ( .ZN(net_19330), .A2(net_19285), .A1(net_19284), .A4(net_13260), .A3(net_5431) );
AOI22_X2 inst_20054 ( .A1(net_6682), .B1(net_6525), .ZN(net_3699), .B2(net_3278), .A2(net_1476) );
INV_X4 inst_16676 ( .A(net_15649), .ZN(net_1613) );
INV_X2 inst_18718 ( .ZN(net_11912), .A(net_8159) );
INV_X4 inst_14089 ( .A(net_6205), .ZN(net_6204) );
INV_X4 inst_18070 ( .A(net_20871), .ZN(net_814) );
INV_X2 inst_18438 ( .ZN(net_19408), .A(net_13612) );
AOI21_X2 inst_20867 ( .ZN(net_8595), .B1(net_8594), .B2(net_4901), .A(net_127) );
NAND2_X2 inst_8366 ( .ZN(net_17373), .A1(net_17372), .A2(net_17341) );
OAI21_X2 inst_1818 ( .ZN(net_14162), .A(net_14086), .B1(net_11121), .B2(net_10611) );
NAND2_X4 inst_7110 ( .ZN(net_13772), .A1(net_10932), .A2(net_4694) );
INV_X4 inst_18341 ( .ZN(net_20714), .A(net_20711) );
NAND2_X2 inst_10705 ( .A2(net_6126), .ZN(net_6029), .A1(net_6028) );
INV_X4 inst_14706 ( .ZN(net_5910), .A(net_4246) );
NAND2_X2 inst_10264 ( .A1(net_11297), .ZN(net_10178), .A2(net_8050) );
OAI21_X2 inst_1766 ( .ZN(net_14702), .A(net_12885), .B2(net_12062), .B1(net_9823) );
INV_X4 inst_13888 ( .ZN(net_7319), .A(net_7318) );
INV_X2 inst_18897 ( .A(net_7954), .ZN(net_6099) );
NAND2_X2 inst_8216 ( .A1(net_20520), .ZN(net_17840), .A2(net_17807) );
CLKBUF_X2 inst_22496 ( .A(net_22367), .Z(net_22368) );
INV_X4 inst_15398 ( .ZN(net_4870), .A(net_2540) );
NAND2_X2 inst_9639 ( .ZN(net_20817), .A1(net_10395), .A2(net_8375) );
AOI21_X2 inst_20499 ( .B1(net_15524), .ZN(net_14655), .A(net_14289), .B2(net_12092) );
NOR2_X2 inst_4548 ( .ZN(net_6875), .A1(net_5551), .A2(net_1905) );
INV_X4 inst_17679 ( .ZN(net_3904), .A(net_758) );
SDFF_X2 inst_876 ( .Q(net_21215), .SI(net_17041), .SE(net_125), .CK(net_22292), .D(x7527) );
NOR2_X4 inst_2979 ( .ZN(net_9776), .A2(net_6394), .A1(net_4637) );
AOI21_X2 inst_20685 ( .ZN(net_12261), .B1(net_11214), .A(net_9565), .B2(net_8517) );
AND2_X2 inst_21296 ( .A1(net_11970), .A2(net_10655), .ZN(net_10392) );
NOR2_X2 inst_4727 ( .ZN(net_3097), .A2(net_3096), .A1(net_2671) );
INV_X2 inst_19182 ( .A(net_4362), .ZN(net_3770) );
OAI211_X2 inst_2433 ( .ZN(net_15022), .A(net_13753), .B(net_12593), .C2(net_12559), .C1(net_1369) );
NAND2_X2 inst_11665 ( .ZN(net_2393), .A2(net_2317), .A1(net_850) );
NAND2_X2 inst_11751 ( .ZN(net_2115), .A2(net_2114), .A1(net_63) );
OAI211_X2 inst_2480 ( .ZN(net_13496), .C1(net_13495), .C2(net_13494), .A(net_8954), .B(net_6728) );
XNOR2_X2 inst_562 ( .B(net_18141), .ZN(net_679), .A(net_678) );
NAND2_X2 inst_9845 ( .ZN(net_10970), .A2(net_9392), .A1(net_8048) );
NAND2_X2 inst_8917 ( .ZN(net_14961), .A1(net_14055), .A2(net_13645) );
INV_X4 inst_14714 ( .ZN(net_18837), .A(net_18025) );
CLKBUF_X2 inst_22616 ( .A(net_22487), .Z(net_22488) );
NAND3_X2 inst_6385 ( .A2(net_20780), .ZN(net_12020), .A3(net_8051), .A1(net_3366) );
NAND2_X2 inst_11445 ( .ZN(net_5587), .A2(net_3094), .A1(net_2274) );
INV_X4 inst_15006 ( .A(net_11866), .ZN(net_11439) );
NAND2_X4 inst_7615 ( .A2(net_20800), .ZN(net_2294), .A1(net_1344) );
NAND2_X2 inst_8277 ( .ZN(net_17722), .A2(net_17496), .A1(net_17375) );
NOR2_X2 inst_4953 ( .ZN(net_7155), .A1(net_4792), .A2(net_3737) );
INV_X8 inst_12404 ( .ZN(net_3745), .A(net_165) );
NAND2_X2 inst_9589 ( .ZN(net_12311), .A2(net_7557), .A1(net_6295) );
NAND2_X4 inst_7164 ( .ZN(net_12791), .A1(net_9466), .A2(net_9465) );
NOR2_X2 inst_3659 ( .A1(net_14346), .ZN(net_12695), .A2(net_11622) );
CLKBUF_X2 inst_21459 ( .A(net_21330), .Z(net_21331) );
NOR2_X2 inst_3604 ( .A1(net_20512), .ZN(net_12430), .A2(net_9112) );
NAND2_X4 inst_7465 ( .ZN(net_5556), .A1(net_2731), .A2(net_956) );
INV_X4 inst_17028 ( .ZN(net_10096), .A(net_8709) );
OR2_X4 inst_1109 ( .ZN(net_5510), .A2(net_1454), .A1(net_1065) );
NAND3_X2 inst_6487 ( .ZN(net_11176), .A2(net_11175), .A3(net_11174), .A1(net_3894) );
AOI22_X2 inst_20052 ( .A1(net_6636), .ZN(net_3702), .A2(net_2701), .B1(net_1607), .B2(net_1434) );
NAND2_X2 inst_12054 ( .ZN(net_3777), .A1(net_900), .A2(net_297) );
NOR2_X4 inst_3037 ( .ZN(net_6253), .A1(net_3644), .A2(net_1138) );
NAND2_X2 inst_11522 ( .ZN(net_5346), .A1(net_4286), .A2(net_2366) );
INV_X4 inst_14857 ( .ZN(net_3799), .A(net_3798) );
OAI22_X2 inst_1314 ( .B2(net_12478), .ZN(net_7108), .A1(net_6879), .A2(net_5605), .B1(net_5220) );
NAND2_X2 inst_7956 ( .ZN(net_18394), .A2(net_18393), .A1(net_17222) );
OR2_X2 inst_1156 ( .A1(net_14617), .A2(net_8348), .ZN(net_8317) );
NAND3_X4 inst_5533 ( .A3(net_20286), .A1(net_20285), .ZN(net_17653), .A2(net_16191) );
NOR2_X2 inst_3378 ( .A1(net_21196), .A2(net_16560), .ZN(net_16430) );
INV_X4 inst_16458 ( .ZN(net_1690), .A(net_338) );
NAND2_X2 inst_11466 ( .ZN(net_5413), .A1(net_4394), .A2(net_3246) );
NAND3_X2 inst_5993 ( .ZN(net_14529), .A1(net_13391), .A3(net_10423), .A2(net_4679) );
INV_X4 inst_12512 ( .A(net_18633), .ZN(net_18618) );
INV_X4 inst_13676 ( .ZN(net_13641), .A(net_8670) );
INV_X4 inst_14259 ( .A(net_9256), .ZN(net_7293) );
INV_X2 inst_19313 ( .A(net_11204), .ZN(net_2659) );
OAI21_X2 inst_1880 ( .ZN(net_13652), .B1(net_13651), .B2(net_13650), .A(net_8354) );
OAI22_X2 inst_1295 ( .ZN(net_11868), .A1(net_11682), .B1(net_11617), .A2(net_9732), .B2(net_4095) );
INV_X2 inst_19333 ( .ZN(net_2517), .A(net_2516) );
NAND2_X4 inst_7457 ( .A2(net_20535), .A1(net_20298), .ZN(net_3768) );
XNOR2_X2 inst_262 ( .ZN(net_17258), .A(net_17254), .B(net_16627) );
NOR2_X2 inst_3630 ( .ZN(net_12213), .A2(net_10421), .A1(net_4689) );
NOR2_X2 inst_4675 ( .A1(net_20541), .ZN(net_3240), .A2(net_2091) );
NAND2_X2 inst_10333 ( .ZN(net_20029), .A1(net_9510), .A2(net_7583) );
INV_X4 inst_16644 ( .A(net_14764), .ZN(net_12627) );
AOI21_X2 inst_20336 ( .ZN(net_20367), .B1(net_19095), .B2(net_15582), .A(net_13082) );
CLKBUF_X2 inst_21939 ( .A(net_21810), .Z(net_21811) );
SDFF_X2 inst_1035 ( .QN(net_21031), .D(net_724), .SE(net_263), .CK(net_21952), .SI(x2468) );
NAND2_X2 inst_7942 ( .ZN(net_18422), .A2(net_18361), .A1(net_18303) );
INV_X2 inst_18466 ( .ZN(net_12731), .A(net_12730) );
NOR2_X2 inst_3637 ( .A2(net_13823), .ZN(net_12183), .A1(net_8662) );
NAND2_X2 inst_11490 ( .A1(net_20537), .ZN(net_3999), .A2(net_3091) );
INV_X4 inst_17286 ( .ZN(net_2788), .A(net_834) );
OAI21_X2 inst_1883 ( .ZN(net_13535), .B1(net_13534), .B2(net_11553), .A(net_10662) );
NAND2_X4 inst_7240 ( .ZN(net_10433), .A1(net_7000), .A2(net_6951) );
NAND2_X2 inst_9580 ( .ZN(net_12603), .A2(net_10927), .A1(net_4018) );
INV_X4 inst_12863 ( .ZN(net_16999), .A(net_16998) );
AOI21_X2 inst_20693 ( .ZN(net_12202), .B2(net_7823), .B1(net_5873), .A(net_816) );
NOR2_X2 inst_3621 ( .ZN(net_12316), .A1(net_12315), .A2(net_9416) );
SDFF_X2 inst_864 ( .Q(net_21147), .SI(net_17118), .SE(net_125), .CK(net_22151), .D(x3376) );
XNOR2_X2 inst_86 ( .ZN(net_18567), .A(net_18505), .B(net_17817) );
SDFF_X2 inst_949 ( .QN(net_21073), .D(net_479), .SE(net_263), .CK(net_21740), .SI(x1869) );
INV_X4 inst_18306 ( .A(net_20493), .ZN(net_20492) );
NOR2_X4 inst_3283 ( .A1(net_20868), .ZN(net_2133), .A2(net_1284) );
INV_X4 inst_12580 ( .ZN(net_18169), .A(net_18168) );
INV_X4 inst_16195 ( .ZN(net_8952), .A(net_5344) );
INV_X4 inst_15651 ( .ZN(net_4275), .A(net_1646) );
NOR2_X2 inst_3730 ( .ZN(net_12308), .A1(net_10886), .A2(net_9125) );
INV_X4 inst_13294 ( .ZN(net_19065), .A(net_12355) );
NOR2_X2 inst_3598 ( .ZN(net_12554), .A1(net_9737), .A2(net_6759) );
NAND2_X2 inst_10342 ( .ZN(net_11025), .A2(net_4554), .A1(net_1790) );
AOI21_X2 inst_20755 ( .ZN(net_11228), .B2(net_9665), .A(net_6226), .B1(net_761) );
CLKBUF_X2 inst_21683 ( .A(net_21554), .Z(net_21555) );
INV_X4 inst_17237 ( .ZN(net_2074), .A(net_662) );
OAI21_X2 inst_2109 ( .A(net_14070), .ZN(net_10045), .B2(net_6157), .B1(net_4059) );
OAI21_X2 inst_1826 ( .ZN(net_14139), .B1(net_11095), .B2(net_7375), .A(net_1052) );
NAND2_X1 inst_12140 ( .A2(net_20711), .ZN(net_17265), .A1(net_631) );
NAND4_X2 inst_5395 ( .A2(net_20322), .A1(net_20321), .ZN(net_14810), .A4(net_10116), .A3(net_5514) );
OAI21_X2 inst_2020 ( .ZN(net_11343), .B1(net_11209), .A(net_10592), .B2(net_6948) );
NAND3_X2 inst_6192 ( .ZN(net_13316), .A2(net_11902), .A3(net_9862), .A1(net_8407) );
NOR2_X2 inst_4361 ( .ZN(net_5976), .A1(net_5503), .A2(net_3342) );
NOR2_X4 inst_2820 ( .ZN(net_16560), .A1(net_16241), .A2(net_16165) );
INV_X4 inst_13721 ( .A(net_7810), .ZN(net_7809) );
CLKBUF_X2 inst_22417 ( .A(net_22288), .Z(net_22289) );
OAI211_X2 inst_2404 ( .ZN(net_15802), .C1(net_15374), .A(net_15277), .B(net_11513), .C2(net_7778) );
INV_X4 inst_14417 ( .ZN(net_6197), .A(net_3652) );
NAND2_X2 inst_7994 ( .A2(net_18360), .ZN(net_18321), .A1(net_17815) );
INV_X4 inst_14075 ( .ZN(net_7572), .A(net_6224) );
INV_X4 inst_15539 ( .ZN(net_11962), .A(net_2366) );
OAI21_X2 inst_1578 ( .A(net_20888), .B2(net_19585), .B1(net_19584), .ZN(net_16313) );
NAND2_X2 inst_7849 ( .ZN(net_20587), .A2(net_18601), .A1(net_15891) );
CLKBUF_X2 inst_21578 ( .A(net_21425), .Z(net_21450) );
NAND2_X4 inst_7662 ( .A1(net_958), .ZN(net_914), .A2(net_913) );
INV_X4 inst_17714 ( .ZN(net_19376), .A(net_244) );
NAND2_X2 inst_9053 ( .A1(net_15174), .ZN(net_14005), .A2(net_12029) );
NOR2_X2 inst_4612 ( .ZN(net_3720), .A1(net_3719), .A2(net_2172) );
CLKBUF_X2 inst_22242 ( .A(net_22113), .Z(net_22114) );
NAND2_X2 inst_9598 ( .ZN(net_13898), .A1(net_9937), .A2(net_9333) );
INV_X2 inst_19363 ( .ZN(net_2248), .A(net_2247) );
NAND2_X2 inst_11398 ( .ZN(net_3469), .A2(net_2139), .A1(net_874) );
INV_X4 inst_15676 ( .ZN(net_2800), .A(net_1570) );
NAND2_X2 inst_8820 ( .ZN(net_15563), .A2(net_14819), .A1(net_12376) );
INV_X2 inst_18802 ( .ZN(net_7416), .A(net_7415) );
INV_X2 inst_19533 ( .ZN(net_20662), .A(net_1491) );
XNOR2_X2 inst_175 ( .ZN(net_17780), .A(net_17548), .B(net_3375) );
NAND2_X2 inst_11989 ( .ZN(net_1249), .A2(net_657), .A1(net_570) );
AOI21_X2 inst_20617 ( .ZN(net_13547), .A(net_8870), .B2(net_7553), .B1(net_5124) );
NOR2_X2 inst_5010 ( .A2(net_3002), .ZN(net_2769), .A1(net_2490) );
NAND2_X2 inst_10491 ( .ZN(net_20200), .A1(net_11476), .A2(net_4061) );
AOI21_X2 inst_20726 ( .ZN(net_11958), .B1(net_11834), .B2(net_5382), .A(net_2302) );
INV_X2 inst_18596 ( .A(net_12036), .ZN(net_10744) );
INV_X4 inst_15764 ( .A(net_9490), .ZN(net_4468) );
OAI21_X2 inst_1737 ( .ZN(net_15068), .A(net_14483), .B1(net_13500), .B2(net_11768) );
NAND2_X2 inst_10895 ( .A1(net_9438), .ZN(net_5398), .A2(net_5397) );
NOR2_X4 inst_2995 ( .ZN(net_9854), .A1(net_5934), .A2(net_4110) );
NAND2_X2 inst_8594 ( .A2(net_17752), .A1(net_16701), .ZN(net_16691) );
CLKBUF_X2 inst_22641 ( .A(net_22512), .Z(net_22513) );
AOI21_X2 inst_20449 ( .ZN(net_19880), .A(net_15087), .B2(net_12893), .B1(net_10889) );
NAND2_X4 inst_7081 ( .A1(net_19600), .ZN(net_18988), .A2(net_11075) );
NAND4_X2 inst_5513 ( .ZN(net_10763), .A2(net_10762), .A4(net_7145), .A3(net_5607), .A1(net_3832) );
CLKBUF_X2 inst_21745 ( .A(net_21616), .Z(net_21617) );
NOR2_X2 inst_4541 ( .A1(net_20541), .ZN(net_4732), .A2(net_3992) );
INV_X4 inst_14073 ( .A(net_7984), .ZN(net_7575) );
INV_X4 inst_18017 ( .A(net_21228), .ZN(net_16402) );
OR2_X2 inst_1149 ( .ZN(net_9848), .A2(net_9847), .A1(net_2276) );
NAND2_X2 inst_10146 ( .A1(net_10037), .ZN(net_8297), .A2(net_6187) );
INV_X4 inst_14354 ( .ZN(net_5756), .A(net_5274) );
NAND3_X2 inst_5640 ( .ZN(net_17999), .A2(net_17962), .A3(net_17961), .A1(net_17591) );
NAND2_X2 inst_9696 ( .A1(net_12056), .A2(net_10773), .ZN(net_10224) );
NAND2_X2 inst_11475 ( .ZN(net_7113), .A2(net_3129), .A1(net_143) );
NOR2_X2 inst_4719 ( .ZN(net_5305), .A2(net_1858), .A1(net_222) );
INV_X4 inst_15026 ( .ZN(net_15360), .A(net_14363) );
INV_X4 inst_17617 ( .ZN(net_305), .A(net_304) );
AOI21_X2 inst_20706 ( .ZN(net_12112), .B2(net_8010), .A(net_6321), .B1(net_2820) );
NOR2_X2 inst_4353 ( .A2(net_12939), .ZN(net_5615), .A1(net_3143) );
NAND3_X2 inst_6003 ( .ZN(net_14428), .A3(net_12449), .A1(net_7853), .A2(net_3252) );
NAND2_X2 inst_9285 ( .ZN(net_12544), .A2(net_9653), .A1(net_60) );
CLKBUF_X2 inst_21592 ( .A(net_21463), .Z(net_21464) );
NOR2_X2 inst_3934 ( .A1(net_9673), .ZN(net_8705), .A2(net_8704) );
NAND2_X2 inst_9716 ( .ZN(net_10169), .A1(net_10168), .A2(net_7710) );
INV_X4 inst_17602 ( .ZN(net_4208), .A(net_321) );
SDFF_X2 inst_948 ( .QN(net_21088), .SE(net_2426), .D(net_376), .CK(net_21795), .SI(x1603) );
INV_X4 inst_12475 ( .ZN(net_18752), .A(net_18709) );
INV_X4 inst_13302 ( .ZN(net_14216), .A(net_12303) );
CLKBUF_X2 inst_21731 ( .A(net_21602), .Z(net_21603) );
INV_X4 inst_17250 ( .A(net_7450), .ZN(net_2884) );
AOI22_X2 inst_20026 ( .A1(net_10920), .ZN(net_9930), .B2(net_9929), .A2(net_8201), .B1(net_1941) );
CLKBUF_X2 inst_22059 ( .A(net_21930), .Z(net_21931) );
INV_X2 inst_18414 ( .ZN(net_20818), .A(net_15783) );
INV_X4 inst_14795 ( .ZN(net_4000), .A(net_3999) );
AOI21_X2 inst_20962 ( .B1(net_5797), .A(net_5575), .ZN(net_5314), .B2(net_2842) );
NAND3_X2 inst_6644 ( .ZN(net_10227), .A1(net_8751), .A3(net_7900), .A2(net_6736) );
INV_X4 inst_13493 ( .ZN(net_11516), .A(net_9469) );
NAND2_X2 inst_11407 ( .A1(net_6135), .ZN(net_4493), .A2(net_3439) );
INV_X4 inst_16079 ( .A(net_1737), .ZN(net_1549) );
NAND2_X2 inst_11275 ( .A1(net_7962), .ZN(net_3876), .A2(net_3875) );
INV_X4 inst_15892 ( .ZN(net_6963), .A(net_1830) );
NAND2_X2 inst_8039 ( .ZN(net_18253), .A1(net_18252), .A2(net_18251) );
NAND2_X2 inst_11647 ( .A2(net_7077), .ZN(net_2478), .A1(net_2477) );
INV_X4 inst_15579 ( .ZN(net_11446), .A(net_5415) );
NAND4_X2 inst_5444 ( .ZN(net_13881), .A1(net_13880), .A2(net_13879), .A3(net_13878), .A4(net_6450) );
NAND2_X2 inst_9966 ( .ZN(net_20740), .A2(net_8895), .A1(net_1864) );
INV_X4 inst_14671 ( .ZN(net_4320), .A(net_4319) );
CLKBUF_X2 inst_22256 ( .A(net_22127), .Z(net_22128) );
OAI21_X2 inst_2002 ( .A(net_13534), .ZN(net_11646), .B2(net_11023), .B1(net_4618) );
NOR2_X2 inst_4380 ( .A1(net_11087), .ZN(net_5347), .A2(net_5346) );
NAND3_X2 inst_6030 ( .A3(net_19892), .ZN(net_14369), .A1(net_13768), .A2(net_8163) );
CLKBUF_X2 inst_22476 ( .A(net_22347), .Z(net_22348) );
NAND2_X2 inst_8430 ( .ZN(net_19269), .A1(net_17177), .A2(net_17138) );
NAND2_X2 inst_10471 ( .ZN(net_6988), .A2(net_4082), .A1(net_3821) );
AOI21_X2 inst_20684 ( .A(net_12504), .ZN(net_12292), .B1(net_7930), .B2(net_7208) );
XNOR2_X2 inst_608 ( .A(net_21137), .B(net_17774), .ZN(net_7650) );
SDFF_X2 inst_834 ( .Q(net_21190), .SI(net_17506), .SE(net_125), .CK(net_22319), .D(x6350) );
AOI22_X2 inst_20042 ( .ZN(net_7079), .B1(net_7078), .B2(net_7077), .A1(net_5344), .A2(net_4267) );
NAND2_X2 inst_11183 ( .ZN(net_6986), .A1(net_6201), .A2(net_4112) );
INV_X4 inst_16869 ( .ZN(net_8616), .A(net_3049) );
NOR2_X4 inst_2920 ( .ZN(net_8072), .A2(net_8071), .A1(net_6058) );
NAND2_X2 inst_8729 ( .ZN(net_16064), .A2(net_15772), .A1(net_8734) );
AOI21_X2 inst_20607 ( .B1(net_14552), .ZN(net_13750), .A(net_13577), .B2(net_9307) );
SDFF_X2 inst_966 ( .QN(net_21102), .D(net_599), .SE(net_263), .CK(net_21777), .SI(x1362) );
INV_X4 inst_14951 ( .ZN(net_6044), .A(net_3508) );
NOR2_X4 inst_2961 ( .A2(net_11041), .ZN(net_8622), .A1(net_6610) );
NAND2_X4 inst_7189 ( .ZN(net_12124), .A2(net_7798), .A1(net_5387) );
NAND2_X2 inst_8924 ( .ZN(net_14946), .A1(net_14945), .A2(net_13685) );
NAND2_X2 inst_11833 ( .ZN(net_1982), .A1(net_1759), .A2(net_1758) );
OAI211_X2 inst_2506 ( .ZN(net_12765), .A(net_12764), .C1(net_12763), .C2(net_12762), .B(net_8054) );
INV_X4 inst_13214 ( .ZN(net_13639), .A(net_12819) );
NAND3_X2 inst_5836 ( .A3(net_20371), .A2(net_20370), .ZN(net_15511), .A1(net_14638) );
NAND3_X2 inst_5976 ( .ZN(net_14741), .A2(net_14740), .A3(net_12321), .A1(net_6921) );
AOI21_X2 inst_20357 ( .ZN(net_15687), .B1(net_15553), .B2(net_15015), .A(net_14790) );
NAND4_X4 inst_5245 ( .A2(net_20687), .A1(net_20686), .A4(net_18963), .ZN(net_14584), .A3(net_6242) );
NAND3_X4 inst_5575 ( .ZN(net_15771), .A3(net_15129), .A2(net_13340), .A1(net_7294) );
AND3_X2 inst_21140 ( .ZN(net_11250), .A2(net_11249), .A3(net_7037), .A1(net_2790) );
CLKBUF_X2 inst_22719 ( .A(net_22590), .Z(net_22591) );
NOR2_X2 inst_4557 ( .ZN(net_6883), .A2(net_3937), .A1(net_1445) );
AND2_X2 inst_21277 ( .ZN(net_13801), .A1(net_13800), .A2(net_12309) );
NOR2_X2 inst_3607 ( .ZN(net_12426), .A2(net_12425), .A1(net_4772) );
CLKBUF_X2 inst_22233 ( .A(net_22104), .Z(net_22105) );
NAND2_X2 inst_8583 ( .ZN(net_16719), .A2(net_16718), .A1(net_16631) );
NAND2_X2 inst_10498 ( .ZN(net_11374), .A1(net_8037), .A2(net_6944) );
INV_X4 inst_13324 ( .ZN(net_20732), .A(net_10076) );
INV_X4 inst_16395 ( .A(net_2400), .ZN(net_1701) );
AOI21_X2 inst_20574 ( .ZN(net_14131), .B1(net_13448), .B2(net_10624), .A(net_7680) );
NOR2_X4 inst_3160 ( .ZN(net_3912), .A2(net_3244), .A1(net_3070) );
INV_X4 inst_14022 ( .ZN(net_10540), .A(net_8250) );
NOR2_X4 inst_2861 ( .ZN(net_15285), .A2(net_11440), .A1(net_10896) );
INV_X4 inst_14825 ( .ZN(net_6707), .A(net_3773) );
XNOR2_X2 inst_66 ( .ZN(net_18823), .B(net_18753), .A(net_17735) );
NOR2_X2 inst_4814 ( .ZN(net_2580), .A2(net_1484), .A1(net_1018) );
NAND2_X2 inst_11139 ( .ZN(net_4966), .A2(net_4247), .A1(net_222) );
NAND2_X2 inst_11012 ( .ZN(net_11158), .A2(net_4859), .A1(net_3297) );
NAND2_X2 inst_7920 ( .ZN(net_18454), .A2(net_18377), .A1(net_17731) );
NAND2_X2 inst_10604 ( .ZN(net_6614), .A2(net_4705), .A1(net_703) );
NAND2_X2 inst_8807 ( .ZN(net_15622), .A1(net_14961), .A2(net_14703) );
XNOR2_X2 inst_273 ( .ZN(net_17210), .A(net_16830), .B(net_635) );
INV_X8 inst_12297 ( .ZN(net_1751), .A(net_562) );
INV_X4 inst_13443 ( .A(net_9787), .ZN(net_9786) );
CLKBUF_X2 inst_22586 ( .A(net_21782), .Z(net_22458) );
INV_X4 inst_15365 ( .ZN(net_3692), .A(net_2263) );
CLKBUF_X2 inst_21762 ( .A(net_21531), .Z(net_21634) );
CLKBUF_X2 inst_21677 ( .A(net_21514), .Z(net_21549) );
OAI211_X2 inst_2418 ( .ZN(net_15407), .A(net_14387), .C2(net_12824), .B(net_7197), .C1(net_1001) );
XNOR2_X2 inst_366 ( .ZN(net_16851), .A(net_16848), .B(net_13951) );
DFF_X1 inst_19797 ( .D(net_18225), .CK(net_22404), .Q(x790) );
NAND3_X2 inst_6162 ( .A2(net_20350), .A1(net_20349), .ZN(net_13640), .A3(net_11948) );
NAND2_X4 inst_7019 ( .ZN(net_17498), .A1(net_16582), .A2(net_16455) );
CLKBUF_X2 inst_22860 ( .A(net_21812), .Z(net_22732) );
NAND2_X2 inst_9397 ( .ZN(net_11701), .A2(net_9671), .A1(net_7646) );
NAND2_X2 inst_9565 ( .ZN(net_13616), .A2(net_11526), .A1(net_10966) );
INV_X4 inst_12542 ( .ZN(net_18343), .A(net_18342) );
NAND2_X2 inst_7964 ( .ZN(net_18369), .A2(net_18365), .A1(net_17206) );
INV_X4 inst_16845 ( .ZN(net_4481), .A(net_4163) );
INV_X4 inst_16737 ( .ZN(net_10737), .A(net_809) );
NAND2_X4 inst_7313 ( .ZN(net_12011), .A2(net_5353), .A1(net_2996) );
NOR2_X2 inst_4746 ( .ZN(net_7048), .A1(net_3069), .A2(net_3038) );
NAND3_X2 inst_5896 ( .ZN(net_19976), .A3(net_14020), .A1(net_11920), .A2(net_10657) );
NAND2_X2 inst_7950 ( .ZN(net_18401), .A1(net_18276), .A2(net_18235) );
INV_X2 inst_18353 ( .ZN(net_18768), .A(net_18767) );
AOI21_X2 inst_20837 ( .ZN(net_9286), .A(net_9285), .B2(net_4548), .B1(net_2768) );
SDFF_X2 inst_707 ( .Q(net_20954), .SE(net_18859), .SI(net_18822), .D(net_385), .CK(net_22266) );
SDFF_X2 inst_1025 ( .QN(net_20982), .D(net_1900), .SE(net_253), .CK(net_21831), .SI(x3290) );
NOR2_X2 inst_4655 ( .A1(net_7268), .ZN(net_5397), .A2(net_2049) );
NOR2_X2 inst_3670 ( .ZN(net_11519), .A1(net_11518), .A2(net_11454) );
NAND2_X4 inst_7566 ( .A1(net_20538), .ZN(net_2080), .A2(net_1669) );
NAND2_X4 inst_7570 ( .ZN(net_3019), .A2(net_1753), .A1(net_221) );
NAND3_X2 inst_5635 ( .A2(net_20588), .A1(net_20587), .ZN(net_18603), .A3(net_18589) );
NAND2_X2 inst_7834 ( .A1(net_20522), .ZN(net_18634), .A2(net_18633) );
AOI211_X2 inst_21017 ( .ZN(net_15552), .C1(net_15369), .C2(net_14582), .B(net_13760), .A(net_11575) );
NAND3_X4 inst_5542 ( .A3(net_19201), .A1(net_19200), .ZN(net_17040), .A2(net_14351) );
NAND2_X2 inst_8654 ( .A1(net_21159), .ZN(net_16545), .A2(net_16515) );
NAND2_X2 inst_10080 ( .ZN(net_13168), .A1(net_9254), .A2(net_7859) );
INV_X4 inst_16730 ( .ZN(net_2696), .A(net_1050) );
INV_X4 inst_15094 ( .A(net_11770), .ZN(net_3248) );
OAI211_X2 inst_2576 ( .ZN(net_8482), .A(net_8481), .B(net_8480), .C2(net_6495), .C1(net_1425) );
NAND2_X4 inst_7269 ( .ZN(net_7561), .A2(net_6200), .A1(net_3696) );
INV_X4 inst_13654 ( .ZN(net_9646), .A(net_8148) );
INV_X4 inst_13710 ( .ZN(net_11886), .A(net_7859) );
NOR3_X4 inst_2631 ( .ZN(net_14578), .A1(net_12725), .A3(net_11796), .A2(net_11248) );
INV_X4 inst_15988 ( .ZN(net_2503), .A(net_1220) );
AOI21_X2 inst_20404 ( .B2(net_18990), .B1(net_18989), .ZN(net_15349), .A(net_15289) );
NOR2_X2 inst_3810 ( .ZN(net_20626), .A1(net_9834), .A2(net_7444) );
NAND2_X2 inst_8453 ( .ZN(net_17196), .A2(net_16746), .A1(net_16611) );
INV_X4 inst_13261 ( .ZN(net_12687), .A(net_11604) );
NOR2_X2 inst_4523 ( .ZN(net_4086), .A1(net_4085), .A2(net_4084) );
AOI22_X2 inst_20036 ( .B1(net_8521), .ZN(net_7662), .A1(net_7661), .A2(net_3487), .B2(net_2156) );
NAND2_X4 inst_7073 ( .A2(net_20156), .A1(net_20155), .ZN(net_15983) );
CLKBUF_X2 inst_21845 ( .A(net_21716), .Z(net_21717) );
NOR3_X2 inst_2636 ( .ZN(net_19989), .A1(net_16003), .A2(net_12530), .A3(net_11753) );
NAND3_X2 inst_6198 ( .A3(net_19107), .A1(net_19106), .ZN(net_18906), .A2(net_8074) );
INV_X4 inst_18039 ( .A(net_21015), .ZN(net_536) );
NAND2_X4 inst_7186 ( .ZN(net_19369), .A2(net_8833), .A1(net_8832) );
INV_X4 inst_16380 ( .A(net_8629), .ZN(net_3156) );
NAND2_X4 inst_7579 ( .ZN(net_3036), .A1(net_1692), .A2(net_200) );
DFF_X1 inst_19886 ( .D(net_17124), .CK(net_22084), .Q(x511) );
INV_X4 inst_16038 ( .ZN(net_11682), .A(net_6889) );
NAND2_X2 inst_11561 ( .ZN(net_5054), .A1(net_1848), .A2(net_1801) );
INV_X4 inst_14491 ( .ZN(net_14874), .A(net_9993) );
XNOR2_X2 inst_445 ( .B(net_21109), .ZN(net_15295), .A(net_15294) );
INV_X4 inst_12961 ( .A(net_17526), .ZN(net_16535) );
INV_X4 inst_13618 ( .ZN(net_12040), .A(net_8891) );
NAND4_X4 inst_5192 ( .A3(net_19318), .A1(net_19317), .A4(net_19100), .ZN(net_17010), .A2(net_16099) );
NAND2_X2 inst_11566 ( .ZN(net_2799), .A1(net_2798), .A2(net_2797) );
NAND2_X2 inst_11400 ( .ZN(net_3464), .A2(net_3463), .A1(net_809) );
INV_X4 inst_17501 ( .ZN(net_1138), .A(net_107) );
INV_X8 inst_12350 ( .ZN(net_9131), .A(net_307) );
INV_X4 inst_15406 ( .ZN(net_15804), .A(net_14572) );
NOR2_X2 inst_3761 ( .ZN(net_10338), .A1(net_10337), .A2(net_9794) );
NOR2_X2 inst_5089 ( .A2(net_3861), .ZN(net_847), .A1(net_846) );
NAND3_X2 inst_5654 ( .ZN(net_16548), .A3(net_16405), .A2(net_16314), .A1(net_14193) );
NAND2_X2 inst_10138 ( .A2(net_20771), .ZN(net_19293), .A1(net_13556) );
SDFF_X2 inst_853 ( .Q(net_21187), .SI(net_17251), .SE(net_125), .CK(net_22299), .D(x6430) );
NAND3_X2 inst_5864 ( .ZN(net_19714), .A3(net_13731), .A1(net_11309), .A2(net_10364) );
XNOR2_X2 inst_657 ( .ZN(net_351), .A(net_350), .B(net_349) );
NOR2_X2 inst_4550 ( .A2(net_20578), .ZN(net_6918), .A1(net_3356) );
INV_X4 inst_12803 ( .ZN(net_17223), .A(net_17222) );
OAI21_X2 inst_2098 ( .A(net_10175), .ZN(net_10071), .B2(net_9974), .B1(net_4065) );
INV_X4 inst_12465 ( .ZN(net_18791), .A(net_18790) );
OAI21_X2 inst_1921 ( .ZN(net_20746), .A(net_11779), .B2(net_11497), .B1(net_5219) );
INV_X4 inst_17467 ( .ZN(net_6570), .A(net_721) );
INV_X4 inst_12890 ( .A(net_17244), .ZN(net_16967) );
INV_X4 inst_13890 ( .ZN(net_11884), .A(net_10496) );
CLKBUF_X2 inst_21965 ( .A(net_21558), .Z(net_21837) );
INV_X2 inst_19636 ( .A(net_19425), .ZN(net_19424) );
NAND2_X4 inst_6977 ( .ZN(net_17320), .A1(net_16905), .A2(net_16715) );
INV_X2 inst_19568 ( .ZN(net_1758), .A(net_780) );
NOR2_X2 inst_4293 ( .ZN(net_7463), .A1(net_6797), .A2(net_5380) );
INV_X4 inst_13996 ( .A(net_8830), .ZN(net_7470) );
INV_X4 inst_14783 ( .ZN(net_6679), .A(net_4028) );
NAND2_X2 inst_10357 ( .ZN(net_7440), .A1(net_7439), .A2(net_5814) );
INV_X4 inst_14285 ( .ZN(net_7057), .A(net_5627) );
NOR3_X2 inst_2638 ( .ZN(net_16007), .A3(net_15420), .A1(net_15063), .A2(net_13067) );
NAND2_X2 inst_8676 ( .A1(net_19449), .ZN(net_16458), .A2(net_16384) );
DFF_X1 inst_19849 ( .D(net_17221), .CK(net_21345), .Q(x107) );
NOR2_X4 inst_3235 ( .ZN(net_4302), .A1(net_3402), .A2(net_2293) );
INV_X4 inst_14019 ( .A(net_7769), .ZN(net_6297) );
NAND2_X2 inst_8672 ( .ZN(net_20744), .A2(net_16619), .A1(net_16464) );
INV_X4 inst_14680 ( .ZN(net_4308), .A(net_4307) );
INV_X4 inst_12786 ( .ZN(net_17298), .A(net_17297) );
NAND2_X2 inst_9421 ( .A1(net_14867), .A2(net_12957), .ZN(net_11633) );
CLKBUF_X2 inst_21972 ( .A(net_21843), .Z(net_21844) );
NAND2_X2 inst_8711 ( .A1(net_20960), .ZN(net_20728), .A2(net_16056) );
CLKBUF_X2 inst_21435 ( .A(net_21306), .Z(net_21307) );
NAND2_X2 inst_8125 ( .ZN(net_18053), .A2(net_18032), .A1(net_7389) );
SDFF_X2 inst_892 ( .Q(net_21152), .D(net_17002), .SE(net_263), .CK(net_22216), .SI(x5637) );
AOI21_X2 inst_20361 ( .A(net_15666), .ZN(net_15662), .B2(net_14914), .B1(net_13750) );
INV_X4 inst_17175 ( .ZN(net_877), .A(net_602) );
NOR2_X2 inst_4100 ( .A1(net_14186), .A2(net_13456), .ZN(net_7216) );
INV_X4 inst_16053 ( .A(net_1737), .ZN(net_1592) );
INV_X4 inst_17560 ( .ZN(net_15178), .A(net_512) );
OAI21_X2 inst_1803 ( .A(net_15088), .ZN(net_14478), .B2(net_12701), .B1(net_6494) );
NAND2_X4 inst_6987 ( .ZN(net_17607), .A1(net_16860), .A2(net_16690) );
NOR2_X4 inst_2814 ( .ZN(net_17268), .A1(net_16829), .A2(net_16674) );
SDFF_X2 inst_936 ( .QN(net_21086), .D(net_681), .SE(net_263), .CK(net_22605), .SI(x1639) );
NAND2_X2 inst_9819 ( .A1(net_11572), .ZN(net_9648), .A2(net_9647) );
NOR2_X2 inst_3809 ( .ZN(net_9835), .A2(net_7446), .A1(net_6530) );
INV_X4 inst_14957 ( .ZN(net_5739), .A(net_3498) );
CLKBUF_X2 inst_22769 ( .A(net_21921), .Z(net_22641) );
NAND2_X2 inst_11368 ( .ZN(net_3580), .A2(net_3301), .A1(net_2168) );
INV_X4 inst_14896 ( .ZN(net_4567), .A(net_3629) );
NAND2_X2 inst_10315 ( .ZN(net_10156), .A2(net_6578), .A1(net_1910) );
NAND3_X2 inst_6171 ( .A2(net_19845), .ZN(net_13612), .A1(net_12646), .A3(net_9566) );
INV_X4 inst_14236 ( .A(net_8187), .ZN(net_5815) );
INV_X4 inst_15300 ( .ZN(net_2690), .A(net_2689) );
NAND2_X4 inst_6865 ( .ZN(net_18318), .A2(net_18301), .A1(net_17738) );
CLKBUF_X2 inst_22661 ( .A(net_22532), .Z(net_22533) );
INV_X4 inst_12948 ( .A(net_17330), .ZN(net_17107) );
NOR2_X2 inst_3780 ( .ZN(net_10136), .A2(net_10135), .A1(net_6689) );
NOR3_X2 inst_2647 ( .ZN(net_15721), .A1(net_15397), .A3(net_13986), .A2(net_7682) );
NAND2_X2 inst_11305 ( .ZN(net_11077), .A1(net_7872), .A2(net_2819) );
INV_X2 inst_18938 ( .A(net_7596), .ZN(net_5822) );
NAND3_X2 inst_6576 ( .ZN(net_10453), .A3(net_10452), .A2(net_6046), .A1(net_4943) );
INV_X2 inst_19090 ( .ZN(net_4558), .A(net_4557) );
INV_X4 inst_15464 ( .ZN(net_2468), .A(net_2467) );
NOR3_X2 inst_2710 ( .A2(net_14593), .ZN(net_13688), .A1(net_12456), .A3(net_10947) );
NAND3_X4 inst_5629 ( .ZN(net_5140), .A2(net_4324), .A1(net_4038), .A3(net_154) );
NAND2_X2 inst_11959 ( .A2(net_2384), .ZN(net_1388), .A1(net_856) );
OR3_X4 inst_1058 ( .ZN(net_10649), .A1(net_10648), .A2(net_10647), .A3(net_10646) );
CLKBUF_X2 inst_22069 ( .A(net_21940), .Z(net_21941) );
INV_X4 inst_12639 ( .ZN(net_17911), .A(net_17910) );
AOI211_X2 inst_21003 ( .ZN(net_19297), .C1(net_15897), .B(net_15203), .A(net_14386), .C2(net_13928) );
NOR2_X2 inst_3360 ( .ZN(net_17423), .A1(net_17422), .A2(net_17421) );
INV_X4 inst_16441 ( .A(net_1246), .ZN(net_1235) );
NAND3_X1 inst_6821 ( .A2(net_20742), .ZN(net_13882), .A1(net_13864), .A3(net_11181) );
NOR2_X2 inst_4984 ( .ZN(net_3092), .A1(net_1848), .A2(net_1336) );
INV_X2 inst_18539 ( .A(net_11712), .ZN(net_11014) );
CLKBUF_X2 inst_22564 ( .A(net_21582), .Z(net_22436) );
INV_X4 inst_18206 ( .A(net_20973), .ZN(net_856) );
OAI21_X2 inst_1788 ( .ZN(net_14645), .B2(net_11765), .A(net_10683), .B1(net_9916) );
INV_X4 inst_14098 ( .ZN(net_7558), .A(net_6180) );
AOI21_X2 inst_20749 ( .ZN(net_11370), .A(net_8298), .B1(net_7198), .B2(net_4379) );
OAI22_X2 inst_1272 ( .B1(net_21180), .ZN(net_16805), .A2(net_16804), .A1(net_16607), .B2(net_16421) );
INV_X4 inst_17780 ( .ZN(net_624), .A(net_112) );
NOR2_X2 inst_4182 ( .ZN(net_8099), .A2(net_6794), .A1(net_6207) );
INV_X4 inst_14566 ( .A(net_7702), .ZN(net_7583) );
NOR2_X4 inst_2852 ( .A2(net_19755), .A1(net_19754), .ZN(net_19615) );
NAND3_X2 inst_6751 ( .ZN(net_14783), .A1(net_8739), .A2(net_6127), .A3(net_5386) );
INV_X4 inst_17008 ( .ZN(net_1219), .A(net_863) );
AOI21_X2 inst_20954 ( .B1(net_12306), .ZN(net_5340), .B2(net_4180), .A(net_3734) );
INV_X2 inst_18458 ( .ZN(net_13261), .A(net_12251) );
NOR2_X2 inst_3973 ( .ZN(net_8405), .A1(net_8404), .A2(net_8364) );
NAND2_X4 inst_7584 ( .ZN(net_1570), .A2(net_1071), .A1(net_826) );
XNOR2_X2 inst_433 ( .ZN(net_16335), .A(net_16334), .B(net_16091) );
INV_X4 inst_13771 ( .ZN(net_11118), .A(net_7594) );
AOI21_X2 inst_20813 ( .ZN(net_10085), .B1(net_6485), .B2(net_6029), .A(net_333) );
NOR2_X2 inst_4939 ( .ZN(net_20394), .A2(net_2751), .A1(net_1195) );
NAND2_X2 inst_11817 ( .ZN(net_3315), .A1(net_1821), .A2(net_1246) );
INV_X4 inst_13249 ( .ZN(net_20299), .A(net_11804) );
INV_X2 inst_18925 ( .ZN(net_5913), .A(net_5912) );
INV_X4 inst_17605 ( .ZN(net_894), .A(net_314) );
INV_X2 inst_18454 ( .ZN(net_13423), .A(net_13422) );
NAND3_X2 inst_6417 ( .ZN(net_11946), .A1(net_9243), .A3(net_7337), .A2(net_5049) );
NAND2_X2 inst_11312 ( .ZN(net_6721), .A2(net_3781), .A1(net_2557) );
INV_X4 inst_13772 ( .ZN(net_11116), .A(net_9285) );
NAND2_X2 inst_8984 ( .ZN(net_14495), .A2(net_13006), .A1(net_11997) );
INV_X4 inst_16411 ( .ZN(net_13525), .A(net_13452) );
NAND2_X2 inst_11955 ( .ZN(net_1963), .A1(net_261), .A2(net_86) );
NAND2_X2 inst_8638 ( .A1(net_16902), .A2(net_16718), .ZN(net_16581) );
NAND2_X2 inst_9269 ( .A2(net_19464), .ZN(net_14878), .A1(net_13383) );
NAND3_X2 inst_5781 ( .ZN(net_15801), .A2(net_15800), .A3(net_14849), .A1(net_14266) );
AOI211_X2 inst_21041 ( .ZN(net_13485), .C2(net_12436), .A(net_11418), .B(net_10711), .C1(net_4512) );
INV_X4 inst_13476 ( .ZN(net_11712), .A(net_9614) );
INV_X4 inst_14733 ( .A(net_4116), .ZN(net_4115) );
NAND2_X4 inst_7151 ( .ZN(net_12835), .A1(net_8592), .A2(net_8241) );
INV_X4 inst_15325 ( .ZN(net_14395), .A(net_8611) );
INV_X4 inst_17564 ( .A(net_14557), .ZN(net_1000) );
AND3_X4 inst_21113 ( .ZN(net_15675), .A3(net_14984), .A2(net_14740), .A1(net_6272) );
OAI21_X4 inst_1475 ( .B2(net_20452), .B1(net_20451), .ZN(net_19645), .A(net_14568) );
INV_X4 inst_15960 ( .ZN(net_2600), .A(net_2107) );
OAI21_X2 inst_1637 ( .ZN(net_19630), .B2(net_19524), .B1(net_19523), .A(net_15450) );
OAI21_X4 inst_1352 ( .B2(net_19512), .B1(net_19511), .A(net_18601), .ZN(net_18593) );
CLKBUF_X2 inst_22873 ( .A(net_21297), .Z(net_22745) );
INV_X4 inst_17079 ( .ZN(net_3990), .A(net_2230) );
INV_X8 inst_12338 ( .ZN(net_6849), .A(net_572) );
AOI21_X2 inst_20532 ( .ZN(net_14522), .B1(net_12583), .B2(net_10136), .A(net_1030) );
OAI21_X2 inst_2261 ( .A(net_13699), .ZN(net_7166), .B2(net_7120), .B1(net_2324) );
NAND2_X2 inst_9955 ( .A1(net_10061), .ZN(net_8926), .A2(net_6508) );
AND3_X2 inst_21138 ( .ZN(net_19903), .A2(net_13168), .A3(net_13167), .A1(net_6708) );
INV_X2 inst_18374 ( .ZN(net_20230), .A(net_17515) );
INV_X4 inst_14524 ( .ZN(net_9870), .A(net_4771) );
NOR2_X2 inst_3390 ( .ZN(net_16167), .A2(net_15935), .A1(net_10556) );
NAND2_X2 inst_9076 ( .ZN(net_13833), .A1(net_13089), .A2(net_11692) );
INV_X4 inst_15742 ( .ZN(net_3641), .A(net_1950) );
INV_X4 inst_16945 ( .ZN(net_1127), .A(net_917) );
NOR2_X4 inst_2930 ( .ZN(net_19601), .A1(net_7729), .A2(net_4375) );
NAND2_X4 inst_7609 ( .A2(net_1751), .ZN(net_1382), .A1(net_343) );
NAND2_X2 inst_8178 ( .ZN(net_17936), .A2(net_17838), .A1(net_17787) );
CLKBUF_X2 inst_22139 ( .A(net_21365), .Z(net_22011) );
NAND3_X2 inst_5683 ( .ZN(net_16323), .A3(net_16073), .A2(net_13358), .A1(net_11726) );
AOI21_X2 inst_20855 ( .ZN(net_9030), .B1(net_7723), .B2(net_6765), .A(net_862) );
NOR2_X2 inst_4790 ( .ZN(net_2789), .A1(net_2788), .A2(net_2787) );
NOR2_X2 inst_4307 ( .ZN(net_7422), .A1(net_5918), .A2(net_4571) );
NAND2_X2 inst_9851 ( .ZN(net_9528), .A2(net_7575), .A1(net_7394) );
INV_X4 inst_18082 ( .A(net_21006), .ZN(net_1865) );
NOR2_X4 inst_3192 ( .ZN(net_4012), .A2(net_2993), .A1(net_1076) );
NOR2_X2 inst_5006 ( .A1(net_1607), .ZN(net_1305), .A2(net_1304) );
CLKBUF_X2 inst_21864 ( .A(net_21735), .Z(net_21736) );
NAND2_X2 inst_9026 ( .ZN(net_19791), .A1(net_14085), .A2(net_11914) );
INV_X2 inst_18485 ( .ZN(net_12384), .A(net_12383) );
NAND2_X2 inst_9780 ( .A2(net_10647), .A1(net_10395), .ZN(net_9765) );
INV_X2 inst_19078 ( .ZN(net_4597), .A(net_4596) );
INV_X4 inst_13585 ( .ZN(net_10403), .A(net_8913) );
NAND2_X2 inst_11129 ( .ZN(net_10638), .A1(net_9109), .A2(net_4272) );
CLKBUF_X2 inst_22424 ( .A(net_22295), .Z(net_22296) );
NOR2_X2 inst_4246 ( .A2(net_13956), .A1(net_12884), .ZN(net_6494) );
NAND2_X2 inst_9146 ( .A1(net_15360), .ZN(net_13405), .A2(net_10653) );
NOR2_X2 inst_3904 ( .A2(net_10609), .ZN(net_8890), .A1(net_8889) );
DFF_X1 inst_19869 ( .D(net_17096), .CK(net_22798), .Q(x1259) );
NAND2_X2 inst_10634 ( .ZN(net_19276), .A1(net_4418), .A2(net_3059) );
NAND3_X2 inst_6333 ( .A3(net_20267), .A1(net_20266), .ZN(net_19810), .A2(net_10873) );
NAND3_X2 inst_5649 ( .A3(net_20168), .A1(net_20167), .ZN(net_17003), .A2(net_15562) );
OAI21_X4 inst_1393 ( .A(net_20848), .B2(net_19582), .B1(net_19581), .ZN(net_16279) );
NAND3_X2 inst_6276 ( .ZN(net_12906), .A2(net_11874), .A1(net_9883), .A3(net_9337) );
NOR2_X2 inst_3519 ( .ZN(net_13758), .A2(net_12568), .A1(net_81) );
NOR2_X2 inst_4075 ( .ZN(net_7496), .A1(net_7472), .A2(net_2431) );
INV_X4 inst_13402 ( .ZN(net_10425), .A(net_10424) );
INV_X4 inst_16191 ( .ZN(net_1414), .A(net_1413) );
INV_X4 inst_17948 ( .A(net_21011), .ZN(net_578) );
AOI222_X1 inst_20069 ( .ZN(net_11917), .C1(net_11296), .A1(net_7975), .A2(net_7541), .C2(net_5422), .B2(net_4516), .B1(net_1619) );
INV_X4 inst_15720 ( .ZN(net_11485), .A(net_10292) );
INV_X4 inst_16576 ( .ZN(net_9349), .A(net_4931) );
NOR2_X1 inst_5153 ( .A1(net_12363), .ZN(net_7808), .A2(net_7807) );
NAND3_X2 inst_5731 ( .ZN(net_18980), .A1(net_15852), .A3(net_15393), .A2(net_12543) );
INV_X4 inst_14264 ( .A(net_7677), .ZN(net_5725) );
INV_X4 inst_15913 ( .ZN(net_1872), .A(net_1748) );
NAND2_X2 inst_8631 ( .ZN(net_16592), .A1(net_16512), .A2(net_16467) );
INV_X4 inst_13118 ( .A(net_21110), .ZN(net_17091) );
INV_X4 inst_14446 ( .ZN(net_7939), .A(net_4983) );
INV_X2 inst_18610 ( .ZN(net_9701), .A(net_9700) );
NOR2_X2 inst_4791 ( .A1(net_4655), .ZN(net_4096), .A2(net_2781) );
NAND3_X2 inst_6459 ( .ZN(net_11394), .A1(net_11393), .A2(net_9550), .A3(net_6286) );
CLKBUF_X2 inst_22481 ( .A(net_22027), .Z(net_22353) );
NAND2_X2 inst_8007 ( .ZN(net_18302), .A2(net_18301), .A1(net_17627) );
INV_X4 inst_15866 ( .ZN(net_11443), .A(net_3041) );
NOR2_X4 inst_2937 ( .A1(net_11614), .ZN(net_7242), .A2(net_6774) );
NAND2_X4 inst_7244 ( .ZN(net_11640), .A2(net_6995), .A1(net_107) );
CLKBUF_X2 inst_22547 ( .A(net_22418), .Z(net_22419) );
INV_X4 inst_17124 ( .ZN(net_7010), .A(net_777) );
XNOR2_X1 inst_687 ( .B(net_17494), .ZN(net_17032), .A(net_17031) );
NAND2_X2 inst_7864 ( .ZN(net_18557), .A1(net_18504), .A2(net_18220) );
OAI21_X2 inst_2319 ( .ZN(net_5676), .A(net_5675), .B1(net_5674), .B2(net_5673) );
NAND2_X4 inst_7091 ( .A1(net_20660), .ZN(net_19172), .A2(net_14463) );
CLKBUF_X2 inst_22444 ( .A(net_22315), .Z(net_22316) );
CLKBUF_X2 inst_22283 ( .A(net_21565), .Z(net_22155) );
DFF_X1 inst_19865 ( .D(net_17105), .CK(net_22361), .Q(x756) );
NAND4_X2 inst_5519 ( .A2(net_9072), .A4(net_8546), .ZN(net_8487), .A3(net_8486), .A1(net_2946) );
INV_X2 inst_19403 ( .ZN(net_3463), .A(net_2702) );
OAI21_X2 inst_2225 ( .B1(net_20482), .ZN(net_8477), .B2(net_8476), .A(net_5146) );
NAND2_X2 inst_7927 ( .ZN(net_18444), .A2(net_18358), .A1(net_17400) );
INV_X2 inst_19561 ( .ZN(net_831), .A(net_830) );
INV_X4 inst_16523 ( .ZN(net_2076), .A(net_963) );
INV_X4 inst_13805 ( .ZN(net_10952), .A(net_7548) );
INV_X4 inst_17889 ( .A(net_189), .ZN(net_71) );
INV_X4 inst_17428 ( .ZN(net_2179), .A(net_168) );
NOR2_X2 inst_4061 ( .ZN(net_19007), .A1(net_14166), .A2(net_7829) );
OAI211_X2 inst_2513 ( .B(net_13174), .ZN(net_12458), .C1(net_12457), .A(net_7480), .C2(net_6212) );
OAI21_X2 inst_2254 ( .ZN(net_7286), .B2(net_4086), .B1(net_3737), .A(net_2463) );
INV_X4 inst_14690 ( .ZN(net_4453), .A(net_4284) );
DFF_X1 inst_19789 ( .D(net_18657), .CK(net_21625), .Q(x577) );
NAND2_X2 inst_7775 ( .ZN(net_18782), .A2(net_18730), .A1(net_17063) );
INV_X2 inst_18844 ( .A(net_10573), .ZN(net_10124) );
NAND3_X2 inst_6255 ( .A3(net_14844), .ZN(net_13004), .A2(net_12976), .A1(net_9705) );
NAND2_X2 inst_10111 ( .ZN(net_8427), .A2(net_5942), .A1(net_5223) );
INV_X2 inst_19380 ( .ZN(net_2148), .A(net_2147) );
AOI21_X4 inst_20103 ( .ZN(net_19063), .B1(net_16390), .A(net_16315), .B2(net_16140) );
NAND2_X2 inst_9255 ( .ZN(net_12648), .A1(net_12647), .A2(net_12646) );
CLKBUF_X2 inst_22933 ( .A(net_21277), .Z(net_22805) );
INV_X4 inst_16531 ( .ZN(net_2255), .A(net_1178) );
CLKBUF_X2 inst_22387 ( .A(net_22258), .Z(net_22259) );
NAND2_X2 inst_10922 ( .A1(net_9510), .ZN(net_5276), .A2(net_3074) );
INV_X4 inst_12519 ( .ZN(net_19767), .A(net_18539) );
INV_X4 inst_15479 ( .ZN(net_6400), .A(net_2453) );
INV_X4 inst_16640 ( .A(net_1389), .ZN(net_1362) );
AOI21_X2 inst_20612 ( .B1(net_13984), .ZN(net_13671), .A(net_12503), .B2(net_8689) );
CLKBUF_X2 inst_22374 ( .A(net_22245), .Z(net_22246) );
DFF_X1 inst_19842 ( .D(net_17284), .CK(net_22381), .Q(x866) );
NAND2_X2 inst_11755 ( .A1(net_3356), .ZN(net_2105), .A2(net_1045) );
XNOR2_X2 inst_354 ( .B(net_17015), .A(net_16935), .ZN(net_16928) );
INV_X4 inst_13794 ( .ZN(net_10903), .A(net_7561) );
OR2_X2 inst_1145 ( .A1(net_13922), .A2(net_10265), .ZN(net_10115) );
CLKBUF_X2 inst_22779 ( .A(net_22650), .Z(net_22651) );
AOI211_X2 inst_21010 ( .ZN(net_15766), .C1(net_15649), .C2(net_15013), .B(net_13758), .A(net_11223) );
NAND3_X2 inst_6235 ( .ZN(net_13214), .A2(net_13213), .A3(net_13169), .A1(net_8313) );
INV_X4 inst_12859 ( .ZN(net_20668), .A(net_16895) );
INV_X4 inst_15380 ( .A(net_6083), .ZN(net_3369) );
INV_X4 inst_15981 ( .A(net_9421), .ZN(net_9018) );
INV_X2 inst_18545 ( .A(net_11558), .ZN(net_10980) );
AOI21_X2 inst_20529 ( .B1(net_14990), .ZN(net_14526), .B2(net_11709), .A(net_11667) );
INV_X4 inst_14804 ( .ZN(net_14653), .A(net_8264) );
AOI21_X4 inst_20147 ( .B1(net_20112), .ZN(net_20012), .A(net_15449), .B2(net_15356) );
INV_X4 inst_16521 ( .A(net_8067), .ZN(net_7836) );
NAND2_X2 inst_7731 ( .ZN(net_18818), .A2(net_18772), .A1(net_17855) );
INV_X4 inst_16006 ( .A(net_1953), .ZN(net_1658) );
NAND2_X2 inst_8414 ( .ZN(net_17229), .A2(net_17227), .A1(net_833) );
CLKBUF_X2 inst_22596 ( .A(net_22467), .Z(net_22468) );
OAI21_X2 inst_1717 ( .ZN(net_15185), .A(net_14006), .B2(net_13953), .B1(net_8400) );
INV_X2 inst_18359 ( .ZN(net_18408), .A(net_18344) );
INV_X4 inst_15206 ( .A(net_3339), .ZN(net_2902) );
NOR2_X4 inst_2901 ( .ZN(net_19688), .A2(net_7127), .A1(net_5108) );
CLKBUF_X2 inst_22770 ( .A(net_22641), .Z(net_22642) );
AND2_X2 inst_21360 ( .A1(net_1195), .ZN(net_1079), .A2(net_110) );
NAND3_X2 inst_6080 ( .ZN(net_13969), .A1(net_13968), .A2(net_13914), .A3(net_10422) );
SDFF_X2 inst_718 ( .Q(net_20927), .SE(net_18863), .SI(net_18754), .D(net_638), .CK(net_22010) );
INV_X4 inst_17488 ( .ZN(net_783), .A(net_313) );
INV_X4 inst_17707 ( .A(net_242), .ZN(net_209) );
NOR2_X2 inst_4024 ( .ZN(net_9560), .A1(net_8020), .A2(net_8019) );
INV_X4 inst_18254 ( .A(net_21008), .ZN(net_565) );
NAND2_X4 inst_7362 ( .ZN(net_8093), .A1(net_4419), .A2(net_2493) );
NAND2_X2 inst_8100 ( .A2(net_20503), .ZN(net_18120), .A1(net_17136) );
NAND2_X2 inst_9166 ( .ZN(net_13373), .A1(net_11494), .A2(net_10427) );
INV_X2 inst_19506 ( .A(net_1593), .ZN(net_1227) );
NAND3_X4 inst_5585 ( .ZN(net_15444), .A3(net_14399), .A1(net_9205), .A2(net_8464) );
NAND2_X2 inst_8350 ( .ZN(net_17471), .A1(net_17470), .A2(net_17469) );
CLKBUF_X2 inst_22448 ( .A(net_21661), .Z(net_22320) );
INV_X4 inst_17827 ( .A(net_1009), .ZN(net_236) );
OAI21_X2 inst_2147 ( .ZN(net_9744), .B1(net_5143), .B2(net_3594), .A(net_1209) );
INV_X4 inst_13171 ( .ZN(net_14621), .A(net_14122) );
OAI21_X2 inst_2091 ( .ZN(net_10217), .A(net_10216), .B1(net_7425), .B2(net_3817) );
INV_X2 inst_19135 ( .ZN(net_4147), .A(net_4146) );
INV_X2 inst_18423 ( .ZN(net_15265), .A(net_14868) );
NAND2_X2 inst_10733 ( .ZN(net_7888), .A1(net_6635), .A2(net_5780) );
INV_X8 inst_12247 ( .ZN(net_3629), .A(net_2342) );
NAND2_X2 inst_8066 ( .A2(net_20793), .ZN(net_18185), .A1(net_17444) );
NAND3_X2 inst_5863 ( .ZN(net_15338), .A3(net_13732), .A1(net_12535), .A2(net_10372) );
AOI21_X2 inst_20495 ( .ZN(net_14737), .A(net_13059), .B2(net_12220), .B1(net_1296) );
INV_X4 inst_16783 ( .ZN(net_2862), .A(net_1017) );
XNOR2_X2 inst_500 ( .B(net_15588), .ZN(net_9000), .A(net_6459) );
NAND4_X2 inst_5348 ( .ZN(net_20688), .A1(net_14549), .A2(net_14442), .A4(net_13779), .A3(net_8535) );
INV_X4 inst_14403 ( .ZN(net_5691), .A(net_5108) );
XNOR2_X2 inst_550 ( .A(net_21194), .B(net_17534), .ZN(net_811) );
CLKBUF_X2 inst_22760 ( .A(net_22631), .Z(net_22632) );
NAND3_X2 inst_6758 ( .A2(net_12478), .ZN(net_5672), .A3(net_5671), .A1(net_2628) );
INV_X4 inst_16270 ( .A(net_9994), .ZN(net_8252) );
INV_X4 inst_17213 ( .ZN(net_1027), .A(net_700) );
NAND3_X2 inst_5913 ( .A2(net_20833), .A1(net_20832), .ZN(net_15010), .A3(net_11815) );
NAND2_X2 inst_11972 ( .ZN(net_1812), .A2(net_1343), .A1(net_252) );
INV_X4 inst_13610 ( .ZN(net_8434), .A(net_7076) );
NAND2_X2 inst_8311 ( .A2(net_20509), .ZN(net_17584), .A1(net_16994) );
INV_X4 inst_17761 ( .ZN(net_14104), .A(net_14022) );
NAND2_X2 inst_8702 ( .A1(net_20888), .ZN(net_19576), .A2(net_16130) );
INV_X4 inst_15417 ( .ZN(net_3391), .A(net_2518) );
NAND4_X2 inst_5471 ( .ZN(net_13216), .A3(net_12989), .A2(net_11656), .A1(net_8438), .A4(net_7148) );
NOR3_X2 inst_2661 ( .ZN(net_15036), .A1(net_13942), .A2(net_10548), .A3(net_10297) );
NAND2_X2 inst_8237 ( .A1(net_17756), .ZN(net_17750), .A2(net_17109) );
NAND3_X2 inst_6034 ( .ZN(net_14338), .A2(net_14337), .A3(net_14336), .A1(net_7226) );
NOR2_X2 inst_3548 ( .ZN(net_20726), .A1(net_12674), .A2(net_11349) );
INV_X4 inst_15246 ( .ZN(net_2809), .A(net_2808) );
XNOR2_X2 inst_594 ( .A(net_16982), .ZN(net_16093), .B(net_643) );
INV_X4 inst_13848 ( .ZN(net_11757), .A(net_7470) );
NOR2_X2 inst_4435 ( .ZN(net_9890), .A1(net_2646), .A2(net_2592) );
OAI21_X2 inst_2175 ( .ZN(net_8878), .A(net_8854), .B1(net_4775), .B2(net_4121) );
OAI21_X2 inst_1632 ( .ZN(net_16018), .A(net_15684), .B2(net_15442), .B1(net_3158) );
NOR2_X2 inst_4241 ( .ZN(net_20341), .A2(net_6552), .A1(net_4034) );
CLKBUF_X2 inst_22052 ( .A(net_21730), .Z(net_21924) );
SDFF_X2 inst_925 ( .Q(net_21138), .D(net_16528), .SE(net_263), .CK(net_22409), .SI(x3701) );
CLKBUF_X2 inst_22822 ( .A(net_22693), .Z(net_22694) );
OAI21_X2 inst_2193 ( .ZN(net_19894), .B2(net_6365), .B1(net_5369), .A(net_1244) );
NAND2_X2 inst_10302 ( .ZN(net_10210), .A1(net_7870), .A2(net_6197) );
NAND2_X2 inst_8734 ( .ZN(net_16049), .A2(net_15765), .A1(net_15086) );
NAND2_X2 inst_9793 ( .ZN(net_11075), .A1(net_10759), .A2(net_9710) );
NAND3_X2 inst_6147 ( .ZN(net_13683), .A2(net_12313), .A3(net_7830), .A1(net_7073) );
NAND2_X2 inst_8999 ( .ZN(net_19384), .A1(net_14296), .A2(net_14295) );
SDFF_X2 inst_881 ( .Q(net_21179), .SI(net_16962), .SE(net_125), .CK(net_21394), .D(x4545) );
OAI21_X2 inst_1536 ( .A(net_18582), .ZN(net_17944), .B1(net_17786), .B2(net_17685) );
NOR2_X2 inst_3876 ( .ZN(net_9358), .A1(net_9357), .A2(net_8071) );
NAND2_X2 inst_11300 ( .ZN(net_8152), .A2(net_3753), .A1(net_1233) );
NOR2_X2 inst_3848 ( .A2(net_12795), .ZN(net_9557), .A1(net_7725) );
AOI21_X2 inst_20298 ( .ZN(net_16123), .B2(net_15725), .B1(net_15681), .A(net_14489) );
NAND2_X4 inst_7001 ( .A2(net_20454), .A1(net_20453), .ZN(net_17194) );
INV_X8 inst_12175 ( .A(net_18211), .ZN(net_18182) );
INV_X2 inst_19034 ( .ZN(net_4861), .A(net_4860) );
NOR2_X2 inst_3706 ( .ZN(net_19607), .A2(net_9163), .A1(net_8197) );
INV_X4 inst_13979 ( .ZN(net_7882), .A(net_6620) );
NAND2_X2 inst_9219 ( .ZN(net_12983), .A1(net_12310), .A2(net_10322) );
CLKBUF_X2 inst_22534 ( .A(net_21425), .Z(net_22406) );
XNOR2_X2 inst_247 ( .ZN(net_17316), .A(net_17310), .B(net_16097) );
XNOR2_X2 inst_403 ( .B(net_21160), .A(net_16677), .ZN(net_16676) );
NAND3_X2 inst_6089 ( .ZN(net_13945), .A1(net_12741), .A3(net_10250), .A2(net_9224) );
NAND2_X4 inst_7066 ( .A2(net_20864), .A1(net_19174), .ZN(net_16240) );
INV_X4 inst_17727 ( .A(net_3745), .ZN(net_2375) );
INV_X4 inst_15969 ( .ZN(net_2420), .A(net_1233) );
INV_X4 inst_15883 ( .ZN(net_3446), .A(net_621) );
DFF_X2 inst_19772 ( .QN(net_20851), .D(net_18074), .CK(net_22639) );
NOR2_X2 inst_3446 ( .A1(net_15924), .ZN(net_14951), .A2(net_13606) );
NOR3_X2 inst_2728 ( .ZN(net_13245), .A3(net_11754), .A1(net_10529), .A2(net_6141) );
INV_X4 inst_16559 ( .ZN(net_10504), .A(net_9080) );
CLKBUF_X2 inst_22735 ( .A(net_22606), .Z(net_22607) );
OAI21_X2 inst_1588 ( .ZN(net_19365), .A(net_16259), .B2(net_15942), .B1(net_10612) );
INV_X2 inst_18790 ( .A(net_8590), .ZN(net_7481) );
INV_X4 inst_18310 ( .A(net_20506), .ZN(net_20505) );
AND2_X4 inst_21220 ( .ZN(net_6744), .A2(net_5545), .A1(net_3368) );
AOI21_X4 inst_20183 ( .B1(net_19277), .ZN(net_15332), .B2(net_14493), .A(net_6397) );
NAND2_X2 inst_8002 ( .ZN(net_18307), .A1(net_18252), .A2(net_18247) );
INV_X4 inst_14484 ( .A(net_6550), .ZN(net_4868) );
NAND2_X2 inst_10996 ( .ZN(net_4919), .A1(net_4918), .A2(net_4910) );
OAI211_X2 inst_2516 ( .ZN(net_12022), .C1(net_10610), .C2(net_10114), .B(net_6210), .A(net_5811) );
INV_X4 inst_13901 ( .A(net_9374), .ZN(net_8573) );
OAI21_X4 inst_1506 ( .ZN(net_9975), .B1(net_7031), .B2(net_5681), .A(net_117) );
NAND2_X2 inst_9567 ( .A2(net_12436), .A1(net_11468), .ZN(net_10964) );
NAND2_X2 inst_9494 ( .ZN(net_19571), .A1(net_11441), .A2(net_9399) );
INV_X4 inst_15515 ( .ZN(net_11432), .A(net_7193) );
NOR2_X2 inst_3785 ( .ZN(net_14418), .A1(net_11549), .A2(net_10210) );
NAND3_X2 inst_6058 ( .A3(net_20360), .A1(net_20359), .ZN(net_14206), .A2(net_10217) );
NAND2_X4 inst_7541 ( .ZN(net_4908), .A1(net_1876), .A2(net_1848) );
NAND2_X2 inst_10455 ( .ZN(net_7030), .A2(net_3672), .A1(net_3447) );
INV_X4 inst_16987 ( .ZN(net_9080), .A(net_1019) );
INV_X4 inst_15800 ( .A(net_15969), .ZN(net_1890) );
INV_X2 inst_19416 ( .ZN(net_1907), .A(net_1201) );
NAND3_X2 inst_5678 ( .A2(net_20658), .A1(net_20657), .A3(net_20379), .ZN(net_16333) );
INV_X2 inst_19706 ( .A(net_20574), .ZN(net_20573) );
CLKBUF_X2 inst_21414 ( .A(net_21285), .Z(net_21286) );
NAND2_X4 inst_7454 ( .A2(net_20568), .ZN(net_3765), .A1(net_2522) );
OAI21_X4 inst_1361 ( .B2(net_20047), .B1(net_20046), .ZN(net_19884), .A(net_18070) );
CLKBUF_X2 inst_21544 ( .A(net_21415), .Z(net_21416) );
NOR2_X2 inst_3401 ( .ZN(net_15847), .A2(net_15642), .A1(net_14674) );
INV_X4 inst_12949 ( .ZN(net_17104), .A(net_17103) );
INV_X4 inst_13105 ( .ZN(net_19732), .A(net_15604) );
CLKBUF_X2 inst_21750 ( .A(net_21621), .Z(net_21622) );
INV_X4 inst_12688 ( .ZN(net_17693), .A(net_17692) );
NAND2_X4 inst_7525 ( .ZN(net_2647), .A1(net_1638), .A2(net_1264) );
NAND2_X2 inst_11916 ( .ZN(net_7091), .A2(net_1636), .A1(net_1547) );
INV_X8 inst_12439 ( .A(net_20495), .ZN(net_20478) );
OAI21_X2 inst_2208 ( .ZN(net_8534), .A(net_8533), .B2(net_6960), .B1(net_3945) );
NOR2_X2 inst_4463 ( .A1(net_9276), .ZN(net_4536), .A2(net_2740) );
INV_X2 inst_18410 ( .ZN(net_16216), .A(net_16161) );
NAND3_X4 inst_5598 ( .ZN(net_19079), .A3(net_11852), .A2(net_7961), .A1(net_6793) );
NAND2_X2 inst_8789 ( .ZN(net_15748), .A1(net_15666), .A2(net_15388) );
NAND2_X2 inst_10698 ( .ZN(net_13880), .A1(net_7850), .A2(net_6052) );
NAND2_X2 inst_8975 ( .ZN(net_14514), .A1(net_14363), .A2(net_12843) );
CLKBUF_X2 inst_21850 ( .A(net_21721), .Z(net_21722) );
NAND2_X2 inst_7873 ( .ZN(net_18541), .A2(net_18485), .A1(net_18456) );
OAI21_X2 inst_2174 ( .A(net_11771), .ZN(net_8899), .B2(net_5653), .B1(net_2364) );
NAND3_X2 inst_6721 ( .ZN(net_7767), .A1(net_6513), .A3(net_6512), .A2(net_2419) );
NAND2_X2 inst_10779 ( .A1(net_7968), .ZN(net_5603), .A2(net_5602) );
CLKBUF_X2 inst_22416 ( .A(net_21286), .Z(net_22288) );
INV_X4 inst_13089 ( .ZN(net_18875), .A(net_15873) );
NAND2_X4 inst_7702 ( .A2(net_525), .ZN(net_372), .A1(net_160) );
XOR2_X2 inst_14 ( .B(net_21127), .Z(net_17027), .A(net_17025) );
NAND2_X2 inst_7886 ( .ZN(net_18512), .A2(net_18436), .A1(net_17918) );
NAND2_X2 inst_9366 ( .ZN(net_12123), .A2(net_12122), .A1(net_9415) );
NAND2_X4 inst_7172 ( .ZN(net_11425), .A2(net_9397), .A1(net_4783) );
CLKBUF_X2 inst_22716 ( .A(net_22587), .Z(net_22588) );
AND2_X4 inst_21157 ( .ZN(net_19817), .A1(net_14301), .A2(net_12732) );
INV_X4 inst_15774 ( .ZN(net_1918), .A(net_1917) );
INV_X4 inst_15085 ( .ZN(net_4736), .A(net_3260) );
CLKBUF_X2 inst_22646 ( .A(net_22517), .Z(net_22518) );
OAI21_X2 inst_2325 ( .ZN(net_5544), .B1(net_2198), .A(net_1156), .B2(net_1089) );
NAND2_X2 inst_12068 ( .ZN(net_823), .A2(net_252), .A1(net_113) );
INV_X8 inst_12354 ( .ZN(net_1735), .A(net_256) );
OR2_X4 inst_1074 ( .A2(net_11282), .ZN(net_8315), .A1(net_2212) );
NAND2_X2 inst_7983 ( .ZN(net_18334), .A2(net_18328), .A1(net_17649) );
NAND2_X4 inst_7375 ( .ZN(net_5505), .A2(net_4315), .A1(net_154) );
NAND2_X2 inst_10149 ( .A1(net_12363), .ZN(net_8292), .A2(net_6193) );
CLKBUF_X2 inst_21905 ( .A(net_21776), .Z(net_21777) );
AOI21_X2 inst_20911 ( .A(net_10096), .ZN(net_7344), .B2(net_7343), .B1(net_2608) );
INV_X2 inst_19293 ( .ZN(net_2823), .A(net_2822) );
INV_X4 inst_14944 ( .A(net_5786), .ZN(net_3520) );
OAI21_X2 inst_1602 ( .B1(net_16743), .ZN(net_16157), .A(net_15796), .B2(net_15767) );
NAND2_X2 inst_9883 ( .A2(net_13226), .A1(net_10580), .ZN(net_9427) );
NAND2_X2 inst_11100 ( .A1(net_20551), .ZN(net_11656), .A2(net_4339) );
SDFF_X2 inst_969 ( .QN(net_21038), .D(net_716), .SE(net_263), .CK(net_21969), .SI(x2357) );
CLKBUF_X2 inst_21588 ( .A(net_21459), .Z(net_21460) );
INV_X4 inst_14569 ( .A(net_11841), .ZN(net_4552) );
INV_X2 inst_18465 ( .A(net_13820), .ZN(net_12732) );
NAND3_X2 inst_6463 ( .ZN(net_11364), .A3(net_11363), .A2(net_9467), .A1(net_3140) );
NAND2_X2 inst_8567 ( .A1(net_21206), .ZN(net_16741), .A2(net_16543) );
INV_X4 inst_13081 ( .ZN(net_16114), .A(net_16025) );
OAI211_X2 inst_2528 ( .ZN(net_11752), .C1(net_11751), .C2(net_10429), .B(net_10156), .A(net_9606) );
INV_X4 inst_12487 ( .ZN(net_18721), .A(net_18696) );
INV_X4 inst_17534 ( .ZN(net_15827), .A(net_15362) );
NOR2_X2 inst_4917 ( .ZN(net_2564), .A2(net_1886), .A1(net_1712) );
NAND2_X2 inst_9749 ( .A2(net_10609), .ZN(net_10076), .A1(net_5216) );
NAND2_X4 inst_7049 ( .A2(net_19162), .A1(net_19161), .ZN(net_16485) );
NOR2_X2 inst_4227 ( .ZN(net_7845), .A2(net_6632), .A1(net_573) );
CLKBUF_X2 inst_22927 ( .A(net_22768), .Z(net_22799) );
NAND2_X4 inst_6840 ( .A2(net_20033), .A1(net_20032), .ZN(net_18703) );
NAND2_X2 inst_9800 ( .ZN(net_12934), .A1(net_10467), .A2(net_9702) );
INV_X4 inst_16599 ( .ZN(net_1492), .A(net_1135) );
NAND2_X2 inst_10824 ( .ZN(net_11598), .A2(net_5900), .A1(net_5498) );
INV_X2 inst_18478 ( .ZN(net_12623), .A(net_12622) );
INV_X8 inst_12290 ( .ZN(net_9478), .A(net_1085) );
OAI21_X2 inst_2343 ( .B2(net_19417), .B1(net_9571), .ZN(net_4399), .A(net_1717) );
OAI211_X2 inst_2538 ( .B(net_13460), .ZN(net_11184), .C1(net_8877), .A(net_8003), .C2(net_6440) );
NAND2_X2 inst_11500 ( .ZN(net_3962), .A2(net_2965), .A1(net_2668) );
NAND3_X2 inst_5708 ( .A3(net_20813), .A1(net_20812), .ZN(net_19253), .A2(net_15709) );
INV_X8 inst_12303 ( .A(net_1981), .ZN(net_1364) );
INV_X4 inst_16980 ( .ZN(net_3134), .A(net_2292) );
INV_X8 inst_12427 ( .A(net_20951), .ZN(net_766) );
NAND2_X2 inst_11929 ( .A1(net_4394), .ZN(net_2899), .A2(net_225) );
INV_X4 inst_15599 ( .ZN(net_4187), .A(net_2217) );
CLKBUF_X2 inst_22271 ( .A(net_22142), .Z(net_22143) );
INV_X4 inst_12584 ( .ZN(net_19902), .A(net_18143) );
NOR2_X2 inst_4945 ( .A1(net_19426), .ZN(net_3091), .A2(net_61) );
NAND4_X4 inst_5169 ( .A4(net_18928), .A1(net_18927), .ZN(net_17109), .A2(net_16193), .A3(net_11663) );
NAND2_X2 inst_8782 ( .A1(net_21220), .ZN(net_15797), .A2(net_15257) );
INV_X4 inst_15497 ( .A(net_7850), .ZN(net_4348) );
NAND2_X2 inst_9982 ( .A2(net_10604), .ZN(net_8856), .A1(net_5998) );
AOI211_X2 inst_21043 ( .ZN(net_13195), .C1(net_13194), .A(net_12538), .B(net_10339), .C2(net_9435) );
INV_X4 inst_17519 ( .A(net_1848), .ZN(net_404) );
NAND2_X2 inst_10970 ( .A1(net_9571), .ZN(net_4986), .A2(net_4902) );
INV_X4 inst_13908 ( .A(net_7016), .ZN(net_7015) );
OR2_X4 inst_1089 ( .ZN(net_5218), .A2(net_4673), .A1(net_1076) );
NAND2_X2 inst_9720 ( .ZN(net_10159), .A1(net_10158), .A2(net_7706) );
INV_X4 inst_17198 ( .ZN(net_3729), .A(net_308) );
NAND3_X2 inst_6537 ( .A2(net_12245), .A3(net_10643), .ZN(net_10579), .A1(net_4019) );
NAND2_X2 inst_10251 ( .ZN(net_9547), .A1(net_8007), .A2(net_8006) );
NAND3_X2 inst_6430 ( .ZN(net_11914), .A3(net_10343), .A1(net_7056), .A2(net_7002) );
INV_X4 inst_17586 ( .ZN(net_523), .A(net_337) );
NAND2_X4 inst_6932 ( .A2(net_19855), .A1(net_19854), .ZN(net_17642) );
NAND4_X2 inst_5367 ( .A1(net_19975), .ZN(net_15238), .A4(net_13363), .A3(net_12061), .A2(net_11502) );
NAND2_X2 inst_9092 ( .ZN(net_13791), .A1(net_12697), .A2(net_12221) );
CLKBUF_X2 inst_22436 ( .A(net_22307), .Z(net_22308) );
DFF_X1 inst_19809 ( .QN(net_21185), .D(net_18024), .CK(net_22341) );
INV_X4 inst_12614 ( .ZN(net_20420), .A(net_18072) );
INV_X4 inst_17127 ( .ZN(net_1241), .A(net_771) );
OAI21_X2 inst_2046 ( .B2(net_11629), .ZN(net_11156), .B1(net_10447), .A(net_2707) );
AOI21_X2 inst_20316 ( .ZN(net_15964), .B1(net_15574), .B2(net_14453), .A(net_1402) );
NAND3_X2 inst_6041 ( .ZN(net_14313), .A2(net_14312), .A3(net_13199), .A1(net_9495) );
NAND2_X2 inst_12021 ( .ZN(net_1236), .A2(net_596), .A1(net_255) );
NOR2_X2 inst_4129 ( .ZN(net_20603), .A1(net_10550), .A2(net_6962) );
NAND2_X4 inst_7505 ( .ZN(net_2620), .A1(net_2253), .A2(net_2252) );
NAND2_X2 inst_11632 ( .ZN(net_2526), .A2(net_253), .A1(x4706) );
NAND3_X2 inst_6340 ( .A3(net_20319), .ZN(net_12267), .A1(net_12266), .A2(net_11816) );
INV_X2 inst_18453 ( .ZN(net_13428), .A(net_13427) );
CLKBUF_X2 inst_22088 ( .A(net_21959), .Z(net_21960) );
INV_X4 inst_16410 ( .ZN(net_4863), .A(net_3491) );
INV_X4 inst_14176 ( .ZN(net_9348), .A(net_5992) );
INV_X4 inst_15953 ( .ZN(net_2993), .A(net_1338) );
CLKBUF_X2 inst_22551 ( .A(net_21552), .Z(net_22423) );
INV_X4 inst_14835 ( .ZN(net_5520), .A(net_3163) );
INV_X2 inst_19121 ( .ZN(net_4417), .A(net_4416) );
INV_X4 inst_13783 ( .ZN(net_12454), .A(net_7572) );
INV_X4 inst_14224 ( .ZN(net_5841), .A(net_5840) );
INV_X4 inst_15833 ( .ZN(net_3614), .A(net_3287) );
NAND3_X2 inst_6533 ( .ZN(net_10585), .A3(net_7239), .A2(net_6214), .A1(net_5739) );
INV_X4 inst_17510 ( .ZN(net_1798), .A(net_894) );
NOR2_X2 inst_3524 ( .ZN(net_19781), .A1(net_11578), .A2(net_8750) );
NOR2_X2 inst_4479 ( .ZN(net_6585), .A2(net_2705), .A1(net_1438) );
INV_X8 inst_12333 ( .ZN(net_1328), .A(net_511) );
NAND2_X2 inst_7719 ( .ZN(net_18841), .A1(net_18840), .A2(net_18827) );
NAND2_X2 inst_10882 ( .ZN(net_6654), .A2(net_3912), .A1(net_2996) );
NOR2_X2 inst_4782 ( .ZN(net_11217), .A1(net_7780), .A2(net_1973) );
INV_X4 inst_15283 ( .ZN(net_4246), .A(net_2352) );
OAI221_X2 inst_1347 ( .C2(net_13196), .ZN(net_12767), .B2(net_12093), .C1(net_10470), .A(net_8962), .B1(net_8674) );
XNOR2_X2 inst_509 ( .ZN(net_7649), .A(net_7648), .B(net_3348) );
NAND2_X2 inst_11073 ( .ZN(net_8085), .A1(net_4481), .A2(net_3788) );
NOR3_X2 inst_2687 ( .ZN(net_14355), .A2(net_14254), .A1(net_12608), .A3(net_8848) );
NAND2_X2 inst_11473 ( .A2(net_5248), .ZN(net_3139), .A1(net_2467) );
NAND2_X2 inst_11775 ( .ZN(net_2046), .A1(net_1433), .A2(net_1252) );
INV_X2 inst_19545 ( .ZN(net_1256), .A(net_941) );
NAND2_X4 inst_7139 ( .ZN(net_13220), .A1(net_9806), .A2(net_4751) );
NOR3_X4 inst_2622 ( .A3(net_19246), .A1(net_19245), .ZN(net_18897), .A2(net_6532) );
XNOR2_X2 inst_153 ( .ZN(net_17989), .A(net_17878), .B(net_16986) );
NOR2_X2 inst_4856 ( .A1(net_6325), .ZN(net_3210), .A2(net_1812) );
NAND2_X2 inst_9751 ( .ZN(net_10055), .A1(net_10054), .A2(net_6972) );
OAI21_X4 inst_1459 ( .ZN(net_20737), .B2(net_20308), .B1(net_20307), .A(net_15077) );
NOR2_X2 inst_4094 ( .A1(net_9349), .ZN(net_7240), .A2(net_7239) );
NAND2_X2 inst_10483 ( .A1(net_10445), .ZN(net_8876), .A2(net_6948) );
XNOR2_X2 inst_209 ( .ZN(net_17570), .B(net_17380), .A(net_17274) );
NAND3_X2 inst_6068 ( .ZN(net_14128), .A3(net_10555), .A1(net_8866), .A2(net_7195) );
CLKBUF_X2 inst_22441 ( .A(net_22312), .Z(net_22313) );
OAI21_X2 inst_1781 ( .B2(net_19942), .B1(net_19941), .ZN(net_14664), .A(net_14663) );
NAND3_X2 inst_6365 ( .ZN(net_20663), .A3(net_12903), .A1(net_6338), .A2(net_2990) );
INV_X4 inst_16304 ( .A(net_10022), .ZN(net_8751) );
AOI21_X4 inst_20232 ( .ZN(net_13137), .B1(net_12497), .A(net_11045), .B2(net_9833) );
NOR3_X2 inst_2769 ( .A2(net_9506), .ZN(net_9251), .A3(net_9250), .A1(net_2944) );
AOI22_X2 inst_19990 ( .ZN(net_14801), .A2(net_13435), .B2(net_11294), .B1(net_5374), .A1(net_902) );
INV_X2 inst_19259 ( .A(net_15099), .ZN(net_3180) );
INV_X4 inst_17794 ( .ZN(net_3456), .A(net_525) );
INV_X4 inst_17625 ( .ZN(net_14678), .A(net_8596) );
NAND3_X2 inst_6230 ( .ZN(net_20204), .A3(net_12122), .A1(net_8589), .A2(net_6102) );
NAND2_X2 inst_11353 ( .ZN(net_3633), .A2(net_3632), .A1(net_3592) );
INV_X4 inst_15797 ( .ZN(net_1893), .A(net_1892) );
NOR2_X2 inst_3982 ( .ZN(net_8380), .A1(net_7854), .A2(net_6299) );
INV_X2 inst_19421 ( .ZN(net_1839), .A(net_1838) );
NAND3_X2 inst_6482 ( .ZN(net_19797), .A3(net_8988), .A1(net_8178), .A2(net_3265) );
NOR2_X4 inst_3215 ( .ZN(net_3874), .A1(net_3101), .A2(net_2327) );
INV_X4 inst_14273 ( .ZN(net_6260), .A(net_5667) );
INV_X4 inst_18231 ( .A(net_20848), .ZN(net_16394) );
NAND3_X2 inst_5810 ( .A3(net_20824), .A1(net_20823), .ZN(net_15652), .A2(net_9123) );
NAND2_X2 inst_8462 ( .ZN(net_20088), .A1(net_19449), .A2(net_17239) );
CLKBUF_X2 inst_22889 ( .A(net_22760), .Z(net_22761) );
NOR2_X2 inst_4167 ( .ZN(net_6864), .A1(net_6863), .A2(net_5199) );
NAND2_X2 inst_9204 ( .A1(net_14186), .ZN(net_13074), .A2(net_10283) );
CLKBUF_X2 inst_21583 ( .A(net_21454), .Z(net_21455) );
NOR2_X2 inst_4374 ( .ZN(net_6652), .A2(net_5413), .A1(net_1279) );
OAI21_X2 inst_1995 ( .ZN(net_20675), .B1(net_11741), .B2(net_7972), .A(net_7193) );
INV_X4 inst_15031 ( .ZN(net_14551), .A(net_3364) );
AND2_X4 inst_21229 ( .ZN(net_4582), .A1(net_4581), .A2(net_4580) );
NAND2_X2 inst_9145 ( .ZN(net_14847), .A2(net_12241), .A1(net_4700) );
INV_X4 inst_17894 ( .A(net_1339), .ZN(net_1080) );
NAND2_X4 inst_7405 ( .ZN(net_9956), .A1(net_3990), .A2(net_3989) );
CLKBUF_X2 inst_22687 ( .A(net_22558), .Z(net_22559) );
NOR2_X2 inst_3367 ( .ZN(net_16868), .A2(net_16867), .A1(net_7293) );
INV_X4 inst_12736 ( .A(net_17952), .ZN(net_17926) );
XNOR2_X2 inst_568 ( .B(net_16839), .ZN(net_642), .A(net_641) );
XNOR2_X2 inst_523 ( .B(net_5616), .ZN(net_4239), .A(net_1883) );
OAI21_X4 inst_1483 ( .B2(net_19323), .B1(net_19322), .ZN(net_14205), .A(net_7170) );
INV_X4 inst_15445 ( .A(net_16051), .ZN(net_3296) );
INV_X4 inst_17843 ( .ZN(net_1347), .A(net_318) );
NAND2_X2 inst_10202 ( .A1(net_10015), .ZN(net_8123), .A2(net_8122) );
OAI21_X4 inst_1492 ( .ZN(net_12540), .B2(net_10337), .B1(net_9227), .A(net_749) );
INV_X4 inst_18328 ( .ZN(net_20551), .A(net_20548) );
DFF_X1 inst_19810 ( .Q(net_20912), .D(net_18001), .CK(net_21305) );
NOR2_X2 inst_4234 ( .ZN(net_6576), .A1(net_6575), .A2(net_6574) );
NAND3_X2 inst_6722 ( .ZN(net_6508), .A2(net_6492), .A1(net_5232), .A3(net_5081) );
NAND2_X2 inst_11982 ( .ZN(net_1287), .A2(net_659), .A1(net_74) );
CLKBUF_X2 inst_21387 ( .A(net_21258), .Z(net_21259) );
INV_X2 inst_19271 ( .ZN(net_3032), .A(net_3031) );
INV_X2 inst_19061 ( .ZN(net_4693), .A(net_4692) );
INV_X4 inst_16694 ( .ZN(net_10098), .A(net_761) );
NOR2_X4 inst_2898 ( .ZN(net_10872), .A1(net_7493), .A2(net_6877) );
AOI21_X2 inst_20506 ( .ZN(net_14635), .B1(net_14634), .B2(net_12080), .A(net_7689) );
NAND2_X2 inst_8875 ( .A1(net_15607), .ZN(net_15249), .A2(net_14191) );
NAND2_X2 inst_10280 ( .ZN(net_7951), .A2(net_6093), .A1(net_4900) );
CLKBUF_X2 inst_22690 ( .A(net_22416), .Z(net_22562) );
INV_X4 inst_17162 ( .ZN(net_9322), .A(net_308) );
OAI21_X4 inst_1368 ( .B2(net_19444), .ZN(net_17504), .A(net_16955), .B1(net_16945) );
INV_X4 inst_13708 ( .ZN(net_9391), .A(net_7861) );
INV_X4 inst_15665 ( .ZN(net_8311), .A(net_5818) );
NAND2_X4 inst_7282 ( .A1(net_19399), .ZN(net_9321), .A2(net_420) );
CLKBUF_X2 inst_22732 ( .A(net_22603), .Z(net_22604) );
OAI21_X2 inst_2088 ( .ZN(net_10353), .B2(net_6312), .B1(net_5941), .A(net_761) );
NAND3_X2 inst_6775 ( .ZN(net_4703), .A1(net_4702), .A2(net_4701), .A3(net_2439) );
INV_X4 inst_15199 ( .A(net_4136), .ZN(net_2915) );
INV_X2 inst_18565 ( .A(net_12417), .ZN(net_10776) );
INV_X4 inst_17475 ( .ZN(net_3242), .A(net_874) );
INV_X4 inst_16026 ( .ZN(net_9301), .A(net_2974) );
NAND3_X2 inst_6673 ( .ZN(net_7760), .A3(net_5940), .A1(net_5490), .A2(net_2826) );
CLKBUF_X2 inst_22659 ( .A(net_22530), .Z(net_22531) );
OAI21_X4 inst_1379 ( .A(net_20968), .B2(net_20139), .B1(net_20138), .ZN(net_19135) );
AOI211_X2 inst_21021 ( .ZN(net_14997), .A(net_14996), .C2(net_12956), .B(net_12068), .C1(net_3985) );
INV_X8 inst_12326 ( .A(net_973), .ZN(net_898) );
NAND2_X2 inst_9582 ( .ZN(net_10926), .A2(net_9150), .A1(net_8697) );
INV_X4 inst_15739 ( .ZN(net_8700), .A(net_5387) );
NAND2_X4 inst_7691 ( .ZN(net_867), .A2(net_317), .A1(net_205) );
INV_X8 inst_12217 ( .ZN(net_9397), .A(net_6067) );
AOI21_X2 inst_20330 ( .B1(net_20706), .ZN(net_20179), .A(net_10269), .B2(net_1171) );
NAND2_X2 inst_9221 ( .ZN(net_18977), .A2(net_12972), .A1(net_2977) );
INV_X4 inst_15582 ( .A(net_11526), .ZN(net_11236) );
NAND3_X2 inst_6131 ( .ZN(net_13740), .A1(net_12887), .A2(net_11081), .A3(net_10940) );
INV_X4 inst_13643 ( .ZN(net_9678), .A(net_6850) );
CLKBUF_X2 inst_22651 ( .A(net_21551), .Z(net_22523) );
NAND3_X2 inst_5796 ( .ZN(net_15720), .A2(net_15114), .A1(net_15070), .A3(net_14561) );
INV_X4 inst_14229 ( .ZN(net_5831), .A(net_5830) );
CLKBUF_X2 inst_22882 ( .A(net_22753), .Z(net_22754) );
NAND2_X2 inst_9571 ( .ZN(net_10959), .A2(net_10958), .A1(net_10022) );
INV_X4 inst_14654 ( .ZN(net_4367), .A(net_4366) );
INV_X4 inst_14924 ( .ZN(net_19487), .A(net_4930) );
XNOR2_X2 inst_583 ( .B(net_678), .ZN(net_592), .A(net_591) );
OAI21_X2 inst_1904 ( .A(net_13437), .ZN(net_13136), .B2(net_9326), .B1(net_5870) );
INV_X4 inst_13970 ( .A(net_8945), .ZN(net_6681) );
NAND2_X2 inst_10732 ( .ZN(net_7355), .A1(net_5599), .A2(net_4669) );
INV_X4 inst_18156 ( .A(net_20885), .ZN(net_106) );
NOR2_X2 inst_4325 ( .ZN(net_5844), .A1(net_2058), .A2(net_1806) );
NAND2_X2 inst_10932 ( .ZN(net_7333), .A2(net_5210), .A1(net_1091) );
INV_X4 inst_14146 ( .ZN(net_11418), .A(net_7902) );
NAND2_X2 inst_10441 ( .ZN(net_7188), .A1(net_7129), .A2(net_5258) );
NAND2_X4 inst_6913 ( .A2(net_20244), .A1(net_20243), .ZN(net_17859) );
AOI21_X2 inst_20897 ( .ZN(net_7739), .A(net_6936), .B1(net_3414), .B2(net_2714) );
NAND3_X2 inst_6788 ( .ZN(net_8954), .A3(net_3836), .A2(net_3789), .A1(net_2245) );
INV_X4 inst_17583 ( .ZN(net_6968), .A(net_3682) );
INV_X4 inst_14346 ( .ZN(net_8408), .A(net_5336) );
NAND2_X2 inst_7709 ( .A1(net_20007), .ZN(net_18857), .A2(net_17038) );
NOR2_X2 inst_4863 ( .ZN(net_4169), .A1(net_2994), .A2(net_1113) );
NOR2_X2 inst_4910 ( .ZN(net_1938), .A2(net_1937), .A1(net_225) );
INV_X4 inst_12513 ( .A(net_18633), .ZN(net_18620) );
INV_X4 inst_14667 ( .ZN(net_18864), .A(net_18025) );
NAND2_X2 inst_12113 ( .A1(net_513), .A2(net_322), .ZN(net_237) );
INV_X4 inst_14985 ( .ZN(net_20031), .A(net_3405) );
AOI21_X2 inst_20383 ( .ZN(net_15505), .B1(net_15334), .B2(net_14528), .A(net_11381) );
NAND2_X2 inst_9811 ( .ZN(net_9677), .A1(net_9676), .A2(net_9675) );
INV_X4 inst_14504 ( .ZN(net_6507), .A(net_5312) );
INV_X4 inst_17523 ( .A(net_606), .ZN(net_400) );
NAND2_X2 inst_8693 ( .A1(net_21236), .ZN(net_16361), .A2(net_16201) );
NAND3_X2 inst_6025 ( .ZN(net_14374), .A3(net_14316), .A2(net_9479), .A1(net_8603) );
INV_X4 inst_17330 ( .A(net_10714), .ZN(net_7801) );
OAI21_X2 inst_2289 ( .ZN(net_6522), .A(net_6521), .B2(net_6520), .B1(net_303) );
CLKBUF_X2 inst_22084 ( .A(net_21542), .Z(net_21956) );
INV_X2 inst_18850 ( .ZN(net_8765), .A(net_6608) );
AND2_X4 inst_21247 ( .ZN(net_9250), .A2(net_2118), .A1(net_143) );
INV_X2 inst_19277 ( .A(net_3758), .ZN(net_2969) );
NOR3_X2 inst_2750 ( .ZN(net_12263), .A2(net_12262), .A1(net_9034), .A3(net_5126) );
CLKBUF_X2 inst_21923 ( .A(net_21794), .Z(net_21795) );
OAI21_X4 inst_1467 ( .A(net_20889), .ZN(net_20164), .B2(net_12901), .B1(net_11429) );
NAND3_X2 inst_5800 ( .ZN(net_19871), .A1(net_15332), .A2(net_15116), .A3(net_14574) );
CLKBUF_X2 inst_22016 ( .A(net_21887), .Z(net_21888) );
DFF_X1 inst_19876 ( .D(net_17026), .CK(net_21331), .Q(x151) );
INV_X4 inst_14313 ( .ZN(net_6766), .A(net_5700) );
NAND3_X2 inst_5772 ( .ZN(net_15894), .A2(net_15402), .A3(net_15373), .A1(net_11514) );
NAND2_X2 inst_10258 ( .ZN(net_13580), .A1(net_11466), .A2(net_7995) );
CLKBUF_X2 inst_21686 ( .A(net_21557), .Z(net_21558) );
NAND2_X2 inst_10803 ( .A1(net_6207), .ZN(net_5546), .A2(net_5545) );
INV_X4 inst_14102 ( .ZN(net_10598), .A(net_7947) );
AND2_X2 inst_21331 ( .A2(net_11253), .A1(net_5486), .ZN(net_5191) );
NAND3_X2 inst_6317 ( .ZN(net_12567), .A2(net_12566), .A1(net_11808), .A3(net_9115) );
INV_X4 inst_13227 ( .A(net_14825), .ZN(net_13594) );
NOR2_X4 inst_2834 ( .ZN(net_19035), .A2(net_15128), .A1(net_13342) );
INV_X4 inst_15067 ( .ZN(net_6592), .A(net_1910) );
INV_X4 inst_17653 ( .ZN(net_3542), .A(net_321) );
INV_X4 inst_16064 ( .ZN(net_7751), .A(net_1575) );
AOI21_X2 inst_20385 ( .ZN(net_15498), .B2(net_14529), .B1(net_13525), .A(net_9731) );
NAND2_X2 inst_8130 ( .A2(net_20912), .ZN(net_18044), .A1(net_16274) );
OAI21_X2 inst_1513 ( .ZN(net_18580), .B2(net_18554), .B1(net_18025), .A(net_12083) );
NAND2_X2 inst_9864 ( .ZN(net_9491), .A1(net_9490), .A2(net_6162) );
NAND2_X2 inst_11756 ( .ZN(net_6107), .A1(net_2493), .A2(net_2104) );
AND2_X2 inst_21281 ( .ZN(net_13145), .A2(net_11274), .A1(net_1070) );
NAND2_X2 inst_10916 ( .ZN(net_11759), .A1(net_5344), .A2(net_5343) );
NOR2_X2 inst_4080 ( .ZN(net_7358), .A2(net_7357), .A1(net_5600) );
NAND2_X4 inst_7667 ( .ZN(net_1284), .A2(net_258), .A1(net_92) );
NAND2_X2 inst_10846 ( .ZN(net_15567), .A1(net_9638), .A2(net_5468) );
OAI21_X2 inst_1545 ( .B1(net_20525), .ZN(net_17868), .A(net_17624), .B2(net_17623) );
INV_X4 inst_12750 ( .ZN(net_17600), .A(net_17414) );
NOR2_X4 inst_3338 ( .ZN(net_1596), .A1(net_915), .A2(net_162) );
AOI21_X2 inst_20828 ( .ZN(net_9862), .B1(net_9861), .B2(net_5977), .A(net_3483) );
AOI21_X2 inst_20972 ( .A(net_7106), .ZN(net_4668), .B1(net_4621), .B2(net_2685) );
AOI21_X2 inst_20791 ( .ZN(net_10542), .B2(net_9822), .B1(net_8710), .A(net_6838) );
XNOR2_X2 inst_406 ( .A(net_16650), .ZN(net_16649), .B(net_16648) );
NOR2_X2 inst_4579 ( .A2(net_20786), .ZN(net_5366), .A1(net_1574) );
NAND3_X2 inst_5933 ( .ZN(net_19652), .A2(net_12692), .A1(net_10359), .A3(net_10024) );
INV_X4 inst_14696 ( .ZN(net_10580), .A(net_4267) );
CLKBUF_X2 inst_22404 ( .A(net_21522), .Z(net_22276) );
INV_X4 inst_13818 ( .A(net_9625), .ZN(net_9178) );
XNOR2_X2 inst_328 ( .B(net_21112), .ZN(net_17310), .A(net_16979) );
INV_X2 inst_19446 ( .ZN(net_1624), .A(net_1623) );
INV_X2 inst_18677 ( .ZN(net_8815), .A(net_8814) );
NOR2_X2 inst_4217 ( .ZN(net_8675), .A1(net_6947), .A2(net_6632) );
NAND2_X2 inst_8496 ( .ZN(net_17227), .A2(net_16555), .A1(net_16446) );
SDFF_X2 inst_818 ( .Q(net_21169), .SI(net_17674), .SE(net_125), .CK(net_22167), .D(x4916) );
INV_X8 inst_12373 ( .ZN(net_826), .A(net_132) );
INV_X4 inst_18336 ( .A(net_20582), .ZN(net_20581) );
INV_X4 inst_18229 ( .A(net_20946), .ZN(net_75) );
NAND2_X2 inst_9902 ( .ZN(net_10884), .A1(net_10831), .A2(net_9363) );
AOI22_X2 inst_19970 ( .ZN(net_15693), .A1(net_15369), .B1(net_15202), .A2(net_15004), .B2(net_12506) );
INV_X4 inst_16959 ( .ZN(net_15343), .A(net_14153) );
NAND2_X4 inst_7561 ( .ZN(net_3162), .A1(net_1692), .A2(net_1024) );
NAND2_X2 inst_9825 ( .ZN(net_20083), .A1(net_9632), .A2(net_9631) );
NAND2_X2 inst_10172 ( .ZN(net_10310), .A1(net_8220), .A2(net_6778) );
NOR2_X4 inst_3274 ( .ZN(net_3090), .A2(net_1733), .A1(net_1348) );
INV_X4 inst_13920 ( .A(net_8758), .ZN(net_8655) );
NAND2_X2 inst_11776 ( .A1(net_3707), .A2(net_2252), .ZN(net_2040) );
INV_X4 inst_12643 ( .ZN(net_17901), .A(net_17900) );
INV_X4 inst_17011 ( .ZN(net_1661), .A(net_867) );
NAND2_X2 inst_9178 ( .ZN(net_13340), .A1(net_10930), .A2(net_10561) );
INV_X4 inst_17207 ( .ZN(net_3310), .A(net_874) );
CLKBUF_X2 inst_22369 ( .A(net_22240), .Z(net_22241) );
INV_X2 inst_19205 ( .ZN(net_5887), .A(net_4319) );
NAND2_X2 inst_10066 ( .ZN(net_8668), .A1(net_8667), .A2(net_6754) );
NAND2_X2 inst_8360 ( .ZN(net_17424), .A1(net_17422), .A2(net_17421) );
INV_X2 inst_19151 ( .A(net_7104), .ZN(net_4059) );
NAND3_X2 inst_6442 ( .ZN(net_11804), .A2(net_9335), .A1(net_8135), .A3(net_7929) );
INV_X4 inst_15622 ( .ZN(net_2748), .A(net_1671) );
CLKBUF_X2 inst_21530 ( .A(net_21401), .Z(net_21402) );
INV_X4 inst_16850 ( .ZN(net_4931), .A(net_535) );
NAND2_X4 inst_7146 ( .A2(net_19254), .ZN(net_12861), .A1(net_9709) );
INV_X4 inst_16056 ( .ZN(net_2146), .A(net_1315) );
SDFF_X2 inst_906 ( .Q(net_21232), .SI(net_16849), .SE(net_125), .CK(net_22422), .D(x6936) );
NOR2_X2 inst_4276 ( .A1(net_9109), .A2(net_6231), .ZN(net_6118) );
INV_X4 inst_17293 ( .ZN(net_2388), .A(net_258) );
NAND4_X4 inst_5222 ( .A2(net_18951), .A1(net_18950), .ZN(net_16341), .A4(net_16182), .A3(net_15736) );
AOI21_X2 inst_20882 ( .ZN(net_8268), .B1(net_7750), .A(net_6639), .B2(net_2954) );
INV_X4 inst_16478 ( .ZN(net_2219), .A(net_1207) );
NOR2_X2 inst_5098 ( .A2(net_3919), .ZN(net_797), .A1(net_86) );
INV_X4 inst_13600 ( .ZN(net_8730), .A(net_8729) );
OAI211_X2 inst_2598 ( .C2(net_6495), .ZN(net_5249), .B(net_5248), .A(net_3550), .C1(net_1047) );
OAI22_X4 inst_1248 ( .A1(net_19490), .ZN(net_14991), .A2(net_14990), .B1(net_13848), .B2(net_3666) );
DFF_X1 inst_19800 ( .D(net_18193), .CK(net_21999), .Q(x1134) );
INV_X2 inst_18626 ( .ZN(net_9549), .A(net_9548) );
AOI21_X2 inst_20779 ( .A(net_15113), .B2(net_12838), .ZN(net_10566), .B1(net_10565) );
NOR2_X2 inst_3998 ( .A1(net_8722), .ZN(net_8229), .A2(net_8228) );
INV_X4 inst_18124 ( .A(net_21240), .ZN(net_170) );
INV_X2 inst_18867 ( .ZN(net_6285), .A(net_6284) );
NAND2_X2 inst_9035 ( .ZN(net_14063), .A1(net_13651), .A2(net_11833) );
INV_X2 inst_18779 ( .ZN(net_7525), .A(net_7524) );
NOR2_X2 inst_4300 ( .ZN(net_7444), .A1(net_5950), .A2(net_5891) );
NAND2_X4 inst_7645 ( .ZN(net_1700), .A2(net_836), .A1(net_387) );
NAND2_X2 inst_12000 ( .ZN(net_6537), .A1(net_3748), .A2(net_170) );
INV_X4 inst_16221 ( .ZN(net_14500), .A(net_238) );
XNOR2_X2 inst_183 ( .A(net_17777), .ZN(net_17765), .B(net_17129) );
NAND2_X2 inst_7748 ( .ZN(net_18780), .A1(net_18731), .A2(net_18706) );
NAND3_X2 inst_6703 ( .A3(net_9073), .ZN(net_7350), .A2(net_4896), .A1(net_4327) );
NAND2_X2 inst_8471 ( .A1(net_21143), .ZN(net_17017), .A2(net_16811) );
CLKBUF_X2 inst_22819 ( .A(net_22268), .Z(net_22691) );
INV_X4 inst_15822 ( .ZN(net_5797), .A(net_1870) );
CLKBUF_X2 inst_22809 ( .A(net_22680), .Z(net_22681) );
INV_X2 inst_19467 ( .ZN(net_8488), .A(net_3908) );
INV_X4 inst_17266 ( .ZN(net_2292), .A(net_1645) );
NAND2_X2 inst_8081 ( .ZN(net_19002), .A2(net_18128), .A1(net_18096) );
CLKBUF_X2 inst_22915 ( .A(net_22786), .Z(net_22787) );
OAI21_X2 inst_1848 ( .ZN(net_14016), .B1(net_11145), .B2(net_8506), .A(net_829) );
CLKBUF_X2 inst_21735 ( .A(net_21554), .Z(net_21607) );
AOI21_X4 inst_20199 ( .B1(net_18977), .ZN(net_15049), .B2(net_15048), .A(net_9588) );
INV_X4 inst_12694 ( .ZN(net_17641), .A(net_17640) );
NOR2_X2 inst_4451 ( .ZN(net_4759), .A2(net_4758), .A1(net_4457) );
XNOR2_X2 inst_487 ( .ZN(net_9713), .B(net_9712), .A(net_5732) );
CLKBUF_X2 inst_21403 ( .A(net_21274), .Z(net_21275) );
NAND2_X2 inst_11338 ( .A1(net_5149), .A2(net_3695), .ZN(net_3684) );
INV_X4 inst_14540 ( .ZN(net_9619), .A(net_4659) );
INV_X4 inst_17810 ( .ZN(net_10087), .A(net_1470) );
NAND4_X2 inst_5315 ( .A4(net_20456), .A1(net_20455), .ZN(net_15780), .A3(net_13943), .A2(net_13799) );
INV_X4 inst_13696 ( .ZN(net_12475), .A(net_7927) );
INV_X4 inst_17376 ( .ZN(net_15077), .A(net_14308) );
OAI21_X2 inst_2133 ( .ZN(net_9991), .A(net_8457), .B1(net_6257), .B2(net_4313) );
OAI21_X2 inst_2163 ( .ZN(net_9081), .A(net_9080), .B1(net_8587), .B2(net_7250) );
INV_X4 inst_17882 ( .A(net_2274), .ZN(net_1509) );
INV_X2 inst_19011 ( .ZN(net_5012), .A(net_5011) );
NAND2_X2 inst_9947 ( .ZN(net_12129), .A1(net_8961), .A2(net_7800) );
NAND3_X2 inst_6051 ( .ZN(net_14238), .A2(net_14237), .A3(net_13561), .A1(net_12601) );
NOR2_X2 inst_4668 ( .ZN(net_9949), .A1(net_5308), .A2(net_2975) );
NAND4_X2 inst_5497 ( .ZN(net_11913), .A4(net_11912), .A2(net_5348), .A3(net_4712), .A1(net_4160) );
OAI21_X2 inst_1861 ( .ZN(net_13797), .A(net_12546), .B2(net_11125), .B1(net_10907) );
AOI21_X2 inst_20396 ( .B2(net_19705), .B1(net_19704), .ZN(net_15449), .A(net_881) );
NOR2_X2 inst_3570 ( .A2(net_12726), .ZN(net_12725), .A1(net_11909) );
NAND2_X2 inst_9133 ( .ZN(net_13518), .A1(net_13517), .A2(net_10800) );
NAND2_X4 inst_7598 ( .A1(net_1630), .ZN(net_1457), .A2(net_1456) );
NOR2_X2 inst_4835 ( .A1(net_5277), .ZN(net_3015), .A2(net_1652) );
INV_X4 inst_15050 ( .ZN(net_6459), .A(net_3321) );
NOR2_X4 inst_2857 ( .ZN(net_11818), .A2(net_8827), .A1(net_7231) );
NAND2_X2 inst_8667 ( .A1(net_21148), .A2(net_16774), .ZN(net_16473) );
INV_X4 inst_15116 ( .A(net_14186), .ZN(net_4154) );
OAI21_X2 inst_1585 ( .A(net_20944), .ZN(net_16263), .B2(net_15931), .B1(net_14189) );
NAND2_X2 inst_10754 ( .ZN(net_7499), .A2(net_5933), .A1(net_90) );
NAND2_X2 inst_11412 ( .ZN(net_4984), .A1(net_4502), .A2(net_3905) );
CLKBUF_X2 inst_22867 ( .A(net_22738), .Z(net_22739) );
OAI21_X2 inst_1873 ( .ZN(net_13704), .A(net_13703), .B1(net_13702), .B2(net_12336) );
NAND2_X2 inst_11965 ( .A1(net_2012), .ZN(net_1857), .A2(net_1787) );
NAND2_X2 inst_7854 ( .A1(net_20703), .ZN(net_18579), .A2(net_18478) );
NAND3_X2 inst_6135 ( .ZN(net_13729), .A2(net_13728), .A3(net_12311), .A1(net_11853) );
NAND2_X2 inst_11765 ( .A1(net_20859), .ZN(net_2713), .A2(net_2079) );
NAND4_X2 inst_5263 ( .A2(net_20594), .A1(net_20593), .ZN(net_19878), .A4(net_15391), .A3(net_10014) );
NOR2_X4 inst_3114 ( .ZN(net_4844), .A2(net_4025), .A1(net_4024) );
NOR2_X2 inst_3577 ( .ZN(net_12703), .A2(net_12422), .A1(net_9432) );
CLKBUF_X2 inst_22323 ( .A(net_22194), .Z(net_22195) );
NAND2_X2 inst_9451 ( .ZN(net_13705), .A1(net_11907), .A2(net_11516) );
INV_X4 inst_15035 ( .ZN(net_4588), .A(net_3359) );
NOR2_X2 inst_4754 ( .ZN(net_5373), .A2(net_3014), .A1(net_3013) );
INV_X4 inst_17711 ( .ZN(net_206), .A(net_205) );
NAND2_X2 inst_10216 ( .ZN(net_12095), .A2(net_8044), .A1(net_7975) );
NAND2_X2 inst_11554 ( .ZN(net_4949), .A2(net_2844), .A1(net_1755) );
NOR2_X2 inst_4680 ( .A1(net_10886), .ZN(net_3223), .A2(net_3217) );
NAND3_X2 inst_6589 ( .ZN(net_10041), .A3(net_9900), .A2(net_6629), .A1(net_5187) );
INV_X4 inst_16216 ( .ZN(net_2410), .A(net_2073) );
CLKBUF_X2 inst_22610 ( .A(net_22481), .Z(net_22482) );
INV_X4 inst_16952 ( .ZN(net_15198), .A(net_909) );
INV_X4 inst_14759 ( .ZN(net_5123), .A(net_4062) );
OAI21_X2 inst_1727 ( .B2(net_20610), .B1(net_20609), .ZN(net_15090), .A(net_12203) );
OAI21_X2 inst_1753 ( .B2(net_20599), .B1(net_20598), .A(net_15550), .ZN(net_14795) );
OR2_X2 inst_1166 ( .A1(net_7116), .ZN(net_7053), .A2(net_7052) );
XNOR2_X2 inst_116 ( .B(net_20761), .ZN(net_18488), .A(net_18323) );
NAND4_X2 inst_5498 ( .ZN(net_11903), .A3(net_11902), .A4(net_10354), .A2(net_5360), .A1(net_4147) );
NAND3_X2 inst_6559 ( .A3(net_20697), .ZN(net_20339), .A1(net_10567), .A2(net_6304) );
INV_X4 inst_15183 ( .ZN(net_5403), .A(net_4287) );
NAND2_X2 inst_10142 ( .A1(net_11466), .ZN(net_8313), .A2(net_8312) );
NOR2_X2 inst_4087 ( .A1(net_10709), .A2(net_9061), .ZN(net_8808) );
XNOR2_X2 inst_471 ( .ZN(net_11892), .A(net_11891), .B(net_2437) );
NAND2_X2 inst_10680 ( .ZN(net_7548), .A2(net_6153), .A1(net_5120) );
NAND2_X2 inst_12104 ( .ZN(net_460), .A2(net_459), .A1(net_334) );
NAND3_X2 inst_6557 ( .ZN(net_10509), .A3(net_6803), .A2(net_5069), .A1(net_2256) );
NAND2_X2 inst_11081 ( .ZN(net_8560), .A2(net_4448), .A1(net_90) );
INV_X4 inst_18349 ( .A(net_20791), .ZN(net_20790) );
SDFF_X2 inst_896 ( .Q(net_21230), .SI(net_16767), .SE(net_125), .CK(net_22141), .D(x7000) );
INV_X8 inst_12315 ( .ZN(net_20676), .A(net_996) );
NAND2_X2 inst_9276 ( .A1(net_13343), .ZN(net_12598), .A2(net_10814) );
INV_X4 inst_14552 ( .ZN(net_5842), .A(net_4590) );
NAND2_X2 inst_9317 ( .ZN(net_12344), .A1(net_9516), .A2(net_9170) );
INV_X4 inst_15021 ( .A(net_10930), .ZN(net_3376) );
NAND2_X4 inst_7445 ( .ZN(net_4360), .A1(net_3090), .A2(net_874) );
NAND2_X2 inst_8577 ( .ZN(net_19681), .A1(net_16727), .A2(net_16524) );
AND3_X2 inst_21133 ( .ZN(net_13686), .A3(net_12314), .A1(net_9958), .A2(net_8560) );
OAI211_X2 inst_2557 ( .C1(net_12067), .A(net_11290), .ZN(net_9948), .B(net_9947), .C2(net_7780) );
NAND2_X4 inst_7438 ( .ZN(net_3323), .A1(net_2140), .A2(net_193) );
INV_X4 inst_15639 ( .ZN(net_3339), .A(net_2130) );
NOR2_X4 inst_3319 ( .ZN(net_1119), .A1(net_958), .A2(net_459) );
INV_X4 inst_15718 ( .ZN(net_3673), .A(net_2787) );
NOR2_X2 inst_4621 ( .A1(net_5797), .ZN(net_3612), .A2(net_3318) );
NAND2_X2 inst_11519 ( .ZN(net_8494), .A2(net_2967), .A1(net_112) );
INV_X4 inst_17262 ( .ZN(net_4726), .A(net_2585) );
OAI211_X2 inst_2550 ( .ZN(net_10817), .A(net_10816), .B(net_10815), .C2(net_4640), .C1(net_3193) );
AOI22_X2 inst_19972 ( .A1(net_15747), .ZN(net_15689), .B1(net_15360), .A2(net_15050), .B2(net_12576) );
INV_X2 inst_18826 ( .ZN(net_12144), .A(net_6821) );
INV_X4 inst_14966 ( .ZN(net_4490), .A(net_2927) );
INV_X4 inst_16301 ( .ZN(net_14981), .A(net_828) );
CLKBUF_X2 inst_21855 ( .A(net_21726), .Z(net_21727) );
NAND2_X4 inst_7559 ( .A2(net_2384), .ZN(net_2033), .A1(net_1711) );
NOR2_X2 inst_4281 ( .ZN(net_10996), .A2(net_6098), .A1(net_5869) );
INV_X4 inst_16425 ( .ZN(net_1707), .A(net_1568) );
OAI21_X2 inst_2142 ( .B1(net_10898), .ZN(net_9946), .B2(net_9945), .A(net_5542) );
AOI21_X2 inst_20671 ( .ZN(net_12856), .B2(net_12804), .B1(net_9006), .A(net_7012) );
INV_X4 inst_12810 ( .A(net_17554), .ZN(net_17466) );
CLKBUF_X2 inst_22227 ( .A(net_21682), .Z(net_22099) );
INV_X4 inst_18021 ( .A(net_20933), .ZN(net_83) );
NOR2_X2 inst_5110 ( .A2(net_20868), .A1(net_2585), .ZN(net_985) );
NAND3_X2 inst_6817 ( .ZN(net_8987), .A3(net_2283), .A2(net_193), .A1(net_175) );
INV_X2 inst_19021 ( .ZN(net_9983), .A(net_6883) );
NOR2_X2 inst_4458 ( .ZN(net_4646), .A2(net_1875), .A1(net_340) );
NAND2_X2 inst_9407 ( .ZN(net_19053), .A1(net_11678), .A2(net_11677) );
INV_X4 inst_14055 ( .A(net_8066), .ZN(net_7612) );
NAND4_X4 inst_5184 ( .A4(net_19060), .A1(net_19059), .ZN(net_17103), .A3(net_14469), .A2(net_13804) );
NAND2_X2 inst_10518 ( .ZN(net_19323), .A1(net_6874), .A2(net_3417) );
CLKBUF_X2 inst_21807 ( .A(net_21270), .Z(net_21679) );
INV_X4 inst_15767 ( .A(net_14430), .ZN(net_11771) );
XNOR2_X2 inst_547 ( .B(net_9712), .ZN(net_725), .A(net_724) );
NAND2_X2 inst_9107 ( .ZN(net_20631), .A1(net_13544), .A2(net_11557) );
INV_X4 inst_16399 ( .A(net_6131), .ZN(net_4156) );
CLKBUF_X2 inst_22248 ( .A(net_22119), .Z(net_22120) );
OAI21_X2 inst_1607 ( .A(net_16368), .ZN(net_16146), .B1(net_15751), .B2(net_15528) );
NAND2_X2 inst_11847 ( .A1(net_3852), .A2(net_1970), .ZN(net_1709) );
NAND2_X2 inst_10367 ( .A1(net_9490), .ZN(net_7408), .A2(net_4572) );
NAND2_X2 inst_11623 ( .ZN(net_5639), .A1(net_4253), .A2(net_3246) );
CLKBUF_X2 inst_22065 ( .A(net_21903), .Z(net_21937) );
OAI21_X2 inst_1854 ( .ZN(net_13997), .A(net_13996), .B1(net_12939), .B2(net_11280) );
NAND2_X2 inst_9002 ( .ZN(net_14285), .A2(net_13487), .A1(net_458) );
INV_X4 inst_12676 ( .ZN(net_17737), .A(net_17736) );
INV_X2 inst_19288 ( .A(net_7395), .ZN(net_2874) );
OAI21_X2 inst_1710 ( .ZN(net_15197), .B1(net_14054), .A(net_12133), .B2(net_10753) );
NAND3_X2 inst_5922 ( .ZN(net_20846), .A3(net_13109), .A2(net_12099), .A1(net_6680) );
NAND2_X4 inst_7295 ( .ZN(net_10523), .A1(net_5573), .A2(net_2909) );
INV_X2 inst_18748 ( .ZN(net_10111), .A(net_8622) );
OAI211_X2 inst_2407 ( .ZN(net_15599), .A(net_14909), .B(net_12626), .C2(net_9304), .C1(net_5186) );
NOR2_X2 inst_4884 ( .ZN(net_4083), .A2(net_2164), .A1(net_1154) );
INV_X4 inst_13814 ( .ZN(net_7533), .A(net_7532) );
NOR2_X4 inst_3142 ( .ZN(net_3714), .A2(net_3713), .A1(net_3501) );
NAND2_X4 inst_7516 ( .ZN(net_3790), .A2(net_1295), .A1(net_938) );
AND2_X2 inst_21289 ( .ZN(net_12173), .A1(net_12172), .A2(net_12171) );
SDFF_X2 inst_753 ( .Q(net_20938), .SE(net_18837), .SI(net_18530), .D(net_11890), .CK(net_21675) );
NAND2_X2 inst_9647 ( .ZN(net_10374), .A1(net_10373), .A2(net_10372) );
NOR2_X2 inst_3427 ( .ZN(net_20418), .A2(net_15066), .A1(net_10868) );
NAND4_X2 inst_5486 ( .ZN(net_12400), .A3(net_8073), .A1(net_6834), .A2(net_6753), .A4(net_5749) );
NAND3_X2 inst_6262 ( .ZN(net_12988), .A3(net_12987), .A2(net_9087), .A1(net_8152) );
NAND3_X2 inst_5768 ( .ZN(net_20340), .A1(net_15223), .A3(net_15172), .A2(net_12152) );
NAND2_X4 inst_6946 ( .ZN(net_20461), .A1(net_17183), .A2(net_17057) );
OAI21_X2 inst_1954 ( .ZN(net_12541), .B1(net_8175), .B2(net_7356), .A(net_1811) );
CLKBUF_X2 inst_22836 ( .A(net_22707), .Z(net_22708) );
INV_X4 inst_16484 ( .ZN(net_1791), .A(net_1755) );
NOR2_X2 inst_3941 ( .A1(net_14078), .A2(net_8769), .ZN(net_8648) );
NAND2_X2 inst_7815 ( .ZN(net_18678), .A2(net_18638), .A1(net_18622) );
INV_X4 inst_13543 ( .ZN(net_20036), .A(net_9199) );
NAND2_X2 inst_10588 ( .A2(net_12935), .A1(net_7427), .ZN(net_6659) );
INV_X4 inst_12746 ( .ZN(net_18718), .A(net_17427) );
NOR2_X2 inst_3858 ( .ZN(net_11510), .A2(net_9467), .A1(net_6092) );
NAND2_X4 inst_7014 ( .A2(net_19668), .A1(net_19667), .ZN(net_17175) );
INV_X4 inst_13129 ( .ZN(net_19599), .A(net_14898) );
INV_X4 inst_13949 ( .ZN(net_6767), .A(net_6766) );
INV_X4 inst_13008 ( .ZN(net_16438), .A(net_16437) );
NAND2_X4 inst_7342 ( .ZN(net_6020), .A1(net_4863), .A2(net_2611) );
NOR2_X2 inst_5105 ( .ZN(net_5959), .A2(net_761), .A1(net_572) );
NAND2_X2 inst_8818 ( .ZN(net_15578), .A2(net_14848), .A1(net_13699) );
INV_X2 inst_19057 ( .ZN(net_4721), .A(net_4720) );
INV_X2 inst_18990 ( .ZN(net_5090), .A(net_5089) );
INV_X4 inst_12725 ( .ZN(net_17521), .A(net_17520) );
DFF_X1 inst_19908 ( .D(net_16781), .CK(net_21811), .Q(x1314) );
NOR2_X2 inst_3561 ( .ZN(net_12977), .A2(net_10287), .A1(net_7627) );
AOI21_X2 inst_20645 ( .ZN(net_13144), .B2(net_9554), .B1(net_2928), .A(net_1471) );
AOI221_X2 inst_20083 ( .B1(net_16051), .ZN(net_15972), .C1(net_15971), .C2(net_15323), .B2(net_13692), .A(net_7765) );
NAND2_X4 inst_7233 ( .A1(net_20477), .ZN(net_8520), .A2(net_7124) );
INV_X4 inst_17773 ( .ZN(net_6863), .A(net_4478) );
INV_X4 inst_14286 ( .A(net_7309), .ZN(net_5610) );
INV_X4 inst_18009 ( .A(net_21192), .ZN(net_11872) );
NOR2_X4 inst_3046 ( .ZN(net_6180), .A2(net_5043), .A1(net_5042) );
INV_X4 inst_16511 ( .ZN(net_5776), .A(net_143) );
NAND2_X2 inst_8751 ( .A1(net_21220), .ZN(net_15947), .A2(net_15551) );
NOR2_X2 inst_4644 ( .A2(net_4230), .ZN(net_3386), .A1(net_955) );
NOR2_X2 inst_4844 ( .ZN(net_5683), .A1(net_4773), .A2(net_2294) );
INV_X4 inst_14994 ( .ZN(net_6295), .A(net_3397) );
NOR2_X2 inst_3757 ( .ZN(net_10360), .A2(net_9394), .A1(net_7321) );
SDFF_X2 inst_917 ( .Q(net_21164), .D(net_16507), .SE(net_253), .CK(net_21640), .SI(x5145) );
NOR2_X2 inst_3712 ( .ZN(net_10997), .A2(net_10996), .A1(net_9165) );
OAI21_X2 inst_1743 ( .ZN(net_14975), .A(net_14974), .B1(net_14813), .B2(net_7329) );
AND2_X4 inst_21263 ( .ZN(net_3282), .A2(net_90), .A1(net_81) );
NAND2_X2 inst_11713 ( .ZN(net_2705), .A2(net_2365), .A1(net_2274) );
INV_X4 inst_13403 ( .ZN(net_10422), .A(net_10421) );
XNOR2_X2 inst_215 ( .ZN(net_17538), .A(net_17537), .B(net_6373) );
NOR2_X2 inst_5022 ( .ZN(net_1189), .A2(net_920), .A1(net_122) );
NOR3_X4 inst_2624 ( .A3(net_19664), .A1(net_19663), .ZN(net_19600), .A2(net_10881) );
INV_X2 inst_18524 ( .A(net_11688), .ZN(net_11131) );
AOI21_X4 inst_20175 ( .ZN(net_20221), .B2(net_14621), .B1(net_13557), .A(net_10122) );
NAND3_X2 inst_6258 ( .ZN(net_12997), .A2(net_12248), .A1(net_11359), .A3(net_10911) );
NAND2_X4 inst_7550 ( .ZN(net_2499), .A2(net_1784), .A1(net_1783) );
NAND2_X2 inst_11293 ( .ZN(net_6632), .A2(net_3819), .A1(net_1228) );
INV_X4 inst_17089 ( .ZN(net_1293), .A(net_364) );
INV_X4 inst_17060 ( .ZN(net_1515), .A(net_133) );
INV_X4 inst_15848 ( .ZN(net_2732), .A(net_1833) );
NAND2_X2 inst_8912 ( .ZN(net_14970), .A2(net_13743), .A1(net_13569) );
INV_X4 inst_17901 ( .A(net_20889), .ZN(net_178) );
NOR2_X2 inst_4819 ( .A1(net_6599), .ZN(net_5184), .A2(net_1767) );
CLKBUF_X2 inst_22167 ( .A(net_21992), .Z(net_22039) );
INV_X4 inst_15437 ( .ZN(net_3197), .A(net_1685) );
INV_X4 inst_17544 ( .ZN(net_3014), .A(net_1376) );
INV_X4 inst_16927 ( .ZN(net_11186), .A(net_8707) );
NOR2_X2 inst_4774 ( .ZN(net_2927), .A2(net_2038), .A1(net_252) );
INV_X4 inst_12997 ( .A(net_16801), .ZN(net_16628) );
NAND2_X2 inst_8622 ( .A1(net_21174), .A2(net_20527), .ZN(net_16604) );
INV_X4 inst_18060 ( .A(net_20998), .ZN(net_1948) );
INV_X8 inst_12401 ( .A(net_1271), .ZN(net_256) );
INV_X4 inst_17454 ( .A(net_9617), .ZN(net_8709) );
INV_X4 inst_18300 ( .A(net_20478), .ZN(net_20477) );
INV_X4 inst_14632 ( .ZN(net_4388), .A(net_4387) );
INV_X2 inst_18876 ( .ZN(net_6206), .A(net_6205) );
NOR2_X2 inst_4016 ( .ZN(net_20081), .A2(net_7163), .A1(net_2355) );
INV_X2 inst_19227 ( .A(net_5131), .ZN(net_3408) );
NOR2_X4 inst_2914 ( .ZN(net_13904), .A2(net_9917), .A1(net_6175) );
NAND2_X4 inst_7648 ( .ZN(net_19222), .A2(net_206), .A1(net_65) );
CLKBUF_X2 inst_22136 ( .A(net_22007), .Z(net_22008) );
NOR2_X4 inst_3294 ( .ZN(net_1638), .A2(net_773), .A1(net_129) );
NOR3_X2 inst_2741 ( .ZN(net_12755), .A1(net_10196), .A3(net_9597), .A2(net_6555) );
NAND2_X2 inst_11825 ( .A1(net_20875), .ZN(net_3290), .A2(net_1787) );
INV_X4 inst_15262 ( .A(net_5621), .ZN(net_2771) );
NAND2_X2 inst_11966 ( .ZN(net_3082), .A1(net_227), .A2(net_187) );
CLKBUF_X2 inst_22365 ( .A(net_22236), .Z(net_22237) );
OAI21_X2 inst_1522 ( .ZN(net_18143), .A(net_18090), .B1(net_18089), .B2(net_5616) );
INV_X4 inst_14380 ( .ZN(net_11347), .A(net_6980) );
NAND2_X1 inst_12135 ( .ZN(net_17558), .A1(net_17557), .A2(net_17232) );
AND4_X2 inst_21108 ( .A3(net_11748), .ZN(net_11730), .A1(net_11729), .A2(net_11728), .A4(net_11727) );
NAND2_X2 inst_11455 ( .ZN(net_4962), .A2(net_3234), .A1(net_1224) );
INV_X4 inst_13955 ( .ZN(net_6756), .A(net_6755) );
INV_X4 inst_16931 ( .ZN(net_10093), .A(net_6877) );
INV_X2 inst_18964 ( .ZN(net_5406), .A(net_5405) );
NAND2_X2 inst_8645 ( .A1(net_20216), .A2(net_16612), .ZN(net_16568) );
INV_X4 inst_16566 ( .ZN(net_1953), .A(net_1162) );
NAND3_X2 inst_5761 ( .ZN(net_15967), .A3(net_15618), .A2(net_12349), .A1(net_9792) );
NAND2_X4 inst_6964 ( .ZN(net_17427), .A2(net_17053), .A1(net_16916) );
INV_X2 inst_19660 ( .A(net_20440), .ZN(net_20439) );
INV_X4 inst_12520 ( .ZN(net_18521), .A(net_18494) );
INV_X4 inst_12809 ( .ZN(net_17307), .A(net_17209) );
NAND2_X2 inst_9528 ( .A1(net_11757), .ZN(net_11121), .A2(net_6293) );
NAND2_X2 inst_11889 ( .ZN(net_2082), .A2(net_1640), .A1(net_955) );
NAND3_X2 inst_5691 ( .ZN(net_16271), .A2(net_15979), .A3(net_15839), .A1(net_5363) );
NAND2_X2 inst_7902 ( .ZN(net_18480), .A2(net_18376), .A1(net_17726) );
SDFF_X2 inst_861 ( .Q(net_21229), .SI(net_17171), .SE(net_125), .CK(net_22154), .D(x7042) );
NAND2_X2 inst_8392 ( .ZN(net_17280), .A2(net_17017), .A1(net_16871) );
INV_X2 inst_18937 ( .ZN(net_5825), .A(net_5824) );
NAND2_X4 inst_7431 ( .ZN(net_10236), .A1(net_3955), .A2(net_1698) );
NAND2_X2 inst_11549 ( .ZN(net_3596), .A2(net_2416), .A1(net_936) );
AOI21_X2 inst_20602 ( .A(net_15205), .ZN(net_13834), .B2(net_10967), .B1(net_4480) );
NOR2_X4 inst_2990 ( .ZN(net_10337), .A2(net_8369), .A1(net_5659) );
NAND2_X4 inst_7495 ( .A2(net_2950), .ZN(net_2342), .A1(net_1733) );
OAI22_X2 inst_1283 ( .B1(net_15481), .ZN(net_15118), .A2(net_13247), .B2(net_10474), .A1(net_5186) );
INV_X4 inst_17345 ( .ZN(net_5594), .A(net_703) );
INV_X4 inst_18299 ( .A(net_20478), .ZN(net_20474) );
NAND2_X2 inst_11225 ( .ZN(net_3956), .A2(net_3955), .A1(net_703) );
INV_X4 inst_17232 ( .ZN(net_2319), .A(net_1148) );
NAND2_X2 inst_10625 ( .A1(net_8543), .ZN(net_6562), .A2(net_6561) );
NOR2_X2 inst_4290 ( .ZN(net_6035), .A2(net_6034), .A1(net_2280) );
INV_X4 inst_18050 ( .A(net_20897), .ZN(net_47) );
INV_X4 inst_16796 ( .ZN(net_5217), .A(net_1357) );
INV_X4 inst_12594 ( .ZN(net_18158), .A(net_18106) );
NAND2_X2 inst_11027 ( .A1(net_5241), .ZN(net_4777), .A2(net_3405) );
INV_X4 inst_15104 ( .ZN(net_3931), .A(net_3762) );
AOI211_X2 inst_21038 ( .ZN(net_14091), .B(net_12965), .C2(net_10432), .A(net_10133), .C1(net_3277) );
INV_X4 inst_17918 ( .A(net_20879), .ZN(net_220) );
NAND2_X2 inst_10238 ( .A1(net_9083), .ZN(net_8038), .A2(net_5145) );
INV_X4 inst_16321 ( .A(net_9339), .ZN(net_4113) );
NAND4_X4 inst_5195 ( .ZN(net_17760), .A1(net_16322), .A4(net_16194), .A2(net_15680), .A3(net_12211) );
INV_X4 inst_14701 ( .A(net_13565), .ZN(net_4452) );
INV_X4 inst_18002 ( .A(net_21063), .ZN(net_520) );
INV_X2 inst_19044 ( .ZN(net_4757), .A(net_4756) );
NOR2_X2 inst_3462 ( .ZN(net_14676), .A1(net_14675), .A2(net_13254) );
INV_X4 inst_16353 ( .ZN(net_8160), .A(net_6221) );
NOR2_X2 inst_4254 ( .A2(net_7672), .ZN(net_6335), .A1(net_6334) );
NAND2_X2 inst_8288 ( .ZN(net_17620), .A2(net_17532), .A1(net_812) );
NOR2_X2 inst_4330 ( .ZN(net_9855), .A2(net_4575), .A1(net_761) );
NAND2_X2 inst_10031 ( .ZN(net_19643), .A1(net_8734), .A2(net_8733) );
NAND2_X2 inst_11925 ( .A2(net_6563), .ZN(net_2247), .A1(net_1451) );
INV_X4 inst_14220 ( .ZN(net_7374), .A(net_5847) );
INV_X2 inst_19085 ( .ZN(net_4576), .A(net_4575) );
INV_X8 inst_12204 ( .ZN(net_11020), .A(net_7590) );
NAND2_X2 inst_9388 ( .ZN(net_20672), .A1(net_9447), .A2(net_7326) );
NOR3_X2 inst_2754 ( .ZN(net_11761), .A1(net_9582), .A3(net_7945), .A2(net_7793) );
SDFF_X2 inst_794 ( .Q(net_20883), .SE(net_18847), .SI(net_18009), .D(net_585), .CK(net_21798) );
INV_X4 inst_14577 ( .ZN(net_7488), .A(net_4218) );
INV_X4 inst_17864 ( .ZN(net_214), .A(net_102) );
NAND2_X4 inst_7354 ( .ZN(net_7472), .A1(net_2641), .A2(net_1645) );
CLKBUF_X2 inst_22312 ( .A(net_22183), .Z(net_22184) );
AOI21_X2 inst_20524 ( .ZN(net_14558), .B1(net_14557), .B2(net_11966), .A(net_7181) );
INV_X4 inst_17663 ( .ZN(net_375), .A(net_253) );
NAND2_X2 inst_12049 ( .A2(net_4718), .ZN(net_1145), .A1(net_934) );
NOR3_X2 inst_2759 ( .ZN(net_11213), .A2(net_11212), .A3(net_11211), .A1(net_7796) );
INV_X4 inst_17378 ( .ZN(net_1195), .A(net_234) );
NAND2_X2 inst_12092 ( .ZN(net_1031), .A1(net_664), .A2(net_625) );
CLKBUF_X2 inst_21728 ( .A(net_21272), .Z(net_21600) );
NAND2_X2 inst_8256 ( .A2(net_17852), .ZN(net_17698), .A1(net_17697) );
NAND2_X2 inst_11165 ( .A1(net_8205), .ZN(net_4176), .A2(net_4175) );
OAI211_X2 inst_2423 ( .ZN(net_15231), .B(net_14142), .C1(net_13871), .A(net_13486), .C2(net_12869) );
INV_X4 inst_16131 ( .ZN(net_2747), .A(net_1479) );
AOI21_X2 inst_20345 ( .A(net_20856), .B2(net_19870), .B1(net_19869), .ZN(net_15760) );
INV_X2 inst_19316 ( .A(net_3501), .ZN(net_2633) );
SDFF_X2 inst_996 ( .QN(net_21032), .D(net_505), .SE(net_263), .CK(net_21958), .SI(x2457) );
NAND2_X2 inst_10963 ( .ZN(net_8233), .A2(net_4632), .A1(net_4288) );
NAND3_X2 inst_5889 ( .ZN(net_15226), .A1(net_14648), .A2(net_13523), .A3(net_13430) );
INV_X4 inst_16230 ( .ZN(net_9401), .A(net_7870) );
NAND2_X2 inst_12074 ( .A2(net_3491), .ZN(net_1234), .A1(net_194) );
OAI21_X2 inst_1527 ( .ZN(net_18024), .B1(net_18003), .B2(net_17943), .A(net_2023) );
NAND3_X2 inst_6142 ( .A2(net_14874), .ZN(net_13712), .A3(net_11049), .A1(net_8251) );
SDFF_X2 inst_740 ( .Q(net_20929), .SE(net_18577), .SI(net_18532), .D(net_577), .CK(net_21442) );
NOR2_X2 inst_4189 ( .ZN(net_13776), .A1(net_6207), .A2(net_5147) );
NAND2_X2 inst_7803 ( .ZN(net_18697), .A2(net_18696), .A1(net_17389) );
INV_X4 inst_17324 ( .A(net_15108), .ZN(net_12916) );
NAND3_X2 inst_6803 ( .A3(net_3385), .ZN(net_3267), .A1(net_2757), .A2(net_986) );
OAI21_X2 inst_1937 ( .ZN(net_12917), .A(net_12916), .B1(net_12915), .B2(net_9585) );
INV_X4 inst_15756 ( .A(net_9514), .ZN(net_5246) );
XNOR2_X2 inst_611 ( .A(net_21164), .B(net_16794), .ZN(net_1516) );
NOR2_X2 inst_4405 ( .ZN(net_6262), .A1(net_3553), .A2(net_3174) );
NAND2_X2 inst_10550 ( .ZN(net_11594), .A2(net_5687), .A1(net_4288) );
OAI211_X2 inst_2487 ( .ZN(net_13250), .A(net_10617), .B(net_9133), .C2(net_5583), .C1(net_1066) );
CLKBUF_X2 inst_22439 ( .A(net_22310), .Z(net_22311) );
INV_X8 inst_12417 ( .A(net_21212), .ZN(net_16743) );
CLKBUF_X2 inst_21496 ( .A(net_21367), .Z(net_21368) );
INV_X4 inst_12462 ( .ZN(net_18828), .A(net_18827) );
INV_X4 inst_12549 ( .ZN(net_18339), .A(net_18283) );
INV_X4 inst_16622 ( .ZN(net_8490), .A(net_983) );
NAND2_X2 inst_7802 ( .ZN(net_18698), .A2(net_18696), .A1(net_17084) );
INV_X4 inst_15856 ( .ZN(net_1942), .A(net_1814) );
XNOR2_X2 inst_490 ( .ZN(net_9241), .A(net_9240), .B(net_4492) );
INV_X2 inst_19685 ( .A(net_20527), .ZN(net_20526) );
AOI21_X2 inst_20930 ( .B1(net_7912), .ZN(net_7070), .B2(net_3848), .A(net_1371) );
CLKBUF_X2 inst_22794 ( .A(net_22665), .Z(net_22666) );
NAND2_X4 inst_7305 ( .ZN(net_6762), .A1(net_5478), .A2(net_232) );
CLKBUF_X2 inst_22217 ( .A(net_22073), .Z(net_22089) );
NAND2_X2 inst_8375 ( .A1(net_20067), .A2(net_17363), .ZN(net_17356) );
INV_X4 inst_13378 ( .ZN(net_13608), .A(net_10871) );
OAI21_X2 inst_2218 ( .B2(net_9072), .ZN(net_8516), .A(net_8515), .B1(net_6698) );
CLKBUF_X2 inst_22079 ( .A(net_21581), .Z(net_21951) );
OAI22_X2 inst_1309 ( .ZN(net_8984), .A1(net_8983), .A2(net_8982), .B1(net_8981), .B2(net_8980) );
INV_X2 inst_18396 ( .ZN(net_20167), .A(net_16427) );
INV_X4 inst_15045 ( .ZN(net_3578), .A(net_3328) );
NOR2_X2 inst_3803 ( .ZN(net_9853), .A2(net_9463), .A1(net_6328) );
NOR2_X2 inst_4938 ( .ZN(net_2971), .A1(net_1148), .A2(net_1127) );
INV_X4 inst_15049 ( .ZN(net_20825), .A(net_3811) );
INV_X4 inst_16103 ( .A(net_5201), .ZN(net_4018) );
NOR2_X4 inst_3183 ( .ZN(net_5478), .A1(net_4014), .A2(net_955) );
NAND2_X2 inst_10242 ( .ZN(net_8024), .A1(net_7677), .A2(net_5679) );
INV_X4 inst_13234 ( .ZN(net_13475), .A(net_12443) );
INV_X4 inst_15095 ( .ZN(net_13095), .A(net_10191) );
NAND2_X2 inst_10860 ( .ZN(net_5444), .A2(net_5443), .A1(net_628) );
INV_X4 inst_16498 ( .ZN(net_7950), .A(net_4250) );
INV_X2 inst_19079 ( .ZN(net_4595), .A(net_4594) );
INV_X4 inst_13301 ( .ZN(net_13553), .A(net_12319) );
NOR2_X2 inst_4312 ( .A1(net_9342), .ZN(net_7411), .A2(net_5874) );
NAND2_X2 inst_11256 ( .ZN(net_5643), .A1(net_4918), .A2(net_3384) );
INV_X4 inst_12950 ( .ZN(net_17066), .A(net_17048) );
NAND4_X2 inst_5328 ( .ZN(net_19077), .A3(net_15457), .A1(net_15075), .A4(net_12165), .A2(net_10118) );
NAND2_X2 inst_8410 ( .A1(net_19435), .ZN(net_17360), .A2(net_17234) );
NAND3_X2 inst_6226 ( .ZN(net_13235), .A3(net_13234), .A1(net_9850), .A2(net_5412) );
INV_X4 inst_13161 ( .ZN(net_14815), .A(net_14233) );
INV_X2 inst_18782 ( .ZN(net_7508), .A(net_7507) );
XNOR2_X2 inst_300 ( .ZN(net_17117), .B(net_16646), .A(net_16629) );
INV_X4 inst_15407 ( .A(net_7394), .ZN(net_6528) );
OR2_X2 inst_1226 ( .A2(net_6387), .ZN(net_2312), .A1(net_2311) );
CLKBUF_X2 inst_21702 ( .A(net_21312), .Z(net_21574) );
NAND3_X2 inst_5964 ( .ZN(net_14785), .A1(net_13324), .A3(net_13273), .A2(net_8459) );
INV_X4 inst_17836 ( .ZN(net_253), .A(net_125) );
XNOR2_X2 inst_446 ( .ZN(net_14918), .B(net_14917), .A(net_12876) );
NAND2_X2 inst_8802 ( .ZN(net_20388), .A2(net_19280), .A1(net_19279) );
INV_X4 inst_15619 ( .ZN(net_5260), .A(net_2160) );
INV_X4 inst_15949 ( .ZN(net_1851), .A(net_1712) );
AOI21_X2 inst_20907 ( .ZN(net_7687), .B2(net_6176), .B1(net_3273), .A(net_1648) );
NOR2_X2 inst_4923 ( .A2(net_3830), .ZN(net_1824), .A1(net_1353) );
INV_X2 inst_18689 ( .ZN(net_8607), .A(net_7180) );
NOR2_X2 inst_3533 ( .ZN(net_13551), .A2(net_10944), .A1(net_4133) );
SDFF_X2 inst_824 ( .Q(net_21173), .SI(net_17575), .SE(net_125), .CK(net_22444), .D(x4781) );
INV_X4 inst_15996 ( .ZN(net_14458), .A(net_11776) );
NAND2_X2 inst_7839 ( .A2(net_18640), .ZN(net_18623), .A1(net_16634) );
INV_X4 inst_12897 ( .ZN(net_16950), .A(net_16787) );
NAND2_X2 inst_10393 ( .A1(net_13762), .A2(net_12035), .ZN(net_7304) );
INV_X4 inst_14678 ( .ZN(net_20335), .A(net_4309) );
INV_X4 inst_16135 ( .ZN(net_5714), .A(net_4179) );
NAND3_X2 inst_6600 ( .ZN(net_9892), .A2(net_9692), .A1(net_6136), .A3(net_4501) );
NAND2_X2 inst_9007 ( .A1(net_14755), .ZN(net_14278), .A2(net_13549) );
INV_X4 inst_13691 ( .ZN(net_12777), .A(net_7944) );
NOR2_X2 inst_3750 ( .A1(net_11406), .ZN(net_10423), .A2(net_10189) );
NAND2_X2 inst_11173 ( .ZN(net_7062), .A2(net_3012), .A1(net_399) );
INV_X4 inst_15286 ( .ZN(net_4837), .A(net_2019) );
AOI21_X2 inst_20668 ( .ZN(net_20114), .A(net_13032), .B1(net_12910), .B2(net_9442) );
NOR2_X2 inst_4056 ( .ZN(net_7839), .A1(net_7838), .A2(net_4699) );
NOR2_X2 inst_4401 ( .ZN(net_19204), .A2(net_12500), .A1(net_761) );
NOR2_X2 inst_3430 ( .ZN(net_15319), .A2(net_14372), .A1(net_11129) );
NAND2_X2 inst_10388 ( .A1(net_14751), .ZN(net_10749), .A2(net_7320) );
CLKBUF_X2 inst_21692 ( .A(net_21563), .Z(net_21564) );
AOI21_X2 inst_20841 ( .A(net_11311), .ZN(net_9269), .B2(net_4558), .B1(net_3020) );
INV_X2 inst_19694 ( .ZN(net_20547), .A(net_20545) );
CLKBUF_X2 inst_22196 ( .A(net_22067), .Z(net_22068) );
INV_X4 inst_13368 ( .A(net_12987), .ZN(net_10908) );
CLKBUF_X2 inst_22360 ( .A(net_22231), .Z(net_22232) );
NAND4_X2 inst_5462 ( .ZN(net_13327), .A1(net_13326), .A2(net_12903), .A4(net_12902), .A3(net_10754) );
NOR2_X2 inst_3439 ( .ZN(net_15199), .A1(net_15198), .A2(net_14556) );
INV_X4 inst_17159 ( .ZN(net_7075), .A(net_5448) );
INV_X4 inst_13968 ( .ZN(net_7966), .A(net_5430) );
NAND4_X2 inst_5412 ( .ZN(net_14587), .A2(net_12439), .A3(net_11282), .A1(net_11140), .A4(net_10001) );
NAND2_X2 inst_8308 ( .ZN(net_19666), .A2(net_17586), .A1(net_17534) );
CLKBUF_X2 inst_22609 ( .A(net_22480), .Z(net_22481) );
NAND2_X2 inst_10901 ( .ZN(net_14921), .A1(net_5448), .A2(net_5373) );
NAND2_X2 inst_10014 ( .ZN(net_10272), .A1(net_9260), .A2(net_8158) );
CLKBUF_X2 inst_22798 ( .A(net_21398), .Z(net_22670) );
INV_X8 inst_12459 ( .ZN(net_20805), .A(net_20802) );
NAND3_X2 inst_6601 ( .ZN(net_9889), .A3(net_6198), .A2(net_6024), .A1(net_4972) );
NAND2_X2 inst_8520 ( .A2(net_20501), .A1(net_17029), .ZN(net_16908) );
AOI21_X2 inst_20939 ( .A(net_6922), .ZN(net_6460), .B1(net_6459), .B2(net_6444) );
OAI21_X2 inst_1571 ( .B1(net_16644), .ZN(net_16388), .A(net_16207), .B2(net_16189) );
INV_X4 inst_15540 ( .A(net_15684), .ZN(net_3164) );
NAND2_X2 inst_12009 ( .ZN(net_9276), .A1(net_1574), .A2(net_824) );
INV_X4 inst_17446 ( .ZN(net_15370), .A(net_15108) );
NAND2_X2 inst_8214 ( .ZN(net_17846), .A2(net_17845), .A1(net_17831) );
OAI21_X4 inst_1402 ( .A(net_20864), .B2(net_19478), .B1(net_19477), .ZN(net_16232) );
NAND3_X2 inst_6511 ( .ZN(net_10778), .A3(net_10777), .A1(net_8296), .A2(net_6874) );
NAND2_X2 inst_11246 ( .ZN(net_8988), .A2(net_3924), .A1(net_721) );
DFF_X1 inst_19811 ( .Q(net_20880), .D(net_18002), .CK(net_22816) );
NOR2_X4 inst_3106 ( .A1(net_19462), .ZN(net_7008), .A2(net_2744) );
NAND3_X2 inst_6810 ( .A1(net_6812), .ZN(net_5585), .A2(net_2948), .A3(net_913) );
INV_X2 inst_18586 ( .ZN(net_10277), .A(net_10276) );
NAND2_X4 inst_6843 ( .ZN(net_20473), .A1(net_18644), .A2(net_18635) );
INV_X4 inst_13379 ( .ZN(net_10868), .A(net_10867) );
INV_X4 inst_17366 ( .ZN(net_7473), .A(net_120) );
NAND3_X2 inst_6270 ( .A2(net_14545), .ZN(net_12956), .A3(net_11622), .A1(net_6823) );
NAND4_X2 inst_5453 ( .ZN(net_13464), .A3(net_13147), .A4(net_11918), .A2(net_9135), .A1(net_5615) );
NAND4_X2 inst_5405 ( .ZN(net_14656), .A2(net_12044), .A3(net_10745), .A4(net_8011), .A1(net_7169) );
NAND2_X2 inst_8810 ( .ZN(net_20037), .A1(net_15833), .A2(net_14924) );
INV_X4 inst_13317 ( .ZN(net_11592), .A(net_11591) );
OAI211_X2 inst_2503 ( .ZN(net_12780), .C2(net_12738), .A(net_11697), .B(net_11554), .C1(net_7394) );
NAND2_X4 inst_7193 ( .ZN(net_11826), .A1(net_7455), .A2(net_5456) );
INV_X4 inst_15347 ( .A(net_16287), .ZN(net_2594) );
NOR2_X2 inst_4877 ( .ZN(net_2201), .A1(net_1784), .A2(net_1756) );
NAND4_X2 inst_5420 ( .ZN(net_14383), .A4(net_14210), .A2(net_11423), .A3(net_9517), .A1(net_8705) );
NAND2_X2 inst_9994 ( .ZN(net_20399), .A1(net_8839), .A2(net_6490) );
CLKBUF_X2 inst_22955 ( .A(net_21567), .Z(net_22827) );
XNOR2_X2 inst_94 ( .ZN(net_18550), .A(net_18449), .B(net_17923) );
AOI221_X2 inst_20081 ( .ZN(net_19963), .B1(net_16051), .C1(net_16050), .C2(net_15367), .B2(net_14772), .A(net_14412) );
INV_X2 inst_19308 ( .ZN(net_6471), .A(net_2055) );
NAND2_X2 inst_10946 ( .ZN(net_5134), .A2(net_3559), .A1(net_1160) );
AOI21_X2 inst_20494 ( .ZN(net_14739), .B1(net_14738), .B2(net_12237), .A(net_9117) );
AOI21_X2 inst_20674 ( .B1(net_19419), .ZN(net_12572), .B2(net_12516), .A(net_1889) );
INV_X2 inst_18489 ( .ZN(net_13406), .A(net_12350) );
INV_X4 inst_14615 ( .ZN(net_13246), .A(net_9033) );
INV_X4 inst_17314 ( .ZN(net_2976), .A(net_165) );
NAND2_X2 inst_11858 ( .ZN(net_2011), .A1(net_1708), .A2(net_1207) );
INV_X4 inst_13060 ( .ZN(net_16353), .A(net_16301) );
XNOR2_X2 inst_591 ( .B(net_16648), .ZN(net_564), .A(net_563) );
XNOR2_X2 inst_424 ( .B(net_21164), .A(net_16506), .ZN(net_16504) );
NOR2_X2 inst_4345 ( .A2(net_12954), .ZN(net_5638), .A1(net_4146) );
AOI21_X2 inst_20488 ( .ZN(net_14770), .B2(net_13225), .A(net_11542), .B1(net_816) );
INV_X4 inst_15504 ( .A(net_4018), .ZN(net_2419) );
INV_X4 inst_15338 ( .ZN(net_13355), .A(net_11909) );
INV_X2 inst_18721 ( .ZN(net_8127), .A(net_8126) );
NAND2_X2 inst_10428 ( .A1(net_8685), .ZN(net_7218), .A2(net_6744) );
INV_X4 inst_17624 ( .ZN(net_2071), .A(net_1861) );
NOR2_X2 inst_4417 ( .ZN(net_8285), .A2(net_5537), .A1(net_4934) );
NAND2_X2 inst_10784 ( .A1(net_9968), .ZN(net_5592), .A2(net_4277) );
NAND2_X2 inst_8320 ( .ZN(net_20244), .A2(net_17552), .A1(net_17522) );
CLKBUF_X2 inst_21477 ( .A(net_21294), .Z(net_21349) );
DFF_X2 inst_19780 ( .D(net_5267), .Q(net_26), .CK(net_21507) );
INV_X2 inst_19699 ( .A(net_20561), .ZN(net_20560) );
INV_X2 inst_19391 ( .ZN(net_2081), .A(net_2080) );
NAND3_X2 inst_5727 ( .ZN(net_19177), .A1(net_15851), .A3(net_15138), .A2(net_7139) );
INV_X4 inst_14012 ( .ZN(net_9693), .A(net_8195) );
NAND2_X2 inst_11861 ( .ZN(net_6485), .A2(net_5259), .A1(net_1495) );
NAND2_X4 inst_6853 ( .A1(net_20320), .ZN(net_18482), .A2(net_17730) );
NOR3_X2 inst_2706 ( .ZN(net_13907), .A1(net_11950), .A3(net_10219), .A2(net_7546) );
INV_X4 inst_16389 ( .ZN(net_5439), .A(net_5097) );
XNOR2_X2 inst_476 ( .ZN(net_11881), .A(net_11880), .B(net_1862) );
NAND2_X2 inst_8640 ( .ZN(net_16578), .A1(net_16577), .A2(net_16576) );
NOR2_X2 inst_3742 ( .ZN(net_10666), .A1(net_8735), .A2(net_7344) );
NAND3_X2 inst_6684 ( .A2(net_12564), .ZN(net_7715), .A3(net_7714), .A1(net_3698) );
NAND2_X2 inst_10249 ( .ZN(net_14193), .A1(net_8674), .A2(net_8013) );
OAI211_X2 inst_2499 ( .C1(net_15297), .ZN(net_12863), .A(net_11102), .B(net_8645), .C2(net_7739) );
INV_X4 inst_16150 ( .ZN(net_15374), .A(net_14548) );
XOR2_X2 inst_20 ( .A(net_21127), .B(net_16887), .Z(net_16878) );
NAND2_X2 inst_11542 ( .ZN(net_2914), .A2(net_2913), .A1(net_85) );
INV_X4 inst_18222 ( .A(net_20881), .ZN(net_126) );
AOI22_X2 inst_20049 ( .ZN(net_3708), .A1(net_3707), .B1(net_3456), .A2(net_3192), .B2(net_2321) );
NAND2_X2 inst_10007 ( .ZN(net_12151), .A2(net_10475), .A1(net_8802) );
DFF_X1 inst_19906 ( .D(net_16800), .CK(net_21816), .Q(x1322) );
NAND3_X4 inst_5549 ( .A3(net_20332), .A1(net_20331), .ZN(net_16996), .A2(net_16078) );
INV_X4 inst_13421 ( .ZN(net_10228), .A(net_10227) );
NOR2_X2 inst_4994 ( .ZN(net_5309), .A1(net_1397), .A2(net_865) );
INV_X4 inst_15387 ( .ZN(net_15270), .A(net_8732) );
XNOR2_X2 inst_576 ( .ZN(net_617), .A(net_616), .B(net_615) );
INV_X4 inst_13590 ( .ZN(net_8860), .A(net_7304) );
INV_X4 inst_14477 ( .A(net_6588), .ZN(net_4893) );
INV_X4 inst_14398 ( .A(net_6837), .ZN(net_6157) );
NAND2_X2 inst_10131 ( .ZN(net_10314), .A1(net_6613), .A2(net_5426) );
NAND2_X2 inst_10182 ( .ZN(net_10186), .A1(net_8186), .A2(net_4970) );
INV_X4 inst_17970 ( .A(net_21018), .ZN(net_574) );
NAND2_X2 inst_10376 ( .A1(net_18025), .ZN(net_7390), .A2(net_416) );
INV_X4 inst_16629 ( .ZN(net_14630), .A(net_14174) );
NOR2_X4 inst_3055 ( .ZN(net_6143), .A2(net_4989), .A1(net_2585) );
NOR2_X4 inst_2876 ( .A2(net_14904), .ZN(net_10324), .A1(net_10323) );
INV_X4 inst_16516 ( .A(net_11297), .ZN(net_1663) );
INV_X4 inst_16371 ( .ZN(net_6947), .A(net_4792) );
SDFF_X2 inst_976 ( .QN(net_21042), .D(net_384), .SE(net_263), .CK(net_22522), .SI(x2280) );
INV_X4 inst_17150 ( .ZN(net_11296), .A(net_3148) );
NAND2_X2 inst_9919 ( .A1(net_9693), .ZN(net_9281), .A2(net_3642) );
INV_X4 inst_17610 ( .A(net_6692), .ZN(net_1020) );
OAI22_X2 inst_1279 ( .ZN(net_16077), .B1(net_16076), .A2(net_15556), .B2(net_14540), .A1(net_4466) );
NAND2_X4 inst_7027 ( .ZN(net_17232), .A1(net_16586), .A2(net_16458) );
NAND3_X2 inst_6562 ( .A2(net_11165), .ZN(net_10485), .A3(net_10484), .A1(net_4786) );
INV_X4 inst_16437 ( .ZN(net_4621), .A(net_1241) );
INV_X4 inst_16554 ( .A(net_3777), .ZN(net_2177) );
NAND2_X4 inst_7474 ( .ZN(net_3416), .A2(net_1527), .A1(net_504) );
INV_X4 inst_13011 ( .ZN(net_16729), .A(net_16574) );
INV_X4 inst_13280 ( .ZN(net_20686), .A(net_11169) );
INV_X4 inst_13287 ( .ZN(net_13566), .A(net_12413) );
AND2_X4 inst_21192 ( .ZN(net_20819), .A1(net_14538), .A2(net_7259) );
NAND2_X2 inst_8025 ( .ZN(net_18270), .A2(net_18265), .A1(net_17185) );
NAND2_X2 inst_11036 ( .A2(net_20469), .ZN(net_11338), .A1(net_3748) );
NAND2_X2 inst_7723 ( .ZN(net_18835), .A2(net_18791), .A1(net_17841) );
AND3_X2 inst_21152 ( .A2(net_10714), .A3(net_6696), .ZN(net_2061), .A1(net_2060) );
INV_X4 inst_18145 ( .A(net_20911), .ZN(net_646) );
NOR2_X2 inst_3414 ( .ZN(net_20182), .A2(net_15096), .A1(net_13771) );
NOR2_X2 inst_3399 ( .ZN(net_18910), .A2(net_15439), .A1(net_15326) );
CLKBUF_X2 inst_22785 ( .A(net_22656), .Z(net_22657) );
INV_X4 inst_17223 ( .A(net_14600), .ZN(net_13517) );
NOR2_X2 inst_4495 ( .ZN(net_6600), .A1(net_4270), .A2(net_4269) );
OAI21_X4 inst_1432 ( .B2(net_20760), .B1(net_20759), .ZN(net_16019), .A(net_15681) );
NAND3_X2 inst_5667 ( .ZN(net_16389), .A2(net_16209), .A3(net_16072), .A1(net_13352) );
NAND2_X1 inst_12159 ( .ZN(net_1973), .A2(net_1689), .A1(net_165) );
NOR2_X4 inst_3084 ( .A1(net_20465), .ZN(net_4375), .A2(net_4374) );
INV_X2 inst_19006 ( .A(net_6846), .ZN(net_5023) );
NAND2_X2 inst_11739 ( .ZN(net_5280), .A1(net_2178), .A2(net_2177) );
INV_X4 inst_15562 ( .ZN(net_4439), .A(net_2307) );
INV_X4 inst_16344 ( .ZN(net_2242), .A(net_971) );
OAI211_X2 inst_2464 ( .ZN(net_14112), .C2(net_13203), .C1(net_10512), .B(net_10460), .A(net_6785) );
NAND2_X2 inst_9790 ( .ZN(net_9740), .A1(net_9739), .A2(net_9738) );
NAND2_X2 inst_8776 ( .ZN(net_15817), .A2(net_15364), .A1(net_14730) );
NAND2_X2 inst_9433 ( .A1(net_12878), .ZN(net_11596), .A2(net_5407) );
NAND2_X2 inst_11197 ( .A1(net_20476), .ZN(net_6989), .A2(net_2447) );
INV_X4 inst_14432 ( .A(net_5029), .ZN(net_5027) );
INV_X4 inst_16347 ( .ZN(net_8741), .A(net_8644) );
NOR2_X2 inst_4010 ( .ZN(net_8077), .A1(net_8076), .A2(net_8075) );
INV_X4 inst_15373 ( .ZN(net_13375), .A(net_6993) );
NOR2_X4 inst_3328 ( .ZN(net_1025), .A2(net_513), .A1(net_322) );
NAND2_X2 inst_9677 ( .ZN(net_20826), .A1(net_9727), .A2(net_9669) );
INV_X4 inst_13254 ( .ZN(net_20014), .A(net_11703) );
NAND2_X2 inst_8399 ( .ZN(net_17394), .A1(net_16956), .A2(net_16790) );
OR2_X4 inst_1111 ( .ZN(net_4838), .A2(net_3120), .A1(net_86) );
INV_X4 inst_14495 ( .ZN(net_6018), .A(net_4843) );
DFF_X1 inst_19873 ( .D(net_17021), .CK(net_22543), .Q(x122) );
INV_X4 inst_17925 ( .A(net_20993), .ZN(net_1862) );
INV_X16 inst_19740 ( .ZN(net_1630), .A(net_875) );
NOR3_X2 inst_2658 ( .ZN(net_18926), .A1(net_14360), .A3(net_14034), .A2(net_4235) );
NAND2_X2 inst_9122 ( .ZN(net_15314), .A1(net_14055), .A2(net_12341) );
CLKBUF_X2 inst_21959 ( .A(net_21830), .Z(net_21831) );
NAND2_X2 inst_11496 ( .ZN(net_11279), .A1(net_5448), .A2(net_3084) );
CLKBUF_X2 inst_22469 ( .A(net_22340), .Z(net_22341) );
XNOR2_X2 inst_480 ( .ZN(net_11864), .A(net_11863), .B(net_2132) );
AOI211_X4 inst_20989 ( .C2(net_20291), .C1(net_20290), .ZN(net_16135), .B(net_15759), .A(net_14418) );
NOR2_X2 inst_4631 ( .ZN(net_20020), .A1(net_3002), .A2(net_2566) );
NOR2_X4 inst_2986 ( .ZN(net_7521), .A1(net_6077), .A2(net_4158) );
OAI21_X2 inst_2206 ( .B1(net_11221), .A(net_10590), .ZN(net_8536), .B2(net_6946) );
NAND2_X2 inst_8074 ( .A2(net_18162), .ZN(net_18161), .A1(net_17456) );
NOR3_X2 inst_2792 ( .ZN(net_4505), .A1(net_4503), .A2(net_1740), .A3(net_222) );
INV_X4 inst_13597 ( .ZN(net_8767), .A(net_7274) );
INV_X4 inst_17053 ( .ZN(net_10521), .A(net_6314) );
SDFF_X2 inst_739 ( .Q(net_20968), .D(net_18551), .SE(net_18025), .SI(net_561), .CK(net_22755) );
AND2_X2 inst_21309 ( .A2(net_12838), .A1(net_11708), .ZN(net_8935) );
INV_X4 inst_18111 ( .A(net_21039), .ZN(net_461) );
XOR2_X2 inst_46 ( .A(net_21117), .Z(net_480), .B(net_479) );
NAND3_X2 inst_6637 ( .A2(net_11162), .ZN(net_8972), .A3(net_8971), .A1(net_4404) );
OAI211_X2 inst_2537 ( .ZN(net_20450), .C2(net_12640), .C1(net_11236), .A(net_7596), .B(net_6060) );
INV_X4 inst_15530 ( .ZN(net_10993), .A(net_8068) );
INV_X4 inst_16862 ( .ZN(net_10512), .A(net_6743) );
OR2_X4 inst_1126 ( .ZN(net_6334), .A2(net_2274), .A1(net_308) );
INV_X8 inst_12361 ( .ZN(net_3491), .A(net_965) );
INV_X4 inst_16180 ( .ZN(net_11550), .A(net_1657) );
NOR2_X2 inst_3470 ( .A1(net_15681), .ZN(net_14489), .A2(net_12745) );
INV_X4 inst_13065 ( .ZN(net_16380), .A(net_16339) );
SDFF_X2 inst_796 ( .Q(net_20915), .SE(net_18847), .SI(net_18007), .D(net_730), .CK(net_21276) );
INV_X4 inst_14135 ( .ZN(net_9660), .A(net_6093) );
INV_X4 inst_16253 ( .A(net_3836), .ZN(net_1911) );
NAND2_X2 inst_11727 ( .ZN(net_3179), .A1(net_2230), .A2(net_1212) );
CLKBUF_X2 inst_21425 ( .A(net_21296), .Z(net_21297) );
NAND3_X2 inst_6699 ( .ZN(net_20698), .A1(net_7396), .A2(net_7395), .A3(net_2058) );
NAND2_X4 inst_7628 ( .A1(net_1662), .ZN(net_1544), .A2(net_1216) );
INV_X4 inst_15030 ( .ZN(net_13752), .A(net_13444) );
OAI21_X4 inst_1499 ( .ZN(net_11319), .A(net_11318), .B2(net_11317), .B1(net_9647) );
NOR2_X4 inst_2972 ( .ZN(net_9812), .A1(net_3991), .A2(net_3333) );
NAND2_X2 inst_9470 ( .ZN(net_13766), .A2(net_10871), .A1(net_5499) );
INV_X4 inst_15554 ( .A(net_3292), .ZN(net_2558) );
NAND2_X2 inst_9293 ( .ZN(net_20599), .A1(net_12409), .A2(net_12408) );
INV_X8 inst_12345 ( .ZN(net_4737), .A(net_4208) );
NOR2_X4 inst_3297 ( .ZN(net_1679), .A2(net_1027), .A1(net_938) );
NAND3_X2 inst_5931 ( .ZN(net_14928), .A2(net_14927), .A1(net_13631), .A3(net_12494) );
NAND4_X2 inst_5429 ( .ZN(net_14114), .A4(net_11312), .A2(net_8436), .A1(net_8379), .A3(net_8288) );
INV_X2 inst_18823 ( .A(net_9099), .ZN(net_6892) );
INV_X4 inst_12556 ( .ZN(net_18363), .A(net_18315) );
NOR2_X2 inst_4423 ( .ZN(net_6114), .A2(net_4849), .A1(net_1102) );
NAND2_X2 inst_10438 ( .A1(net_11443), .A2(net_7235), .ZN(net_7195) );
INV_X4 inst_13384 ( .ZN(net_13716), .A(net_10769) );
NAND2_X2 inst_11880 ( .ZN(net_3020), .A2(net_1619), .A1(net_1190) );
NOR2_X2 inst_4342 ( .ZN(net_7608), .A2(net_3308), .A1(net_409) );
INV_X4 inst_15691 ( .A(net_2044), .ZN(net_2025) );
NAND2_X2 inst_8664 ( .A1(net_21171), .ZN(net_16477), .A2(net_16476) );
NAND2_X2 inst_10398 ( .ZN(net_12105), .A2(net_7283), .A1(net_5733) );
INV_X4 inst_12887 ( .ZN(net_16970), .A(net_16813) );
NOR2_X2 inst_4339 ( .ZN(net_5690), .A1(net_5689), .A2(net_4217) );
NOR2_X2 inst_5060 ( .ZN(net_10377), .A1(net_7268), .A2(net_47) );
INV_X4 inst_17666 ( .ZN(net_2557), .A(net_900) );
INV_X4 inst_14187 ( .ZN(net_8003), .A(net_5981) );
OAI21_X4 inst_1421 ( .B2(net_19078), .B1(net_19077), .A(net_16187), .ZN(net_16109) );
INV_X2 inst_18909 ( .ZN(net_6038), .A(net_6037) );
INV_X4 inst_16836 ( .ZN(net_1563), .A(net_982) );
NOR2_X2 inst_4262 ( .ZN(net_6232), .A2(net_6231), .A1(net_874) );
INV_X4 inst_12819 ( .ZN(net_17193), .A(net_17192) );
NAND2_X2 inst_8298 ( .ZN(net_17605), .A2(net_17414), .A1(net_17412) );
INV_X4 inst_12607 ( .A(net_18083), .ZN(net_18082) );
NAND2_X2 inst_10406 ( .A1(net_20120), .ZN(net_7267), .A2(net_120) );
INV_X4 inst_16283 ( .ZN(net_1455), .A(net_1029) );
CLKBUF_X2 inst_21599 ( .A(net_21383), .Z(net_21471) );
INV_X4 inst_17797 ( .ZN(net_861), .A(net_130) );
INV_X4 inst_17436 ( .A(net_1980), .ZN(net_1619) );
INV_X4 inst_13882 ( .A(net_14348), .ZN(net_8978) );
NOR2_X2 inst_3664 ( .ZN(net_11561), .A1(net_11560), .A2(net_9584) );
NAND2_X2 inst_9688 ( .ZN(net_20673), .A2(net_10245), .A1(net_9169) );
CLKBUF_X2 inst_22893 ( .A(net_22764), .Z(net_22765) );
NAND2_X2 inst_9961 ( .ZN(net_8908), .A2(net_8213), .A1(net_6188) );
NAND3_X2 inst_6011 ( .ZN(net_14422), .A1(net_13473), .A3(net_9998), .A2(net_4044) );
NAND2_X2 inst_10536 ( .ZN(net_6809), .A2(net_6808), .A1(net_5935) );
INV_X2 inst_18437 ( .ZN(net_14311), .A(net_13844) );
INV_X4 inst_17412 ( .A(net_14563), .ZN(net_1006) );
NOR2_X2 inst_3486 ( .ZN(net_14292), .A1(net_14291), .A2(net_13370) );
NAND2_X2 inst_8833 ( .ZN(net_15503), .A2(net_15137), .A1(net_7135) );
INV_X4 inst_13246 ( .ZN(net_12981), .A(net_12048) );
INV_X4 inst_13961 ( .ZN(net_13146), .A(net_6744) );
NAND2_X2 inst_9636 ( .ZN(net_13125), .A1(net_10386), .A2(net_8357) );
INV_X2 inst_19384 ( .ZN(net_2134), .A(net_2133) );
NAND2_X2 inst_8970 ( .ZN(net_14520), .A1(net_14078), .A2(net_12868) );
NAND2_X2 inst_12099 ( .ZN(net_514), .A2(net_513), .A1(net_88) );
INV_X4 inst_13358 ( .ZN(net_12360), .A(net_10954) );
INV_X4 inst_13769 ( .A(net_9610), .ZN(net_7603) );
INV_X2 inst_18987 ( .ZN(net_5117), .A(net_5116) );
NAND3_X2 inst_6628 ( .A3(net_14921), .ZN(net_9038), .A2(net_9037), .A1(net_5617) );
INV_X4 inst_17257 ( .ZN(net_3426), .A(net_2094) );
NAND2_X4 inst_7621 ( .ZN(net_1310), .A1(net_967), .A2(net_207) );
NAND2_X2 inst_10029 ( .ZN(net_20091), .A1(net_15191), .A2(net_8737) );
INV_X4 inst_13877 ( .A(net_7561), .ZN(net_7373) );
XNOR2_X2 inst_230 ( .ZN(net_17454), .A(net_17033), .B(net_283) );
NAND3_X2 inst_5903 ( .ZN(net_15131), .A3(net_13396), .A2(net_11568), .A1(net_9641) );
INV_X4 inst_18022 ( .A(net_20862), .ZN(net_317) );
INV_X2 inst_18982 ( .ZN(net_5143), .A(net_5142) );
INV_X4 inst_16668 ( .ZN(net_1082), .A(net_1081) );
NAND2_X2 inst_10089 ( .A1(net_12885), .ZN(net_8624), .A2(net_7925) );
AOI221_X2 inst_20092 ( .B1(net_15955), .ZN(net_14822), .C1(net_14593), .C2(net_13197), .B2(net_12239), .A(net_11958) );
INV_X4 inst_17337 ( .ZN(net_3748), .A(net_90) );
OAI21_X2 inst_1893 ( .ZN(net_13366), .A(net_10688), .B1(net_9852), .B2(net_8514) );
NOR2_X2 inst_5101 ( .A2(net_20495), .ZN(net_772), .A1(net_115) );
NOR2_X2 inst_4728 ( .A1(net_20488), .ZN(net_3555), .A2(net_3095) );
INV_X4 inst_16074 ( .ZN(net_2481), .A(net_1554) );
AOI222_X2 inst_20064 ( .ZN(net_13672), .A2(net_11510), .C1(net_9378), .B2(net_4663), .C2(net_4069), .B1(net_3906), .A1(net_81) );
NAND3_X2 inst_6480 ( .ZN(net_11248), .A2(net_11247), .A3(net_9838), .A1(net_2799) );
NAND2_X2 inst_8325 ( .A1(net_20775), .ZN(net_17553), .A2(net_17231) );
NOR2_X2 inst_4385 ( .A2(net_20795), .ZN(net_7818), .A1(net_5435) );
AOI21_X4 inst_20193 ( .ZN(net_15137), .B2(net_13325), .A(net_8277), .B1(net_1889) );
AOI22_X4 inst_19955 ( .B2(net_20936), .ZN(net_19020), .A2(net_18601), .A1(net_16333), .B1(net_15923) );
INV_X4 inst_16841 ( .ZN(net_15012), .A(net_7071) );
NOR2_X2 inst_4606 ( .ZN(net_3747), .A2(net_2543), .A1(net_2339) );
INV_X2 inst_18986 ( .ZN(net_5119), .A(net_5118) );
CLKBUF_X2 inst_22510 ( .A(net_21660), .Z(net_22382) );
INV_X4 inst_17782 ( .ZN(net_2214), .A(net_194) );
INV_X2 inst_18472 ( .ZN(net_12680), .A(net_12679) );
XNOR2_X2 inst_452 ( .ZN(net_14415), .B(net_14414), .A(net_11873) );
INV_X4 inst_14375 ( .ZN(net_19210), .A(net_5176) );
INV_X2 inst_18603 ( .ZN(net_9788), .A(net_9787) );
INV_X4 inst_17088 ( .ZN(net_8543), .A(net_877) );
NAND2_X2 inst_10338 ( .A2(net_9698), .A1(net_8961), .ZN(net_7554) );
NAND2_X2 inst_9392 ( .ZN(net_11711), .A2(net_11710), .A1(net_8938) );
INV_X2 inst_19381 ( .A(net_2781), .ZN(net_2145) );
NAND2_X2 inst_8397 ( .ZN(net_17398), .A1(net_16978), .A2(net_16826) );
AOI22_X1 inst_20059 ( .B2(net_3134), .ZN(net_2628), .A1(net_2627), .A2(net_2365), .B1(net_1798) );
NOR2_X4 inst_3061 ( .ZN(net_8070), .A1(net_4950), .A2(net_1566) );
INV_X4 inst_13146 ( .ZN(net_15053), .A(net_14620) );
CLKBUF_X2 inst_22210 ( .A(net_22081), .Z(net_22082) );
NOR2_X2 inst_4144 ( .ZN(net_6913), .A2(net_6883), .A1(net_4869) );
INV_X4 inst_14000 ( .A(net_7937), .ZN(net_7656) );
INV_X4 inst_17953 ( .A(net_21021), .ZN(net_443) );
INV_X4 inst_17710 ( .A(net_20851), .ZN(net_640) );
NAND2_X2 inst_10254 ( .ZN(net_10155), .A2(net_8175), .A1(net_4762) );
SDFF_X2 inst_728 ( .Q(net_20877), .SE(net_18584), .SI(net_18567), .D(net_3582), .CK(net_21919) );
NAND2_X2 inst_11180 ( .A2(net_4136), .ZN(net_4121), .A1(net_2065) );
INV_X4 inst_14308 ( .A(net_10562), .ZN(net_5502) );
NAND2_X2 inst_10372 ( .ZN(net_12507), .A1(net_10031), .A2(net_4576) );
NOR2_X4 inst_3121 ( .ZN(net_6443), .A2(net_4374), .A1(net_3970) );
NOR3_X2 inst_2780 ( .A3(net_8870), .A1(net_8395), .ZN(net_6532), .A2(net_1070) );
AND3_X4 inst_21117 ( .ZN(net_13606), .A2(net_13605), .A3(net_13532), .A1(net_9497) );
INV_X4 inst_15034 ( .A(net_5488), .ZN(net_4898) );
NAND3_X2 inst_6655 ( .ZN(net_8496), .A2(net_8495), .A3(net_8494), .A1(net_5337) );
CLKBUF_X2 inst_21798 ( .A(net_21669), .Z(net_21670) );
INV_X2 inst_18957 ( .ZN(net_5514), .A(net_5513) );
NOR2_X2 inst_4152 ( .A1(net_8709), .ZN(net_6901), .A2(net_5079) );
INV_X4 inst_16325 ( .A(net_7010), .ZN(net_5009) );
AOI21_X4 inst_20121 ( .B1(net_19590), .ZN(net_19067), .B2(net_16214), .A(net_15464) );
NAND2_X2 inst_11031 ( .ZN(net_10255), .A1(net_4762), .A2(net_3499) );
NOR2_X4 inst_2844 ( .ZN(net_14250), .A1(net_12610), .A2(net_11271) );
INV_X2 inst_19178 ( .ZN(net_3795), .A(net_3794) );
OAI211_X2 inst_2492 ( .ZN(net_13158), .C1(net_13157), .C2(net_13156), .A(net_11744), .B(net_8673) );
INV_X4 inst_17046 ( .ZN(net_3900), .A(net_1547) );
AOI21_X2 inst_20603 ( .ZN(net_13760), .B2(net_10951), .A(net_8559), .B1(net_2785) );
NOR2_X2 inst_3582 ( .A1(net_12870), .ZN(net_12682), .A2(net_12681) );
INV_X4 inst_15571 ( .ZN(net_14966), .A(net_14636) );
NOR2_X2 inst_3480 ( .ZN(net_14379), .A1(net_14378), .A2(net_12929) );
INV_X4 inst_14125 ( .ZN(net_7532), .A(net_6121) );
INV_X4 inst_18114 ( .A(net_21098), .ZN(net_719) );
NAND2_X2 inst_11721 ( .A2(net_3045), .ZN(net_2817), .A1(net_2246) );
AOI21_X2 inst_20442 ( .B1(net_15245), .ZN(net_15123), .B2(net_13216), .A(net_12134) );
INV_X2 inst_19662 ( .A(net_20467), .ZN(net_20466) );
CLKBUF_X2 inst_22490 ( .A(net_21533), .Z(net_22362) );
NAND3_X2 inst_5705 ( .A3(net_20013), .A1(net_20012), .ZN(net_16204), .A2(net_14876) );
NAND2_X2 inst_10879 ( .A2(net_12915), .ZN(net_11800), .A1(net_5415) );
CLKBUF_X2 inst_21875 ( .A(net_21746), .Z(net_21747) );
INV_X4 inst_15314 ( .ZN(net_3424), .A(net_2647) );
NAND2_X4 inst_7638 ( .A2(net_1328), .ZN(net_1150), .A1(net_570) );
INV_X4 inst_14776 ( .ZN(net_7723), .A(net_5433) );
NAND2_X4 inst_7093 ( .A2(net_20841), .A1(net_20840), .ZN(net_19358) );
NAND2_X2 inst_11017 ( .A2(net_6053), .ZN(net_5968), .A1(net_5448) );
NOR2_X2 inst_4818 ( .A1(net_3780), .ZN(net_2560), .A2(net_2559) );
NAND2_X2 inst_10381 ( .A1(net_18025), .ZN(net_7385), .A2(net_441) );
AOI211_X2 inst_21009 ( .ZN(net_15776), .B(net_15126), .C2(net_12909), .A(net_8716), .C1(net_5166) );
AOI21_X2 inst_20458 ( .B1(net_15121), .ZN(net_15038), .B2(net_12951), .A(net_10990) );
SDFF_X2 inst_974 ( .QN(net_21013), .D(net_799), .SE(net_263), .CK(net_22729), .SI(x2809) );
AOI21_X2 inst_20584 ( .ZN(net_14034), .A(net_14033), .B1(net_13121), .B2(net_7251) );
DFF_X1 inst_19826 ( .D(net_17678), .CK(net_22117), .Q(x361) );
CLKBUF_X2 inst_22168 ( .A(net_22039), .Z(net_22040) );
INV_X4 inst_17685 ( .ZN(net_930), .A(net_330) );
INV_X2 inst_18700 ( .ZN(net_8302), .A(net_8301) );
CLKBUF_X2 inst_21736 ( .A(net_21607), .Z(net_21608) );
INV_X2 inst_19590 ( .A(net_333), .ZN(net_296) );
SDFF_X2 inst_1001 ( .QN(net_21005), .D(net_2095), .SE(net_263), .CK(net_21890), .SI(x2978) );
AOI21_X2 inst_20520 ( .ZN(net_14564), .B1(net_14563), .B2(net_11976), .A(net_10088) );
INV_X4 inst_17281 ( .ZN(net_639), .A(net_227) );
NAND3_X2 inst_5825 ( .ZN(net_15566), .A2(net_15565), .A1(net_14815), .A3(net_12493) );
NOR2_X4 inst_3033 ( .ZN(net_9832), .A2(net_5169), .A1(net_5131) );
NOR2_X4 inst_2925 ( .ZN(net_11741), .A1(net_10144), .A2(net_7886) );
NAND2_X2 inst_7843 ( .ZN(net_19765), .A2(net_18620), .A1(net_16411) );
NAND2_X2 inst_10537 ( .ZN(net_8771), .A1(net_8724), .A2(net_6842) );
CLKBUF_X2 inst_21456 ( .A(net_21327), .Z(net_21328) );
OAI21_X2 inst_1828 ( .A(net_15362), .ZN(net_14138), .B2(net_10464), .B1(net_9908) );
NAND2_X2 inst_9510 ( .ZN(net_11266), .A2(net_8193), .A1(net_4335) );
NOR2_X2 inst_3388 ( .ZN(net_16189), .A2(net_16016), .A1(net_7931) );
NOR2_X2 inst_3735 ( .ZN(net_10727), .A2(net_10708), .A1(net_5122) );
NAND2_X2 inst_11238 ( .ZN(net_3938), .A2(net_2748), .A1(net_955) );
NAND4_X2 inst_5311 ( .ZN(net_19030), .A4(net_15090), .A1(net_15069), .A3(net_13266), .A2(net_13041) );
NOR3_X2 inst_2675 ( .ZN(net_14803), .A2(net_14802), .A3(net_13424), .A1(net_5191) );
INV_X4 inst_18115 ( .A(net_21005), .ZN(net_2095) );
XNOR2_X2 inst_141 ( .ZN(net_18173), .A(net_18095), .B(net_9173) );
OAI211_X2 inst_2520 ( .ZN(net_11875), .B(net_11874), .C1(net_9487), .A(net_6810), .C2(net_4645) );
NAND2_X2 inst_10578 ( .ZN(net_8702), .A2(net_6594), .A1(net_5984) );
AOI21_X2 inst_20329 ( .ZN(net_15828), .B1(net_15827), .B2(net_15273), .A(net_14931) );
XNOR2_X2 inst_571 ( .ZN(net_633), .A(net_632), .B(net_631) );
INV_X4 inst_16405 ( .ZN(net_8839), .A(net_906) );
NAND3_X2 inst_6007 ( .A2(net_20827), .A1(net_20826), .A3(net_20237), .ZN(net_19957) );
OAI21_X2 inst_1974 ( .ZN(net_12198), .A(net_8596), .B2(net_7799), .B1(net_4536) );
OAI21_X2 inst_2017 ( .ZN(net_11367), .A(net_11366), .B1(net_11365), .B2(net_7006) );
OR2_X2 inst_1154 ( .A2(net_12233), .ZN(net_10350), .A1(net_8981) );
INV_X4 inst_14901 ( .ZN(net_5895), .A(net_3606) );
INV_X4 inst_16267 ( .ZN(net_2305), .A(net_1672) );
NAND2_X2 inst_7728 ( .ZN(net_18826), .A1(net_18792), .A2(net_18774) );
INV_X8 inst_12413 ( .A(net_20941), .ZN(net_1271) );
NAND2_X2 inst_9584 ( .ZN(net_10921), .A1(net_10920), .A2(net_10919) );
CLKBUF_X2 inst_22132 ( .A(net_21746), .Z(net_22004) );
INV_X4 inst_16339 ( .ZN(net_1799), .A(net_1753) );
NAND2_X4 inst_7224 ( .ZN(net_11091), .A1(net_5839), .A2(net_4253) );
XNOR2_X2 inst_469 ( .ZN(net_12269), .B(net_12268), .A(net_7652) );
NAND2_X4 inst_7468 ( .ZN(net_4387), .A1(net_2668), .A2(net_391) );
NAND2_X2 inst_8598 ( .A1(net_21166), .A2(net_19448), .ZN(net_19262) );
NAND2_X4 inst_7133 ( .ZN(net_14541), .A1(net_9615), .A2(net_8311) );
NAND2_X4 inst_6837 ( .A2(net_18723), .ZN(net_18719), .A1(net_18718) );
INV_X4 inst_15013 ( .ZN(net_14755), .A(net_10141) );
INV_X4 inst_16919 ( .ZN(net_1135), .A(net_936) );
NAND2_X2 inst_8866 ( .ZN(net_15326), .A2(net_14501), .A1(net_10859) );
DFF_X1 inst_19928 ( .D(net_2525), .CK(net_22765), .Q(x1330) );
NAND3_X2 inst_6642 ( .ZN(net_8946), .A3(net_8945), .A1(net_5428), .A2(net_3549) );
NAND3_X2 inst_6507 ( .ZN(net_10793), .A3(net_10792), .A1(net_5647), .A2(net_3363) );
OAI21_X2 inst_2339 ( .ZN(net_4679), .B2(net_3675), .B1(net_3538), .A(net_2121) );
INV_X2 inst_18911 ( .A(net_8187), .ZN(net_6032) );
INV_X8 inst_12300 ( .ZN(net_4042), .A(net_950) );
AOI21_X2 inst_20581 ( .B2(net_20641), .B1(net_20640), .ZN(net_14077), .A(net_10686) );
INV_X2 inst_18692 ( .A(net_10655), .ZN(net_8375) );
NAND2_X2 inst_11603 ( .A1(net_3491), .ZN(net_2653), .A2(net_2413) );
OR2_X2 inst_1216 ( .ZN(net_12500), .A2(net_2940), .A1(net_2076) );
NAND2_X2 inst_8260 ( .ZN(net_17689), .A2(net_17665), .A1(net_17399) );
NAND3_X2 inst_6697 ( .ZN(net_7666), .A3(net_7665), .A2(net_6130), .A1(net_2812) );
INV_X4 inst_15544 ( .ZN(net_9925), .A(net_6626) );
INV_X4 inst_17019 ( .A(net_13089), .ZN(net_852) );
SDFF_X2 inst_952 ( .QN(net_21090), .SE(net_17277), .D(net_676), .CK(net_21787), .SI(x1551) );
INV_X2 inst_18833 ( .ZN(net_6771), .A(net_6770) );
INV_X4 inst_16069 ( .ZN(net_2442), .A(net_1239) );
NAND3_X2 inst_5972 ( .ZN(net_19511), .A1(net_14149), .A3(net_13060), .A2(net_8652) );
AOI211_X2 inst_21069 ( .ZN(net_7699), .B(net_6433), .C2(net_4624), .A(net_4508), .C1(net_2107) );
NAND2_X4 inst_7254 ( .A1(net_19816), .ZN(net_8029), .A2(net_6736) );
CLKBUF_X2 inst_22912 ( .A(net_22783), .Z(net_22784) );
AOI21_X2 inst_20338 ( .B1(net_15831), .ZN(net_15792), .B2(net_14810), .A(net_11905) );
CLKBUF_X2 inst_21680 ( .A(net_21551), .Z(net_21552) );
INV_X4 inst_14710 ( .ZN(net_20647), .A(net_5370) );
SDFF_X2 inst_721 ( .Q(net_20905), .SE(net_18858), .SI(net_18587), .D(net_11881), .CK(net_21869) );
NAND2_X2 inst_11135 ( .ZN(net_6591), .A2(net_2308), .A1(net_222) );
NAND2_X4 inst_7211 ( .ZN(net_11878), .A2(net_7892), .A1(net_7790) );
NAND2_X2 inst_10838 ( .ZN(net_8886), .A1(net_5479), .A2(net_4053) );
CLKBUF_X2 inst_22576 ( .A(net_22447), .Z(net_22448) );
CLKBUF_X2 inst_22715 ( .A(net_22586), .Z(net_22587) );
CLKBUF_X2 inst_21953 ( .A(net_21824), .Z(net_21825) );
NOR2_X4 inst_3009 ( .ZN(net_8080), .A1(net_3476), .A2(net_270) );
OAI21_X4 inst_1366 ( .B1(net_21113), .ZN(net_17843), .B2(net_17675), .A(net_17583) );
INV_X4 inst_13667 ( .ZN(net_11959), .A(net_8062) );
INV_X4 inst_13079 ( .ZN(net_16190), .A(net_16120) );
AOI21_X4 inst_20253 ( .B2(net_20441), .ZN(net_6501), .B1(net_1569), .A(net_196) );
INV_X4 inst_17675 ( .A(net_255), .ZN(net_241) );
CLKBUF_X2 inst_22235 ( .A(net_22106), .Z(net_22107) );
OAI21_X2 inst_1915 ( .A(net_15077), .ZN(net_13064), .B1(net_11534), .B2(net_5809) );
NOR3_X2 inst_2794 ( .A2(net_9387), .ZN(net_3445), .A1(net_2427), .A3(net_1004) );
OAI22_X2 inst_1254 ( .A2(net_17876), .B2(net_17875), .ZN(net_17833), .A1(net_8997), .B1(net_5724) );
NAND2_X4 inst_7111 ( .A2(net_20551), .ZN(net_13768), .A1(net_10872) );
NOR2_X2 inst_3553 ( .ZN(net_13060), .A2(net_12308), .A1(net_10232) );
INV_X4 inst_14031 ( .ZN(net_7628), .A(net_6277) );
INV_X4 inst_14412 ( .A(net_6862), .ZN(net_5094) );
CLKBUF_X2 inst_22247 ( .A(net_21300), .Z(net_22119) );
OAI21_X2 inst_1811 ( .ZN(net_19674), .B2(net_12250), .A(net_10683), .B1(net_8092) );
NOR2_X2 inst_4544 ( .ZN(net_11113), .A1(net_4711), .A2(net_4041) );
NAND2_X2 inst_11147 ( .ZN(net_5275), .A1(net_4481), .A2(net_2688) );
NAND2_X2 inst_11351 ( .ZN(net_4871), .A1(net_3645), .A2(net_2537) );
INV_X4 inst_14479 ( .ZN(net_5823), .A(net_3519) );
CLKBUF_X2 inst_21884 ( .A(net_21510), .Z(net_21756) );
NAND2_X2 inst_10801 ( .ZN(net_10534), .A2(net_5553), .A1(net_2585) );
NAND2_X4 inst_7054 ( .A2(net_19356), .A1(net_19355), .ZN(net_16451) );
INV_X4 inst_18075 ( .A(net_20886), .ZN(net_203) );
INV_X4 inst_14834 ( .ZN(net_4853), .A(net_3037) );
AOI22_X2 inst_20028 ( .ZN(net_9927), .A1(net_9926), .B1(net_9925), .A2(net_8207), .B2(net_3443) );
NAND2_X2 inst_8826 ( .A1(net_20165), .ZN(net_19598), .A2(net_15697) );
XNOR2_X2 inst_163 ( .ZN(net_17898), .A(net_17770), .B(net_679) );
NAND2_X2 inst_9156 ( .A1(net_13416), .ZN(net_13387), .A2(net_10441) );
CLKBUF_X2 inst_21779 ( .A(net_21650), .Z(net_21651) );
XNOR2_X2 inst_394 ( .ZN(net_16765), .A(net_16764), .B(net_14918) );
NAND2_X2 inst_8455 ( .ZN(net_17185), .A2(net_16741), .A1(net_16600) );
CLKBUF_X2 inst_21756 ( .A(net_21627), .Z(net_21628) );
NAND2_X2 inst_11619 ( .ZN(net_5189), .A1(net_2917), .A2(net_2842) );
INV_X2 inst_18978 ( .ZN(net_5159), .A(net_5158) );
INV_X4 inst_17678 ( .ZN(net_1660), .A(net_307) );
INV_X4 inst_16268 ( .ZN(net_1488), .A(net_1348) );
OAI21_X2 inst_1814 ( .ZN(net_14172), .B2(net_10697), .B1(net_9753), .A(net_816) );
AOI22_X2 inst_19957 ( .ZN(net_16349), .B1(net_16287), .A2(net_16104), .A1(net_15369), .B2(net_14985) );
NOR2_X2 inst_4470 ( .ZN(net_4426), .A1(net_3890), .A2(net_3486) );
INV_X4 inst_17392 ( .A(net_2094), .ZN(net_818) );
NAND2_X2 inst_10875 ( .A1(net_10512), .A2(net_5436), .ZN(net_5425) );
XNOR2_X2 inst_361 ( .A(net_20213), .B(net_17247), .ZN(net_16884) );
CLKBUF_X2 inst_22645 ( .A(net_22157), .Z(net_22517) );
CLKBUF_X2 inst_22173 ( .A(net_22044), .Z(net_22045) );
AOI21_X2 inst_20347 ( .A(net_21236), .ZN(net_15757), .B2(net_15021), .B1(net_12183) );
NAND2_X2 inst_11358 ( .ZN(net_3616), .A2(net_3467), .A1(net_1757) );
AOI21_X2 inst_20734 ( .B1(net_12298), .ZN(net_11738), .B2(net_11737), .A(net_9182) );
NOR2_X2 inst_3400 ( .ZN(net_15849), .A2(net_15421), .A1(net_15199) );
NAND2_X2 inst_8127 ( .A2(net_20912), .ZN(net_18052), .A1(net_15896) );
CLKBUF_X2 inst_22464 ( .A(net_22335), .Z(net_22336) );
NAND2_X1 inst_12134 ( .ZN(net_18189), .A1(net_18183), .A2(net_2400) );
NAND2_X2 inst_8082 ( .ZN(net_19001), .A2(net_18153), .A1(net_18118) );
INV_X2 inst_19056 ( .ZN(net_4725), .A(net_4724) );
NAND2_X2 inst_11008 ( .ZN(net_19332), .A2(net_4877), .A1(net_3297) );
INV_X4 inst_14852 ( .A(net_5419), .ZN(net_4818) );
SDFF_X2 inst_786 ( .Q(net_20945), .SE(net_18804), .SI(net_18039), .D(net_480), .CK(net_21282) );
XOR2_X2 inst_2 ( .Z(net_18194), .B(net_18093), .A(net_1943) );
NAND2_X2 inst_11003 ( .A1(net_9325), .ZN(net_4887), .A2(net_2706) );
CLKBUF_X2 inst_21981 ( .A(net_21852), .Z(net_21853) );
AOI22_X2 inst_19985 ( .ZN(net_15204), .A1(net_14600), .A2(net_14114), .B2(net_11291), .B1(net_5372) );
SDFF_X2 inst_888 ( .Q(net_21135), .SI(net_16881), .SE(net_125), .CK(net_21647), .D(x3791) );
INV_X2 inst_19688 ( .A(net_20533), .ZN(net_20532) );
OAI21_X2 inst_1769 ( .B2(net_20109), .B1(net_20108), .ZN(net_14696), .A(net_11771) );
INV_X8 inst_12306 ( .ZN(net_1669), .A(net_760) );
NAND3_X2 inst_5999 ( .ZN(net_14434), .A1(net_12721), .A3(net_12548), .A2(net_11618) );
NOR2_X2 inst_3625 ( .ZN(net_13577), .A1(net_12658), .A2(net_9157) );
INV_X2 inst_19356 ( .ZN(net_2360), .A(net_2359) );
NAND3_X2 inst_6598 ( .A3(net_20333), .ZN(net_9901), .A1(net_9900), .A2(net_4024) );
NAND3_X2 inst_5979 ( .ZN(net_14606), .A1(net_13249), .A2(net_13196), .A3(net_12788) );
INV_X4 inst_15896 ( .ZN(net_15694), .A(net_14694) );
NAND2_X2 inst_7817 ( .ZN(net_18672), .A1(net_18636), .A2(net_18621) );
OAI211_X2 inst_2581 ( .ZN(net_7674), .A(net_6332), .B(net_3794), .C2(net_1875), .C1(net_1032) );
NOR2_X2 inst_4110 ( .ZN(net_7086), .A1(net_4317), .A2(net_4254) );
OAI21_X2 inst_2164 ( .A(net_15499), .ZN(net_9029), .B2(net_9028), .B1(net_5409) );
INV_X4 inst_17112 ( .A(net_15113), .ZN(net_15107) );
INV_X4 inst_16618 ( .ZN(net_8330), .A(net_5766) );
NAND2_X4 inst_7198 ( .ZN(net_12099), .A2(net_8250), .A1(net_143) );
INV_X4 inst_13208 ( .ZN(net_13726), .A(net_12985) );
NOR2_X2 inst_4392 ( .ZN(net_20398), .A1(net_12295), .A2(net_5198) );
NAND2_X2 inst_11696 ( .A1(net_4052), .ZN(net_2772), .A2(net_2317) );
NAND2_X2 inst_11093 ( .A2(net_20579), .ZN(net_5442), .A1(net_4737) );
NOR2_X2 inst_4915 ( .ZN(net_2575), .A2(net_1905), .A1(net_167) );
NAND2_X2 inst_8590 ( .A1(net_17091), .A2(net_16935), .ZN(net_16710) );
INV_X4 inst_14424 ( .ZN(net_6184), .A(net_5047) );
INV_X4 inst_15758 ( .A(net_15842), .ZN(net_1930) );
NAND2_X2 inst_8530 ( .ZN(net_20063), .A1(net_17019), .A2(net_16866) );
NAND2_X2 inst_9655 ( .ZN(net_10344), .A2(net_10343), .A1(net_4004) );
CLKBUF_X2 inst_22632 ( .A(net_22503), .Z(net_22504) );
NAND2_X2 inst_11245 ( .A2(net_5579), .A1(net_4794), .ZN(net_3925) );
INV_X4 inst_16276 ( .ZN(net_8328), .A(net_70) );
INV_X4 inst_16926 ( .ZN(net_10515), .A(net_8664) );
INV_X4 inst_17385 ( .ZN(net_3645), .A(net_252) );
NOR2_X2 inst_3385 ( .ZN(net_20287), .A2(net_16157), .A1(net_16155) );
OAI21_X2 inst_1572 ( .A(net_20960), .B2(net_20162), .B1(net_20161), .ZN(net_16358) );
CLKBUF_X2 inst_22511 ( .A(net_22382), .Z(net_22383) );
NAND2_X2 inst_11753 ( .ZN(net_4219), .A2(net_1136), .A1(net_447) );
NOR2_X2 inst_4906 ( .A2(net_4773), .ZN(net_3472), .A1(net_3184) );
INV_X4 inst_16550 ( .A(net_2744), .ZN(net_1409) );
INV_X4 inst_14932 ( .ZN(net_7755), .A(net_3541) );
CLKBUF_X2 inst_21960 ( .A(net_21601), .Z(net_21832) );
INV_X4 inst_14815 ( .ZN(net_9738), .A(net_3936) );
AND2_X4 inst_21183 ( .ZN(net_18959), .A1(net_15694), .A2(net_11546) );
INV_X4 inst_15634 ( .ZN(net_3439), .A(net_3122) );
INV_X4 inst_14026 ( .ZN(net_11124), .A(net_8120) );
NAND2_X2 inst_10221 ( .ZN(net_8084), .A2(net_4614), .A1(net_866) );
NOR2_X2 inst_4978 ( .ZN(net_3087), .A2(net_1542), .A1(net_170) );
INV_X2 inst_18608 ( .ZN(net_11489), .A(net_10221) );
NAND2_X2 inst_7875 ( .ZN(net_18537), .A1(net_18484), .A2(net_18455) );
INV_X2 inst_18787 ( .ZN(net_9167), .A(net_7497) );
INV_X2 inst_19418 ( .ZN(net_1880), .A(net_1879) );
NAND2_X2 inst_9721 ( .ZN(net_19815), .A2(net_10155), .A1(net_7084) );
AND2_X4 inst_21191 ( .A1(net_13192), .ZN(net_10748), .A2(net_10747) );
NAND2_X2 inst_12048 ( .ZN(net_6495), .A1(net_508), .A2(net_222) );
NOR2_X2 inst_4367 ( .A1(net_6849), .ZN(net_6093), .A2(net_5490) );
NAND2_X2 inst_10346 ( .ZN(net_11012), .A1(net_5157), .A2(net_4539) );
NAND2_X2 inst_7712 ( .ZN(net_18853), .A2(net_18828), .A1(net_17922) );
OAI21_X2 inst_1731 ( .ZN(net_15081), .B2(net_12863), .B1(net_8012), .A(net_1915) );
INV_X2 inst_19327 ( .ZN(net_5195), .A(net_2564) );
INV_X4 inst_16631 ( .ZN(net_7078), .A(net_1110) );
AND2_X2 inst_21310 ( .ZN(net_8715), .A1(net_8714), .A2(net_8713) );
NAND2_X2 inst_7960 ( .ZN(net_18388), .A2(net_18351), .A1(net_17267) );
NOR2_X4 inst_2960 ( .ZN(net_7879), .A1(net_6613), .A2(net_6612) );
OAI21_X2 inst_1909 ( .ZN(net_13092), .A(net_13091), .B2(net_9708), .B1(net_6816) );
INV_X4 inst_16674 ( .ZN(net_15121), .A(net_843) );
NAND3_X2 inst_6616 ( .ZN(net_9068), .A1(net_8091), .A3(net_6966), .A2(net_5994) );
NOR2_X2 inst_4318 ( .ZN(net_9354), .A1(net_7487), .A2(net_3556) );
NAND2_X2 inst_11080 ( .ZN(net_10608), .A1(net_4457), .A2(net_3969) );
NAND2_X2 inst_11669 ( .ZN(net_3191), .A1(net_2331), .A2(net_367) );
NAND2_X2 inst_7991 ( .ZN(net_18323), .A2(net_18270), .A1(net_18230) );
NAND2_X2 inst_9063 ( .ZN(net_13990), .A1(net_13544), .A2(net_11992) );
CLKBUF_X2 inst_22843 ( .A(net_22714), .Z(net_22715) );
NAND2_X4 inst_7455 ( .ZN(net_3764), .A2(net_2981), .A1(net_874) );
NAND2_X2 inst_8443 ( .ZN(net_20158), .A1(net_19441), .A2(net_16451) );
INV_X4 inst_16047 ( .ZN(net_2676), .A(net_1690) );
NOR2_X4 inst_3161 ( .ZN(net_4102), .A1(net_3242), .A2(net_3159) );
INV_X4 inst_14908 ( .ZN(net_6040), .A(net_2391) );
NAND2_X2 inst_10032 ( .ZN(net_10198), .A1(net_8732), .A2(net_8731) );
NAND2_X2 inst_11462 ( .ZN(net_3190), .A1(net_1341), .A2(net_1312) );
NOR2_X4 inst_2816 ( .ZN(net_16786), .A1(net_16419), .A2(net_16369) );
XNOR2_X2 inst_276 ( .B(net_21182), .ZN(net_17188), .A(net_17187) );
INV_X2 inst_18640 ( .ZN(net_12859), .A(net_9380) );
INV_X4 inst_13380 ( .ZN(net_12241), .A(net_10787) );
INV_X2 inst_19337 ( .ZN(net_3269), .A(net_2469) );
NOR2_X2 inst_3339 ( .ZN(net_20691), .A2(net_18824), .A1(net_17164) );
NOR2_X2 inst_3791 ( .ZN(net_10079), .A1(net_6681), .A2(net_6335) );
INV_X2 inst_19296 ( .ZN(net_2805), .A(net_2804) );
CLKBUF_X2 inst_21673 ( .A(net_21544), .Z(net_21545) );
NAND4_X2 inst_5297 ( .ZN(net_19519), .A4(net_15352), .A1(net_15068), .A3(net_14405), .A2(net_13755) );
XNOR2_X2 inst_91 ( .ZN(net_18554), .A(net_18464), .B(net_18300) );
CLKBUF_X2 inst_22119 ( .A(net_21768), .Z(net_21991) );
OAI21_X2 inst_1762 ( .ZN(net_14707), .A(net_14706), .B1(net_12757), .B2(net_12162) );
OAI21_X2 inst_2023 ( .A(net_13544), .ZN(net_11328), .B2(net_6974), .B1(net_5559) );
NOR3_X2 inst_2779 ( .ZN(net_7372), .A2(net_4428), .A1(net_3314), .A3(net_1247) );
NAND3_X2 inst_6508 ( .ZN(net_10791), .A3(net_10790), .A2(net_6663), .A1(net_5634) );
NOR2_X2 inst_4919 ( .A2(net_7156), .ZN(net_1882), .A1(net_1337) );
INV_X4 inst_13250 ( .ZN(net_12793), .A(net_11797) );
INV_X1 inst_19758 ( .A(net_7009), .ZN(net_5164) );
NAND2_X4 inst_7424 ( .A1(net_19175), .ZN(net_5894), .A2(net_2292) );
NOR2_X2 inst_4715 ( .A1(net_4037), .ZN(net_3137), .A2(net_2210) );
INV_X4 inst_17622 ( .A(net_20897), .ZN(net_14483) );
INV_X2 inst_18625 ( .ZN(net_9556), .A(net_9555) );
INV_X2 inst_19703 ( .A(net_20567), .ZN(net_20566) );
NAND3_X2 inst_6648 ( .ZN(net_8558), .A2(net_6742), .A3(net_4397), .A1(net_3826) );
NAND2_X2 inst_11897 ( .ZN(net_2396), .A2(net_1083), .A1(net_880) );
INV_X4 inst_14079 ( .ZN(net_9437), .A(net_6220) );
INV_X4 inst_16398 ( .ZN(net_13495), .A(net_11461) );
NAND2_X2 inst_8851 ( .ZN(net_19915), .A2(net_14701), .A1(net_14513) );
CLKBUF_X2 inst_21721 ( .A(net_21592), .Z(net_21593) );
NAND2_X2 inst_8075 ( .A2(net_20794), .ZN(net_18160), .A1(net_17443) );
INV_X4 inst_17394 ( .A(net_1922), .ZN(net_1356) );
CLKBUF_X2 inst_22143 ( .A(net_21901), .Z(net_22015) );
NAND3_X2 inst_6415 ( .A3(net_19896), .ZN(net_11949), .A1(net_11948), .A2(net_10618) );
NAND2_X2 inst_11187 ( .ZN(net_5311), .A2(net_3861), .A1(net_2889) );
NAND4_X4 inst_5161 ( .A4(net_18953), .A1(net_18952), .ZN(net_18107), .A3(net_14943), .A2(net_12173) );
INV_X2 inst_18803 ( .A(net_9509), .ZN(net_7413) );
INV_X2 inst_18813 ( .A(net_9764), .ZN(net_7316) );
INV_X4 inst_16754 ( .A(net_10417), .ZN(net_1810) );
NAND2_X2 inst_7984 ( .A2(net_18339), .ZN(net_18333), .A1(net_17157) );
NAND3_X2 inst_6489 ( .A2(net_11811), .ZN(net_11170), .A3(net_8919), .A1(net_3885) );
XNOR2_X2 inst_266 ( .ZN(net_17252), .A(net_16754), .B(net_147) );
OAI21_X2 inst_2051 ( .ZN(net_10851), .A(net_7593), .B2(net_4854), .B1(net_1731) );
NAND2_X2 inst_9288 ( .ZN(net_12529), .A1(net_12528), .A2(net_9331) );
NAND2_X2 inst_8382 ( .ZN(net_17342), .A2(net_17341), .A1(net_17078) );
INV_X2 inst_18766 ( .ZN(net_7602), .A(net_7601) );
CLKBUF_X2 inst_21767 ( .A(net_21638), .Z(net_21639) );
INV_X4 inst_17276 ( .ZN(net_13437), .A(net_278) );
OR2_X2 inst_1198 ( .A1(net_8563), .A2(net_6439), .ZN(net_3855) );
XNOR2_X2 inst_171 ( .A(net_17876), .ZN(net_17821), .B(net_17820) );
INV_X4 inst_17835 ( .ZN(net_327), .A(net_279) );
INV_X2 inst_19543 ( .ZN(net_19844), .A(net_4093) );
NAND2_X2 inst_10950 ( .ZN(net_5105), .A2(net_5104), .A1(net_1983) );
XNOR2_X2 inst_374 ( .B(net_21160), .ZN(net_16990), .A(net_16843) );
INV_X4 inst_18023 ( .A(net_21075), .ZN(net_568) );
XNOR2_X2 inst_103 ( .ZN(net_18532), .A(net_18423), .B(net_17569) );
INV_X4 inst_12832 ( .ZN(net_17137), .A(net_17136) );
INV_X4 inst_14864 ( .ZN(net_6695), .A(net_3764) );
NOR2_X2 inst_3690 ( .ZN(net_20110), .A2(net_9589), .A1(net_6915) );
INV_X4 inst_17372 ( .ZN(net_911), .A(net_703) );
NAND2_X2 inst_10763 ( .A1(net_7659), .ZN(net_5647), .A2(net_5646) );
NAND3_X2 inst_6353 ( .A3(net_12284), .ZN(net_12098), .A1(net_8164), .A2(net_6340) );
NAND3_X2 inst_6061 ( .ZN(net_14184), .A3(net_14183), .A1(net_6400), .A2(net_2542) );
NAND2_X2 inst_11716 ( .ZN(net_9085), .A1(net_4715), .A2(net_3208) );
NAND2_X2 inst_9905 ( .ZN(net_11437), .A2(net_9363), .A1(net_731) );
NOR2_X2 inst_3738 ( .ZN(net_10717), .A1(net_10716), .A2(net_10715) );
NOR2_X4 inst_2855 ( .ZN(net_12615), .A1(net_12614), .A2(net_10274) );
NAND2_X2 inst_8247 ( .ZN(net_17716), .A2(net_17715), .A1(net_17046) );
AND4_X2 inst_21107 ( .A1(net_13164), .A3(net_12800), .ZN(net_11732), .A4(net_11731), .A2(net_11040) );
NAND3_X2 inst_6749 ( .A2(net_7844), .ZN(net_5796), .A3(net_3062), .A1(net_2022) );
NAND2_X2 inst_10097 ( .ZN(net_13171), .A2(net_7882), .A1(net_7253) );
CLKBUF_X2 inst_22018 ( .A(net_21264), .Z(net_21890) );
INV_X2 inst_19202 ( .ZN(net_6071), .A(net_3568) );
OAI21_X2 inst_2058 ( .ZN(net_10703), .A(net_10702), .B1(net_10701), .B2(net_6903) );
SDFF_X2 inst_809 ( .Q(net_20848), .SE(net_18804), .SI(net_17949), .D(net_390), .CK(net_22607) );
INV_X2 inst_19107 ( .A(net_7714), .ZN(net_4488) );
INV_X4 inst_16609 ( .A(net_9571), .ZN(net_6346) );
NOR2_X2 inst_3675 ( .ZN(net_11471), .A2(net_11470), .A1(net_8188) );
INV_X4 inst_15821 ( .ZN(net_4491), .A(net_1871) );
NAND2_X2 inst_7816 ( .ZN(net_18662), .A1(net_18661), .A2(net_17436) );
OAI211_X2 inst_2562 ( .C1(net_10659), .ZN(net_9908), .C2(net_8901), .A(net_5794), .B(net_3921) );
INV_X4 inst_14245 ( .ZN(net_5774), .A(net_5242) );
SDFF_X2 inst_1022 ( .QN(net_21078), .D(net_378), .SE(net_263), .CK(net_22563), .SI(x1747) );
INV_X4 inst_13925 ( .A(net_14384), .ZN(net_8642) );
INV_X4 inst_15054 ( .ZN(net_19671), .A(net_3312) );
NAND2_X2 inst_9248 ( .ZN(net_12670), .A1(net_12669), .A2(net_10985) );
CLKBUF_X2 inst_21409 ( .A(net_21280), .Z(net_21281) );
AND2_X2 inst_21270 ( .ZN(net_19021), .A2(net_12729), .A1(net_12680) );
INV_X4 inst_16876 ( .ZN(net_1173), .A(net_308) );
NAND2_X2 inst_10416 ( .A1(net_9921), .ZN(net_7243), .A2(net_7203) );
NAND3_X2 inst_6241 ( .ZN(net_13193), .A2(net_13192), .A3(net_12168), .A1(net_7209) );
NOR2_X2 inst_3906 ( .ZN(net_13823), .A1(net_13700), .A2(net_8876) );
NAND2_X2 inst_8928 ( .ZN(net_14862), .A2(net_14093), .A1(net_11674) );
NAND2_X2 inst_8657 ( .A2(net_19449), .ZN(net_19263), .A1(net_16759) );
INV_X2 inst_19187 ( .ZN(net_3722), .A(net_3721) );
NAND2_X2 inst_9322 ( .ZN(net_12327), .A1(net_12326), .A2(net_9067) );
INV_X4 inst_15103 ( .A(net_11432), .ZN(net_9263) );
NAND2_X2 inst_10665 ( .ZN(net_9795), .A2(net_6346), .A1(net_6255) );
INV_X4 inst_16804 ( .ZN(net_9324), .A(net_3886) );
NOR2_X4 inst_2915 ( .ZN(net_10284), .A2(net_8190), .A1(net_8189) );
INV_X4 inst_17387 ( .ZN(net_8224), .A(net_895) );
NOR2_X4 inst_3296 ( .A1(net_2788), .ZN(net_2141), .A2(net_85) );
CLKBUF_X2 inst_22852 ( .A(net_21423), .Z(net_22724) );
INV_X4 inst_18129 ( .A(net_21082), .ZN(net_473) );
NAND3_X2 inst_6148 ( .ZN(net_19776), .A3(net_12742), .A2(net_10959), .A1(net_8606) );
NAND2_X2 inst_9135 ( .ZN(net_13470), .A2(net_10670), .A1(net_3968) );
INV_X4 inst_14792 ( .ZN(net_4005), .A(net_4004) );
NAND3_X2 inst_6379 ( .ZN(net_12034), .A3(net_12033), .A2(net_4298), .A1(net_3528) );
XNOR2_X2 inst_532 ( .A(net_15957), .ZN(net_2401), .B(net_2400) );
NOR2_X4 inst_3164 ( .A2(net_20868), .ZN(net_3202), .A1(net_3111) );
NOR2_X4 inst_2965 ( .A1(net_9692), .ZN(net_7821), .A2(net_6570) );
OAI211_X4 inst_2382 ( .ZN(net_14135), .C1(net_12231), .C2(net_9896), .B(net_7980), .A(net_7089) );
INV_X8 inst_12228 ( .ZN(net_5176), .A(net_3202) );
NOR2_X4 inst_2969 ( .ZN(net_11151), .A1(net_6394), .A2(net_5357) );
AOI211_X2 inst_21076 ( .C1(net_12238), .ZN(net_7352), .B(net_7351), .A(net_7080), .C2(net_4357) );
NOR2_X4 inst_3314 ( .A2(net_1533), .ZN(net_1162), .A1(net_700) );
CLKBUF_X2 inst_21600 ( .A(net_21471), .Z(net_21472) );
INV_X4 inst_14854 ( .A(net_3822), .ZN(net_3821) );
INV_X4 inst_15891 ( .ZN(net_13080), .A(net_1777) );
NOR2_X2 inst_4037 ( .A1(net_13785), .ZN(net_7931), .A2(net_7930) );
INV_X4 inst_15294 ( .ZN(net_5170), .A(net_2090) );
INV_X4 inst_13277 ( .ZN(net_12451), .A(net_11176) );
OAI221_X4 inst_1327 ( .B1(net_20042), .ZN(net_14758), .B2(net_14185), .C1(net_14175), .C2(net_10527), .A(net_7349) );
NAND2_X2 inst_12073 ( .ZN(net_1250), .A2(net_958), .A1(net_459) );
INV_X4 inst_13566 ( .ZN(net_10711), .A(net_9137) );
NAND2_X2 inst_10598 ( .ZN(net_11964), .A2(net_4813), .A1(net_4250) );
NAND2_X2 inst_11715 ( .A1(net_3493), .ZN(net_3149), .A2(net_1151) );
INV_X4 inst_16423 ( .ZN(net_2073), .A(net_1251) );
INV_X4 inst_16683 ( .A(net_13514), .ZN(net_8128) );
INV_X2 inst_19647 ( .A(net_19449), .ZN(net_19448) );
INV_X4 inst_17969 ( .A(net_21126), .ZN(net_604) );
INV_X4 inst_16943 ( .A(net_4111), .ZN(net_1634) );
NAND3_X2 inst_6066 ( .ZN(net_14136), .A3(net_10725), .A2(net_9530), .A1(net_7064) );
OAI22_X2 inst_1255 ( .B1(net_21146), .ZN(net_17664), .A2(net_17383), .B2(net_17382), .A1(net_16982) );
NAND2_X2 inst_9844 ( .ZN(net_11547), .A1(net_9541), .A2(net_6199) );
CLKBUF_X2 inst_22553 ( .A(net_22424), .Z(net_22425) );
NAND2_X2 inst_9279 ( .ZN(net_12588), .A1(net_10920), .A2(net_10852) );
OAI21_X2 inst_1791 ( .A(net_15071), .ZN(net_14614), .B2(net_11821), .B1(net_9261) );
NOR2_X2 inst_3420 ( .A1(net_15842), .ZN(net_15575), .A2(net_14805) );
NAND2_X2 inst_8834 ( .ZN(net_15493), .A2(net_14906), .A1(net_13190) );
AOI21_X2 inst_20774 ( .A(net_13554), .B2(net_10762), .ZN(net_10628), .B1(net_10627) );
NOR2_X2 inst_5064 ( .ZN(net_983), .A2(net_212), .A1(net_123) );
INV_X8 inst_12341 ( .ZN(net_996), .A(net_273) );
NAND2_X2 inst_11827 ( .ZN(net_3159), .A1(net_2746), .A2(net_299) );
XNOR2_X2 inst_528 ( .A(net_16839), .ZN(net_3348), .B(net_3347) );
DFF_X2 inst_19767 ( .QN(net_20859), .D(net_18869), .CK(net_22056) );
NAND2_X2 inst_9360 ( .ZN(net_19702), .A2(net_9892), .A1(net_6963) );
AOI21_X2 inst_20827 ( .ZN(net_9865), .B1(net_8179), .B2(net_6507), .A(net_2719) );
NAND2_X2 inst_9782 ( .ZN(net_11632), .A1(net_8273), .A2(net_6258) );
INV_X4 inst_13574 ( .ZN(net_10705), .A(net_9125) );
INV_X4 inst_16244 ( .ZN(net_2952), .A(net_1367) );
INV_X4 inst_17065 ( .ZN(net_5479), .A(net_4264) );
INV_X4 inst_13173 ( .ZN(net_14393), .A(net_13935) );
NOR2_X2 inst_4957 ( .ZN(net_2359), .A1(net_1634), .A2(net_1633) );
SDFF_X2 inst_846 ( .Q(net_21184), .SI(net_17314), .SE(net_125), .CK(net_22309), .D(x6521) );
NAND2_X2 inst_11377 ( .ZN(net_6384), .A2(net_3406), .A1(net_1647) );
NAND3_X2 inst_5925 ( .A3(net_20015), .A1(net_20014), .ZN(net_14979), .A2(net_4682) );
AOI221_X4 inst_20072 ( .C1(net_19867), .ZN(net_19060), .C2(net_15995), .B2(net_13741), .A(net_13261), .B1(net_12001) );
OAI21_X2 inst_1734 ( .ZN(net_15072), .A(net_15071), .B1(net_13506), .B2(net_8966) );
NAND2_X4 inst_7036 ( .ZN(net_16557), .A2(net_16556), .A1(net_16489) );
INV_X4 inst_17976 ( .A(net_21159), .ZN(net_349) );
NOR2_X2 inst_4646 ( .ZN(net_6948), .A2(net_3940), .A1(net_1102) );
CLKBUF_X2 inst_22340 ( .A(net_22211), .Z(net_22212) );
CLKBUF_X2 inst_21951 ( .A(net_21822), .Z(net_21823) );
DFF_X1 inst_19847 ( .D(net_17190), .CK(net_22110), .Q(x413) );
AND2_X4 inst_21258 ( .ZN(net_2718), .A2(net_193), .A1(net_109) );
DFF_X1 inst_19899 ( .D(net_16884), .CK(net_21586), .Q(x610) );
NOR2_X2 inst_3354 ( .ZN(net_17786), .A2(net_17639), .A1(net_17119) );
INV_X4 inst_17887 ( .ZN(net_261), .A(net_72) );
NOR2_X2 inst_4993 ( .ZN(net_2840), .A2(net_901), .A1(net_225) );
CLKBUF_X2 inst_21914 ( .A(net_21407), .Z(net_21786) );
NAND2_X2 inst_9500 ( .ZN(net_11398), .A1(net_11397), .A2(net_6322) );
NAND2_X2 inst_8199 ( .ZN(net_17884), .A1(net_17863), .A2(net_17802) );
DFF_X1 inst_19840 ( .D(net_17285), .CK(net_21988), .Q(x975) );
INV_X4 inst_17215 ( .A(net_816), .ZN(net_696) );
NOR2_X2 inst_3927 ( .A2(net_10762), .A1(net_10141), .ZN(net_8746) );
NOR3_X2 inst_2718 ( .ZN(net_13329), .A2(net_11450), .A1(net_10903), .A3(net_7330) );
DFF_X1 inst_19857 ( .D(net_17142), .CK(net_21755), .Q(x55) );
XNOR2_X2 inst_58 ( .ZN(net_18843), .A(net_18799), .B(net_17646) );
NOR2_X2 inst_3633 ( .ZN(net_19199), .A2(net_12196), .A1(net_7234) );
NAND2_X2 inst_9574 ( .A1(net_14085), .ZN(net_10953), .A2(net_10557) );
NAND2_X2 inst_11653 ( .A2(net_7078), .ZN(net_6429), .A1(net_3385) );
NAND2_X2 inst_9775 ( .ZN(net_9790), .A1(net_9041), .A2(net_4105) );
INV_X4 inst_13792 ( .A(net_7564), .ZN(net_7563) );
AOI21_X2 inst_20490 ( .ZN(net_14765), .B1(net_14764), .B2(net_13204), .A(net_11484) );
CLKBUF_X2 inst_22351 ( .A(net_22222), .Z(net_22223) );
OAI21_X4 inst_1469 ( .ZN(net_20682), .B2(net_20134), .B1(net_20133), .A(net_15044) );
INV_X2 inst_18806 ( .ZN(net_7405), .A(net_7404) );
INV_X2 inst_19315 ( .ZN(net_2652), .A(net_2651) );
NAND2_X2 inst_10295 ( .ZN(net_10117), .A1(net_7901), .A2(net_6217) );
NAND2_X2 inst_12056 ( .ZN(net_892), .A1(net_807), .A2(net_598) );
AOI21_X2 inst_20702 ( .ZN(net_12134), .A(net_12133), .B2(net_8390), .B1(net_5334) );
INV_X4 inst_16156 ( .ZN(net_7538), .A(net_1458) );
INV_X4 inst_17949 ( .A(net_21163), .ZN(net_636) );
INV_X4 inst_12878 ( .ZN(net_20285), .A(net_16708) );
INV_X4 inst_16918 ( .ZN(net_8293), .A(net_242) );
NAND3_X2 inst_5690 ( .A3(net_19551), .A1(net_19550), .ZN(net_16272), .A2(net_15978) );
NAND2_X2 inst_9592 ( .A1(net_13569), .ZN(net_10857), .A2(net_7361) );
NAND4_X2 inst_5288 ( .ZN(net_15940), .A1(net_15265), .A4(net_14789), .A3(net_13311), .A2(net_12940) );
INV_X4 inst_18302 ( .A(net_20486), .ZN(net_20482) );
OAI211_X2 inst_2424 ( .ZN(net_15225), .C1(net_15224), .C2(net_13329), .A(net_8531), .B(net_8266) );
INV_X4 inst_15860 ( .ZN(net_8232), .A(net_1810) );
NOR2_X2 inst_4517 ( .A1(net_4799), .A2(net_4162), .ZN(net_4153) );
INV_X4 inst_13719 ( .ZN(net_11784), .A(net_7821) );
NOR2_X4 inst_3144 ( .ZN(net_4869), .A2(net_4026), .A1(net_809) );
INV_X4 inst_13386 ( .ZN(net_14183), .A(net_10761) );
CLKBUF_X2 inst_22304 ( .A(net_21679), .Z(net_22176) );
NAND3_X2 inst_6124 ( .ZN(net_13749), .A3(net_13669), .A1(net_11133), .A2(net_5063) );
CLKBUF_X2 inst_22590 ( .A(net_21672), .Z(net_22462) );
CLKBUF_X2 inst_21443 ( .A(net_21251), .Z(net_21315) );
NAND2_X2 inst_11530 ( .ZN(net_5317), .A1(net_2913), .A2(net_1455) );
NOR2_X2 inst_3666 ( .ZN(net_12655), .A1(net_11866), .A2(net_10970) );
SDFF_X2 inst_993 ( .QN(net_21030), .SE(net_17277), .D(net_586), .CK(net_22725), .SI(x2481) );
INV_X4 inst_14882 ( .ZN(net_12283), .A(net_3671) );
NAND4_X4 inst_5177 ( .ZN(net_16663), .A1(net_16352), .A4(net_16313), .A3(net_15992), .A2(net_10820) );
CLKBUF_X2 inst_21667 ( .A(net_21531), .Z(net_21539) );
NAND3_X2 inst_6407 ( .ZN(net_11966), .A1(net_9963), .A3(net_9376), .A2(net_9039) );
INV_X4 inst_14590 ( .A(net_9626), .ZN(net_4461) );
INV_X4 inst_17137 ( .A(net_7230), .ZN(net_1197) );
INV_X4 inst_17034 ( .A(net_3047), .ZN(net_842) );
NAND2_X4 inst_7264 ( .ZN(net_7631), .A2(net_6200), .A1(net_3033) );
INV_X4 inst_13855 ( .A(net_9356), .ZN(net_9138) );
INV_X4 inst_16646 ( .ZN(net_2235), .A(net_1096) );
NAND3_X4 inst_5535 ( .A3(net_20195), .A1(net_20194), .ZN(net_17337), .A2(net_16040) );
XNOR2_X2 inst_630 ( .B(net_21173), .ZN(net_15959), .A(net_726) );
INV_X2 inst_19466 ( .ZN(net_3169), .A(net_1453) );
NAND4_X2 inst_5268 ( .A4(net_19829), .A1(net_19828), .ZN(net_16140), .A3(net_15187), .A2(net_14877) );
NAND2_X2 inst_11796 ( .A1(net_7890), .ZN(net_4351), .A2(net_1121) );
CLKBUF_X2 inst_21935 ( .A(net_21763), .Z(net_21807) );
NAND2_X2 inst_9662 ( .ZN(net_10326), .A1(net_10325), .A2(net_7749) );
OAI22_X2 inst_1273 ( .B1(net_21155), .ZN(net_16776), .A1(net_16775), .B2(net_16774), .A2(net_16412) );
XNOR2_X2 inst_512 ( .ZN(net_6373), .A(net_6372), .B(net_2555) );
NAND2_X2 inst_11337 ( .A1(net_5246), .ZN(net_3689), .A2(net_3688) );
INV_X4 inst_12791 ( .ZN(net_17283), .A(net_17282) );
NOR2_X2 inst_4966 ( .ZN(net_6299), .A2(net_1705), .A1(net_1114) );
INV_X4 inst_14307 ( .ZN(net_20606), .A(net_11822) );
INV_X8 inst_12278 ( .ZN(net_2117), .A(net_929) );
INV_X4 inst_15308 ( .ZN(net_3681), .A(net_1938) );
OAI21_X2 inst_2151 ( .ZN(net_9307), .A(net_9306), .B1(net_8490), .B2(net_3591) );
NOR2_X4 inst_3054 ( .ZN(net_6144), .A1(net_4991), .A2(net_3185) );
AND2_X4 inst_21266 ( .ZN(net_1174), .A2(net_221), .A1(net_168) );
DFF_X1 inst_19850 ( .D(net_17188), .CK(net_22376), .Q(x876) );
INV_X4 inst_15450 ( .ZN(net_2728), .A(net_2492) );
NAND2_X2 inst_11744 ( .ZN(net_4337), .A1(net_3311), .A2(net_2144) );
NOR2_X2 inst_4764 ( .ZN(net_3775), .A2(net_3221), .A1(net_2985) );
AND3_X4 inst_21114 ( .A2(net_14533), .ZN(net_14344), .A3(net_13078), .A1(net_12621) );
AOI21_X4 inst_20224 ( .ZN(net_14037), .B1(net_13938), .B2(net_10145), .A(net_9976) );
INV_X2 inst_18750 ( .ZN(net_7831), .A(net_7830) );
INV_X4 inst_13271 ( .ZN(net_12527), .A(net_12526) );
INV_X4 inst_15755 ( .ZN(net_10114), .A(net_7528) );
NOR2_X2 inst_3772 ( .ZN(net_13072), .A1(net_10285), .A2(net_10284) );
NOR2_X2 inst_4210 ( .ZN(net_8684), .A1(net_6647), .A2(net_6646) );
OAI21_X2 inst_2043 ( .ZN(net_11190), .B1(net_11189), .A(net_5398), .B2(net_5069) );
SDFF_X2 inst_960 ( .QN(net_21068), .D(net_415), .SE(net_263), .CK(net_21731), .SI(x1948) );
INV_X4 inst_16051 ( .A(net_8720), .ZN(net_5818) );
OAI211_X2 inst_2411 ( .ZN(net_15523), .C1(net_15522), .A(net_14867), .B(net_14655), .C2(net_12860) );
XOR2_X2 inst_38 ( .A(net_21199), .Z(net_649), .B(net_648) );
NOR4_X2 inst_2601 ( .ZN(net_12143), .A4(net_12142), .A2(net_7820), .A1(net_6769), .A3(net_6012) );
XNOR2_X2 inst_381 ( .B(net_21108), .ZN(net_17168), .A(net_16802) );
INV_X4 inst_14846 ( .ZN(net_4829), .A(net_3845) );
NAND2_X2 inst_9448 ( .A1(net_12764), .ZN(net_11529), .A2(net_10243) );
NOR2_X2 inst_3837 ( .ZN(net_9686), .A1(net_8254), .A2(net_7482) );
NAND2_X4 inst_6876 ( .A2(net_20280), .A1(net_20279), .ZN(net_18242) );
CLKBUF_X2 inst_22864 ( .A(net_21402), .Z(net_22736) );
NAND2_X4 inst_7577 ( .A2(net_2283), .ZN(net_2265), .A1(net_1299) );
NAND2_X2 inst_10355 ( .ZN(net_7456), .A1(net_7455), .A2(net_7454) );
INV_X4 inst_13108 ( .ZN(net_15704), .A(net_15495) );
NAND2_X2 inst_8068 ( .ZN(net_20616), .A1(net_18182), .A2(net_18143) );
AOI21_X2 inst_20906 ( .ZN(net_7693), .B2(net_4638), .B1(net_3575), .A(net_2743) );
NAND4_X2 inst_5496 ( .ZN(net_11951), .A2(net_10131), .A4(net_8063), .A3(net_7795), .A1(net_4347) );
INV_X4 inst_18135 ( .A(net_20894), .ZN(net_162) );
NAND3_X2 inst_6002 ( .ZN(net_14429), .A1(net_12717), .A3(net_11336), .A2(net_8786) );
INV_X4 inst_13880 ( .A(net_9586), .ZN(net_9203) );
NAND2_X2 inst_10228 ( .ZN(net_8058), .A1(net_7812), .A2(net_6128) );
INV_X4 inst_14599 ( .ZN(net_5737), .A(net_4450) );
AOI22_X2 inst_20041 ( .B1(net_20560), .A1(net_13076), .ZN(net_7107), .B2(net_7106), .A2(net_4339) );
INV_X4 inst_15008 ( .ZN(net_9692), .A(net_2586) );
NAND4_X2 inst_5503 ( .A3(net_11959), .A4(net_11855), .ZN(net_11806), .A1(net_11805), .A2(net_5491) );
NOR2_X2 inst_4597 ( .A1(net_9148), .ZN(net_7068), .A2(net_2602) );
OR2_X2 inst_1188 ( .A2(net_4963), .A1(net_4520), .ZN(net_4519) );
CLKBUF_X2 inst_22186 ( .A(net_22057), .Z(net_22058) );
INV_X4 inst_14579 ( .ZN(net_4523), .A(net_4522) );
AOI21_X2 inst_20797 ( .B2(net_12248), .ZN(net_10418), .A(net_10417), .B1(net_2010) );
INV_X4 inst_13462 ( .ZN(net_11518), .A(net_10245) );
NAND2_X2 inst_9960 ( .ZN(net_20175), .A2(net_8912), .A1(net_6203) );
NAND2_X4 inst_6957 ( .ZN(net_20762), .A2(net_19398), .A1(net_19397) );
NAND2_X4 inst_7184 ( .ZN(net_10735), .A1(net_9162), .A2(net_8160) );
NAND2_X2 inst_8966 ( .ZN(net_14620), .A1(net_14619), .A2(net_13388) );
NOR2_X2 inst_3873 ( .ZN(net_18990), .A1(net_9368), .A2(net_6684) );
NAND2_X2 inst_8363 ( .A1(net_21147), .ZN(net_17377), .A2(net_17376) );
INV_X2 inst_19017 ( .ZN(net_4982), .A(net_4981) );
AOI211_X2 inst_21058 ( .C1(net_11494), .ZN(net_11199), .C2(net_11198), .A(net_9897), .B(net_3032) );
CLKBUF_X2 inst_22391 ( .A(net_21309), .Z(net_22263) );
INV_X4 inst_16290 ( .A(net_12307), .ZN(net_1335) );
AOI21_X2 inst_20266 ( .B2(net_20912), .ZN(net_18063), .B1(net_16205), .A(net_12121) );
XNOR2_X2 inst_387 ( .B(net_17366), .ZN(net_16781), .A(net_16780) );
INV_X2 inst_18370 ( .ZN(net_17531), .A(net_17424) );
NOR2_X2 inst_4601 ( .ZN(net_6564), .A1(net_4481), .A2(net_3762) );
INV_X4 inst_15416 ( .ZN(net_14509), .A(net_2520) );
INV_X4 inst_14769 ( .ZN(net_9988), .A(net_4053) );
CLKBUF_X2 inst_22092 ( .A(net_21407), .Z(net_21964) );
INV_X4 inst_12784 ( .ZN(net_17301), .A(net_17300) );
INV_X2 inst_18757 ( .A(net_13442), .ZN(net_7641) );
INV_X2 inst_18711 ( .A(net_10493), .ZN(net_8230) );
OAI21_X2 inst_2129 ( .ZN(net_9998), .A(net_9997), .B1(net_9801), .B2(net_4836) );
NAND2_X2 inst_8801 ( .A1(net_16030), .ZN(net_15661), .A2(net_15315) );
NAND3_X2 inst_5750 ( .ZN(net_16006), .A3(net_15624), .A2(net_14940), .A1(net_12682) );
INV_X2 inst_18714 ( .ZN(net_8210), .A(net_8209) );
INV_X4 inst_16422 ( .A(net_12363), .ZN(net_11482) );
NAND2_X2 inst_11273 ( .ZN(net_3887), .A1(net_3886), .A2(net_2081) );
OR2_X2 inst_1181 ( .ZN(net_4790), .A2(net_4789), .A1(net_612) );
INV_X1 inst_19760 ( .A(net_4075), .ZN(net_2826) );
CLKBUF_X2 inst_21509 ( .A(net_21380), .Z(net_21381) );
INV_X4 inst_18223 ( .A(net_20929), .ZN(net_910) );
NAND2_X2 inst_8986 ( .A1(net_15628), .ZN(net_14485), .A2(net_12906) );
NAND3_X2 inst_6165 ( .A2(net_14211), .ZN(net_13634), .A1(net_12344), .A3(net_8768) );
NOR2_X2 inst_5045 ( .ZN(net_1078), .A2(net_870), .A1(net_61) );
CLKBUF_X2 inst_22566 ( .A(net_22249), .Z(net_22438) );
INV_X4 inst_17863 ( .ZN(net_942), .A(net_89) );
OAI21_X2 inst_1548 ( .ZN(net_17734), .B2(net_17651), .A(net_17481), .B1(net_17480) );
INV_X4 inst_15916 ( .ZN(net_9014), .A(net_4907) );
INV_X4 inst_17100 ( .A(net_10667), .ZN(net_8286) );
NAND2_X2 inst_9913 ( .ZN(net_11508), .A1(net_10309), .A2(net_7834) );
INV_X4 inst_17607 ( .ZN(net_993), .A(net_311) );
NAND2_X4 inst_7013 ( .A2(net_19639), .A1(net_19638), .ZN(net_17136) );
NAND2_X2 inst_9457 ( .A1(net_12419), .ZN(net_11502), .A2(net_11501) );
INV_X4 inst_14255 ( .ZN(net_7590), .A(net_5092) );
NAND2_X2 inst_10899 ( .ZN(net_6608), .A2(net_6512), .A1(net_5387) );
NAND3_X2 inst_5715 ( .ZN(net_16141), .A3(net_15714), .A2(net_15361), .A1(net_15316) );
NAND2_X2 inst_8470 ( .A1(net_21178), .ZN(net_17018), .A2(net_17011) );
INV_X4 inst_18338 ( .A(net_20585), .ZN(net_20584) );
NAND2_X2 inst_10462 ( .ZN(net_10655), .A1(net_9541), .A2(net_6980) );
NAND2_X2 inst_7799 ( .ZN(net_18700), .A2(net_18690), .A1(net_18684) );
INV_X4 inst_16089 ( .A(net_2331), .ZN(net_2197) );
CLKBUF_X2 inst_22930 ( .A(net_22801), .Z(net_22802) );
NAND2_X2 inst_12018 ( .A1(net_3009), .A2(net_2214), .ZN(net_1063) );
NOR2_X2 inst_5130 ( .A2(net_229), .ZN(net_228), .A1(net_227) );
INV_X4 inst_14629 ( .ZN(net_4626), .A(net_4393) );
INV_X4 inst_15447 ( .A(net_3351), .ZN(net_2777) );
NAND4_X2 inst_5489 ( .A1(net_13497), .ZN(net_12285), .A2(net_12284), .A3(net_12283), .A4(net_12282) );
INV_X4 inst_16765 ( .ZN(net_9754), .A(net_3297) );
INV_X2 inst_19207 ( .ZN(net_3529), .A(net_3528) );
NAND2_X2 inst_7765 ( .ZN(net_18764), .A2(net_18726), .A1(net_18699) );
INV_X4 inst_16453 ( .ZN(net_3281), .A(net_1226) );
INV_X4 inst_14662 ( .ZN(net_19195), .A(net_15974) );
NAND2_X2 inst_8682 ( .A2(net_16576), .A1(net_16497), .ZN(net_16450) );
NAND2_X2 inst_9760 ( .ZN(net_9852), .A1(net_9849), .A2(net_4745) );
NAND4_X2 inst_5290 ( .A4(net_19712), .A1(net_19711), .ZN(net_19344), .A2(net_12492), .A3(net_12114) );
INV_X4 inst_16468 ( .ZN(net_1632), .A(net_1213) );
NAND2_X2 inst_10239 ( .ZN(net_8036), .A1(net_8035), .A2(net_5967) );
AOI21_X2 inst_20473 ( .ZN(net_14957), .B1(net_13117), .B2(net_12676), .A(net_1132) );
AOI21_X4 inst_20214 ( .B1(net_20355), .ZN(net_14399), .A(net_6734), .B2(net_308) );
NAND2_X2 inst_8585 ( .A2(net_16727), .ZN(net_16715), .A1(net_16663) );
OAI21_X2 inst_2307 ( .A(net_9754), .ZN(net_5765), .B2(net_4145), .B1(net_3243) );
NAND2_X2 inst_11611 ( .ZN(net_8342), .A1(net_7007), .A2(net_2610) );
NOR3_X4 inst_2611 ( .ZN(net_15998), .A3(net_15408), .A1(net_14640), .A2(net_14473) );
INV_X4 inst_13469 ( .ZN(net_12891), .A(net_9669) );
NOR2_X2 inst_5004 ( .ZN(net_10325), .A2(net_6318), .A1(net_1470) );
AOI21_X2 inst_20464 ( .ZN(net_15002), .B1(net_14636), .B2(net_12997), .A(net_7314) );
NAND2_X2 inst_9926 ( .ZN(net_12425), .A1(net_8573), .A2(net_4085) );
INV_X2 inst_19236 ( .ZN(net_3337), .A(net_3336) );
NOR2_X4 inst_2994 ( .A1(net_19483), .ZN(net_9476), .A2(net_955) );
NOR2_X4 inst_3023 ( .ZN(net_8364), .A1(net_6492), .A2(net_3862) );
OR2_X2 inst_1243 ( .ZN(net_1304), .A2(net_268), .A1(net_154) );
INV_X4 inst_13155 ( .ZN(net_14872), .A(net_14332) );
AND3_X2 inst_21147 ( .A3(net_8565), .ZN(net_6405), .A2(net_6404), .A1(net_3701) );
INV_X4 inst_14970 ( .ZN(net_3425), .A(net_3424) );
CLKBUF_X2 inst_21774 ( .A(net_21645), .Z(net_21646) );
NAND2_X2 inst_9512 ( .ZN(net_11188), .A1(net_8196), .A2(net_6614) );
INV_X4 inst_13074 ( .ZN(net_16229), .A(net_16170) );
NAND2_X2 inst_10514 ( .ZN(net_8211), .A1(net_6879), .A2(net_6878) );
INV_X4 inst_14639 ( .ZN(net_4778), .A(net_4381) );
NAND3_X2 inst_5958 ( .ZN(net_14845), .A3(net_14844), .A2(net_13423), .A1(net_7611) );
OR2_X4 inst_1093 ( .A2(net_6971), .ZN(net_4033), .A1(net_4032) );
NAND2_X4 inst_7646 ( .ZN(net_1346), .A2(net_972), .A1(net_935) );
INV_X4 inst_14728 ( .ZN(net_6533), .A(net_4122) );
INV_X2 inst_19624 ( .A(net_20919), .ZN(net_20005) );
CLKBUF_X2 inst_21560 ( .A(net_21431), .Z(net_21432) );
NOR2_X4 inst_3271 ( .ZN(net_2814), .A2(net_1881), .A1(net_1526) );
OAI21_X4 inst_1430 ( .B2(net_19535), .B1(net_19534), .ZN(net_18946), .A(net_16347) );
NAND2_X2 inst_10707 ( .ZN(net_6013), .A2(net_4407), .A1(net_90) );
INV_X4 inst_14516 ( .ZN(net_8002), .A(net_4813) );
CLKBUF_X2 inst_22740 ( .A(net_22611), .Z(net_22612) );
NOR2_X4 inst_3257 ( .A1(net_20868), .ZN(net_2259), .A2(net_2242) );
NAND2_X2 inst_10759 ( .A1(net_8037), .ZN(net_6710), .A2(net_5423) );
INV_X4 inst_14081 ( .ZN(net_13497), .A(net_6218) );
NAND2_X2 inst_11498 ( .A1(net_10183), .ZN(net_3078), .A2(net_2161) );
INV_X4 inst_16543 ( .ZN(net_11549), .A(net_1505) );
CLKBUF_X2 inst_22328 ( .A(net_22199), .Z(net_22200) );
CLKBUF_X2 inst_22316 ( .A(net_21332), .Z(net_22188) );
AOI21_X4 inst_20102 ( .ZN(net_19546), .B1(net_16394), .A(net_16252), .B2(net_16225) );
NAND2_X2 inst_9979 ( .A2(net_10565), .ZN(net_8864), .A1(net_5988) );
SDFF_X2 inst_763 ( .Q(net_20870), .SE(net_18577), .SI(net_18520), .D(net_717), .CK(net_22450) );
OAI21_X2 inst_2330 ( .ZN(net_20149), .A(net_9636), .B2(net_4326), .B1(net_2397) );
NAND2_X4 inst_7377 ( .A1(net_5635), .ZN(net_5457), .A2(net_4287) );
NOR2_X2 inst_3636 ( .ZN(net_20180), .A2(net_12187), .A1(net_8777) );
NAND2_X2 inst_11069 ( .ZN(net_8251), .A2(net_2803), .A1(net_874) );
INV_X4 inst_14018 ( .ZN(net_11181), .A(net_6298) );
INV_X4 inst_13754 ( .A(net_7619), .ZN(net_7618) );
INV_X4 inst_15970 ( .ZN(net_1887), .A(net_1686) );
INV_X4 inst_17185 ( .ZN(net_4264), .A(net_308) );
INV_X2 inst_19514 ( .A(net_1615), .ZN(net_1153) );
XNOR2_X2 inst_537 ( .ZN(net_1512), .A(net_1511), .B(net_959) );
AND3_X4 inst_21125 ( .ZN(net_12057), .A3(net_12056), .A1(net_10641), .A2(net_6835) );
NOR2_X2 inst_5069 ( .ZN(net_4516), .A2(net_949), .A1(net_221) );
CLKBUF_X2 inst_21900 ( .A(net_21771), .Z(net_21772) );
INV_X4 inst_17935 ( .A(net_21064), .ZN(net_530) );
NAND2_X4 inst_7141 ( .ZN(net_12746), .A2(net_9807), .A1(net_9418) );
INV_X4 inst_14977 ( .ZN(net_14972), .A(net_14460) );
INV_X4 inst_15232 ( .ZN(net_3627), .A(net_2837) );
INV_X4 inst_14341 ( .ZN(net_5988), .A(net_5366) );
NAND2_X2 inst_8431 ( .ZN(net_19764), .A2(net_17141), .A1(net_17048) );
NAND2_X2 inst_10786 ( .ZN(net_10595), .A2(net_5590), .A1(net_573) );
NOR2_X2 inst_3950 ( .A1(net_12496), .A2(net_10503), .ZN(net_8612) );
NAND2_X2 inst_8863 ( .ZN(net_15336), .A2(net_14481), .A1(net_10660) );
NOR2_X2 inst_4288 ( .ZN(net_7492), .A2(net_6039), .A1(net_4655) );
SDFF_X2 inst_869 ( .Q(net_21192), .SI(net_17090), .SE(net_125), .CK(net_22297), .D(x6300) );
NAND2_X2 inst_10671 ( .ZN(net_8917), .A1(net_5277), .A2(net_3540) );
NOR3_X2 inst_2646 ( .ZN(net_15778), .A3(net_14763), .A1(net_14633), .A2(net_13782) );
INV_X4 inst_18321 ( .A(net_20535), .ZN(net_20534) );
NAND3_X2 inst_6543 ( .ZN(net_10568), .A3(net_10567), .A1(net_6799), .A2(net_6368) );
INV_X2 inst_18493 ( .ZN(net_14262), .A(net_12324) );
INV_X4 inst_17824 ( .ZN(net_270), .A(net_156) );
INV_X4 inst_13229 ( .ZN(net_13521), .A(net_12512) );
NAND2_X2 inst_9753 ( .ZN(net_10043), .A1(net_10042), .A2(net_6577) );
INV_X4 inst_13649 ( .ZN(net_12063), .A(net_8155) );
NOR2_X4 inst_3267 ( .ZN(net_3513), .A2(net_1981), .A1(net_1586) );
NAND2_X2 inst_9849 ( .A1(net_10395), .ZN(net_9533), .A2(net_9532) );
NOR2_X4 inst_3205 ( .ZN(net_5525), .A1(net_3035), .A2(net_3034) );
INV_X4 inst_14315 ( .ZN(net_6755), .A(net_5474) );
INV_X4 inst_17109 ( .ZN(net_1046), .A(net_278) );
NAND3_X2 inst_6048 ( .ZN(net_14246), .A2(net_13956), .A3(net_13439), .A1(net_8422) );
NAND2_X2 inst_8945 ( .ZN(net_14729), .A2(net_13236), .A1(net_1015) );
XNOR2_X2 inst_612 ( .B(net_5788), .ZN(net_501), .A(net_500) );
INV_X4 inst_12505 ( .ZN(net_18610), .A(net_18609) );
NAND3_X2 inst_6185 ( .ZN(net_13471), .A3(net_9145), .A2(net_7970), .A1(net_7067) );
OAI21_X2 inst_1692 ( .B2(net_19307), .B1(net_19306), .ZN(net_15359), .A(net_12298) );
AOI21_X4 inst_20150 ( .ZN(net_20653), .B2(net_14938), .B1(net_14700), .A(net_8279) );
INV_X4 inst_15875 ( .A(net_5869), .ZN(net_2682) );
INV_X2 inst_19604 ( .A(net_20869), .ZN(net_91) );
NOR2_X2 inst_3986 ( .ZN(net_8323), .A2(net_8322), .A1(net_4552) );
NAND2_X4 inst_7627 ( .ZN(net_7703), .A2(net_353), .A1(net_309) );
INV_X4 inst_13137 ( .ZN(net_15130), .A(net_14746) );
NAND2_X4 inst_7275 ( .ZN(net_11175), .A1(net_4111), .A2(net_3558) );
INV_X4 inst_14328 ( .ZN(net_11974), .A(net_5696) );
NAND2_X2 inst_10819 ( .ZN(net_19997), .A2(net_5752), .A1(net_1777) );
INV_X4 inst_14535 ( .ZN(net_4660), .A(net_4659) );
OAI211_X2 inst_2455 ( .ZN(net_14322), .A(net_14321), .B(net_14320), .C1(net_14319), .C2(net_9020) );
INV_X4 inst_18157 ( .A(net_21034), .ZN(net_518) );
CLKBUF_X2 inst_22345 ( .A(net_22033), .Z(net_22217) );
INV_X4 inst_12923 ( .ZN(net_16813), .A(net_16689) );
NAND2_X2 inst_10575 ( .ZN(net_19940), .A1(net_11786), .A2(net_11317) );
INV_X4 inst_15690 ( .ZN(net_3989), .A(net_2033) );
INV_X4 inst_17570 ( .ZN(net_6525), .A(net_523) );
NAND3_X2 inst_6724 ( .ZN(net_6505), .A2(net_4735), .A3(net_3992), .A1(net_1577) );
NAND2_X2 inst_11581 ( .ZN(net_3341), .A2(net_2726), .A1(net_170) );
AND2_X2 inst_21317 ( .A2(net_9039), .ZN(net_7176), .A1(net_3622) );
NOR2_X2 inst_4828 ( .ZN(net_4236), .A1(net_2485), .A2(net_787) );
INV_X4 inst_18258 ( .A(net_21151), .ZN(net_17247) );
NAND4_X4 inst_5218 ( .A3(net_20304), .A1(net_20303), .ZN(net_17767), .A2(net_16145), .A4(net_16063) );
CLKBUF_X2 inst_22833 ( .A(net_22704), .Z(net_22705) );
NAND4_X2 inst_5389 ( .A4(net_20276), .A1(net_20275), .ZN(net_15009), .A2(net_11250), .A3(net_11024) );
AOI21_X2 inst_20543 ( .ZN(net_14413), .A(net_14412), .B2(net_12562), .B1(net_7077) );
INV_X2 inst_19249 ( .ZN(net_3259), .A(net_3258) );
INV_X4 inst_17152 ( .A(net_3108), .ZN(net_1434) );
SDFF_X2 inst_885 ( .Q(net_21206), .D(net_16936), .SE(net_263), .CK(net_22148), .SI(x5926) );
INV_X4 inst_15995 ( .ZN(net_13938), .A(net_9728) );
INV_X2 inst_18509 ( .ZN(net_11626), .A(net_11625) );
INV_X4 inst_17796 ( .ZN(net_1955), .A(net_131) );
NAND3_X2 inst_5803 ( .ZN(net_15703), .A3(net_15052), .A1(net_13988), .A2(net_5580) );
NAND2_X2 inst_10748 ( .ZN(net_10733), .A2(net_4308), .A1(net_1173) );
INV_X4 inst_18314 ( .ZN(net_20512), .A(net_7637) );
NOR2_X2 inst_3610 ( .ZN(net_12416), .A1(net_8537), .A2(net_7573) );
NOR2_X4 inst_2999 ( .ZN(net_9359), .A2(net_6571), .A1(net_4573) );
INV_X4 inst_13097 ( .ZN(net_20278), .A(net_15737) );
AOI21_X2 inst_20807 ( .ZN(net_10297), .B1(net_6455), .B2(net_6054), .A(net_603) );
NAND2_X2 inst_8351 ( .ZN(net_17468), .A1(net_17303), .A2(net_17293) );
INV_X4 inst_12822 ( .ZN(net_17488), .A(net_17341) );
INV_X2 inst_19244 ( .A(net_11446), .ZN(net_3277) );
NAND2_X2 inst_8188 ( .ZN(net_17906), .A2(net_17798), .A1(net_17717) );
NAND3_X2 inst_5956 ( .ZN(net_14848), .A3(net_14847), .A2(net_11079), .A1(net_7050) );
INV_X4 inst_17750 ( .A(net_1645), .ZN(net_420) );
NAND4_X2 inst_5305 ( .ZN(net_19971), .A4(net_19646), .A1(net_19645), .A3(net_13900), .A2(net_11005) );
NOR2_X2 inst_4156 ( .ZN(net_6891), .A1(net_6807), .A2(net_5439) );
NAND2_X2 inst_9875 ( .A2(net_9854), .ZN(net_9457), .A1(net_3297) );
INV_X4 inst_16896 ( .ZN(net_4794), .A(net_628) );
XNOR2_X2 inst_200 ( .B(net_20713), .ZN(net_17667), .A(net_17662) );
INV_X4 inst_16490 ( .ZN(net_15790), .A(net_15602) );
NAND2_X2 inst_11986 ( .ZN(net_2883), .A2(net_2327), .A1(net_1269) );
INV_X4 inst_17649 ( .ZN(net_721), .A(net_271) );
NOR2_X2 inst_4373 ( .ZN(net_19562), .A1(net_13091), .A2(net_9064) );
NAND2_X2 inst_9198 ( .A1(net_15270), .ZN(net_13088), .A2(net_11235) );
NAND2_X2 inst_9939 ( .ZN(net_9132), .A1(net_9131), .A2(net_7092) );
INV_X2 inst_18463 ( .ZN(net_12736), .A(net_11714) );
INV_X4 inst_16094 ( .ZN(net_9575), .A(net_9109) );
INV_X2 inst_18434 ( .ZN(net_14486), .A(net_14019) );
OAI21_X2 inst_1750 ( .ZN(net_14833), .B2(net_13451), .B1(net_10369), .A(net_750) );
NAND4_X4 inst_5242 ( .ZN(net_20046), .A1(net_14671), .A3(net_14536), .A4(net_13098), .A2(net_7206) );
INV_X2 inst_19264 ( .A(net_4089), .ZN(net_3859) );
NAND2_X2 inst_10155 ( .ZN(net_8269), .A2(net_8195), .A1(net_948) );
CLKBUF_X2 inst_22954 ( .A(net_22825), .Z(net_22826) );
NAND2_X2 inst_7758 ( .ZN(net_18763), .A2(net_18711), .A1(net_18688) );
NAND2_X4 inst_7593 ( .ZN(net_3182), .A2(net_1343), .A1(net_123) );
INV_X4 inst_16185 ( .ZN(net_2436), .A(net_2195) );
NAND2_X2 inst_9569 ( .ZN(net_19004), .A1(net_14075), .A2(net_7600) );
INV_X4 inst_17528 ( .ZN(net_6637), .A(net_4394) );
INV_X8 inst_12294 ( .ZN(net_2283), .A(net_419) );
NOR2_X2 inst_3499 ( .ZN(net_14066), .A2(net_11844), .A1(net_10292) );
SDFF_X2 inst_893 ( .Q(net_21216), .SI(net_17001), .SE(net_125), .CK(net_22284), .D(x7497) );
NAND2_X2 inst_8128 ( .A2(net_20880), .ZN(net_18048), .A1(net_16119) );
INV_X4 inst_15711 ( .ZN(net_19508), .A(net_2726) );
INV_X4 inst_15435 ( .A(net_2979), .ZN(net_2819) );
INV_X2 inst_19671 ( .A(net_20486), .ZN(net_20485) );
INV_X4 inst_17923 ( .A(net_20921), .ZN(net_1021) );
XNOR2_X2 inst_569 ( .ZN(net_638), .A(net_637), .B(net_636) );
NAND2_X2 inst_9209 ( .ZN(net_13050), .A2(net_13049), .A1(net_12991) );
INV_X4 inst_12763 ( .ZN(net_17385), .A(net_17384) );
INV_X4 inst_14730 ( .A(net_5792), .ZN(net_4661) );
INV_X4 inst_15440 ( .ZN(net_3300), .A(net_1642) );
INV_X4 inst_14451 ( .A(net_8476), .ZN(net_4958) );
CLKBUF_X2 inst_21453 ( .A(net_21324), .Z(net_21325) );
INV_X4 inst_12554 ( .A(net_18312), .ZN(net_18248) );
INV_X4 inst_16328 ( .ZN(net_3688), .A(net_1311) );
INV_X2 inst_18555 ( .ZN(net_10885), .A(net_10884) );
NOR2_X2 inst_4220 ( .A1(net_13968), .A2(net_9418), .ZN(net_8649) );
XNOR2_X2 inst_522 ( .ZN(net_5733), .A(net_1656), .B(net_33) );
INV_X2 inst_18658 ( .ZN(net_9207), .A(net_9206) );
NOR2_X2 inst_5040 ( .ZN(net_1094), .A1(net_895), .A2(net_367) );
INV_X2 inst_19172 ( .ZN(net_4817), .A(net_3237) );
NAND2_X2 inst_9037 ( .A1(net_14365), .ZN(net_14061), .A2(net_11829) );
INV_X8 inst_12408 ( .ZN(net_314), .A(net_164) );
INV_X4 inst_14458 ( .A(net_8511), .ZN(net_4946) );
NAND2_X2 inst_9842 ( .ZN(net_12812), .A2(net_7564), .A1(net_6668) );
NOR2_X4 inst_2809 ( .ZN(net_17793), .A1(net_17531), .A2(net_17423) );
NAND2_X2 inst_9654 ( .ZN(net_13980), .A2(net_9771), .A1(net_5432) );
INV_X4 inst_14011 ( .A(net_8197), .ZN(net_6307) );
INV_X4 inst_15147 ( .A(net_3080), .ZN(net_3079) );
INV_X4 inst_12478 ( .ZN(net_18730), .A(net_18703) );
INV_X4 inst_17076 ( .ZN(net_8260), .A(net_904) );
INV_X4 inst_13141 ( .ZN(net_15082), .A(net_14685) );
INV_X4 inst_12797 ( .ZN(net_17267), .A(net_17266) );
INV_X4 inst_18273 ( .A(net_19454), .ZN(net_19453) );
NAND2_X4 inst_6936 ( .A2(net_19764), .A1(net_19763), .ZN(net_17539) );
DFF_X1 inst_19912 ( .D(net_16840), .CK(net_22342), .Q(x844) );
INV_X2 inst_18401 ( .ZN(net_19962), .A(net_16400) );
CLKBUF_X2 inst_22122 ( .A(net_21993), .Z(net_21994) );
INV_X4 inst_17497 ( .ZN(net_2426), .A(net_125) );
NAND2_X4 inst_6911 ( .A2(net_19666), .A1(net_19665), .ZN(net_17890) );
NAND2_X2 inst_9144 ( .A1(net_14085), .ZN(net_13408), .A2(net_10510) );
INV_X2 inst_18662 ( .ZN(net_12505), .A(net_10952) );
NAND2_X2 inst_11131 ( .A2(net_20796), .ZN(net_6603), .A1(net_4268) );
NAND2_X2 inst_8997 ( .ZN(net_14400), .A2(net_13043), .A1(net_10310) );
NAND3_X2 inst_6493 ( .ZN(net_11160), .A2(net_11159), .A3(net_11158), .A1(net_3579) );
INV_X4 inst_14779 ( .ZN(net_6468), .A(net_4045) );
INV_X4 inst_16603 ( .ZN(net_1128), .A(net_1127) );
SDFF_X2 inst_719 ( .Q(net_20957), .SE(net_18804), .SI(net_18735), .D(net_744), .CK(net_22005) );
INV_X4 inst_15699 ( .ZN(net_19175), .A(net_2014) );
NAND2_X2 inst_10195 ( .ZN(net_8140), .A1(net_6316), .A2(net_6294) );
NOR2_X2 inst_4166 ( .ZN(net_6868), .A1(net_6867), .A2(net_5202) );
INV_X4 inst_18182 ( .A(net_21061), .ZN(net_483) );
AOI21_X4 inst_20248 ( .ZN(net_9863), .B1(net_5975), .B2(net_5241), .A(net_2372) );
INV_X4 inst_18234 ( .A(net_20955), .ZN(net_143) );
NOR2_X2 inst_3868 ( .ZN(net_11470), .A1(net_9374), .A2(net_9373) );
NAND2_X2 inst_8695 ( .ZN(net_19186), .A1(net_16357), .A2(net_16204) );
INV_X4 inst_17574 ( .A(net_841), .ZN(net_764) );
OR2_X2 inst_1134 ( .ZN(net_12628), .A1(net_12627), .A2(net_12626) );
AOI21_X2 inst_20315 ( .ZN(net_20327), .B1(net_15974), .B2(net_15591), .A(net_13333) );
AOI22_X2 inst_20046 ( .ZN(net_20125), .B1(net_5239), .A2(net_3911), .B2(net_2158), .A1(net_1091) );
NOR2_X2 inst_3546 ( .ZN(net_13115), .A2(net_13114), .A1(net_10127) );
NAND3_X2 inst_5748 ( .ZN(net_19069), .A1(net_15625), .A3(net_15448), .A2(net_12140) );
OR2_X2 inst_1144 ( .A2(net_11091), .ZN(net_10918), .A1(net_10917) );
NAND4_X4 inst_5165 ( .ZN(net_20220), .A3(net_18897), .A1(net_18896), .A4(net_18050), .A2(net_15832) );
NAND3_X2 inst_6426 ( .ZN(net_11930), .A2(net_11929), .A3(net_8146), .A1(net_3694) );
NAND4_X2 inst_5366 ( .A1(net_19540), .ZN(net_15239), .A4(net_12038), .A3(net_11742), .A2(net_8660) );
NAND3_X4 inst_5551 ( .A3(net_20261), .A1(net_20260), .ZN(net_16766), .A2(net_12272) );
INV_X4 inst_17599 ( .A(net_874), .ZN(net_399) );
OAI211_X2 inst_2568 ( .ZN(net_9034), .C2(net_9033), .C1(net_8674), .A(net_8567), .B(net_3186) );
OAI21_X2 inst_2295 ( .ZN(net_6470), .B1(net_5852), .A(net_5405), .B2(net_4378) );
INV_X4 inst_17168 ( .ZN(net_1017), .A(net_212) );
INV_X4 inst_13021 ( .ZN(net_16564), .A(net_16451) );
AOI21_X2 inst_20437 ( .ZN(net_15155), .A(net_14610), .B1(net_10812), .B2(net_6446) );
INV_X4 inst_17759 ( .ZN(net_14006), .A(net_8596) );
INV_X2 inst_19039 ( .ZN(net_4781), .A(net_4780) );
NOR2_X2 inst_3532 ( .ZN(net_13552), .A2(net_12300), .A1(net_320) );
NOR2_X4 inst_3028 ( .ZN(net_8587), .A1(net_6221), .A2(net_3683) );
NAND2_X2 inst_9190 ( .ZN(net_19520), .A1(net_13122), .A2(net_13121) );
NOR2_X2 inst_3854 ( .A1(net_10930), .ZN(net_9501), .A2(net_9500) );
NAND2_X2 inst_9432 ( .ZN(net_11599), .A1(net_11598), .A2(net_11597) );
NAND2_X2 inst_10881 ( .A1(net_9459), .A2(net_6684), .ZN(net_6664) );
AOI221_X2 inst_20090 ( .C1(net_15369), .B1(net_15369), .ZN(net_15236), .A(net_13701), .B2(net_13200), .C2(net_10782) );
NAND2_X4 inst_7089 ( .A1(net_19025), .ZN(net_15246), .A2(net_15191) );
OAI21_X2 inst_1530 ( .ZN(net_18004), .B1(net_18003), .B2(net_17898), .A(net_2027) );
INV_X4 inst_18004 ( .A(net_21122), .ZN(net_634) );
NAND4_X2 inst_5421 ( .ZN(net_14251), .A4(net_13406), .A3(net_13014), .A1(net_12945), .A2(net_2312) );
INV_X4 inst_17091 ( .ZN(net_14684), .A(net_10699) );
NAND2_X4 inst_7635 ( .ZN(net_2532), .A2(net_1159), .A1(net_1158) );
NAND3_X2 inst_6308 ( .ZN(net_12779), .A2(net_11693), .A3(net_11552), .A1(net_8194) );
NAND2_X2 inst_11599 ( .A1(net_6963), .ZN(net_2664), .A2(net_2663) );
INV_X2 inst_18816 ( .ZN(net_7234), .A(net_7233) );
NAND3_X2 inst_5948 ( .A3(net_20226), .ZN(net_14886), .A1(net_14272), .A2(net_7532) );
NAND2_X2 inst_9340 ( .A1(net_13517), .ZN(net_12212), .A2(net_9948) );
NAND3_X2 inst_6282 ( .ZN(net_12897), .A3(net_9099), .A1(net_7660), .A2(net_7553) );
NAND2_X2 inst_10076 ( .ZN(net_12122), .A1(net_7878), .A2(net_7825) );
NAND2_X2 inst_10955 ( .ZN(net_19748), .A2(net_5088), .A1(net_2044) );
INV_X4 inst_13318 ( .A(net_15457), .ZN(net_11576) );
NAND2_X2 inst_12111 ( .A2(net_325), .ZN(net_302), .A1(net_301) );
CLKBUF_X2 inst_22671 ( .A(net_22542), .Z(net_22543) );
INV_X4 inst_17598 ( .A(net_20851), .ZN(net_733) );
INV_X2 inst_19026 ( .A(net_10426), .ZN(net_4924) );
INV_X4 inst_13876 ( .ZN(net_9158), .A(net_7374) );
INV_X2 inst_18477 ( .ZN(net_12630), .A(net_12629) );
INV_X4 inst_17051 ( .ZN(net_9148), .A(net_4890) );
AND2_X4 inst_21166 ( .ZN(net_20286), .A1(net_14542), .A2(net_13125) );
INV_X4 inst_12586 ( .ZN(net_18136), .A(net_18135) );
NAND3_X2 inst_6244 ( .ZN(net_13175), .A2(net_13174), .A3(net_13173), .A1(net_8677) );
NAND2_X2 inst_8753 ( .A1(net_16357), .ZN(net_15914), .A2(net_15513) );
NOR2_X2 inst_4174 ( .A1(net_9183), .ZN(net_8157), .A2(net_5047) );
INV_X4 inst_17841 ( .A(net_1697), .ZN(net_1461) );
INV_X4 inst_15133 ( .ZN(net_4070), .A(net_2338) );
NAND3_X2 inst_6369 ( .ZN(net_12074), .A1(net_11908), .A3(net_9434), .A2(net_8248) );
OAI211_X2 inst_2502 ( .ZN(net_12785), .C1(net_12784), .B(net_11602), .C2(net_10236), .A(net_7809) );
AOI21_X2 inst_20932 ( .ZN(net_6800), .B2(net_4230), .B1(net_2578), .A(net_1084) );
INV_X4 inst_17473 ( .A(net_20897), .ZN(net_864) );
NAND2_X2 inst_9114 ( .ZN(net_19914), .A1(net_15666), .A2(net_13577) );
NAND2_X2 inst_11233 ( .ZN(net_12025), .A1(net_4074), .A2(net_3945) );
NOR2_X2 inst_3974 ( .ZN(net_8403), .A1(net_8402), .A2(net_8360) );
INV_X4 inst_17425 ( .A(net_761), .ZN(net_495) );
INV_X4 inst_13290 ( .ZN(net_13600), .A(net_12402) );
INV_X4 inst_12601 ( .ZN(net_18129), .A(net_18112) );
XNOR2_X2 inst_213 ( .B(net_21203), .A(net_20071), .ZN(net_17543) );
NAND2_X2 inst_11501 ( .ZN(net_3539), .A2(net_1746), .A1(net_85) );
INV_X4 inst_18167 ( .A(net_21136), .ZN(net_16836) );
INV_X2 inst_18408 ( .ZN(net_19237), .A(net_16296) );
XNOR2_X2 inst_205 ( .ZN(net_17705), .A(net_17413), .B(net_17220) );
OAI21_X2 inst_1645 ( .A(net_16260), .ZN(net_15915), .B2(net_15398), .B1(net_15061) );
NAND2_X2 inst_7904 ( .ZN(net_18477), .A2(net_18400), .A1(net_18338) );
CLKBUF_X2 inst_21532 ( .A(net_21271), .Z(net_21404) );
NOR2_X2 inst_3722 ( .ZN(net_10967), .A2(net_9361), .A1(net_7578) );
NAND2_X2 inst_8043 ( .ZN(net_18236), .A2(net_18218), .A1(net_17806) );
NAND4_X2 inst_5410 ( .ZN(net_14607), .A2(net_12027), .A4(net_9947), .A1(net_9559), .A3(net_6721) );
NOR2_X2 inst_4311 ( .ZN(net_9845), .A1(net_9571), .A2(net_5899) );
INV_X4 inst_15618 ( .ZN(net_3449), .A(net_2163) );
CLKBUF_X2 inst_21993 ( .A(net_21864), .Z(net_21865) );
INV_X4 inst_14469 ( .ZN(net_6055), .A(net_5687) );
INV_X4 inst_14916 ( .ZN(net_4586), .A(net_3567) );
AOI21_X2 inst_20854 ( .A(net_9762), .ZN(net_9044), .B1(net_8982), .B2(net_8951) );
NAND4_X4 inst_5173 ( .ZN(net_20515), .A1(net_16386), .A4(net_16215), .A2(net_15970), .A3(net_13829) );
INV_X4 inst_14117 ( .ZN(net_6145), .A(net_6144) );
INV_X4 inst_15388 ( .ZN(net_3413), .A(net_2550) );
NAND3_X2 inst_6464 ( .ZN(net_11362), .A2(net_11245), .A3(net_11243), .A1(net_5639) );
NOR2_X4 inst_2951 ( .ZN(net_13065), .A1(net_5179), .A2(net_2996) );
NAND2_X2 inst_9176 ( .ZN(net_13344), .A1(net_13343), .A2(net_10456) );
CLKBUF_X2 inst_21557 ( .A(net_21270), .Z(net_21429) );
NOR2_X2 inst_3890 ( .ZN(net_9242), .A1(net_6113), .A2(net_4782) );
CLKBUF_X2 inst_21719 ( .A(net_21590), .Z(net_21591) );
INV_X4 inst_13526 ( .ZN(net_20366), .A(net_9323) );
NAND2_X2 inst_10209 ( .ZN(net_11663), .A1(net_11426), .A2(net_7979) );
OAI211_X2 inst_2535 ( .ZN(net_11252), .A(net_11251), .C1(net_10415), .C2(net_9985), .B(net_5189) );
NOR2_X2 inst_4569 ( .A2(net_4908), .A1(net_4802), .ZN(net_3871) );
INV_X2 inst_18873 ( .ZN(net_6236), .A(net_6235) );
INV_X8 inst_12393 ( .ZN(net_1533), .A(net_938) );
NOR2_X2 inst_4480 ( .A1(net_10292), .ZN(net_5446), .A2(net_4355) );
AOI21_X2 inst_20518 ( .B1(net_14622), .ZN(net_14570), .B2(net_12078), .A(net_8898) );
NAND3_X2 inst_6676 ( .ZN(net_7752), .A2(net_7751), .A3(net_7750), .A1(net_5895) );
NAND2_X2 inst_10723 ( .A1(net_10815), .A2(net_5958), .ZN(net_5876) );
NAND2_X2 inst_9378 ( .ZN(net_11963), .A1(net_11962), .A2(net_9859) );
INV_X4 inst_18058 ( .A(net_20856), .ZN(net_16390) );
INV_X4 inst_17536 ( .A(net_14568), .ZN(net_13058) );
NAND3_X2 inst_5639 ( .A1(net_19493), .ZN(net_18078), .A2(net_18048), .A3(net_13679) );
NOR2_X2 inst_3502 ( .ZN(net_14036), .A2(net_11716), .A1(net_2302) );
NOR2_X2 inst_3473 ( .ZN(net_14453), .A2(net_12779), .A1(net_9629) );
INV_X4 inst_14584 ( .ZN(net_9506), .A(net_4490) );
AND2_X2 inst_21323 ( .A2(net_10426), .ZN(net_6783), .A1(net_6782) );
INV_X4 inst_18160 ( .A(net_21162), .ZN(net_17426) );
NAND3_X2 inst_6018 ( .ZN(net_14385), .A3(net_14384), .A2(net_13620), .A1(net_12895) );
NAND2_X2 inst_9942 ( .ZN(net_12125), .A2(net_7826), .A1(net_3700) );
INV_X4 inst_14644 ( .ZN(net_18577), .A(net_18025) );
NAND2_X2 inst_8502 ( .ZN(net_17063), .A2(net_16606), .A1(net_16472) );
DFF_X1 inst_19791 ( .D(net_18627), .CK(net_22121), .Q(x546) );
INV_X4 inst_17556 ( .ZN(net_5450), .A(net_90) );
NAND3_X2 inst_5822 ( .ZN(net_15584), .A1(net_14958), .A3(net_12736), .A2(net_2963) );
INV_X2 inst_19123 ( .ZN(net_4392), .A(net_4391) );
NAND3_X2 inst_6448 ( .ZN(net_11765), .A2(net_11764), .A3(net_11763), .A1(net_5892) );
INV_X4 inst_16013 ( .ZN(net_20249), .A(net_15790) );
CLKBUF_X2 inst_21492 ( .A(net_21363), .Z(net_21364) );
XNOR2_X2 inst_348 ( .ZN(net_16940), .A(net_16748), .B(net_5738) );
NAND2_X4 inst_7676 ( .ZN(net_815), .A1(net_159), .A2(net_153) );
NAND2_X2 inst_8737 ( .A1(net_16390), .ZN(net_16025), .A2(net_15723) );
NOR2_X2 inst_5123 ( .A2(net_312), .ZN(net_280), .A1(net_279) );
NOR3_X2 inst_2686 ( .ZN(net_14358), .A2(net_14357), .A1(net_12604), .A3(net_10718) );
INV_X4 inst_14911 ( .ZN(net_6126), .A(net_3578) );
CLKBUF_X2 inst_21640 ( .A(net_21511), .Z(net_21512) );
NAND2_X2 inst_10774 ( .ZN(net_10618), .A2(net_7151), .A1(net_6854) );
NOR2_X2 inst_3740 ( .ZN(net_10673), .A1(net_10672), .A2(net_8549) );
OAI21_X2 inst_2293 ( .ZN(net_6496), .B2(net_4664), .A(net_3827), .B1(net_2598) );
NAND2_X2 inst_9600 ( .ZN(net_10758), .A2(net_10757), .A1(net_4288) );
CLKBUF_X2 inst_21816 ( .A(net_21687), .Z(net_21688) );
NAND2_X2 inst_11299 ( .ZN(net_9652), .A1(net_6647), .A2(net_2783) );
INV_X4 inst_18108 ( .A(net_21022), .ZN(net_694) );
XNOR2_X2 inst_645 ( .B(net_516), .ZN(net_393), .A(net_392) );
INV_X4 inst_13299 ( .ZN(net_12329), .A(net_12328) );
INV_X4 inst_15615 ( .A(net_15955), .ZN(net_15818) );
CLKBUF_X2 inst_21710 ( .A(net_21581), .Z(net_21582) );
NOR2_X4 inst_3041 ( .A2(net_20868), .ZN(net_5092), .A1(net_4989) );
INV_X4 inst_14967 ( .ZN(net_4843), .A(net_3430) );
NOR3_X2 inst_2719 ( .ZN(net_13309), .A2(net_11221), .A1(net_10507), .A3(net_7847) );
OAI21_X2 inst_2352 ( .ZN(net_3343), .B1(net_3342), .A(net_2527), .B2(net_1302) );
XNOR2_X2 inst_269 ( .B(net_21181), .A(net_20499), .ZN(net_17219) );
CLKBUF_X2 inst_21907 ( .A(net_21720), .Z(net_21779) );
NAND2_X4 inst_6864 ( .A2(net_19392), .A1(net_19391), .ZN(net_18377) );
INV_X4 inst_17125 ( .ZN(net_775), .A(net_774) );
INV_X4 inst_12534 ( .ZN(net_18381), .A(net_18380) );
INV_X4 inst_14278 ( .A(net_9035), .ZN(net_5656) );
INV_X2 inst_18383 ( .ZN(net_20194), .A(net_16550) );
INV_X4 inst_15947 ( .ZN(net_11536), .A(net_6346) );
INV_X2 inst_19370 ( .ZN(net_2209), .A(net_2208) );
NAND2_X2 inst_9796 ( .A1(net_10449), .ZN(net_9708), .A2(net_9707) );
XNOR2_X2 inst_514 ( .B(net_15585), .ZN(net_5791), .A(net_3422) );
AND2_X4 inst_21212 ( .A1(net_11296), .ZN(net_7826), .A2(net_6572) );
OAI21_X2 inst_1541 ( .ZN(net_17900), .B2(net_17851), .A(net_17696), .B1(net_17695) );
INV_X4 inst_12707 ( .ZN(net_17573), .A(net_17572) );
INV_X4 inst_15867 ( .ZN(net_2042), .A(net_1802) );
NOR2_X2 inst_4236 ( .ZN(net_7828), .A1(net_5308), .A2(net_4817) );
CLKBUF_X2 inst_21378 ( .A(net_21249), .Z(net_21250) );
INV_X2 inst_19437 ( .A(net_8326), .ZN(net_1721) );
CLKBUF_X2 inst_21480 ( .A(net_21351), .Z(net_21352) );
INV_X4 inst_16828 ( .ZN(net_1418), .A(net_830) );
CLKBUF_X2 inst_21518 ( .A(net_21389), .Z(net_21390) );
INV_X4 inst_12952 ( .ZN(net_16698), .A(net_16543) );
AOI21_X2 inst_20514 ( .B1(net_20667), .ZN(net_14604), .A(net_13904), .B2(net_8618) );
INV_X4 inst_14061 ( .A(net_7995), .ZN(net_7604) );
NOR2_X2 inst_4656 ( .A2(net_10672), .ZN(net_3662), .A1(net_3309) );
NAND2_X2 inst_10658 ( .ZN(net_6312), .A2(net_6311), .A1(net_2689) );
INV_X4 inst_14358 ( .ZN(net_5238), .A(net_4199) );
NAND3_X4 inst_5621 ( .ZN(net_19653), .A3(net_9799), .A1(net_9445), .A2(net_7109) );
NAND2_X2 inst_10636 ( .A1(net_13196), .ZN(net_6424), .A2(net_3939) );
NAND2_X2 inst_11585 ( .ZN(net_20589), .A2(net_4343), .A1(net_2710) );
NOR2_X2 inst_3432 ( .ZN(net_19611), .A1(net_15285), .A2(net_14267) );
INV_X4 inst_14047 ( .ZN(net_9500), .A(net_6256) );
INV_X4 inst_15760 ( .A(net_12306), .ZN(net_8611) );
INV_X4 inst_13984 ( .ZN(net_7827), .A(net_6566) );
INV_X4 inst_15211 ( .A(net_4272), .ZN(net_2893) );
NAND2_X2 inst_8959 ( .ZN(net_14710), .A1(net_14709), .A2(net_13290) );
NAND2_X4 inst_6881 ( .ZN(net_18263), .A1(net_18121), .A2(net_18108) );
NOR2_X2 inst_3840 ( .ZN(net_11010), .A2(net_9610), .A1(net_7244) );
AOI22_X2 inst_20005 ( .B1(net_13030), .ZN(net_12929), .A1(net_12928), .A2(net_12927), .B2(net_8813) );
NAND2_X2 inst_8905 ( .ZN(net_15041), .A2(net_14044), .A1(net_6535) );
NAND2_X2 inst_9477 ( .ZN(net_13778), .A1(net_11461), .A2(net_9379) );
INV_X4 inst_13852 ( .ZN(net_9140), .A(net_7466) );
INV_X4 inst_16695 ( .ZN(net_6896), .A(net_5432) );
NAND2_X4 inst_6973 ( .ZN(net_20774), .A2(net_20189), .A1(net_20188) );
AOI21_X2 inst_20710 ( .B2(net_13941), .ZN(net_12073), .B1(net_12072), .A(net_11461) );
NAND4_X2 inst_5333 ( .ZN(net_15555), .A1(net_14650), .A4(net_14531), .A3(net_14391), .A2(net_13356) );
CLKBUF_X2 inst_21574 ( .A(net_21445), .Z(net_21446) );
INV_X4 inst_17553 ( .A(net_657), .ZN(net_366) );
NAND2_X4 inst_7170 ( .A1(net_19984), .ZN(net_12987), .A2(net_6712) );
NOR2_X2 inst_4944 ( .ZN(net_1706), .A2(net_1705), .A1(net_1135) );
INV_X4 inst_13971 ( .ZN(net_7949), .A(net_5420) );
NAND2_X2 inst_10975 ( .ZN(net_13320), .A2(net_4967), .A1(net_170) );
NAND2_X2 inst_10259 ( .A1(net_20532), .ZN(net_15844), .A2(net_7992) );
XNOR2_X2 inst_312 ( .A(net_17092), .ZN(net_17085), .B(net_10805) );
INV_X4 inst_13429 ( .ZN(net_9883), .A(net_8443) );
NAND2_X2 inst_9554 ( .ZN(net_11013), .A1(net_11012), .A2(net_8398) );
INV_X4 inst_17829 ( .ZN(net_293), .A(net_104) );
XNOR2_X2 inst_309 ( .B(net_21163), .A(net_17092), .ZN(net_17089) );
NOR2_X2 inst_3416 ( .ZN(net_15600), .A2(net_14912), .A1(net_12279) );
CLKBUF_X2 inst_22203 ( .A(net_22074), .Z(net_22075) );
INV_X4 inst_13765 ( .ZN(net_10927), .A(net_7606) );
AOI21_X4 inst_20204 ( .B1(net_19924), .ZN(net_19633), .B2(net_14769), .A(net_12355) );
NAND2_X2 inst_9365 ( .A1(net_12944), .ZN(net_12130), .A2(net_12129) );
NAND2_X4 inst_7265 ( .ZN(net_12976), .A1(net_6274), .A2(net_6273) );
NAND2_X2 inst_8038 ( .ZN(net_18254), .A2(net_18175), .A1(net_17286) );
NOR3_X2 inst_2694 ( .ZN(net_14221), .A1(net_12643), .A2(net_9496), .A3(net_7518) );
NAND2_X2 inst_9833 ( .ZN(net_9592), .A1(net_9591), .A2(net_7537) );
INV_X4 inst_15207 ( .ZN(net_5210), .A(net_2901) );
INV_X2 inst_19366 ( .A(net_3038), .ZN(net_2238) );
OAI21_X2 inst_1968 ( .ZN(net_12256), .B1(net_10886), .B2(net_8498), .A(net_7272) );
CLKBUF_X2 inst_22679 ( .A(net_22550), .Z(net_22551) );
INV_X4 inst_12983 ( .A(net_17760), .ZN(net_17625) );
INV_X8 inst_12168 ( .ZN(net_18670), .A(net_18639) );
OAI221_X2 inst_1330 ( .ZN(net_19388), .B2(net_15844), .C1(net_15790), .C2(net_14932), .B1(net_10930), .A(net_9449) );
NAND2_X2 inst_12038 ( .ZN(net_3484), .A1(net_761), .A2(net_107) );
INV_X4 inst_17903 ( .ZN(net_19027), .A(net_1697) );
INV_X4 inst_13728 ( .ZN(net_7779), .A(net_6539) );
INV_X4 inst_13963 ( .ZN(net_8651), .A(net_5444) );
INV_X8 inst_12410 ( .A(net_1733), .ZN(net_965) );
OAI21_X2 inst_1898 ( .A(net_14600), .ZN(net_13358), .B1(net_8862), .B2(net_8572) );
INV_X4 inst_15644 ( .ZN(net_11380), .A(net_9926) );
NAND3_X2 inst_6275 ( .ZN(net_12909), .A1(net_12908), .A3(net_12907), .A2(net_5957) );
OAI21_X2 inst_1714 ( .B2(net_20259), .B1(net_20258), .ZN(net_19239), .A(net_15191) );
NAND2_X2 inst_8551 ( .A1(net_16965), .ZN(net_16791), .A2(net_16497) );
NAND2_X2 inst_9164 ( .ZN(net_13376), .A1(net_13375), .A2(net_10577) );
INV_X4 inst_14630 ( .A(net_4934), .ZN(net_4594) );
NAND2_X2 inst_9428 ( .ZN(net_11615), .A1(net_11614), .A2(net_11038) );
AOI21_X4 inst_20117 ( .B2(net_20904), .ZN(net_20749), .B1(net_20272), .A(net_15241) );
NOR2_X2 inst_4777 ( .ZN(net_11253), .A1(net_8490), .A2(net_2395) );
INV_X4 inst_15789 ( .A(net_13576), .ZN(net_8959) );
NAND2_X2 inst_10762 ( .ZN(net_6714), .A2(net_5515), .A1(net_3187) );
NAND2_X2 inst_10851 ( .A2(net_5709), .ZN(net_5464), .A1(net_154) );
INV_X4 inst_15333 ( .A(net_4151), .ZN(net_2604) );
OAI21_X4 inst_1496 ( .B1(net_20415), .ZN(net_19265), .A(net_14022), .B2(net_12147) );
NAND2_X2 inst_11292 ( .ZN(net_8515), .A1(net_4032), .A2(net_2084) );
NAND2_X2 inst_9091 ( .A1(net_15046), .ZN(net_13793), .A2(net_12560) );
NOR2_X2 inst_4297 ( .ZN(net_5965), .A2(net_4538), .A1(net_1773) );
NAND2_X2 inst_9381 ( .ZN(net_11937), .A2(net_8929), .A1(net_7934) );
INV_X4 inst_13005 ( .A(net_16577), .ZN(net_16443) );
OAI21_X2 inst_1565 ( .ZN(net_16932), .B2(net_16762), .B1(net_16716), .A(net_16454) );
SDFF_X2 inst_924 ( .Q(net_21220), .D(net_16502), .SE(net_263), .CK(net_21520), .SI(x7366) );
AOI22_X2 inst_19961 ( .ZN(net_16192), .A2(net_15870), .A1(net_15369), .B2(net_14317), .B1(net_4364) );
INV_X2 inst_19461 ( .ZN(net_2250), .A(net_1198) );
XNOR2_X2 inst_287 ( .A(net_17170), .ZN(net_17152), .B(net_16921) );
NAND2_X2 inst_10614 ( .ZN(net_8713), .A2(net_6594), .A1(net_1274) );
AOI21_X2 inst_20614 ( .ZN(net_13658), .B2(net_13657), .B1(net_12888), .A(net_6994) );
NAND2_X2 inst_7929 ( .ZN(net_18442), .A2(net_18352), .A1(net_17266) );
INV_X4 inst_16144 ( .ZN(net_3301), .A(net_2135) );
NAND2_X2 inst_12030 ( .A1(net_20865), .A2(net_1959), .ZN(net_1111) );
NOR2_X4 inst_3094 ( .ZN(net_9973), .A1(net_4228), .A2(net_2601) );
INV_X4 inst_16305 ( .ZN(net_3206), .A(net_1326) );
NOR2_X4 inst_2903 ( .ZN(net_10661), .A2(net_9098), .A1(net_5659) );
INV_X4 inst_13830 ( .ZN(net_12530), .A(net_7499) );
NOR2_X2 inst_4045 ( .A2(net_20528), .ZN(net_11733), .A1(net_7232) );
INV_X4 inst_16749 ( .ZN(net_10274), .A(net_749) );
INV_X4 inst_12623 ( .ZN(net_20166), .A(net_17991) );
NOR2_X2 inst_4890 ( .ZN(net_6446), .A2(net_1514), .A1(net_170) );
SDFF_X2 inst_984 ( .QN(net_21037), .D(net_456), .SE(net_263), .CK(net_21963), .SI(x2367) );
NAND3_X2 inst_6734 ( .ZN(net_6477), .A2(net_6476), .A1(net_4197), .A3(net_1553) );
OAI21_X2 inst_2064 ( .ZN(net_10679), .B1(net_9430), .B2(net_5589), .A(net_4264) );
INV_X4 inst_14604 ( .ZN(net_9002), .A(net_5567) );
INV_X2 inst_19267 ( .ZN(net_3081), .A(net_3080) );
INV_X2 inst_18546 ( .ZN(net_10971), .A(net_10970) );
INV_X4 inst_15057 ( .ZN(net_11317), .A(net_3307) );
OAI22_X2 inst_1292 ( .A2(net_12520), .ZN(net_12479), .B2(net_12478), .A1(net_9989), .B1(net_1965) );
INV_X4 inst_15769 ( .A(net_15840), .ZN(net_1923) );
NOR2_X2 inst_5014 ( .ZN(net_13996), .A2(net_1253), .A1(net_855) );
OAI21_X2 inst_1963 ( .ZN(net_12403), .B2(net_7372), .A(net_5872), .B1(net_2211) );
SDFF_X1 inst_1056 ( .QN(net_21080), .D(net_440), .SE(net_263), .CK(net_22634), .SI(x1718) );
NAND2_X2 inst_11818 ( .ZN(net_1820), .A2(net_1789), .A1(net_227) );
INV_X2 inst_18611 ( .ZN(net_11622), .A(net_10284) );
INV_X4 inst_17401 ( .ZN(net_8664), .A(net_60) );
NOR2_X2 inst_4247 ( .ZN(net_7539), .A1(net_6856), .A2(net_6436) );
NOR2_X2 inst_3648 ( .ZN(net_11676), .A2(net_11675), .A1(net_8105) );
INV_X2 inst_19571 ( .ZN(net_756), .A(net_445) );
CLKBUF_X2 inst_21571 ( .A(net_21334), .Z(net_21443) );
INV_X4 inst_14434 ( .A(net_5021), .ZN(net_5020) );
INV_X4 inst_14359 ( .A(net_16054), .ZN(net_9256) );
CLKBUF_X2 inst_22278 ( .A(net_22149), .Z(net_22150) );
NAND3_X2 inst_6524 ( .A2(net_11224), .ZN(net_10622), .A1(net_10593), .A3(net_7848) );
NOR2_X2 inst_4988 ( .A2(net_1934), .ZN(net_1432), .A1(net_308) );
NAND2_X2 inst_11325 ( .A1(net_8160), .ZN(net_6558), .A2(net_2655) );
INV_X4 inst_15074 ( .A(net_3509), .ZN(net_3273) );
INV_X4 inst_14216 ( .A(net_12457), .ZN(net_5865) );
INV_X4 inst_17815 ( .ZN(net_232), .A(net_115) );
AOI21_X2 inst_20818 ( .ZN(net_19747), .B1(net_9322), .B2(net_6269), .A(net_5936) );
NAND2_X2 inst_11677 ( .A1(net_4155), .ZN(net_2351), .A2(net_2350) );
INV_X4 inst_14996 ( .ZN(net_6720), .A(net_3395) );
INV_X4 inst_18170 ( .A(net_20904), .ZN(net_16210) );
NAND2_X2 inst_11559 ( .A2(net_7399), .ZN(net_2830), .A1(net_1532) );
NAND2_X2 inst_10064 ( .ZN(net_13152), .A1(net_8676), .A2(net_8675) );
NAND2_X2 inst_10999 ( .A2(net_4902), .ZN(net_4901), .A1(net_4900) );
CLKBUF_X2 inst_21821 ( .A(net_21428), .Z(net_21693) );
NAND2_X2 inst_9077 ( .ZN(net_13832), .A2(net_12730), .A1(net_1077) );
CLKBUF_X2 inst_21838 ( .A(net_21709), .Z(net_21710) );
NAND2_X2 inst_9023 ( .A1(net_15158), .ZN(net_14156), .A2(net_12274) );
INV_X2 inst_19309 ( .A(net_3884), .ZN(net_2721) );
NAND2_X2 inst_10244 ( .A1(net_13350), .ZN(net_10204), .A2(net_6250) );
INV_X4 inst_12714 ( .ZN(net_17610), .A(net_17550) );
NAND2_X4 inst_7650 ( .A1(net_1581), .ZN(net_1204), .A2(net_795) );
INV_X4 inst_14750 ( .ZN(net_8039), .A(net_5467) );
INV_X4 inst_17876 ( .ZN(net_4850), .A(net_2673) );
NAND2_X2 inst_8296 ( .ZN(net_20595), .A2(net_18684), .A1(net_16684) );
NAND2_X1 inst_12160 ( .A1(net_20477), .ZN(net_1444), .A2(net_1112) );
INV_X8 inst_12246 ( .ZN(net_4109), .A(net_3790) );
OAI21_X2 inst_1590 ( .ZN(net_20294), .A(net_16402), .B2(net_15940), .B1(net_12933) );
INV_X4 inst_17353 ( .ZN(net_5342), .A(net_549) );
NAND2_X4 inst_7591 ( .ZN(net_20802), .A1(net_1513), .A2(net_1026) );
CLKBUF_X2 inst_21801 ( .A(net_21672), .Z(net_21673) );
NAND3_X2 inst_6229 ( .ZN(net_13228), .A3(net_12131), .A2(net_11076), .A1(net_8598) );
NAND2_X2 inst_10648 ( .ZN(net_9829), .A1(net_6358), .A2(net_6357) );
NAND2_X2 inst_10931 ( .A1(net_9367), .ZN(net_5214), .A2(net_2912) );
INV_X4 inst_18093 ( .A(net_20858), .ZN(net_86) );
NAND4_X2 inst_5347 ( .ZN(net_15434), .A1(net_14553), .A4(net_14281), .A3(net_11369), .A2(net_9197) );
OAI21_X2 inst_2318 ( .A(net_12001), .ZN(net_5682), .B2(net_5681), .B1(net_2207) );
XNOR2_X2 inst_399 ( .ZN(net_16702), .A(net_16701), .B(net_16700) );
INV_X8 inst_12433 ( .A(net_20071), .ZN(net_20070) );
NOR2_X2 inst_3957 ( .ZN(net_8597), .A1(net_8596), .A2(net_6517) );
NOR2_X2 inst_4020 ( .ZN(net_9567), .A2(net_8023), .A1(net_1037) );
NAND2_X2 inst_9953 ( .ZN(net_8934), .A1(net_8933), .A2(net_8113) );
INV_X4 inst_13404 ( .ZN(net_13970), .A(net_8934) );
INV_X4 inst_17014 ( .ZN(net_1582), .A(net_192) );
OAI22_X2 inst_1299 ( .ZN(net_11271), .B1(net_11270), .B2(net_11269), .A1(net_9278), .A2(net_5861) );
CLKBUF_X2 inst_21601 ( .A(net_21341), .Z(net_21473) );
NAND3_X2 inst_6450 ( .ZN(net_11760), .A2(net_11759), .A1(net_9580), .A3(net_8571) );
NAND2_X2 inst_8404 ( .A2(net_17498), .ZN(net_17248), .A1(net_17247) );
NAND2_X2 inst_10404 ( .A1(net_11830), .ZN(net_7273), .A2(net_7272) );
INV_X4 inst_13487 ( .ZN(net_11542), .A(net_9523) );
INV_X4 inst_17133 ( .ZN(net_11045), .A(net_4264) );
XNOR2_X2 inst_674 ( .A(net_21156), .B(net_21124), .ZN(net_1674) );
INV_X4 inst_14683 ( .ZN(net_4428), .A(net_4296) );
NAND4_X2 inst_5259 ( .A4(net_20328), .A1(net_20327), .ZN(net_16302), .A2(net_13858), .A3(net_13085) );
NAND4_X2 inst_5518 ( .A1(net_11743), .ZN(net_9886), .A3(net_9885), .A2(net_8714), .A4(net_4824) );
INV_X4 inst_14151 ( .ZN(net_6031), .A(net_6030) );
NAND2_X2 inst_10859 ( .ZN(net_8962), .A1(net_5449), .A2(net_4011) );
OAI21_X2 inst_2253 ( .ZN(net_19506), .A(net_11541), .B2(net_6752), .B1(net_3603) );
INV_X4 inst_13670 ( .ZN(net_8054), .A(net_8053) );
INV_X4 inst_18148 ( .A(net_21078), .ZN(net_378) );
NAND2_X2 inst_10115 ( .ZN(net_8423), .A2(net_7807), .A1(net_7062) );
NAND2_X2 inst_9674 ( .ZN(net_13813), .A1(net_10279), .A2(net_8173) );
INV_X4 inst_16255 ( .ZN(net_1628), .A(net_1355) );
NOR2_X4 inst_2868 ( .ZN(net_14357), .A2(net_11015), .A1(net_7862) );
NAND3_X2 inst_6522 ( .A3(net_12118), .A1(net_11065), .ZN(net_10633), .A2(net_7343) );
INV_X8 inst_12254 ( .ZN(net_3359), .A(net_2281) );
INV_X4 inst_18031 ( .A(net_21172), .ZN(net_17253) );
INV_X4 inst_14549 ( .ZN(net_4607), .A(net_4606) );
INV_X8 inst_12261 ( .ZN(net_3924), .A(net_2568) );
AOI21_X2 inst_20295 ( .B2(net_19914), .B1(net_19913), .A(net_16359), .ZN(net_16153) );
OAI21_X2 inst_1832 ( .B1(net_20205), .ZN(net_14076), .A(net_14075), .B2(net_10352) );
INV_X4 inst_13241 ( .A(net_13589), .ZN(net_13389) );
NOR2_X2 inst_4562 ( .A1(net_20457), .ZN(net_4852), .A2(net_3937) );
XNOR2_X2 inst_640 ( .B(net_16680), .ZN(net_414), .A(net_413) );
INV_X4 inst_15740 ( .A(net_12100), .ZN(net_11654) );
NAND2_X2 inst_9893 ( .ZN(net_11555), .A2(net_7560), .A1(net_7007) );
NAND2_X4 inst_7500 ( .ZN(net_4226), .A2(net_2296), .A1(net_225) );
INV_X4 inst_17785 ( .A(net_855), .ZN(net_449) );
INV_X4 inst_16932 ( .A(net_14945), .ZN(net_12275) );
OAI21_X4 inst_1478 ( .A(net_14678), .ZN(net_14677), .B2(net_11946), .B1(net_11698) );
NAND3_X2 inst_6098 ( .ZN(net_13917), .A3(net_13165), .A1(net_11434), .A2(net_10964) );
INV_X2 inst_18500 ( .ZN(net_12158), .A(net_12157) );
CLKBUF_X2 inst_21832 ( .A(net_21570), .Z(net_21704) );
NAND2_X2 inst_9535 ( .A1(net_15012), .ZN(net_12411), .A2(net_7515) );
INV_X4 inst_17717 ( .A(net_20897), .ZN(net_197) );
NAND2_X2 inst_9085 ( .ZN(net_19579), .A1(net_13811), .A2(net_13810) );
INV_X4 inst_12957 ( .ZN(net_16909), .A(net_16727) );
INV_X4 inst_16661 ( .ZN(net_1538), .A(net_1083) );
NAND3_X2 inst_6075 ( .ZN(net_14107), .A1(net_12299), .A3(net_9081), .A2(net_8885) );
INV_X4 inst_13739 ( .ZN(net_12734), .A(net_7644) );
INV_X4 inst_16977 ( .ZN(net_6696), .A(net_3009) );
INV_X4 inst_16742 ( .ZN(net_19929), .A(net_864) );
OAI21_X2 inst_2089 ( .ZN(net_10308), .B2(net_6283), .B1(net_4850), .A(net_4068) );
INV_X4 inst_15128 ( .ZN(net_3143), .A(net_3142) );
NAND2_X2 inst_11378 ( .ZN(net_3549), .A1(net_3548), .A2(net_1917) );
INV_X4 inst_16775 ( .ZN(net_8629), .A(net_5449) );
OAI21_X2 inst_1679 ( .B1(net_15706), .ZN(net_15488), .B2(net_14569), .A(net_12212) );
INV_X4 inst_16280 ( .ZN(net_4179), .A(net_1341) );
OAI21_X2 inst_2215 ( .ZN(net_8523), .A(net_6863), .B1(net_5575), .B2(net_5366) );
OAI21_X2 inst_1855 ( .ZN(net_20683), .A(net_13554), .B1(net_10926), .B2(net_5718) );
XNOR2_X2 inst_337 ( .B(net_21121), .ZN(net_16986), .A(net_16985) );
NAND2_X2 inst_11564 ( .ZN(net_9632), .A2(net_2952), .A1(net_1487) );
AOI21_X2 inst_20306 ( .B2(net_19857), .B1(net_19856), .A(net_16187), .ZN(net_16070) );
INV_X4 inst_16575 ( .ZN(net_9591), .A(net_112) );
NAND2_X2 inst_11193 ( .ZN(net_5171), .A2(net_4083), .A1(net_573) );
NAND3_X2 inst_6220 ( .ZN(net_13242), .A3(net_12194), .A2(net_9473), .A1(net_8432) );
INV_X4 inst_15355 ( .ZN(net_4967), .A(net_2233) );
INV_X4 inst_13355 ( .A(net_11710), .ZN(net_10983) );
INV_X4 inst_13775 ( .ZN(net_7589), .A(net_7588) );
NAND2_X2 inst_9262 ( .A2(net_12624), .ZN(net_12621), .A1(net_12620) );
INV_X4 inst_17249 ( .ZN(net_863), .A(net_418) );
NAND2_X2 inst_7738 ( .A1(net_18840), .ZN(net_18808), .A2(net_18807) );
INV_X4 inst_18278 ( .A(net_20067), .ZN(net_20066) );
OAI211_X2 inst_2396 ( .ZN(net_16082), .C1(net_16076), .B(net_15554), .C2(net_12938), .A(net_11373) );
CLKBUF_X2 inst_21839 ( .A(net_21710), .Z(net_21711) );
NAND2_X2 inst_10232 ( .ZN(net_8049), .A1(net_8048), .A2(net_7729) );
INV_X4 inst_15704 ( .A(net_7659), .ZN(net_2003) );
INV_X2 inst_19583 ( .A(net_1369), .ZN(net_373) );
NAND2_X2 inst_10281 ( .ZN(net_19857), .A1(net_13023), .A2(net_5656) );
INV_X4 inst_14295 ( .ZN(net_5555), .A(net_5554) );
INV_X2 inst_18589 ( .ZN(net_10199), .A(net_10198) );
INV_X4 inst_14628 ( .ZN(net_20315), .A(net_4396) );
NAND3_X2 inst_5908 ( .ZN(net_15057), .A3(net_12921), .A1(net_11650), .A2(net_11445) );
XNOR2_X2 inst_246 ( .ZN(net_17317), .A(net_17312), .B(net_12268) );
NOR2_X2 inst_4443 ( .ZN(net_4803), .A1(net_4802), .A2(net_4801) );
XNOR2_X2 inst_635 ( .A(net_21200), .B(net_16836), .ZN(net_434) );
INV_X8 inst_12384 ( .ZN(net_289), .A(net_246) );
NAND3_X2 inst_5787 ( .A3(net_19744), .A1(net_19743), .ZN(net_15774), .A2(net_13347) );
CLKBUF_X2 inst_22268 ( .A(net_22139), .Z(net_22140) );
INV_X2 inst_19509 ( .ZN(net_1203), .A(net_216) );
NAND2_X2 inst_8510 ( .ZN(net_16920), .A1(net_16919), .A2(net_16619) );
NAND2_X2 inst_10569 ( .ZN(net_20038), .A1(net_10389), .A2(net_9529) );
INV_X4 inst_16208 ( .ZN(net_10386), .A(net_8252) );
INV_X4 inst_15140 ( .ZN(net_13350), .A(net_3251) );
XNOR2_X2 inst_519 ( .A(net_16265), .ZN(net_6374), .B(net_2401) );
NAND2_X4 inst_7641 ( .A1(net_1331), .ZN(net_1104), .A2(net_108) );
NOR2_X2 inst_3796 ( .ZN(net_10025), .A1(net_6907), .A2(net_6780) );
NAND2_X2 inst_9359 ( .ZN(net_12150), .A2(net_9884), .A1(net_6377) );
INV_X4 inst_12758 ( .ZN(net_17399), .A(net_17398) );
INV_X4 inst_18198 ( .A(net_20972), .ZN(net_225) );
INV_X8 inst_12174 ( .ZN(net_17681), .A(net_17653) );
AOI21_X2 inst_20286 ( .A(net_16404), .ZN(net_16245), .B2(net_15900), .B1(net_10157) );
SDFF_X2 inst_1053 ( .QN(net_21028), .D(net_593), .SE(net_263), .CK(net_21941), .SI(x2531) );
NOR2_X1 inst_5158 ( .ZN(net_971), .A2(net_938), .A1(net_258) );
NAND2_X4 inst_7231 ( .A1(net_20606), .ZN(net_14782), .A2(net_5712) );
INV_X4 inst_17639 ( .ZN(net_5748), .A(net_1435) );
NOR3_X2 inst_2774 ( .A2(net_15636), .A3(net_14083), .A1(net_8495), .ZN(net_7776) );
INV_X4 inst_14673 ( .ZN(net_18862), .A(net_18025) );
AOI21_X2 inst_20922 ( .A(net_15452), .B1(net_11925), .ZN(net_7213), .B2(net_2695) );
INV_X4 inst_17630 ( .ZN(net_288), .A(net_287) );
NAND2_X4 inst_6871 ( .A2(net_20324), .A1(net_20323), .ZN(net_18280) );
INV_X8 inst_12202 ( .ZN(net_12372), .A(net_11015) );
AOI21_X2 inst_20701 ( .A(net_14022), .ZN(net_12135), .B2(net_8386), .B1(net_7786) );
NOR2_X2 inst_4577 ( .ZN(net_4836), .A1(net_3852), .A2(net_3112) );
XNOR2_X2 inst_239 ( .ZN(net_17390), .B(net_17091), .A(net_16928) );
CLKBUF_X2 inst_21641 ( .A(net_21439), .Z(net_21513) );
INV_X2 inst_18449 ( .ZN(net_19672), .A(net_12639) );
INV_X4 inst_18098 ( .A(net_21169), .ZN(net_17774) );
AND2_X4 inst_21232 ( .ZN(net_19801), .A1(net_7836), .A2(net_4169) );
AND4_X4 inst_21093 ( .ZN(net_2525), .A3(net_2524), .A4(net_625), .A2(net_32), .A1(net_25) );
OR2_X2 inst_1193 ( .A2(net_7669), .ZN(net_5212), .A1(net_4783) );
INV_X4 inst_14770 ( .ZN(net_6732), .A(net_4051) );
INV_X4 inst_17703 ( .A(net_6692), .ZN(net_655) );
INV_X4 inst_18248 ( .A(net_21040), .ZN(net_610) );
NAND2_X2 inst_10582 ( .ZN(net_6675), .A1(net_6674), .A2(net_4923) );
INV_X4 inst_15228 ( .ZN(net_4616), .A(net_3449) );
INV_X8 inst_12395 ( .A(net_814), .ZN(net_185) );
NAND3_X2 inst_6091 ( .ZN(net_20258), .A1(net_12450), .A3(net_7130), .A2(net_4048) );
XNOR2_X2 inst_601 ( .B(net_17097), .ZN(net_537), .A(net_536) );
NAND2_X4 inst_7391 ( .A2(net_20859), .ZN(net_6895), .A1(net_4187) );
INV_X4 inst_13709 ( .ZN(net_11898), .A(net_7860) );
CLKBUF_X2 inst_21625 ( .A(net_21496), .Z(net_21497) );
INV_X2 inst_18852 ( .A(net_9075), .ZN(net_6593) );
NAND2_X2 inst_7952 ( .ZN(net_18400), .A2(net_18399), .A1(net_17997) );
NAND2_X2 inst_8097 ( .A2(net_20503), .ZN(net_18123), .A1(net_17290) );
OAI21_X2 inst_1773 ( .B2(net_20022), .B1(net_20021), .ZN(net_14690), .A(net_14689) );
NAND2_X2 inst_10133 ( .ZN(net_20430), .A1(net_11572), .A2(net_5440) );
NAND2_X2 inst_10278 ( .ZN(net_7955), .A2(net_7954), .A1(net_7917) );
OAI21_X2 inst_1583 ( .A(net_20952), .B2(net_19934), .B1(net_19933), .ZN(net_16305) );
SDFF_X2 inst_771 ( .Q(net_20866), .SE(net_18584), .SI(net_18488), .D(net_519), .CK(net_22175) );
NAND3_X2 inst_6325 ( .ZN(net_12512), .A3(net_12511), .A2(net_11391), .A1(net_2918) );
NAND2_X2 inst_11552 ( .ZN(net_20094), .A1(net_2861), .A2(net_2860) );
INV_X4 inst_16002 ( .A(net_9080), .ZN(net_2355) );
INV_X4 inst_15654 ( .ZN(net_3949), .A(net_1377) );
NAND2_X4 inst_7324 ( .ZN(net_8019), .A2(net_5097), .A1(net_4251) );
NAND2_X4 inst_7402 ( .ZN(net_5203), .A2(net_4037), .A1(net_2897) );
NAND2_X2 inst_9334 ( .ZN(net_12296), .A1(net_12295), .A2(net_8957) );
NAND2_X2 inst_8169 ( .A1(net_20107), .ZN(net_17956), .A2(net_17952) );
NAND2_X4 inst_7138 ( .ZN(net_11688), .A1(net_9807), .A2(net_7414) );
INV_X4 inst_12945 ( .ZN(net_16954), .A(net_16631) );
NAND3_X2 inst_5782 ( .ZN(net_15783), .A3(net_14794), .A2(net_13976), .A1(net_13086) );
INV_X4 inst_13873 ( .ZN(net_7423), .A(net_7422) );
CLKBUF_X2 inst_22871 ( .A(net_22742), .Z(net_22743) );
NAND2_X2 inst_10520 ( .ZN(net_10499), .A1(net_6861), .A2(net_6860) );
OAI22_X2 inst_1319 ( .ZN(net_4240), .A2(net_3102), .A1(net_2994), .B2(net_1605), .B1(net_1272) );
XNOR2_X2 inst_358 ( .ZN(net_16889), .A(net_16499), .B(net_158) );
NOR2_X2 inst_4462 ( .ZN(net_4551), .A2(net_4520), .A1(net_1473) );
OAI21_X2 inst_1756 ( .ZN(net_14789), .A(net_14788), .B2(net_13293), .B1(net_6928) );
INV_X4 inst_14037 ( .A(net_9900), .ZN(net_6271) );
INV_X4 inst_17041 ( .ZN(net_1059), .A(net_940) );
NAND3_X2 inst_6766 ( .ZN(net_20120), .A3(net_3903), .A1(net_2923), .A2(net_1637) );
NAND2_X2 inst_8794 ( .A1(net_15897), .ZN(net_15741), .A2(net_15368) );
NAND2_X4 inst_7108 ( .ZN(net_12633), .A1(net_11534), .A2(net_11016) );
NAND2_X2 inst_9309 ( .ZN(net_12364), .A1(net_12363), .A2(net_10769) );
INV_X4 inst_15215 ( .ZN(net_20257), .A(net_3344) );
INV_X4 inst_14177 ( .ZN(net_7464), .A(net_5991) );
XNOR2_X2 inst_655 ( .B(net_15588), .ZN(net_357), .A(net_356) );
NAND3_X2 inst_5914 ( .ZN(net_20586), .A2(net_13507), .A3(net_12793), .A1(net_10396) );
AOI21_X4 inst_20159 ( .ZN(net_15702), .B1(net_15366), .B2(net_15010), .A(net_14309) );
NAND3_X2 inst_5817 ( .A1(net_19953), .ZN(net_15604), .A3(net_12442), .A2(net_5963) );
NAND3_X2 inst_5934 ( .ZN(net_14925), .A3(net_13477), .A1(net_12316), .A2(net_4550) );
NAND2_X2 inst_8422 ( .ZN(net_17297), .A2(net_16923), .A1(net_16744) );
CLKBUF_X2 inst_22102 ( .A(net_21973), .Z(net_21974) );
CLKBUF_X2 inst_22571 ( .A(net_22442), .Z(net_22443) );
CLKBUF_X2 inst_22097 ( .A(net_21493), .Z(net_21969) );
NAND2_X2 inst_9373 ( .A1(net_20399), .ZN(net_12048), .A2(net_6612) );
AOI21_X2 inst_20947 ( .ZN(net_5862), .B1(net_5104), .A(net_4279), .B2(net_1754) );
NAND2_X2 inst_11316 ( .A1(net_5499), .ZN(net_5052), .A2(net_4275) );
NOR2_X2 inst_4438 ( .ZN(net_5906), .A2(net_4828), .A1(net_628) );
NAND3_X2 inst_6662 ( .A3(net_13968), .ZN(net_8450), .A2(net_6588), .A1(net_4195) );
INV_X2 inst_19557 ( .A(net_3704), .ZN(net_844) );
NAND2_X2 inst_8800 ( .ZN(net_20155), .A1(net_15969), .A2(net_15337) );
NAND3_X2 inst_6303 ( .ZN(net_12801), .A2(net_12800), .A1(net_10921), .A3(net_8137) );
NAND3_X4 inst_5623 ( .ZN(net_19650), .A3(net_19333), .A2(net_11159), .A1(net_10026) );
CLKBUF_X2 inst_21672 ( .A(net_21258), .Z(net_21544) );
CLKBUF_X2 inst_22857 ( .A(net_22728), .Z(net_22729) );
NAND2_X2 inst_9669 ( .A2(net_11822), .ZN(net_10312), .A1(net_8336) );
NAND2_X2 inst_11996 ( .ZN(net_5775), .A1(net_1741), .A2(net_465) );
XOR2_X2 inst_41 ( .A(net_21135), .Z(net_585), .B(net_584) );
NAND2_X2 inst_11516 ( .A1(net_3063), .ZN(net_2995), .A2(net_1838) );
AOI21_X2 inst_20408 ( .ZN(net_15330), .A(net_14802), .B1(net_14552), .B2(net_13720) );
NAND2_X2 inst_11743 ( .ZN(net_5240), .A1(net_1027), .A2(net_985) );
INV_X4 inst_12569 ( .A(net_18202), .ZN(net_18201) );
INV_X2 inst_18445 ( .ZN(net_13624), .A(net_12766) );
OAI21_X2 inst_1989 ( .B1(net_13274), .ZN(net_12029), .A(net_12028), .B2(net_11845) );
NAND2_X2 inst_11868 ( .ZN(net_1646), .A1(net_1645), .A2(net_1644) );
INV_X4 inst_13260 ( .ZN(net_19709), .A(net_11608) );
XNOR2_X2 inst_152 ( .ZN(net_17982), .B(net_17906), .A(net_17499) );
NAND2_X2 inst_9694 ( .ZN(net_10230), .A1(net_10229), .A2(net_8052) );
NAND3_X4 inst_5609 ( .ZN(net_19298), .A3(net_10492), .A2(net_7955), .A1(net_5489) );
NAND2_X2 inst_11111 ( .A1(net_9450), .ZN(net_8915), .A2(net_4321) );
NAND2_X4 inst_6944 ( .ZN(net_19010), .A1(net_18313), .A2(net_17235) );
INV_X8 inst_12314 ( .ZN(net_1783), .A(net_786) );
INV_X2 inst_18763 ( .ZN(net_7625), .A(net_7624) );
NAND3_X2 inst_6388 ( .ZN(net_12012), .A3(net_12011), .A2(net_11397), .A1(net_5150) );
OAI21_X4 inst_1400 ( .ZN(net_20729), .B2(net_20341), .B1(net_20340), .A(net_16242) );
INV_X4 inst_14374 ( .ZN(net_6290), .A(net_5178) );
NAND4_X4 inst_5233 ( .A1(net_18929), .ZN(net_18882), .A3(net_12232), .A2(net_9602), .A4(net_5801) );
XNOR2_X2 inst_89 ( .ZN(net_18563), .A(net_18496), .B(net_17821) );
AOI21_X2 inst_20279 ( .A(net_16644), .ZN(net_16303), .B2(net_16012), .B1(net_15483) );
OAI21_X2 inst_1520 ( .ZN(net_18380), .A(net_18233), .B2(net_18232), .B1(net_17187) );
OAI21_X2 inst_1535 ( .A(net_18582), .ZN(net_17945), .B2(net_17789), .B1(net_17688) );
INV_X4 inst_13609 ( .ZN(net_8437), .A(net_7083) );
INV_X4 inst_14112 ( .ZN(net_9709), .A(net_6155) );
INV_X2 inst_19419 ( .ZN(net_3914), .A(net_3068) );
SDFF_X2 inst_788 ( .Q(net_20884), .SE(net_18862), .SI(net_18034), .D(net_492), .CK(net_21802) );
INV_X4 inst_15525 ( .ZN(net_3632), .A(net_2395) );
NAND2_X4 inst_7526 ( .ZN(net_3762), .A2(net_2744), .A1(net_817) );
INV_X4 inst_13391 ( .ZN(net_10724), .A(net_10723) );
INV_X4 inst_17174 ( .ZN(net_4357), .A(net_734) );
NAND3_X2 inst_5990 ( .ZN(net_14534), .A2(net_14533), .A1(net_13373), .A3(net_12028) );
NAND4_X2 inst_5407 ( .ZN(net_20365), .A2(net_18895), .A1(net_18894), .A3(net_14642), .A4(net_6224) );
OAI21_X2 inst_1579 ( .A(net_20856), .B2(net_19683), .B1(net_19682), .ZN(net_16312) );
INV_X4 inst_13482 ( .ZN(net_9564), .A(net_9563) );
XNOR2_X2 inst_193 ( .ZN(net_17678), .A(net_17336), .B(net_324) );
INV_X4 inst_14568 ( .ZN(net_5824), .A(net_4555) );
INV_X4 inst_16153 ( .ZN(net_2981), .A(net_1263) );
CLKBUF_X2 inst_22637 ( .A(net_22508), .Z(net_22509) );
INV_X4 inst_17541 ( .ZN(net_6606), .A(net_381) );
NAND2_X2 inst_11704 ( .ZN(net_2932), .A1(net_2300), .A2(net_1142) );
CLKBUF_X2 inst_21543 ( .A(net_21414), .Z(net_21415) );
OAI21_X2 inst_1709 ( .ZN(net_19231), .A(net_14203), .B2(net_13981), .B1(net_6628) );
INV_X16 inst_19732 ( .A(net_1630), .ZN(net_1442) );
INV_X4 inst_16583 ( .ZN(net_1427), .A(net_1418) );
INV_X4 inst_15358 ( .A(net_5852), .ZN(net_3422) );
AOI21_X2 inst_20664 ( .A(net_15186), .ZN(net_12924), .B2(net_12923), .B1(net_12035) );
INV_X4 inst_17600 ( .A(net_20868), .ZN(net_663) );
NAND2_X4 inst_7531 ( .ZN(net_1957), .A1(net_1956), .A2(net_1803) );
OAI21_X2 inst_2202 ( .ZN(net_20600), .B1(net_8553), .B2(net_6998), .A(net_6867) );
CLKBUF_X2 inst_22781 ( .A(net_22652), .Z(net_22653) );
CLKBUF_X2 inst_21485 ( .A(net_21356), .Z(net_21357) );
NAND2_X2 inst_11673 ( .ZN(net_5623), .A1(net_4253), .A2(net_2358) );
INV_X2 inst_19218 ( .ZN(net_19646), .A(net_3473) );
NOR2_X4 inst_3180 ( .A1(net_20868), .ZN(net_3132), .A2(net_3131) );
NAND2_X2 inst_7969 ( .ZN(net_18362), .A2(net_18248), .A1(net_17301) );
AND4_X4 inst_21086 ( .ZN(net_16482), .A4(net_16179), .A2(net_15909), .A1(net_15536), .A3(net_14822) );
NOR2_X2 inst_4737 ( .ZN(net_3922), .A2(net_3075), .A1(net_3063) );
NAND2_X2 inst_9965 ( .A1(net_12295), .ZN(net_8897), .A2(net_8896) );
NOR2_X4 inst_2987 ( .ZN(net_7507), .A2(net_6078), .A1(net_6077) );
NAND2_X2 inst_10618 ( .A2(net_20782), .ZN(net_12177), .A1(net_6586) );
INV_X4 inst_15162 ( .ZN(net_5165), .A(net_3024) );
NAND2_X2 inst_11645 ( .ZN(net_5621), .A1(net_3915), .A2(net_1142) );
INV_X2 inst_19303 ( .ZN(net_2764), .A(net_2763) );
NAND3_X2 inst_5884 ( .ZN(net_15242), .A3(net_14172), .A2(net_13531), .A1(net_12913) );
NAND2_X2 inst_11853 ( .ZN(net_3253), .A1(net_1655), .A2(net_1389) );
CLKBUF_X2 inst_21595 ( .A(net_21466), .Z(net_21467) );
NAND2_X2 inst_11170 ( .ZN(net_7052), .A1(net_4340), .A2(net_2239) );
CLKBUF_X2 inst_22153 ( .A(net_22024), .Z(net_22025) );
CLKBUF_X2 inst_22002 ( .A(net_21873), .Z(net_21874) );
INV_X4 inst_12874 ( .ZN(net_16947), .A(net_16946) );
INV_X2 inst_19311 ( .ZN(net_2706), .A(net_2705) );
OAI211_X2 inst_2473 ( .ZN(net_13662), .A(net_11244), .B(net_10902), .C1(net_9502), .C2(net_3178) );
NAND2_X4 inst_7125 ( .ZN(net_12665), .A2(net_10903), .A1(net_9925) );
INV_X4 inst_17361 ( .ZN(net_2202), .A(net_149) );
NOR2_X2 inst_4516 ( .A1(net_10962), .ZN(net_5221), .A2(net_4908) );
INV_X8 inst_12442 ( .A(net_20940), .ZN(net_20495) );
INV_X4 inst_13952 ( .ZN(net_8681), .A(net_6765) );
CLKBUF_X2 inst_21707 ( .A(net_21396), .Z(net_21579) );
NOR2_X4 inst_2864 ( .ZN(net_20028), .A1(net_7467), .A2(net_3298) );
NOR2_X2 inst_3476 ( .ZN(net_14445), .A1(net_14444), .A2(net_13037) );
INV_X4 inst_14645 ( .ZN(net_4637), .A(net_4373) );
NOR2_X2 inst_3789 ( .ZN(net_19171), .A2(net_6337), .A1(net_5416) );
INV_X4 inst_15001 ( .A(net_14605), .ZN(net_11645) );
NAND2_X4 inst_7096 ( .ZN(net_18883), .A1(net_13064), .A2(net_8718) );
INV_X4 inst_16127 ( .ZN(net_1482), .A(net_1481) );
XNOR2_X2 inst_367 ( .ZN(net_16850), .A(net_16846), .B(net_7648) );
SDFF_X2 inst_957 ( .QN(net_21058), .D(net_477), .SE(net_253), .CK(net_21734), .SI(x2087) );
NAND2_X2 inst_11589 ( .A1(net_2727), .ZN(net_2695), .A2(net_2694) );
DFF_X1 inst_19816 ( .D(net_17833), .CK(net_22812), .Q(x1283) );
OAI21_X2 inst_1871 ( .ZN(net_13710), .A(net_13709), .B2(net_11737), .B1(net_11072) );
INV_X2 inst_19451 ( .ZN(net_2988), .A(net_2293) );
INV_X4 inst_16653 ( .ZN(net_2164), .A(net_1092) );
NAND3_X2 inst_6460 ( .ZN(net_11392), .A2(net_11391), .A3(net_11347), .A1(net_11251) );
OAI21_X2 inst_2300 ( .ZN(net_6416), .A(net_6415), .B1(net_6379), .B2(net_4092) );
NAND2_X4 inst_7552 ( .A1(net_3456), .ZN(net_2017), .A2(net_1764) );
NAND2_X2 inst_10800 ( .ZN(net_5561), .A2(net_5560), .A1(net_154) );
CLKBUF_X2 inst_22240 ( .A(net_22111), .Z(net_22112) );
INV_X2 inst_18666 ( .A(net_11021), .ZN(net_9176) );
SDFF_X2 inst_745 ( .Q(net_20961), .SE(net_18804), .SI(net_18548), .D(net_534), .CK(net_22181) );
NAND2_X2 inst_11694 ( .A2(net_2683), .ZN(net_2320), .A1(net_2319) );
NAND2_X4 inst_7024 ( .ZN(net_17353), .A1(net_16557), .A2(net_16448) );
AOI21_X2 inst_20556 ( .ZN(net_14281), .B1(net_13984), .B2(net_13589), .A(net_8302) );
NAND2_X2 inst_11622 ( .ZN(net_5044), .A1(net_2013), .A2(net_1360) );
CLKBUF_X2 inst_22840 ( .A(net_21415), .Z(net_22712) );
CLKBUF_X2 inst_22487 ( .A(net_22358), .Z(net_22359) );
OAI21_X2 inst_2032 ( .ZN(net_11310), .B2(net_9774), .B1(net_9673), .A(net_2574) );
NOR2_X2 inst_4113 ( .ZN(net_7066), .A1(net_7065), .A2(net_4148) );
XNOR2_X2 inst_80 ( .B(net_21163), .ZN(net_18660), .A(net_18610) );
NAND2_X4 inst_7698 ( .ZN(net_503), .A2(net_220), .A1(net_118) );
SDFF_X2 inst_836 ( .Q(net_21238), .SI(net_17503), .SE(net_125), .CK(net_21559), .D(x6740) );
NAND2_X2 inst_8821 ( .ZN(net_15560), .A2(net_14832), .A1(net_11847) );
NAND2_X2 inst_9521 ( .ZN(net_11139), .A2(net_11138), .A1(net_7638) );
NAND3_X2 inst_6564 ( .A3(net_19753), .ZN(net_10482), .A2(net_8162), .A1(net_6779) );
NAND2_X2 inst_10771 ( .A1(net_14865), .ZN(net_6723), .A2(net_5629) );
NAND2_X2 inst_9562 ( .ZN(net_12374), .A1(net_11020), .A2(net_6999) );
CLKBUF_X2 inst_22255 ( .A(net_22091), .Z(net_22127) );
XNOR2_X2 inst_241 ( .B(net_21181), .ZN(net_17379), .A(net_17378) );
AOI21_X2 inst_20641 ( .ZN(net_13230), .B1(net_10937), .B2(net_10041), .A(net_7598) );
NOR2_X2 inst_5120 ( .A2(net_513), .ZN(net_298), .A1(net_108) );
NOR2_X2 inst_4409 ( .ZN(net_6218), .A1(net_4840), .A2(net_2807) );
DFF_X2 inst_19776 ( .D(net_5773), .Q(net_28), .CK(net_22272) );
INV_X4 inst_16957 ( .ZN(net_7850), .A(net_388) );
NOR2_X2 inst_4934 ( .ZN(net_2479), .A2(net_1741), .A1(net_123) );
INV_X4 inst_14705 ( .ZN(net_5174), .A(net_3145) );
INV_X4 inst_16356 ( .ZN(net_8961), .A(net_8376) );
INV_X4 inst_15384 ( .ZN(net_3365), .A(net_2723) );
NAND3_X2 inst_6690 ( .ZN(net_7706), .A3(net_7705), .A1(net_4656), .A2(net_3017) );
AOI21_X2 inst_20669 ( .B1(net_13070), .ZN(net_12894), .A(net_11266), .B2(net_8688) );
NOR2_X2 inst_3918 ( .ZN(net_10288), .A1(net_8800), .A2(net_8192) );
INV_X4 inst_13491 ( .A(net_11717), .ZN(net_9484) );
INV_X4 inst_14142 ( .ZN(net_8475), .A(net_6068) );
INV_X4 inst_15534 ( .A(net_9183), .ZN(net_7872) );
NOR3_X2 inst_2758 ( .ZN(net_11222), .A2(net_11221), .A3(net_11220), .A1(net_7792) );
NOR2_X2 inst_4504 ( .A1(net_12004), .ZN(net_4243), .A2(net_2983) );
OR2_X4 inst_1116 ( .ZN(net_10886), .A2(net_955), .A1(net_115) );
NAND2_X2 inst_7947 ( .ZN(net_18407), .A2(net_18342), .A1(net_18337) );
INV_X4 inst_18311 ( .ZN(net_20506), .A(net_20504) );
NOR2_X2 inst_3753 ( .ZN(net_10394), .A1(net_10393), .A2(net_6652) );
NAND3_X4 inst_5545 ( .ZN(net_17006), .A3(net_16364), .A1(net_16320), .A2(net_15682) );
NAND2_X2 inst_12050 ( .ZN(net_929), .A2(net_928), .A1(net_459) );
CLKBUF_X2 inst_22279 ( .A(net_22150), .Z(net_22151) );
AOI21_X2 inst_20628 ( .ZN(net_13430), .B1(net_10216), .A(net_10084), .B2(net_9047) );
INV_X4 inst_16393 ( .ZN(net_1831), .A(net_864) );
INV_X4 inst_17858 ( .ZN(net_889), .A(net_108) );
NAND2_X2 inst_11555 ( .ZN(net_3721), .A1(net_2841), .A2(net_2840) );
INV_X4 inst_17363 ( .ZN(net_7465), .A(net_761) );
NAND3_X2 inst_6394 ( .ZN(net_12002), .A2(net_11717), .A1(net_7447), .A3(net_6709) );
NOR2_X4 inst_3136 ( .A2(net_20568), .ZN(net_6662), .A1(net_3797) );
XNOR2_X2 inst_402 ( .A(net_19432), .ZN(net_16679), .B(net_11888) );
NAND2_X2 inst_10962 ( .A1(net_9785), .ZN(net_8228), .A2(net_4641) );
INV_X4 inst_16084 ( .A(net_5479), .ZN(net_1927) );
CLKBUF_X2 inst_22039 ( .A(net_21288), .Z(net_21911) );
NAND2_X2 inst_11259 ( .ZN(net_11240), .A1(net_4305), .A2(net_3911) );
INV_X4 inst_13025 ( .A(net_16476), .ZN(net_16441) );
NAND3_X2 inst_5832 ( .A3(net_18874), .ZN(net_15515), .A1(net_14131), .A2(net_13518) );
INV_X4 inst_12815 ( .ZN(net_17300), .A(net_17198) );
NAND2_X4 inst_7350 ( .ZN(net_7877), .A1(net_4821), .A2(net_3505) );
OAI22_X2 inst_1288 ( .ZN(net_12886), .A1(net_12885), .B1(net_12884), .B2(net_12883), .A2(net_12844) );
NOR2_X2 inst_3844 ( .ZN(net_11571), .A2(net_9586), .A1(net_6702) );
INV_X2 inst_19128 ( .ZN(net_4283), .A(net_4282) );
NAND2_X4 inst_7610 ( .ZN(net_2462), .A2(net_200), .A1(net_63) );
NAND2_X2 inst_11329 ( .ZN(net_6122), .A2(net_3736), .A1(net_2171) );
SDFF_X2 inst_1033 ( .QN(net_21053), .D(net_616), .SE(net_263), .CK(net_22495), .SI(x2149) );
NAND2_X2 inst_11845 ( .ZN(net_2492), .A2(net_2384), .A1(net_367) );
NOR2_X2 inst_4673 ( .A1(net_3458), .ZN(net_3243), .A2(net_2167) );
AOI21_X2 inst_20732 ( .ZN(net_11742), .B2(net_11741), .B1(net_11572), .A(net_6117) );
INV_X4 inst_14201 ( .ZN(net_5955), .A(net_5954) );
CLKBUF_X2 inst_21520 ( .A(net_21379), .Z(net_21392) );
INV_X2 inst_19081 ( .ZN(net_4587), .A(net_4586) );
INV_X4 inst_16138 ( .ZN(net_1473), .A(net_1472) );
NAND3_X4 inst_5582 ( .A2(net_19813), .A1(net_19812), .ZN(net_15530), .A3(net_14719) );
OAI221_X2 inst_1348 ( .ZN(net_12239), .B1(net_12238), .C1(net_10947), .A(net_10126), .B2(net_7026), .C2(net_4363) );
NAND4_X2 inst_5427 ( .A3(net_20029), .A1(net_20028), .ZN(net_19389), .A2(net_10314), .A4(net_10017) );
OAI21_X2 inst_1748 ( .ZN(net_14941), .A(net_14820), .B2(net_12683), .B1(net_9143) );
INV_X4 inst_15686 ( .ZN(net_2905), .A(net_1649) );
NAND2_X4 inst_7356 ( .ZN(net_8393), .A1(net_3489), .A2(net_2274) );
NAND2_X2 inst_11423 ( .A1(net_7917), .ZN(net_3363), .A2(net_3362) );
DFF_X1 inst_19879 ( .D(net_17128), .CK(net_22538), .Q(x23) );
CLKBUF_X2 inst_21968 ( .A(net_21397), .Z(net_21840) );
NAND3_X4 inst_5565 ( .ZN(net_15986), .A3(net_15619), .A1(net_14842), .A2(net_14727) );
NAND2_X2 inst_11684 ( .ZN(net_13002), .A1(net_4286), .A2(net_2340) );
INV_X4 inst_14781 ( .ZN(net_14141), .A(net_4034) );
NAND2_X2 inst_11864 ( .A1(net_2919), .A2(net_2190), .ZN(net_1654) );
NAND2_X2 inst_8637 ( .A1(net_20527), .A2(net_16612), .ZN(net_16582) );
NAND2_X2 inst_9712 ( .ZN(net_10177), .A1(net_7618), .A2(net_6766) );
NAND2_X2 inst_10145 ( .ZN(net_20742), .A1(net_11182), .A2(net_6202) );
INV_X4 inst_14058 ( .ZN(net_9640), .A(net_6248) );
INV_X4 inst_18211 ( .A(net_21204), .ZN(net_17262) );
NAND2_X2 inst_9216 ( .ZN(net_12998), .A2(net_11385), .A1(net_6839) );
INV_X4 inst_16439 ( .ZN(net_1780), .A(net_63) );
INV_X2 inst_19004 ( .ZN(net_7930), .A(net_6730) );
NAND2_X2 inst_11088 ( .ZN(net_4912), .A2(net_4315), .A1(net_70) );
AOI22_X2 inst_20032 ( .ZN(net_8960), .A1(net_8959), .B2(net_8958), .A2(net_5408), .B1(net_4151) );
AOI21_X4 inst_20095 ( .ZN(net_18915), .B2(net_18601), .A(net_18594), .B1(net_16302) );
NAND2_X2 inst_12046 ( .ZN(net_1081), .A1(net_938), .A2(net_258) );
NAND3_X2 inst_6397 ( .ZN(net_11993), .A3(net_11924), .A2(net_5898), .A1(net_3358) );
NAND2_X4 inst_7337 ( .ZN(net_6049), .A1(net_4902), .A2(net_3865) );
OAI211_X2 inst_2461 ( .B(net_14337), .ZN(net_14150), .C2(net_9207), .C1(net_5282), .A(net_4905) );
INV_X2 inst_18420 ( .ZN(net_15623), .A(net_15384) );
AOI21_X2 inst_20934 ( .B1(net_7121), .ZN(net_6542), .B2(net_6541), .A(net_5184) );
NAND2_X2 inst_8814 ( .ZN(net_19596), .A2(net_14887), .A1(net_12357) );
SDFF_X2 inst_732 ( .Q(net_20941), .SE(net_18862), .SI(net_18563), .D(net_6549), .CK(net_22758) );
INV_X8 inst_12183 ( .ZN(net_17244), .A(net_16656) );
INV_X4 inst_13044 ( .ZN(net_18954), .A(net_16373) );
NAND2_X2 inst_8023 ( .A2(net_18280), .ZN(net_18275), .A1(net_17630) );
NAND3_X2 inst_5968 ( .ZN(net_14775), .A3(net_13417), .A2(net_12301), .A1(net_11639) );
XNOR2_X2 inst_79 ( .ZN(net_18664), .A(net_18614), .B(net_17777) );
NAND2_X2 inst_11250 ( .ZN(net_8467), .A2(net_5284), .A1(net_2709) );
NAND2_X2 inst_8930 ( .ZN(net_20354), .A1(net_15742), .A2(net_13602) );
NOR3_X2 inst_2654 ( .ZN(net_15474), .A3(net_14534), .A2(net_10148), .A1(net_5152) );
NAND2_X4 inst_7088 ( .ZN(net_19357), .A2(net_14487), .A1(net_14249) );
INV_X4 inst_16526 ( .ZN(net_9366), .A(net_4799) );
INV_X4 inst_16691 ( .ZN(net_13999), .A(net_8260) );
CLKBUF_X2 inst_22409 ( .A(net_22280), .Z(net_22281) );
CLKBUF_X2 inst_22499 ( .A(net_22370), .Z(net_22371) );
NAND2_X2 inst_11662 ( .A1(net_4711), .ZN(net_4345), .A2(net_2412) );
CLKBUF_X2 inst_21986 ( .A(net_21408), .Z(net_21858) );
NAND2_X2 inst_8838 ( .ZN(net_15473), .A2(net_14850), .A1(net_12154) );
NAND2_X2 inst_11962 ( .A2(net_20480), .ZN(net_1383), .A1(net_294) );
NAND2_X2 inst_7895 ( .ZN(net_18489), .A2(net_18446), .A1(net_17951) );
NOR2_X2 inst_4413 ( .A1(net_5157), .ZN(net_5045), .A2(net_5044) );
INV_X4 inst_16293 ( .ZN(net_10225), .A(net_761) );
CLKBUF_X2 inst_21749 ( .A(net_21525), .Z(net_21621) );
INV_X4 inst_17938 ( .A(net_21221), .ZN(net_130) );
NOR2_X4 inst_2975 ( .A2(net_8369), .ZN(net_7591), .A1(net_3970) );
OAI21_X2 inst_1741 ( .ZN(net_15028), .A(net_15027), .B2(net_12749), .B1(net_9264) );
NAND3_X4 inst_5594 ( .ZN(net_15011), .A2(net_12687), .A3(net_11769), .A1(net_5592) );
OAI21_X2 inst_1658 ( .ZN(net_15787), .B2(net_14781), .B1(net_6296), .A(net_1774) );
NAND3_X2 inst_6515 ( .A3(net_11915), .ZN(net_10653), .A1(net_10609), .A2(net_3995) );
INV_X4 inst_14991 ( .A(net_15974), .ZN(net_13827) );
NAND2_X2 inst_9003 ( .ZN(net_14283), .A2(net_13595), .A1(net_11345) );
NOR2_X2 inst_4267 ( .ZN(net_6167), .A2(net_6166), .A1(net_3759) );
NOR2_X2 inst_3965 ( .ZN(net_8420), .A1(net_7059), .A2(net_4731) );
INV_X2 inst_19291 ( .ZN(net_2865), .A(net_2864) );
CLKBUF_X2 inst_22494 ( .A(net_22365), .Z(net_22366) );
INV_X4 inst_12829 ( .ZN(net_20633), .A(net_17141) );
XNOR2_X2 inst_440 ( .A(net_21207), .B(net_16857), .ZN(net_16090) );
DFF_X1 inst_19872 ( .D(net_17030), .CK(net_22356), .Q(x745) );
INV_X2 inst_18963 ( .ZN(net_5408), .A(net_5407) );
INV_X4 inst_14386 ( .ZN(net_8191), .A(net_5147) );
DFF_X2 inst_19783 ( .D(net_14378), .QN(net_29), .CK(net_22186) );
AND3_X4 inst_21128 ( .A1(net_11426), .A2(net_8700), .ZN(net_7186), .A3(net_5780) );
NOR2_X2 inst_4927 ( .A1(net_20495), .ZN(net_2926), .A2(net_1785) );
OAI21_X2 inst_1887 ( .ZN(net_13503), .A(net_10659), .B2(net_9074), .B1(net_7017) );
INV_X4 inst_15287 ( .ZN(net_9282), .A(net_2777) );
INV_X4 inst_15423 ( .ZN(net_3299), .A(net_3111) );
NAND2_X2 inst_11708 ( .ZN(net_12887), .A1(net_8462), .A2(net_1223) );
INV_X4 inst_15108 ( .ZN(net_3840), .A(net_3210) );
AOI21_X4 inst_20189 ( .B1(net_19298), .ZN(net_19050), .A(net_10680), .B2(net_816) );
NOR2_X2 inst_3579 ( .A1(net_14357), .ZN(net_12688), .A2(net_12386) );
INV_X2 inst_19537 ( .A(net_2244), .ZN(net_969) );
INV_X4 inst_16560 ( .A(net_13343), .ZN(net_8889) );
INV_X4 inst_16537 ( .ZN(net_1819), .A(net_1075) );
NAND3_X2 inst_5688 ( .ZN(net_16295), .A1(net_16024), .A3(net_16017), .A2(net_15639) );
CLKBUF_X2 inst_22297 ( .A(net_22168), .Z(net_22169) );
OAI21_X2 inst_1672 ( .ZN(net_15601), .B1(net_15542), .B2(net_14259), .A(net_5324) );
INV_X4 inst_16921 ( .ZN(net_5766), .A(net_624) );
INV_X4 inst_13705 ( .ZN(net_9407), .A(net_7869) );
NAND2_X2 inst_8625 ( .ZN(net_16600), .A1(net_16599), .A2(net_16577) );
NAND2_X2 inst_12120 ( .A2(net_20538), .ZN(net_1369), .A1(net_146) );
INV_X4 inst_17661 ( .ZN(net_895), .A(net_257) );
OAI21_X2 inst_2015 ( .ZN(net_11375), .A(net_11374), .B1(net_10587), .B2(net_5855) );
INV_X4 inst_18110 ( .A(net_20862), .ZN(net_64) );
NAND2_X2 inst_12108 ( .ZN(net_335), .A2(net_272), .A1(net_64) );
AOI21_X2 inst_20433 ( .ZN(net_15171), .B1(net_14643), .B2(net_13893), .A(net_7983) );
NOR2_X2 inst_3937 ( .ZN(net_13184), .A2(net_8942), .A1(net_8674) );
NOR2_X4 inst_2970 ( .ZN(net_7643), .A1(net_5322), .A2(net_4917) );
INV_X4 inst_14488 ( .ZN(net_6014), .A(net_4851) );
NAND2_X2 inst_11950 ( .A1(net_1823), .ZN(net_1419), .A2(net_1418) );
DFF_X2 inst_19777 ( .QN(net_21107), .D(net_5717), .CK(net_22461) );
NAND2_X2 inst_10942 ( .ZN(net_6821), .A2(net_5575), .A1(net_5157) );
CLKBUF_X2 inst_21733 ( .A(net_21604), .Z(net_21605) );
NAND2_X2 inst_8278 ( .A2(net_19932), .A1(net_19931), .ZN(net_17631) );
NAND2_X2 inst_9281 ( .ZN(net_12585), .A2(net_9507), .A1(net_6955) );
NOR2_X2 inst_4085 ( .ZN(net_13186), .A2(net_10306), .A1(net_5186) );
INV_X4 inst_16360 ( .ZN(net_4401), .A(net_143) );
CLKBUF_X2 inst_22178 ( .A(net_22049), .Z(net_22050) );
INV_X2 inst_18576 ( .ZN(net_10487), .A(net_8974) );
INV_X4 inst_14719 ( .ZN(net_8939), .A(net_8581) );
INV_X4 inst_18194 ( .A(net_20956), .ZN(net_252) );
INV_X4 inst_17058 ( .ZN(net_6924), .A(net_5450) );
INV_X4 inst_13183 ( .ZN(net_14259), .A(net_13706) );
NOR2_X2 inst_4990 ( .A1(net_20495), .ZN(net_1417), .A2(net_1168) );
NAND3_X2 inst_5664 ( .ZN(net_16400), .A3(net_16258), .A2(net_15544), .A1(net_10809) );
NAND2_X2 inst_10317 ( .ZN(net_12225), .A2(net_5353), .A1(net_1067) );
INV_X8 inst_12285 ( .ZN(net_2139), .A(net_753) );
CLKBUF_X2 inst_22389 ( .A(net_22260), .Z(net_22261) );
NAND2_X2 inst_9442 ( .ZN(net_18981), .A1(net_11553), .A2(net_11552) );
NAND2_X2 inst_11090 ( .ZN(net_6430), .A2(net_3771), .A1(net_3148) );
AOI21_X2 inst_20484 ( .ZN(net_14836), .B2(net_13466), .B1(net_12595), .A(net_10683) );
SDFF_X2 inst_815 ( .Q(net_21129), .SI(net_17773), .SE(net_125), .CK(net_21416), .D(x4041) );
AND2_X4 inst_21178 ( .A1(net_11644), .ZN(net_11636), .A2(net_11635) );
OAI21_X2 inst_2165 ( .A(net_12133), .ZN(net_9026), .B2(net_7235), .B1(net_5684) );
INV_X4 inst_15433 ( .ZN(net_10389), .A(net_9023) );
NOR2_X4 inst_3081 ( .ZN(net_7729), .A1(net_4409), .A2(net_131) );
AOI21_X2 inst_20605 ( .ZN(net_13756), .B2(net_11101), .B1(net_2620), .A(net_1998) );
NAND4_X4 inst_5187 ( .A4(net_18942), .A1(net_18941), .ZN(net_17526), .A2(net_16343), .A3(net_14255) );
NAND2_X2 inst_12096 ( .A2(net_20851), .ZN(net_554), .A1(net_214) );
INV_X2 inst_19376 ( .A(net_2189), .ZN(net_2169) );
NAND2_X2 inst_8227 ( .A2(net_17797), .ZN(net_17795), .A1(net_17200) );
INV_X4 inst_16330 ( .ZN(net_1768), .A(net_1308) );
NAND2_X4 inst_7006 ( .ZN(net_20097), .A2(net_19459), .A1(net_16969) );
NAND2_X2 inst_8888 ( .ZN(net_15142), .A2(net_14094), .A1(net_11668) );
AOI21_X2 inst_20579 ( .ZN(net_14100), .B1(net_11451), .B2(net_10651), .A(net_10388) );
OAI21_X2 inst_2108 ( .ZN(net_19951), .B1(net_10046), .A(net_7252), .B2(net_4667) );
NOR2_X2 inst_3572 ( .ZN(net_12723), .A2(net_10935), .A1(net_7015) );
NAND2_X2 inst_7761 ( .ZN(net_18755), .A2(net_18705), .A1(net_18685) );
INV_X8 inst_12178 ( .ZN(net_17363), .A(net_17236) );
NAND2_X2 inst_11177 ( .A1(net_5244), .ZN(net_5206), .A2(net_4138) );
XNOR2_X2 inst_413 ( .A(net_16569), .ZN(net_16547), .B(net_11884) );
NOR2_X2 inst_5094 ( .ZN(net_2096), .A1(net_809), .A2(net_85) );
CLKBUF_X2 inst_21563 ( .A(net_21335), .Z(net_21435) );
NAND2_X2 inst_8118 ( .A2(net_18089), .ZN(net_18088), .A1(net_17371) );
NAND3_X2 inst_6623 ( .A3(net_19305), .ZN(net_9050), .A1(net_6758), .A2(net_4776) );
SDFF_X2 inst_859 ( .Q(net_21172), .SI(net_17173), .SE(net_125), .CK(net_22155), .D(x4815) );
INV_X4 inst_13446 ( .ZN(net_11108), .A(net_8305) );
NOR2_X4 inst_3323 ( .A2(net_20901), .ZN(net_1644), .A1(net_163) );
INV_X4 inst_12634 ( .ZN(net_18687), .A(net_17919) );
CLKBUF_X2 inst_21870 ( .A(net_21337), .Z(net_21742) );
INV_X4 inst_17448 ( .A(net_2224), .ZN(net_922) );
INV_X4 inst_13013 ( .ZN(net_16874), .A(net_16762) );
INV_X2 inst_18391 ( .ZN(net_16629), .A(net_16628) );
INV_X2 inst_19394 ( .ZN(net_19529), .A(net_2026) );
CLKBUF_X2 inst_21411 ( .A(net_21272), .Z(net_21283) );
NAND3_X2 inst_5938 ( .ZN(net_14919), .A1(net_13625), .A2(net_10774), .A3(net_9075) );
AOI21_X2 inst_20722 ( .ZN(net_11978), .A(net_10006), .B2(net_7715), .B1(net_3802) );
INV_X4 inst_13061 ( .ZN(net_16352), .A(net_16300) );
NAND3_X2 inst_5736 ( .ZN(net_19363), .A3(net_19304), .A1(net_19303), .A2(net_11232) );
OAI21_X2 inst_1691 ( .B2(net_20383), .B1(net_20382), .ZN(net_15365), .A(net_15301) );
INV_X4 inst_15626 ( .ZN(net_4203), .A(net_2149) );
AOI21_X2 inst_20752 ( .ZN(net_11349), .B1(net_11348), .B2(net_11347), .A(net_11148) );
NAND2_X2 inst_9019 ( .A1(net_15833), .ZN(net_14173), .A2(net_12244) );
NAND2_X2 inst_11156 ( .A1(net_9418), .ZN(net_4195), .A2(net_3302) );
CLKBUF_X2 inst_21479 ( .A(net_21324), .Z(net_21351) );
AOI21_X2 inst_20378 ( .ZN(net_15562), .B1(net_15561), .B2(net_14435), .A(net_6657) );
AOI21_X2 inst_20675 ( .ZN(net_12531), .B2(net_12530), .A(net_11207), .B1(net_81) );
INV_X4 inst_15413 ( .ZN(net_15166), .A(net_14009) );
NOR2_X2 inst_3688 ( .ZN(net_11412), .A1(net_9570), .A2(net_9287) );
NAND2_X2 inst_7716 ( .ZN(net_18846), .A1(net_18812), .A2(net_18795) );
NAND4_X2 inst_5476 ( .A3(net_12968), .ZN(net_12905), .A2(net_11895), .A4(net_5178), .A1(net_3425) );
AND3_X2 inst_21134 ( .A3(net_13941), .ZN(net_13262), .A2(net_12762), .A1(net_10516) );
NAND3_X2 inst_5776 ( .ZN(net_15872), .A3(net_15365), .A2(net_14729), .A1(net_13711) );
INV_X2 inst_18863 ( .ZN(net_6293), .A(net_6292) );
NAND2_X1 inst_12149 ( .A2(net_17767), .ZN(net_16432), .A1(net_6548) );
CLKBUF_X2 inst_22109 ( .A(net_21980), .Z(net_21981) );
NAND2_X2 inst_10186 ( .ZN(net_8178), .A1(net_7822), .A2(net_7057) );
INV_X4 inst_13124 ( .ZN(net_15403), .A(net_15146) );
XNOR2_X2 inst_560 ( .B(net_17534), .ZN(net_682), .A(net_681) );
NAND2_X2 inst_11167 ( .A1(net_11062), .ZN(net_4173), .A2(net_4172) );
NAND4_X2 inst_5393 ( .ZN(net_14827), .A4(net_13365), .A3(net_11778), .A1(net_9786), .A2(net_9059) );
NAND4_X4 inst_5199 ( .A4(net_19146), .A1(net_19145), .ZN(net_16780), .A3(net_13374), .A2(net_12178) );
NAND2_X2 inst_9729 ( .A1(net_12330), .ZN(net_10118), .A2(net_8000) );
INV_X4 inst_12953 ( .ZN(net_16901), .A(net_16732) );
NAND2_X4 inst_7479 ( .ZN(net_4991), .A1(net_1764), .A2(net_1446) );
NOR2_X2 inst_4809 ( .ZN(net_10459), .A1(net_2646), .A2(net_2645) );
OAI21_X2 inst_1802 ( .ZN(net_14479), .B1(net_12461), .B2(net_11438), .A(net_652) );
CLKBUF_X2 inst_21390 ( .A(net_21261), .Z(net_21262) );
NAND2_X2 inst_10260 ( .ZN(net_10265), .A2(net_3421), .A1(net_1076) );
NAND2_X4 inst_6851 ( .A2(net_20721), .A1(net_20720), .ZN(net_18500) );
NOR2_X4 inst_2982 ( .ZN(net_9699), .A2(net_3970), .A1(net_1931) );
INV_X4 inst_15444 ( .ZN(net_3509), .A(net_2499) );
NAND2_X2 inst_11837 ( .A1(net_20851), .ZN(net_2386), .A2(net_1625) );
NOR2_X2 inst_3359 ( .A2(net_20207), .ZN(net_17486), .A1(net_17485) );
NAND2_X2 inst_10100 ( .ZN(net_20360), .A1(net_10216), .A2(net_7030) );
CLKBUF_X2 inst_22290 ( .A(net_21697), .Z(net_22162) );
INV_X2 inst_18974 ( .ZN(net_5213), .A(net_5212) );
NAND2_X4 inst_7491 ( .ZN(net_2699), .A2(net_2402), .A1(net_1269) );
INV_X4 inst_14338 ( .ZN(net_5382), .A(net_5381) );
NOR2_X2 inst_4418 ( .ZN(net_4996), .A1(net_4995), .A2(net_3596) );
XNOR2_X2 inst_96 ( .ZN(net_18548), .A(net_18445), .B(net_17379) );
NOR2_X2 inst_4346 ( .ZN(net_20756), .A1(net_5637), .A2(net_3362) );
NAND2_X2 inst_8564 ( .A1(net_21180), .ZN(net_16745), .A2(net_16576) );
INV_X2 inst_18705 ( .ZN(net_8259), .A(net_8258) );
INV_X4 inst_17156 ( .ZN(net_1246), .A(net_857) );
NAND2_X2 inst_11205 ( .ZN(net_4043), .A1(net_4042), .A2(net_3924) );
NAND2_X2 inst_9330 ( .ZN(net_14210), .A1(net_10815), .A2(net_9139) );
INV_X2 inst_19388 ( .A(net_3177), .ZN(net_2088) );
INV_X2 inst_18687 ( .ZN(net_8662), .A(net_8661) );
INV_X4 inst_17616 ( .A(net_20875), .ZN(net_381) );
NAND2_X2 inst_10912 ( .A1(net_12100), .ZN(net_5354), .A2(net_5353) );
INV_X4 inst_15558 ( .ZN(net_7147), .A(net_2068) );
INV_X4 inst_14575 ( .ZN(net_7454), .A(net_4537) );
INV_X4 inst_15937 ( .ZN(net_2917), .A(net_1723) );
OAI211_X2 inst_2436 ( .ZN(net_15004), .C2(net_13747), .B(net_12778), .C1(net_10011), .A(net_9906) );
INV_X16 inst_19736 ( .ZN(net_1981), .A(net_412) );
NOR2_X4 inst_2832 ( .A2(net_19938), .A1(net_19937), .ZN(net_19550) );
INV_X2 inst_19168 ( .ZN(net_13201), .A(net_5423) );
CLKBUF_X2 inst_22703 ( .A(net_22574), .Z(net_22575) );
XNOR2_X2 inst_603 ( .B(net_17253), .ZN(net_531), .A(net_530) );
XNOR2_X2 inst_291 ( .B(net_21168), .ZN(net_17134), .A(net_16974) );
CLKBUF_X2 inst_22148 ( .A(net_21285), .Z(net_22020) );
NAND2_X2 inst_9488 ( .A1(net_13375), .ZN(net_11445), .A2(net_11444) );
AND2_X4 inst_21185 ( .A2(net_12804), .ZN(net_11447), .A1(net_11446) );
INV_X4 inst_15521 ( .ZN(net_2737), .A(net_2399) );
INV_X8 inst_12213 ( .ZN(net_9618), .A(net_6233) );
INV_X4 inst_16569 ( .ZN(net_2060), .A(net_606) );
AND2_X2 inst_21347 ( .A2(net_2891), .ZN(net_2662), .A1(net_1901) );
AND4_X2 inst_21102 ( .ZN(net_12465), .A4(net_12025), .A3(net_10580), .A2(net_10208), .A1(net_3221) );
INV_X2 inst_18709 ( .A(net_8655), .ZN(net_8239) );
INV_X4 inst_16846 ( .ZN(net_14769), .A(net_1030) );
INV_X4 inst_16688 ( .A(net_3900), .ZN(net_3812) );
NAND2_X4 inst_6849 ( .A2(net_20936), .ZN(net_18591), .A1(net_15769) );
NAND2_X2 inst_10310 ( .ZN(net_9383), .A2(net_7851), .A1(net_7850) );
NAND2_X2 inst_9110 ( .ZN(net_14858), .A1(net_14264), .A2(net_12410) );
NAND3_X2 inst_6512 ( .A3(net_12902), .ZN(net_10755), .A2(net_10754), .A1(net_3726) );
NAND2_X4 inst_6925 ( .A2(net_19048), .A1(net_19047), .ZN(net_17744) );
NAND2_X2 inst_7745 ( .ZN(net_18792), .A2(net_18761), .A1(net_17564) );
INV_X2 inst_19239 ( .ZN(net_3313), .A(net_3312) );
AOI21_X2 inst_20976 ( .A(net_20486), .ZN(net_4217), .B2(net_4216), .B1(net_3543) );
OAI21_X2 inst_1807 ( .ZN(net_14469), .B1(net_12935), .B2(net_12518), .A(net_8839) );
NAND2_X2 inst_8600 ( .A2(net_21134), .ZN(net_19142), .A1(net_16675) );
NAND2_X4 inst_7236 ( .ZN(net_8368), .A1(net_7010), .A2(net_7009) );
NAND2_X2 inst_9989 ( .ZN(net_13800), .A2(net_6969), .A1(net_3383) );
SDFF_X2 inst_913 ( .Q(net_21128), .D(net_16678), .SE(net_263), .CK(net_21522), .SI(x4099) );
INV_X8 inst_12274 ( .ZN(net_9514), .A(net_5439) );
INV_X4 inst_12712 ( .A(net_17777), .ZN(net_17746) );
INV_X4 inst_18267 ( .A(net_19444), .ZN(net_19443) );
INV_X4 inst_16434 ( .ZN(net_9459), .A(net_2828) );
INV_X4 inst_15999 ( .ZN(net_15681), .A(net_15110) );
INV_X4 inst_17567 ( .ZN(net_2280), .A(net_612) );
INV_X4 inst_18120 ( .A(net_21142), .ZN(net_17015) );
INV_X4 inst_15188 ( .A(net_7712), .ZN(net_4666) );
INV_X4 inst_15502 ( .ZN(net_3761), .A(net_2421) );
NAND3_X2 inst_6633 ( .ZN(net_8989), .A2(net_8988), .A3(net_8987), .A1(net_5729) );
NAND2_X2 inst_10322 ( .ZN(net_9327), .A1(net_7812), .A2(net_7811) );
NAND2_X2 inst_12004 ( .ZN(net_1609), .A2(net_1174), .A1(net_873) );
NAND2_X2 inst_9298 ( .ZN(net_12394), .A1(net_12393), .A2(net_12342) );
NAND2_X2 inst_11214 ( .ZN(net_4006), .A2(net_2817), .A1(net_1884) );
OAI211_X2 inst_2483 ( .ZN(net_13482), .B(net_13481), .C2(net_11357), .A(net_10724), .C1(net_3369) );
OAI21_X4 inst_1414 ( .A(net_20904), .ZN(net_20390), .B2(net_19031), .B1(net_19030) );
NAND2_X4 inst_7624 ( .A2(net_2001), .A1(net_1344), .ZN(net_1268) );
INV_X4 inst_16101 ( .ZN(net_15955), .A(net_14630) );
INV_X4 inst_17658 ( .ZN(net_14308), .A(net_261) );
NAND2_X2 inst_8451 ( .ZN(net_17206), .A2(net_16751), .A1(net_16616) );
NOR2_X2 inst_3994 ( .ZN(net_8271), .A2(net_6094), .A1(net_6026) );
XNOR2_X2 inst_449 ( .B(net_21108), .A(net_17262), .ZN(net_14851) );
CLKBUF_X2 inst_22665 ( .A(net_22536), .Z(net_22537) );
CLKBUF_X2 inst_22603 ( .A(net_22474), .Z(net_22475) );
NAND2_X2 inst_10797 ( .A1(net_8041), .ZN(net_7289), .A2(net_3935) );
CLKBUF_X2 inst_22815 ( .A(net_22607), .Z(net_22687) );
NAND2_X2 inst_10354 ( .ZN(net_13412), .A1(net_7465), .A2(net_4579) );
NOR3_X2 inst_2790 ( .ZN(net_4510), .A1(net_2491), .A3(net_2025), .A2(net_1173) );
OAI21_X2 inst_2138 ( .ZN(net_13167), .A(net_9254), .B1(net_6395), .B2(net_5683) );
NAND2_X4 inst_7152 ( .ZN(net_10987), .A1(net_8588), .A2(net_7886) );
NAND3_X4 inst_5599 ( .ZN(net_14580), .A3(net_11818), .A2(net_10278), .A1(net_8327) );
INV_X4 inst_16823 ( .A(net_7455), .ZN(net_5432) );
INV_X2 inst_19209 ( .ZN(net_3522), .A(net_3521) );
NAND3_X2 inst_6593 ( .ZN(net_9953), .A2(net_5315), .A3(net_4721), .A1(net_3209) );
NAND2_X2 inst_11417 ( .ZN(net_7380), .A2(net_3766), .A1(net_409) );
NAND3_X2 inst_6055 ( .ZN(net_14230), .A2(net_13608), .A1(net_13400), .A3(net_11606) );
INV_X4 inst_13362 ( .ZN(net_12345), .A(net_10936) );
NOR2_X4 inst_3249 ( .ZN(net_3077), .A1(net_2328), .A2(net_2099) );
NOR2_X2 inst_4935 ( .ZN(net_10168), .A2(net_9342), .A1(net_609) );
INV_X4 inst_17505 ( .ZN(net_9461), .A(net_690) );
NAND2_X2 inst_8961 ( .A1(net_20897), .ZN(net_14698), .A2(net_13218) );
NAND2_X4 inst_7498 ( .ZN(net_3112), .A1(net_2327), .A2(net_1216) );
CLKBUF_X2 inst_21852 ( .A(net_21640), .Z(net_21724) );
NAND2_X2 inst_9860 ( .A1(net_20549), .ZN(net_9497), .A2(net_9496) );
INV_X8 inst_12420 ( .A(net_20892), .ZN(net_1733) );
INV_X4 inst_13369 ( .ZN(net_12322), .A(net_10906) );
NAND2_X2 inst_11044 ( .A1(net_8276), .ZN(net_4719), .A2(net_3931) );
INV_X4 inst_12973 ( .ZN(net_17233), .A(net_16512) );
CLKBUF_X2 inst_22501 ( .A(net_21540), .Z(net_22373) );
INV_X2 inst_19103 ( .A(net_6243), .ZN(net_4500) );
NAND2_X2 inst_8201 ( .ZN(net_17878), .A2(net_17755), .A1(net_17661) );
NOR2_X2 inst_3614 ( .ZN(net_12381), .A2(net_12380), .A1(net_10740) );
NAND2_X2 inst_8893 ( .A1(net_20699), .ZN(net_15112), .A2(net_14022) );
INV_X2 inst_18672 ( .ZN(net_9123), .A(net_9122) );
INV_X4 inst_16224 ( .ZN(net_9260), .A(net_1478) );
INV_X4 inst_12776 ( .ZN(net_17322), .A(net_17321) );
XNOR2_X2 inst_588 ( .B(net_17494), .ZN(net_569), .A(net_568) );
NAND2_X2 inst_10752 ( .ZN(net_5699), .A2(net_5474), .A1(net_3760) );
NAND2_X2 inst_10394 ( .A1(net_14337), .ZN(net_7303), .A2(net_7302) );
NAND2_X2 inst_11411 ( .ZN(net_4560), .A1(net_2096), .A2(net_2048) );
INV_X4 inst_16488 ( .ZN(net_12179), .A(net_10091) );
INV_X4 inst_17296 ( .ZN(net_5205), .A(net_809) );
AOI211_X2 inst_21051 ( .ZN(net_12420), .C1(net_12419), .C2(net_8449), .B(net_7433), .A(net_5997) );
INV_X4 inst_14015 ( .ZN(net_7638), .A(net_6303) );
NAND2_X2 inst_10329 ( .ZN(net_7724), .A2(net_7723), .A1(net_4525) );
NAND2_X2 inst_9405 ( .ZN(net_20276), .A1(net_11682), .A2(net_11136) );
INV_X4 inst_16557 ( .ZN(net_2350), .A(net_1168) );
INV_X2 inst_19063 ( .A(net_6807), .ZN(net_4650) );
NAND2_X2 inst_11060 ( .ZN(net_4603), .A1(net_2588), .A2(net_2449) );
NOR2_X2 inst_4752 ( .A1(net_20568), .ZN(net_3848), .A2(net_3065) );
OAI21_X4 inst_1356 ( .ZN(net_20391), .A(net_18176), .B2(net_17479), .B1(net_17361) );
INV_X4 inst_12913 ( .ZN(net_16853), .A(net_16683) );
CLKBUF_X2 inst_22613 ( .A(net_22484), .Z(net_22485) );
NAND3_X2 inst_6447 ( .ZN(net_11768), .A2(net_11767), .A3(net_11766), .A1(net_2972) );
NOR3_X4 inst_2628 ( .ZN(net_15037), .A3(net_12818), .A1(net_12724), .A2(net_12591) );
CLKBUF_X2 inst_22076 ( .A(net_21947), .Z(net_21948) );
OAI21_X2 inst_2196 ( .A(net_10569), .ZN(net_8577), .B1(net_4016), .B2(net_3769) );
INV_X4 inst_14159 ( .ZN(net_9570), .A(net_7885) );
NAND2_X2 inst_7754 ( .ZN(net_18770), .A2(net_18746), .A1(net_18724) );
NAND2_X4 inst_7145 ( .ZN(net_12878), .A1(net_9750), .A2(net_9478) );
INV_X4 inst_14083 ( .ZN(net_7567), .A(net_6216) );
AOI21_X2 inst_20418 ( .ZN(net_15262), .B2(net_13897), .A(net_11515), .B1(net_11407) );
INV_X2 inst_19497 ( .ZN(net_1723), .A(net_835) );
SDFF_X2 inst_1045 ( .QN(net_21046), .D(net_354), .SE(net_263), .CK(net_22485), .SI(x2240) );
INV_X4 inst_18054 ( .A(net_21147), .ZN(net_437) );
INV_X4 inst_18042 ( .A(net_20946), .ZN(net_48) );
XNOR2_X2 inst_252 ( .ZN(net_17309), .A(net_17308), .B(net_9239) );
SDFF_X2 inst_865 ( .Q(net_21158), .D(net_17094), .SE(net_263), .CK(net_21470), .SI(x5409) );
SDFF_X2 inst_956 ( .QN(net_21011), .D(net_578), .SE(net_263), .CK(net_22735), .SI(x2855) );
NAND2_X2 inst_10959 ( .A2(net_19461), .ZN(net_8244), .A1(net_6177) );
INV_X4 inst_17269 ( .ZN(net_4211), .A(net_154) );
INV_X2 inst_18827 ( .A(net_11830), .ZN(net_6804) );
NAND2_X2 inst_10177 ( .A1(net_8748), .ZN(net_8198), .A2(net_8197) );
NOR2_X2 inst_4684 ( .ZN(net_3845), .A2(net_3065), .A1(net_655) );
INV_X4 inst_12757 ( .ZN(net_17401), .A(net_17400) );
XNOR2_X2 inst_484 ( .ZN(net_10802), .A(net_10801), .B(net_5793) );
INV_X4 inst_16041 ( .ZN(net_16011), .A(net_1613) );
AOI22_X2 inst_19977 ( .ZN(net_15483), .A2(net_14608), .B1(net_13565), .B2(net_13548), .A1(net_2072) );
NOR2_X2 inst_4474 ( .A1(net_9276), .ZN(net_4981), .A2(net_4118) );
NAND2_X2 inst_9272 ( .ZN(net_12602), .A2(net_10846), .A1(net_8618) );
INV_X4 inst_15902 ( .ZN(net_16281), .A(net_449) );
CLKBUF_X2 inst_22752 ( .A(net_22475), .Z(net_22624) );
XOR2_X2 inst_32 ( .A(net_21127), .Z(net_730), .B(net_729) );
NAND2_X2 inst_9129 ( .A1(net_14171), .ZN(net_13529), .A2(net_10794) );
OAI21_X2 inst_1821 ( .ZN(net_14157), .A(net_12325), .B2(net_10553), .B1(net_10031) );
CLKBUF_X2 inst_22472 ( .A(net_22343), .Z(net_22344) );
INV_X4 inst_16316 ( .ZN(net_1749), .A(net_299) );
NAND2_X4 inst_7271 ( .A1(net_20440), .ZN(net_9631), .A2(net_4810) );
AND2_X4 inst_21198 ( .A1(net_10325), .ZN(net_10110), .A2(net_7666) );
XNOR2_X2 inst_616 ( .ZN(net_490), .A(net_489), .B(net_488) );
NAND2_X2 inst_10683 ( .A1(net_20561), .ZN(net_6134), .A2(net_6042) );
INV_X4 inst_18293 ( .A(net_20438), .ZN(net_20437) );
NAND4_X2 inst_5381 ( .ZN(net_15051), .A2(net_12977), .A4(net_12513), .A1(net_11058), .A3(net_5949) );
AOI21_X2 inst_20560 ( .ZN(net_14255), .B2(net_14254), .A(net_11399), .B1(net_5750) );
OAI21_X2 inst_1784 ( .B2(net_19981), .B1(net_19980), .ZN(net_14658), .A(net_14657) );
INV_X2 inst_18670 ( .ZN(net_12342), .A(net_10240) );
CLKBUF_X2 inst_21636 ( .A(net_21332), .Z(net_21508) );
CLKBUF_X2 inst_21474 ( .A(net_21251), .Z(net_21346) );
NAND2_X2 inst_8040 ( .ZN(net_18250), .A1(net_18178), .A2(net_18154) );
CLKBUF_X2 inst_21802 ( .A(net_21673), .Z(net_21674) );
INV_X4 inst_16402 ( .ZN(net_15864), .A(net_15020) );
OAI21_X2 inst_2071 ( .ZN(net_20123), .A(net_14092), .B1(net_11476), .B2(net_6438) );
INV_X4 inst_14921 ( .A(net_4821), .ZN(net_4573) );
OAI21_X4 inst_1427 ( .ZN(net_16033), .B2(net_15497), .A(net_13666), .B1(net_588) );
NAND2_X2 inst_10421 ( .A1(net_13091), .ZN(net_7226), .A2(net_5522) );
NAND2_X2 inst_9183 ( .ZN(net_19707), .A1(net_10694), .A2(net_10169) );
NAND2_X4 inst_7259 ( .A1(net_19553), .ZN(net_7908), .A2(net_6692) );
NAND2_X2 inst_10056 ( .ZN(net_13165), .A1(net_9461), .A2(net_8688) );
AND2_X4 inst_21224 ( .ZN(net_19679), .A2(net_9819), .A1(net_8785) );
INV_X4 inst_17346 ( .A(net_2585), .ZN(net_777) );
NOR2_X2 inst_4662 ( .A1(net_14038), .A2(net_7002), .ZN(net_3285) );
INV_X4 inst_14296 ( .ZN(net_6871), .A(net_5549) );
XNOR2_X2 inst_87 ( .ZN(net_18566), .A(net_18500), .B(net_17768) );
INV_X4 inst_17704 ( .ZN(net_937), .A(net_215) );
INV_X4 inst_16172 ( .ZN(net_15699), .A(net_10891) );
NOR2_X4 inst_2918 ( .ZN(net_19779), .A2(net_8090), .A1(net_6045) );
NAND2_X2 inst_10036 ( .ZN(net_13231), .A2(net_10695), .A1(net_8328) );
NOR3_X2 inst_2721 ( .ZN(net_13255), .A1(net_10588), .A3(net_8566), .A2(net_8030) );
NAND2_X2 inst_9576 ( .ZN(net_10946), .A1(net_10945), .A2(net_7360) );
NOR2_X4 inst_3074 ( .ZN(net_10072), .A2(net_2514), .A1(net_399) );
SDFF_X2 inst_800 ( .Q(net_20951), .SE(net_18581), .SI(net_17982), .D(net_407), .CK(net_21268) );
NAND4_X2 inst_5281 ( .ZN(net_20758), .A2(net_20038), .A1(net_20037), .A4(net_15600), .A3(net_6677) );
XOR2_X2 inst_10 ( .A(net_21126), .B(net_17086), .Z(net_17073) );
NAND2_X2 inst_9925 ( .A2(net_20777), .A1(net_20465), .ZN(net_9228) );
NAND2_X2 inst_7770 ( .A2(net_20210), .ZN(net_18743), .A1(net_17080) );
NOR2_X2 inst_4337 ( .ZN(net_5697), .A2(net_5696), .A1(net_3232) );
INV_X4 inst_15550 ( .ZN(net_14241), .A(net_11430) );
NAND2_X2 inst_10475 ( .ZN(net_10606), .A2(net_8541), .A1(net_6982) );
NAND2_X2 inst_7981 ( .ZN(net_18338), .A2(net_18337), .A1(net_17998) );
INV_X4 inst_13555 ( .ZN(net_12408), .A(net_9161) );
NAND4_X2 inst_5459 ( .ZN(net_13413), .A3(net_13412), .A1(net_12500), .A4(net_9590), .A2(net_7158) );
INV_X4 inst_13186 ( .ZN(net_14225), .A(net_13622) );
CLKBUF_X2 inst_22106 ( .A(net_21977), .Z(net_21978) );
NAND2_X2 inst_9867 ( .A2(net_12757), .ZN(net_9488), .A1(net_9487) );
INV_X4 inst_18281 ( .A(net_20076), .ZN(net_20073) );
CLKBUF_X2 inst_21511 ( .A(net_21382), .Z(net_21383) );
NAND2_X2 inst_10090 ( .A1(net_9681), .ZN(net_8623), .A2(net_7923) );
INV_X4 inst_16623 ( .ZN(net_5845), .A(net_3174) );
NAND2_X2 inst_11961 ( .ZN(net_2645), .A2(net_1418), .A1(net_1385) );
INV_X4 inst_16443 ( .A(net_6812), .ZN(net_4751) );
INV_X2 inst_18368 ( .ZN(net_17723), .A(net_17722) );
NAND3_X2 inst_6700 ( .A1(net_14337), .A3(net_8696), .ZN(net_7361), .A2(net_6885) );
INV_X4 inst_14462 ( .ZN(net_6085), .A(net_4939) );
INV_X4 inst_16078 ( .ZN(net_11472), .A(net_6316) );
NOR2_X2 inst_4731 ( .A1(net_20548), .ZN(net_3974), .A2(net_2650) );
AOI21_X2 inst_20380 ( .B1(net_15955), .ZN(net_15558), .A(net_14388), .B2(net_14194) );
OAI22_X2 inst_1276 ( .A2(net_17290), .B2(net_17177), .ZN(net_16621), .A1(net_13655), .B1(net_8738) );
XNOR2_X2 inst_256 ( .B(net_21134), .ZN(net_17288), .A(net_17287) );
NAND3_X2 inst_6205 ( .ZN(net_13293), .A3(net_8817), .A1(net_8745), .A2(net_8654) );
OAI21_X2 inst_1902 ( .A(net_14006), .ZN(net_13328), .B1(net_9105), .B2(net_5566) );
NAND2_X2 inst_9180 ( .ZN(net_13334), .A2(net_10741), .A1(net_8576) );
INV_X4 inst_16518 ( .ZN(net_1743), .A(net_755) );
NAND2_X2 inst_8626 ( .A1(net_21165), .ZN(net_20743), .A2(net_16605) );
NAND2_X2 inst_9635 ( .ZN(net_13127), .A1(net_12542), .A2(net_9808) );
DFF_X1 inst_19829 ( .D(net_17525), .CK(net_21995), .Q(x936) );
NOR2_X2 inst_5052 ( .ZN(net_6449), .A1(net_1155), .A2(net_429) );
INV_X4 inst_16874 ( .ZN(net_10031), .A(net_3814) );
AOI21_X2 inst_20399 ( .ZN(net_15412), .B1(net_15411), .B2(net_14383), .A(net_6748) );
NAND3_X2 inst_6038 ( .ZN(net_14326), .A3(net_13209), .A2(net_11473), .A1(net_9534) );
INV_X4 inst_13791 ( .ZN(net_9043), .A(net_7564) );
NOR2_X2 inst_3978 ( .ZN(net_8392), .A2(net_8391), .A1(net_8389) );
NAND3_X2 inst_6106 ( .ZN(net_13896), .A3(net_13053), .A2(net_9716), .A1(net_8599) );
NAND2_X2 inst_11264 ( .A1(net_10667), .A2(net_4192), .ZN(net_3897) );
NAND2_X2 inst_9354 ( .ZN(net_12164), .A2(net_12163), .A1(net_10328) );
NAND2_X2 inst_10042 ( .ZN(net_19777), .A2(net_8712), .A1(net_7622) );
NAND2_X2 inst_10214 ( .ZN(net_19544), .A1(net_8088), .A2(net_8087) );
OAI21_X2 inst_2078 ( .ZN(net_10556), .A(net_10002), .B2(net_6405), .B1(net_3663) );
NAND2_X2 inst_9161 ( .ZN(net_13380), .A1(net_12551), .A2(net_10439) );
NAND3_X2 inst_6555 ( .A3(net_20125), .ZN(net_19965), .A1(net_10523), .A2(net_7558) );
AOI21_X4 inst_20219 ( .ZN(net_14118), .B1(net_13512), .A(net_11071), .B2(net_10443) );
INV_X2 inst_18773 ( .ZN(net_20266), .A(net_9540) );
INV_X4 inst_17422 ( .ZN(net_2563), .A(net_955) );
OAI21_X4 inst_1462 ( .ZN(net_19532), .B2(net_19127), .B1(net_19126), .A(net_238) );
NAND2_X2 inst_8509 ( .A1(net_21212), .ZN(net_20404), .A2(net_16922) );
OAI21_X2 inst_2273 ( .A(net_10930), .ZN(net_7137), .B2(net_7136), .B1(net_4316) );
AND2_X4 inst_21241 ( .ZN(net_11220), .A2(net_5269), .A1(net_859) );
DFF_X1 inst_19835 ( .D(net_17417), .CK(net_22804), .Q(x1215) );
NAND2_X2 inst_9138 ( .ZN(net_13441), .A2(net_13367), .A1(net_13213) );
NAND3_X2 inst_6391 ( .ZN(net_12003), .A3(net_11340), .A2(net_7440), .A1(net_7040) );
INV_X4 inst_13944 ( .ZN(net_8111), .A(net_6803) );
OAI21_X2 inst_2003 ( .ZN(net_11619), .A(net_9861), .B2(net_7526), .B1(net_3959) );
INV_X4 inst_15954 ( .ZN(net_2113), .A(net_1707) );
NAND3_X2 inst_6100 ( .ZN(net_13908), .A1(net_12054), .A2(net_11031), .A3(net_10064) );
NAND3_X2 inst_6084 ( .ZN(net_13960), .A3(net_11177), .A1(net_9385), .A2(net_3616) );
NAND4_X2 inst_5430 ( .A2(net_19689), .A1(net_19688), .ZN(net_14110), .A4(net_10969), .A3(net_4887) );
CLKBUF_X2 inst_21859 ( .A(net_21338), .Z(net_21731) );
NOR2_X2 inst_5119 ( .ZN(net_299), .A1(net_162), .A2(net_137) );
NOR2_X2 inst_4963 ( .A2(net_20860), .ZN(net_1603), .A1(net_1602) );
NOR3_X2 inst_2787 ( .ZN(net_5577), .A1(net_5576), .A2(net_5402), .A3(net_4014) );
NAND3_X4 inst_5612 ( .ZN(net_20451), .A3(net_8921), .A2(net_8082), .A1(net_8042) );
INV_X4 inst_13638 ( .A(net_10530), .ZN(net_8188) );
INV_X8 inst_12455 ( .A(net_20766), .ZN(net_20765) );
NAND2_X2 inst_9386 ( .ZN(net_11935), .A1(net_9454), .A2(net_7328) );
NAND2_X2 inst_11074 ( .A1(net_8618), .ZN(net_4480), .A2(net_2009) );
NOR4_X2 inst_2599 ( .ZN(net_15722), .A1(net_15150), .A4(net_13845), .A2(net_11403), .A3(net_10132) );
INV_X4 inst_16062 ( .ZN(net_4098), .A(net_1580) );
NAND3_X2 inst_6254 ( .ZN(net_13008), .A3(net_13007), .A2(net_11353), .A1(net_9094) );
CLKBUF_X2 inst_22191 ( .A(net_22062), .Z(net_22063) );
INV_X4 inst_18286 ( .A(net_20210), .ZN(net_20208) );
NOR2_X2 inst_3971 ( .A1(net_9250), .ZN(net_8407), .A2(net_8366) );
NAND2_X2 inst_11573 ( .A2(net_7399), .ZN(net_6776), .A1(net_1696) );
NAND2_X2 inst_9858 ( .ZN(net_9503), .A1(net_9502), .A2(net_6066) );
INV_X2 inst_18772 ( .ZN(net_7569), .A(net_7568) );
INV_X4 inst_13596 ( .A(net_11882), .ZN(net_8774) );
INV_X4 inst_18013 ( .A(net_20979), .ZN(net_2432) );
OR2_X4 inst_1123 ( .ZN(net_2221), .A2(net_252), .A1(net_143) );
INV_X4 inst_18028 ( .A(net_21137), .ZN(net_17422) );
NAND2_X2 inst_8747 ( .ZN(net_19581), .A1(net_15825), .A2(net_15377) );
INV_X4 inst_13383 ( .A(net_12962), .ZN(net_10770) );
INV_X4 inst_17256 ( .ZN(net_3054), .A(net_2629) );
NAND2_X2 inst_11763 ( .ZN(net_4041), .A1(net_1823), .A2(net_783) );
CLKBUF_X2 inst_22254 ( .A(net_22125), .Z(net_22126) );
NAND2_X4 inst_7169 ( .ZN(net_12900), .A1(net_7308), .A2(net_874) );
INV_X4 inst_16429 ( .ZN(net_4301), .A(net_2996) );
NAND2_X2 inst_8061 ( .ZN(net_18197), .A2(net_18130), .A1(net_18113) );
OAI21_X2 inst_1628 ( .ZN(net_20650), .B2(net_15443), .B1(net_14080), .A(net_588) );
NAND2_X4 inst_6844 ( .ZN(net_18723), .A1(net_18643), .A2(net_18631) );
DFF_X1 inst_19804 ( .D(net_18173), .CK(net_22822), .Q(x1087) );
INV_X4 inst_17506 ( .A(net_1299), .ZN(net_857) );
NAND2_X2 inst_9640 ( .ZN(net_10391), .A2(net_9821), .A1(net_7204) );
NOR2_X2 inst_4840 ( .ZN(net_3944), .A2(net_2369), .A1(net_168) );
XNOR2_X2 inst_225 ( .ZN(net_17503), .A(net_17502), .B(net_13282) );
INV_X4 inst_12530 ( .ZN(net_18412), .A(net_18411) );
INV_X4 inst_14261 ( .ZN(net_14348), .A(net_4350) );
INV_X4 inst_17832 ( .ZN(net_12133), .A(net_10216) );
NOR2_X2 inst_5020 ( .A1(net_1415), .ZN(net_1199), .A2(net_922) );
NAND2_X2 inst_9030 ( .A1(net_15573), .ZN(net_14073), .A2(net_11896) );
NAND2_X4 inst_7349 ( .ZN(net_7833), .A2(net_4093), .A1(net_3340) );
INV_X4 inst_14808 ( .A(net_9493), .ZN(net_3971) );
XNOR2_X2 inst_508 ( .ZN(net_7651), .A(net_7650), .B(net_3437) );
NOR2_X2 inst_4888 ( .A1(net_6091), .ZN(net_3959), .A2(net_2110) );
NAND2_X2 inst_8150 ( .ZN(net_18014), .A2(net_17966), .A1(net_17937) );
CLKBUF_X2 inst_21699 ( .A(net_21486), .Z(net_21571) );
INV_X4 inst_12611 ( .A(net_18147), .ZN(net_18101) );
XNOR2_X2 inst_590 ( .A(net_16648), .B(net_16646), .ZN(net_1676) );
OAI211_X2 inst_2553 ( .ZN(net_10498), .B(net_8793), .A(net_5177), .C1(net_3400), .C2(net_2929) );
INV_X2 inst_18427 ( .ZN(net_20724), .A(net_14508) );
INV_X8 inst_12209 ( .ZN(net_9496), .A(net_4812) );
INV_X4 inst_12671 ( .ZN(net_17759), .A(net_17758) );
INV_X4 inst_13051 ( .ZN(net_16383), .A(net_16382) );
INV_X4 inst_13897 ( .ZN(net_7179), .A(net_5693) );
AOI21_X2 inst_20491 ( .ZN(net_14756), .B1(net_14755), .B2(net_12289), .A(net_8268) );
NOR2_X2 inst_4531 ( .ZN(net_4443), .A1(net_4228), .A2(net_4022) );
OR2_X4 inst_1105 ( .ZN(net_2249), .A2(net_1602), .A1(net_1058) );
NOR3_X2 inst_2746 ( .A1(net_20184), .ZN(net_12577), .A3(net_7852), .A2(net_7146) );
INV_X4 inst_14746 ( .ZN(net_7343), .A(net_4277) );
INV_X4 inst_14387 ( .A(net_8035), .ZN(net_5145) );
NAND2_X4 inst_6961 ( .A2(net_20089), .A1(net_20088), .ZN(net_17439) );
NAND2_X2 inst_8200 ( .A1(net_20634), .ZN(net_17883), .A2(net_17437) );
XNOR2_X2 inst_330 ( .ZN(net_17002), .A(net_17000), .B(net_12264) );
INV_X4 inst_13345 ( .ZN(net_11071), .A(net_11070) );
INV_X4 inst_13558 ( .ZN(net_12405), .A(net_9158) );
AOI21_X4 inst_20116 ( .ZN(net_19613), .B2(net_16005), .A(net_15200), .B1(net_1052) );
NOR2_X2 inst_4305 ( .ZN(net_9460), .A1(net_4569), .A2(net_154) );
NAND2_X2 inst_12101 ( .A2(net_874), .ZN(net_487), .A1(net_251) );
INV_X4 inst_13546 ( .A(net_11918), .ZN(net_10761) );
NAND2_X2 inst_8786 ( .ZN(net_15754), .A1(net_15753), .A2(net_15160) );
NOR2_X2 inst_3566 ( .ZN(net_12828), .A2(net_10311), .A1(net_4425) );
INV_X4 inst_13864 ( .A(net_9496), .ZN(net_7457) );
NAND2_X2 inst_11803 ( .A2(net_19418), .ZN(net_1909), .A1(net_107) );
AOI211_X2 inst_21031 ( .B(net_15202), .ZN(net_14386), .A(net_13785), .C2(net_11628), .C1(net_10010) );
INV_X4 inst_15455 ( .ZN(net_15876), .A(net_15694) );
CLKBUF_X2 inst_22943 ( .A(net_22814), .Z(net_22815) );
AOI211_X2 inst_21074 ( .B(net_8563), .ZN(net_7682), .C2(net_7681), .A(net_4453), .C1(net_2773) );
INV_X4 inst_16108 ( .ZN(net_2831), .A(net_1499) );
OR2_X2 inst_1232 ( .ZN(net_12930), .A2(net_7325), .A1(net_126) );
INV_X4 inst_14431 ( .A(net_5029), .ZN(net_5028) );
INV_X4 inst_16562 ( .ZN(net_13198), .A(net_10592) );
INV_X2 inst_18968 ( .A(net_15519), .ZN(net_5294) );
SDFF_X2 inst_758 ( .Q(net_20933), .SE(net_18576), .SI(net_18525), .D(net_444), .CK(net_21434) );
INV_X4 inst_17915 ( .ZN(net_251), .A(net_120) );
OAI21_X2 inst_2146 ( .B1(net_10714), .ZN(net_9864), .B2(net_8833), .A(net_2711) );
INV_X4 inst_13332 ( .ZN(net_13012), .A(net_11134) );
NAND2_X2 inst_8543 ( .A2(net_17126), .ZN(net_16817), .A1(net_16636) );
NOR2_X2 inst_3437 ( .ZN(net_15253), .A2(net_14736), .A1(net_2594) );
INV_X4 inst_13425 ( .A(net_10995), .ZN(net_10785) );
NAND3_X2 inst_6813 ( .A2(net_4394), .ZN(net_3000), .A3(net_2384), .A1(net_135) );
INV_X4 inst_17777 ( .ZN(net_2493), .A(net_1509) );
NAND3_X2 inst_5764 ( .A1(net_19591), .ZN(net_18996), .A3(net_11865), .A2(net_3735) );
NAND2_X4 inst_7442 ( .A1(net_20875), .ZN(net_4784), .A2(net_3192) );
OAI21_X2 inst_1953 ( .ZN(net_12552), .A(net_12551), .B2(net_7523), .B1(net_4764) );
NOR2_X2 inst_4570 ( .ZN(net_20782), .A1(net_2794), .A2(net_940) );
NOR2_X4 inst_3016 ( .ZN(net_6843), .A2(net_3918), .A1(net_2274) );
OAI21_X2 inst_1958 ( .ZN(net_19738), .A(net_9128), .B2(net_8833), .B1(net_6696) );
INV_X4 inst_14050 ( .ZN(net_9822), .A(net_6252) );
INV_X2 inst_18639 ( .ZN(net_9382), .A(net_9381) );
NAND2_X4 inst_6885 ( .A1(net_20505), .ZN(net_18146), .A2(net_17177) );
NOR2_X4 inst_3240 ( .ZN(net_4180), .A2(net_2258), .A1(net_131) );
NAND2_X2 inst_9403 ( .ZN(net_11685), .A2(net_11068), .A1(net_6190) );
AOI21_X2 inst_20821 ( .A(net_13781), .ZN(net_10003), .B2(net_10002), .B1(net_8189) );
INV_X4 inst_17201 ( .ZN(net_4685), .A(net_706) );
INV_X4 inst_16950 ( .ZN(net_5572), .A(net_912) );
INV_X2 inst_19022 ( .ZN(net_12317), .A(net_6616) );
XNOR2_X2 inst_111 ( .ZN(net_18539), .A(net_18384), .B(net_18210) );
INV_X4 inst_13196 ( .ZN(net_14040), .A(net_13376) );
AOI21_X2 inst_20394 ( .ZN(net_15460), .B1(net_14459), .B2(net_14452), .A(net_11407) );
OAI21_X2 inst_1723 ( .B2(net_19469), .B1(net_19468), .ZN(net_15094), .A(net_14472) );
NOR2_X4 inst_3278 ( .ZN(net_3061), .A1(net_1630), .A2(net_1303) );
NAND2_X2 inst_11425 ( .ZN(net_4422), .A1(net_3719), .A2(net_3120) );
NOR2_X2 inst_5145 ( .ZN(net_664), .A2(net_26), .A1(net_25) );
NAND2_X2 inst_11296 ( .ZN(net_11746), .A1(net_3812), .A2(net_3811) );
INV_X4 inst_16703 ( .A(net_11189), .ZN(net_9638) );
INV_X4 inst_13407 ( .ZN(net_10359), .A(net_8882) );
INV_X2 inst_19433 ( .A(net_12203), .ZN(net_1744) );
INV_X4 inst_17906 ( .ZN(net_792), .A(net_466) );
SDFF_X2 inst_978 ( .QN(net_21084), .D(net_527), .SE(net_263), .CK(net_22589), .SI(x1662) );
INV_X4 inst_14757 ( .A(net_13375), .ZN(net_13026) );
NOR2_X4 inst_2955 ( .ZN(net_8708), .A1(net_6812), .A2(net_5174) );
INV_X4 inst_13506 ( .ZN(net_9415), .A(net_9414) );
NOR2_X2 inst_3926 ( .A2(net_11589), .A1(net_10142), .ZN(net_8747) );
NAND2_X4 inst_7293 ( .ZN(net_7337), .A2(net_5575), .A1(net_809) );
INV_X4 inst_16515 ( .ZN(net_2232), .A(net_947) );
INV_X4 inst_13160 ( .ZN(net_14819), .A(net_14239) );
INV_X4 inst_17765 ( .A(net_874), .ZN(net_454) );
CLKBUF_X2 inst_22337 ( .A(net_21696), .Z(net_22209) );
NAND2_X2 inst_9745 ( .ZN(net_15800), .A1(net_14367), .A2(net_11150) );
INV_X4 inst_18295 ( .A(net_20441), .ZN(net_20440) );
INV_X2 inst_19030 ( .A(net_9692), .ZN(net_8076) );
XNOR2_X2 inst_495 ( .B(net_16599), .ZN(net_9007), .A(net_9006) );
INV_X4 inst_14366 ( .ZN(net_8197), .A(net_5781) );
INV_X4 inst_15041 ( .ZN(net_4408), .A(net_3340) );
NAND3_X2 inst_6437 ( .ZN(net_11827), .A2(net_11826), .A1(net_7456), .A3(net_6786) );
OAI21_X2 inst_1864 ( .ZN(net_13777), .B1(net_13776), .B2(net_11026), .A(net_449) );
NAND2_X2 inst_9632 ( .ZN(net_10408), .A1(net_10407), .A2(net_10406) );
NOR2_X4 inst_3224 ( .ZN(net_5114), .A1(net_3070), .A2(net_252) );
INV_X4 inst_16626 ( .A(net_9966), .ZN(net_9083) );
NAND2_X2 inst_10887 ( .ZN(net_5740), .A2(net_5343), .A1(net_998) );
CLKBUF_X2 inst_22073 ( .A(net_21944), .Z(net_21945) );
INV_X2 inst_18534 ( .ZN(net_11074), .A(net_11073) );
CLKBUF_X2 inst_21629 ( .A(net_21377), .Z(net_21501) );
NAND2_X2 inst_7917 ( .ZN(net_18456), .A2(net_18385), .A1(net_17814) );
CLKBUF_X2 inst_22028 ( .A(net_21899), .Z(net_21900) );
INV_X4 inst_12616 ( .ZN(net_18065), .A(net_18057) );
INV_X4 inst_15826 ( .A(net_9401), .ZN(net_4512) );
INV_X4 inst_16852 ( .ZN(net_3836), .A(net_2539) );
INV_X4 inst_13305 ( .A(net_13399), .ZN(net_12195) );
NAND2_X4 inst_7286 ( .A1(net_20335), .ZN(net_10790), .A2(net_5476) );
INV_X4 inst_12644 ( .ZN(net_17888), .A(net_17887) );
NAND2_X2 inst_8914 ( .ZN(net_14968), .A1(net_14706), .A2(net_13749) );
INV_X4 inst_18150 ( .A(net_21165), .ZN(net_16464) );
NOR2_X4 inst_2893 ( .ZN(net_10932), .A1(net_9445), .A2(net_547) );
NAND2_X2 inst_9497 ( .ZN(net_15595), .A1(net_14365), .A2(net_11479) );
AOI21_X2 inst_20953 ( .B1(net_9342), .ZN(net_5341), .A(net_4172), .B2(net_2227) );
NAND3_X2 inst_6727 ( .A1(net_20795), .ZN(net_6493), .A2(net_6492), .A3(net_6491) );
INV_X8 inst_12447 ( .ZN(net_20535), .A(net_20529) );
CLKBUF_X2 inst_21580 ( .A(net_21451), .Z(net_21452) );
NAND2_X2 inst_7937 ( .ZN(net_18431), .A2(net_18370), .A1(net_18316) );
NAND3_X2 inst_6347 ( .ZN(net_12235), .A3(net_9975), .A2(net_9695), .A1(net_8297) );
CLKBUF_X2 inst_22627 ( .A(net_22498), .Z(net_22499) );
OAI21_X4 inst_1453 ( .A(net_15353), .ZN(net_15352), .B2(net_13677), .B1(net_10095) );
INV_X4 inst_12466 ( .ZN(net_19955), .A(net_18789) );
NAND2_X2 inst_8871 ( .A1(net_15699), .ZN(net_15288), .A2(net_14251) );
INV_X4 inst_17961 ( .A(net_20946), .ZN(net_70) );
NOR2_X4 inst_3007 ( .ZN(net_9285), .A2(net_5754), .A1(net_3333) );
INV_X4 inst_18344 ( .A(net_20772), .ZN(net_20771) );
INV_X4 inst_15081 ( .A(net_6404), .ZN(net_3638) );
NOR2_X2 inst_4185 ( .A1(net_11214), .ZN(net_8055), .A2(net_4818) );
AOI21_X2 inst_20504 ( .B1(net_14751), .ZN(net_14639), .B2(net_12086), .A(net_5264) );
NAND3_X2 inst_6358 ( .ZN(net_18912), .A2(net_10681), .A1(net_9230), .A3(net_7861) );
NOR2_X2 inst_3512 ( .ZN(net_13826), .A1(net_13444), .A2(net_12577) );
NAND2_X2 inst_11018 ( .A2(net_12262), .ZN(net_5967), .A1(net_3900) );
NAND2_X2 inst_11485 ( .ZN(net_11805), .A1(net_6682), .A2(net_3088) );
NAND2_X2 inst_10738 ( .ZN(net_14544), .A1(net_8190), .A2(net_6960) );
NAND3_X2 inst_5632 ( .ZN(net_18793), .A2(net_18777), .A3(net_18776), .A1(net_17722) );
INV_X4 inst_14839 ( .ZN(net_13878), .A(net_5384) );
OR2_X2 inst_1206 ( .ZN(net_5853), .A2(net_3389), .A1(net_90) );
INV_X4 inst_15778 ( .ZN(net_8991), .A(net_2420) );
INV_X4 inst_15270 ( .ZN(net_3537), .A(net_2046) );
NAND3_X2 inst_6773 ( .ZN(net_5141), .A2(net_3758), .A1(net_2654), .A3(net_893) );
INV_X4 inst_15485 ( .ZN(net_2443), .A(net_2442) );
NAND2_X4 inst_7075 ( .A2(net_19629), .A1(net_19628), .ZN(net_19115) );
NAND2_X2 inst_10328 ( .ZN(net_7732), .A1(net_7731), .A2(net_3008) );
NOR2_X2 inst_3466 ( .ZN(net_19184), .A2(net_13244), .A1(net_8129) );
NAND2_X2 inst_8106 ( .ZN(net_18113), .A2(net_18112), .A1(net_16683) );
NAND2_X2 inst_8358 ( .A2(net_17607), .ZN(net_17449), .A1(net_17448) );
INV_X4 inst_13907 ( .ZN(net_8895), .A(net_7016) );
NOR2_X2 inst_4800 ( .ZN(net_3877), .A2(net_2992), .A1(net_143) );
NOR2_X2 inst_4394 ( .A1(net_8836), .ZN(net_5196), .A2(net_5195) );
INV_X4 inst_15684 ( .A(net_3459), .ZN(net_2632) );
NAND2_X2 inst_11303 ( .ZN(net_4771), .A2(net_3866), .A1(net_3789) );
INV_X4 inst_12631 ( .ZN(net_18840), .A(net_17922) );
INV_X4 inst_13086 ( .ZN(net_16028), .A(net_15916) );
OAI21_X4 inst_1487 ( .ZN(net_14798), .B1(net_12428), .B2(net_8575), .A(net_4931) );
CLKBUF_X2 inst_21410 ( .A(net_21281), .Z(net_21282) );
NAND2_X2 inst_7807 ( .ZN(net_18686), .A2(net_18665), .A1(net_17076) );
NAND2_X4 inst_7246 ( .ZN(net_8811), .A2(net_6854), .A1(net_6853) );
OAI21_X2 inst_1933 ( .B1(net_15375), .ZN(net_12933), .A(net_12932), .B2(net_9268) );
INV_X4 inst_13169 ( .ZN(net_14625), .A(net_14127) );
NAND2_X4 inst_7511 ( .A2(net_19347), .ZN(net_3977), .A1(net_2950) );
INV_X2 inst_18996 ( .ZN(net_5068), .A(net_5067) );
NAND2_X2 inst_12025 ( .ZN(net_2978), .A2(net_344), .A1(net_211) );
NOR2_X2 inst_4320 ( .A2(net_5894), .ZN(net_5870), .A1(net_5869) );
CLKBUF_X2 inst_21540 ( .A(net_21396), .Z(net_21412) );
INV_X2 inst_19493 ( .A(net_2497), .ZN(net_1294) );
CLKBUF_X2 inst_22517 ( .A(net_22388), .Z(net_22389) );
INV_X4 inst_16120 ( .ZN(net_19254), .A(net_2627) );
INV_X4 inst_16031 ( .ZN(net_2494), .A(net_1628) );
NAND2_X4 inst_7572 ( .ZN(net_4014), .A1(net_1403), .A2(net_1271) );
NAND3_X2 inst_6313 ( .ZN(net_12740), .A3(net_11120), .A1(net_6072), .A2(net_5538) );
NAND2_X4 inst_7680 ( .A2(net_1271), .ZN(net_1168), .A1(net_795) );
INV_X4 inst_16810 ( .A(net_3115), .ZN(net_2948) );
INV_X4 inst_18101 ( .A(net_21226), .ZN(net_189) );
INV_X4 inst_15516 ( .ZN(net_3144), .A(net_2405) );
INV_X4 inst_14228 ( .A(net_5833), .ZN(net_5832) );
INV_X4 inst_14316 ( .ZN(net_9028), .A(net_5471) );
INV_X4 inst_14182 ( .ZN(net_12795), .A(net_7833) );
NOR2_X2 inst_4771 ( .ZN(net_6376), .A2(net_2964), .A1(net_2113) );
INV_X4 inst_16986 ( .ZN(net_881), .A(net_333) );
INV_X4 inst_16375 ( .ZN(net_15731), .A(net_15107) );
NAND2_X4 inst_7695 ( .ZN(net_803), .A2(net_246), .A1(net_73) );
NOR2_X2 inst_4669 ( .ZN(net_3930), .A1(net_3254), .A2(net_3253) );
INV_X4 inst_15091 ( .A(net_5674), .ZN(net_4312) );
AOI21_X2 inst_20889 ( .ZN(net_7789), .B1(net_7432), .B2(net_6369), .A(net_6349) );
INV_X4 inst_15476 ( .ZN(net_3954), .A(net_2428) );
NAND2_X2 inst_8016 ( .ZN(net_18282), .A2(net_18261), .A1(net_17996) );
NAND2_X2 inst_8707 ( .ZN(net_16284), .A2(net_16149), .A1(net_16069) );
INV_X4 inst_13204 ( .ZN(net_13857), .A(net_13172) );
INV_X4 inst_15191 ( .ZN(net_5200), .A(net_2257) );
INV_X8 inst_12230 ( .ZN(net_7124), .A(net_3643) );
INV_X4 inst_15650 ( .ZN(net_3771), .A(net_3019) );
SDFF_X2 inst_1017 ( .QN(net_21077), .D(net_589), .SE(net_253), .CK(net_22568), .SI(x1765) );
CLKBUF_X2 inst_21881 ( .A(net_21752), .Z(net_21753) );
INV_X4 inst_13802 ( .A(net_9710), .ZN(net_7551) );
XNOR2_X2 inst_281 ( .ZN(net_17169), .A(net_17168), .B(net_1510) );
CLKBUF_X2 inst_21663 ( .A(net_21534), .Z(net_21535) );
NAND3_X2 inst_6336 ( .ZN(net_12443), .A2(net_12442), .A3(net_12236), .A1(net_2059) );
NAND2_X2 inst_10306 ( .ZN(net_9398), .A1(net_6982), .A2(net_4927) );
NAND2_X4 inst_7062 ( .A2(net_20856), .A1(net_19109), .ZN(net_18917) );
OAI21_X2 inst_1836 ( .A(net_15659), .ZN(net_14044), .B1(net_11520), .B2(net_8746) );
INV_X4 inst_18103 ( .A(net_21176), .ZN(net_16842) );
NAND2_X4 inst_7005 ( .ZN(net_17184), .A1(net_16722), .A2(net_16567) );
CLKBUF_X2 inst_21715 ( .A(net_21366), .Z(net_21587) );
NOR2_X2 inst_4274 ( .A1(net_9571), .ZN(net_7536), .A2(net_4543) );
NOR2_X2 inst_4250 ( .ZN(net_6390), .A1(net_3747), .A2(net_3139) );
OAI21_X2 inst_2170 ( .ZN(net_8928), .A(net_7153), .B2(net_6144), .B1(net_2896) );
CLKBUF_X2 inst_21895 ( .A(net_21766), .Z(net_21767) );
NAND2_X4 inst_7414 ( .ZN(net_8580), .A2(net_4481), .A1(net_3761) );
INV_X4 inst_13322 ( .ZN(net_11449), .A(net_11448) );
INV_X4 inst_15490 ( .A(net_15955), .ZN(net_2434) );
CLKBUF_X2 inst_22924 ( .A(net_22795), .Z(net_22796) );
NOR2_X4 inst_2946 ( .ZN(net_8231), .A2(net_7414), .A1(net_4998) );
NAND2_X2 inst_9940 ( .ZN(net_10681), .A2(net_8518), .A1(net_8304) );
INV_X4 inst_14149 ( .ZN(net_9683), .A(net_6046) );
INV_X4 inst_16415 ( .ZN(net_2634), .A(net_1256) );
INV_X4 inst_15234 ( .ZN(net_4181), .A(net_4027) );
INV_X4 inst_13827 ( .ZN(net_13164), .A(net_9363) );
NAND2_X2 inst_10828 ( .ZN(net_6786), .A1(net_4183), .A2(net_4057) );
INV_X2 inst_18932 ( .ZN(net_5849), .A(net_5848) );
NOR2_X4 inst_3211 ( .A1(net_20490), .ZN(net_5419), .A2(net_3023) );
NAND2_X2 inst_10364 ( .ZN(net_10838), .A1(net_9461), .A2(net_7392) );
INV_X4 inst_12702 ( .A(net_18252), .ZN(net_18205) );
NAND2_X4 inst_7270 ( .ZN(net_12738), .A1(net_5964), .A2(net_809) );
DFF_X1 inst_19903 ( .D(net_16964), .CK(net_22073), .Q(x339) );
NAND2_X2 inst_10906 ( .ZN(net_5794), .A1(net_3574), .A2(net_1126) );
INV_X4 inst_14803 ( .ZN(net_6676), .A(net_6674) );
AOI21_X2 inst_20850 ( .B2(net_14384), .ZN(net_9088), .B1(net_9087), .A(net_81) );
INV_X2 inst_18415 ( .ZN(net_15857), .A(net_15705) );
OAI211_X2 inst_2386 ( .C1(net_16743), .ZN(net_16399), .C2(net_16167), .A(net_15910), .B(net_15235) );
INV_X4 inst_13846 ( .ZN(net_11464), .A(net_7474) );
NOR2_X2 inst_4103 ( .A2(net_12805), .ZN(net_7208), .A1(net_7207) );
OAI22_X2 inst_1267 ( .B1(net_21187), .ZN(net_17098), .A1(net_17097), .B2(net_16576), .A2(net_16536) );
OAI21_X4 inst_1507 ( .ZN(net_10777), .B2(net_7120), .B1(net_5689), .A(net_673) );
INV_X4 inst_15276 ( .ZN(net_5055), .A(net_2748) );
INV_X2 inst_19116 ( .ZN(net_6242), .A(net_4443) );
INV_X2 inst_19091 ( .A(net_6153), .ZN(net_4556) );
NAND2_X4 inst_7301 ( .ZN(net_10247), .A1(net_9514), .A2(net_5534) );
CLKBUF_X2 inst_22034 ( .A(net_21905), .Z(net_21906) );
CLKBUF_X2 inst_22693 ( .A(net_22564), .Z(net_22565) );
NAND2_X4 inst_7260 ( .ZN(net_7883), .A2(net_6135), .A1(net_4823) );
NOR2_X2 inst_3786 ( .A1(net_13093), .ZN(net_10100), .A2(net_9548) );
CLKBUF_X2 inst_22725 ( .A(net_22596), .Z(net_22597) );
CLKBUF_X2 inst_21584 ( .A(net_21455), .Z(net_21456) );
INV_X4 inst_14960 ( .ZN(net_5935), .A(net_3489) );
NAND2_X4 inst_7367 ( .ZN(net_6837), .A2(net_4242), .A1(net_3713) );
NOR2_X2 inst_3404 ( .ZN(net_15812), .A2(net_15263), .A1(net_3552) );
AND2_X2 inst_21301 ( .ZN(net_14416), .A2(net_11753), .A1(net_10447) );
NAND2_X2 inst_7878 ( .ZN(net_18528), .A2(net_18462), .A1(net_17701) );
NAND4_X2 inst_5351 ( .ZN(net_19534), .A1(net_14673), .A3(net_14542), .A4(net_13102), .A2(net_11483) );
XNOR2_X2 inst_542 ( .ZN(net_794), .A(net_793), .B(net_792) );
XNOR2_X2 inst_128 ( .ZN(net_18342), .B(net_18197), .A(net_16838) );
CLKBUF_X2 inst_22114 ( .A(net_21985), .Z(net_21986) );
INV_X4 inst_13589 ( .ZN(net_8888), .A(net_7310) );
INV_X2 inst_18946 ( .ZN(net_8033), .A(net_6662) );
INV_X4 inst_14172 ( .ZN(net_18964), .A(net_8830) );
INV_X4 inst_14322 ( .ZN(net_5456), .A(net_5455) );
INV_X4 inst_13100 ( .ZN(net_15829), .A(net_15658) );
AOI21_X4 inst_20210 ( .ZN(net_20431), .B1(net_19528), .B2(net_14568), .A(net_11420) );
INV_X4 inst_13222 ( .ZN(net_13625), .A(net_12767) );
INV_X4 inst_15252 ( .ZN(net_4785), .A(net_2512) );
NOR2_X2 inst_4000 ( .ZN(net_9700), .A2(net_6867), .A1(net_6173) );
AOI211_X2 inst_21026 ( .ZN(net_14589), .C1(net_12916), .A(net_12228), .C2(net_11339), .B(net_8557) );
INV_X4 inst_13625 ( .ZN(net_14321), .A(net_8324) );
AOI21_X4 inst_20244 ( .B2(net_11702), .ZN(net_10081), .B1(net_5678), .A(net_1030) );
NOR2_X4 inst_3218 ( .A2(net_4374), .ZN(net_2754), .A1(net_2753) );
NAND2_X4 inst_6904 ( .ZN(net_17921), .A2(net_17751), .A1(net_17657) );
NAND2_X2 inst_9345 ( .ZN(net_20302), .A1(net_15245), .A2(net_8909) );
NAND2_X2 inst_8137 ( .ZN(net_18031), .A1(net_18013), .A2(net_17988) );
CLKBUF_X2 inst_22280 ( .A(net_21780), .Z(net_22152) );
NAND3_X2 inst_5723 ( .ZN(net_16130), .A2(net_15663), .A1(net_15592), .A3(net_14833) );
NOR2_X4 inst_2958 ( .A2(net_8748), .ZN(net_8064), .A1(net_5660) );
CLKBUF_X2 inst_22656 ( .A(net_22424), .Z(net_22528) );
XOR2_X2 inst_24 ( .B(net_21138), .A(net_16530), .Z(net_16528) );
OR2_X2 inst_1209 ( .ZN(net_3222), .A2(net_3221), .A1(net_944) );
INV_X4 inst_16832 ( .ZN(net_15833), .A(net_15452) );
NAND2_X2 inst_8190 ( .ZN(net_17897), .A2(net_17791), .A1(net_17689) );
OAI21_X2 inst_1611 ( .A(net_16359), .ZN(net_16113), .B1(net_15656), .B2(net_14761) );
NOR2_X2 inst_4469 ( .ZN(net_5927), .A1(net_4464), .A2(net_2835) );
NAND3_X2 inst_6779 ( .ZN(net_4504), .A1(net_4503), .A2(net_4502), .A3(net_1871) );
INV_X4 inst_12764 ( .ZN(net_17383), .A(net_17382) );
CLKBUF_X2 inst_22128 ( .A(net_21848), .Z(net_22000) );
AOI21_X2 inst_20914 ( .A(net_10956), .B2(net_10635), .ZN(net_7336), .B1(net_3659) );
CLKBUF_X2 inst_22804 ( .A(net_22675), .Z(net_22676) );
NAND2_X2 inst_8730 ( .ZN(net_16063), .A1(net_15924), .A2(net_15771) );
NAND2_X2 inst_8466 ( .ZN(net_17049), .A2(net_17048), .A1(net_16696) );
NAND3_X2 inst_5849 ( .ZN(net_15432), .A3(net_14325), .A2(net_13328), .A1(net_12587) );
INV_X4 inst_17005 ( .A(net_14027), .ZN(net_10536) );
OAI21_X2 inst_1663 ( .ZN(net_15755), .A(net_15411), .B2(net_15056), .B1(net_11431) );
CLKBUF_X2 inst_22461 ( .A(net_22332), .Z(net_22333) );
NOR3_X2 inst_2714 ( .ZN(net_13510), .A2(net_13509), .A3(net_12353), .A1(net_10866) );
INV_X4 inst_13223 ( .ZN(net_13623), .A(net_12765) );
NAND2_X4 inst_7099 ( .ZN(net_19400), .A1(net_13560), .A2(net_11869) );
AND2_X2 inst_21348 ( .ZN(net_2643), .A1(net_2642), .A2(net_1486) );
INV_X4 inst_13036 ( .A(net_16774), .ZN(net_16411) );
INV_X2 inst_19524 ( .ZN(net_4747), .A(net_1518) );
NAND2_X2 inst_7962 ( .ZN(net_18371), .A2(net_18319), .A1(net_17432) );
INV_X4 inst_15730 ( .ZN(net_12864), .A(net_9438) );
CLKBUF_X2 inst_21978 ( .A(net_21849), .Z(net_21850) );
INV_X4 inst_16029 ( .ZN(net_2163), .A(net_1632) );
INV_X4 inst_15420 ( .A(net_3710), .ZN(net_2596) );
NAND2_X2 inst_11285 ( .ZN(net_5312), .A1(net_3924), .A2(net_3844) );
NAND2_X2 inst_10713 ( .A1(net_9591), .ZN(net_5953), .A2(net_5952) );
INV_X4 inst_14928 ( .ZN(net_13472), .A(net_3555) );
INV_X4 inst_15088 ( .ZN(net_3643), .A(net_3256) );
INV_X2 inst_18929 ( .ZN(net_5882), .A(net_5881) );
INV_X4 inst_16228 ( .ZN(net_11426), .A(net_6635) );
AND2_X2 inst_21328 ( .ZN(net_5966), .A1(net_4770), .A2(net_2758) );
NAND3_X2 inst_6021 ( .A3(net_20734), .A1(net_20733), .ZN(net_19080), .A2(net_10635) );
SDFF_X2 inst_820 ( .Q(net_21233), .SI(net_17670), .SE(net_125), .CK(net_22241), .D(x6912) );
AND2_X2 inst_21286 ( .ZN(net_12713), .A1(net_12712), .A2(net_10856) );
XNOR2_X2 inst_157 ( .ZN(net_17983), .A(net_17858), .B(net_17690) );
OAI21_X4 inst_1441 ( .B2(net_20385), .B1(net_20384), .ZN(net_15811), .A(net_15810) );
NOR2_X4 inst_2929 ( .ZN(net_9332), .A1(net_7815), .A2(net_6354) );
NAND2_X1 inst_12154 ( .A2(net_8333), .ZN(net_8307), .A1(net_8306) );
NOR2_X2 inst_3443 ( .ZN(net_15032), .A2(net_13908), .A1(net_10892) );
INV_X16 inst_19743 ( .A(net_879), .ZN(net_875) );
CLKBUF_X2 inst_21927 ( .A(net_21696), .Z(net_21799) );
NAND3_X2 inst_6159 ( .A1(net_20079), .A3(net_19560), .ZN(net_13646), .A2(net_10567) );
NOR2_X2 inst_4287 ( .ZN(net_6047), .A2(net_5329), .A1(net_4052) );
NAND2_X2 inst_10986 ( .ZN(net_8096), .A2(net_3601), .A1(net_526) );
NAND4_X2 inst_5491 ( .ZN(net_12247), .A3(net_12246), .A2(net_8458), .A1(net_7188), .A4(net_5768) );
OAI21_X2 inst_2177 ( .B2(net_19327), .B1(net_9999), .ZN(net_8872), .A(net_8741) );
INV_X4 inst_16963 ( .ZN(net_8037), .A(net_2976) );
NAND2_X2 inst_9588 ( .ZN(net_12314), .A2(net_7461), .A1(net_6924) );
NAND2_X4 inst_7447 ( .A1(net_19964), .ZN(net_6488), .A2(net_3107) );
NAND2_X2 inst_8348 ( .ZN(net_17476), .A2(net_17321), .A1(net_17071) );
INV_X4 inst_17549 ( .ZN(net_1776), .A(net_154) );
NOR2_X2 inst_3410 ( .ZN(net_15726), .A2(net_15180), .A1(net_14069) );
NAND4_X2 inst_5339 ( .A2(net_20681), .A1(net_20680), .A3(net_20496), .ZN(net_19234), .A4(net_12617) );
NAND2_X2 inst_11506 ( .A1(net_20488), .ZN(net_4828), .A2(net_3053) );
INV_X4 inst_13478 ( .ZN(net_9609), .A(net_9608) );
INV_X4 inst_13216 ( .ZN(net_13637), .A(net_12810) );
INV_X4 inst_17227 ( .A(net_9581), .ZN(net_5735) );
XOR2_X2 inst_17 ( .B(net_21170), .Z(net_17020), .A(net_17019) );
CLKBUF_X2 inst_21539 ( .A(net_21410), .Z(net_21411) );
NAND2_X2 inst_10105 ( .ZN(net_11849), .A1(net_8485), .A2(net_6184) );
AOI21_X2 inst_20341 ( .B1(net_20336), .ZN(net_15765), .A(net_12164), .B2(net_2573) );
NAND2_X2 inst_7838 ( .ZN(net_18625), .A2(net_18605), .A1(net_615) );
XNOR2_X2 inst_249 ( .ZN(net_17314), .A(net_16988), .B(net_188) );
CLKBUF_X2 inst_22800 ( .A(net_22671), .Z(net_22672) );
OAI21_X2 inst_2234 ( .ZN(net_7764), .B2(net_7663), .A(net_6261), .B1(net_3704) );
INV_X8 inst_12407 ( .ZN(net_808), .A(net_598) );
NAND3_X2 inst_6251 ( .ZN(net_13011), .A3(net_13010), .A1(net_9717), .A2(net_7338) );
CLKBUF_X2 inst_22828 ( .A(net_22699), .Z(net_22700) );
AOI21_X2 inst_20291 ( .ZN(net_16191), .B1(net_15969), .B2(net_15868), .A(net_15577) );
INV_X2 inst_18879 ( .ZN(net_6194), .A(net_6193) );
INV_X4 inst_14509 ( .ZN(net_7846), .A(net_4824) );
NAND4_X4 inst_5204 ( .A3(net_18985), .A1(net_18984), .ZN(net_16571), .A4(net_16246), .A2(net_15661) );
OAI21_X4 inst_1480 ( .ZN(net_19622), .A(net_14029), .B2(net_11590), .B1(net_8828) );
INV_X2 inst_18905 ( .A(net_7989), .ZN(net_6057) );
INV_X4 inst_17461 ( .ZN(net_8502), .A(net_4718) );
NAND2_X2 inst_10676 ( .ZN(net_9714), .A1(net_6201), .A2(net_6200) );
INV_X4 inst_14121 ( .A(net_7939), .ZN(net_7541) );
INV_X4 inst_15305 ( .A(net_10989), .ZN(net_6363) );
INV_X2 inst_18856 ( .ZN(net_6339), .A(net_6338) );
INV_X4 inst_17334 ( .ZN(net_15372), .A(net_855) );
INV_X4 inst_15708 ( .A(net_2687), .ZN(net_1988) );
INV_X4 inst_17173 ( .ZN(net_940), .A(net_85) );
INV_X8 inst_12359 ( .A(net_20876), .ZN(net_412) );
NAND2_X4 inst_7409 ( .A1(net_19348), .ZN(net_4926), .A2(net_367) );
NAND3_X2 inst_6472 ( .ZN(net_11289), .A2(net_9553), .A3(net_6674), .A1(net_2823) );
NAND2_X2 inst_10504 ( .ZN(net_8274), .A2(net_6917), .A1(net_6896) );
INV_X2 inst_18450 ( .ZN(net_13488), .A(net_12462) );
INV_X4 inst_16704 ( .A(net_3713), .ZN(net_3322) );
XNOR2_X2 inst_664 ( .A(net_21181), .B(net_21117), .ZN(net_254) );
NAND2_X2 inst_11638 ( .ZN(net_2512), .A2(net_1667), .A1(net_85) );
INV_X4 inst_13977 ( .ZN(net_8602), .A(net_8560) );
NAND2_X2 inst_10486 ( .ZN(net_6937), .A2(net_6936), .A1(net_1663) );
INV_X4 inst_12485 ( .ZN(net_18734), .A(net_18675) );
INV_X4 inst_14262 ( .ZN(net_8098), .A(net_5732) );
NAND2_X2 inst_9911 ( .ZN(net_11459), .A2(net_9496), .A1(net_9324) );
CLKBUF_X2 inst_22643 ( .A(net_22514), .Z(net_22515) );
OAI21_X2 inst_1918 ( .A(net_14605), .ZN(net_13041), .B2(net_12934), .B1(net_6811) );
NAND2_X2 inst_9466 ( .ZN(net_13693), .A1(net_11485), .A2(net_11484) );
INV_X4 inst_14500 ( .ZN(net_13762), .A(net_4836) );
INV_X4 inst_17441 ( .ZN(net_8181), .A(net_5748) );
INV_X4 inst_16590 ( .ZN(net_19516), .A(net_1303) );
INV_X4 inst_15394 ( .A(net_4026), .ZN(net_3570) );
NOR2_X2 inst_4064 ( .ZN(net_7796), .A2(net_7795), .A1(net_60) );
NOR2_X2 inst_4427 ( .ZN(net_6095), .A1(net_5557), .A2(net_4949) );
INV_X4 inst_15806 ( .A(net_3347), .ZN(net_2571) );
INV_X4 inst_12543 ( .ZN(net_18395), .A(net_18330) );
CLKBUF_X2 inst_22050 ( .A(net_21921), .Z(net_21922) );
NOR2_X2 inst_4635 ( .ZN(net_3502), .A1(net_3501), .A2(net_1323) );
NOR2_X2 inst_3839 ( .ZN(net_9655), .A2(net_9654), .A1(net_6032) );
AOI21_X2 inst_20531 ( .ZN(net_14524), .B1(net_14515), .B2(net_11704), .A(net_11670) );
NAND2_X2 inst_7862 ( .ZN(net_18560), .A2(net_18522), .A1(net_18495) );
OAI211_X4 inst_2368 ( .C2(net_20880), .ZN(net_18072), .B(net_18047), .C1(net_16203), .A(net_14470) );
NOR3_X2 inst_2735 ( .ZN(net_12806), .A2(net_12805), .A3(net_12804), .A1(net_8262) );
NOR2_X4 inst_2934 ( .ZN(net_12525), .A2(net_5842), .A1(net_732) );
NOR3_X2 inst_2767 ( .ZN(net_9871), .A2(net_9870), .A3(net_4881), .A1(net_3018) );
OAI21_X4 inst_1370 ( .B1(net_20068), .ZN(net_17214), .A(net_16572), .B2(net_16571) );
OAI211_X2 inst_2512 ( .C2(net_20780), .B(net_13762), .ZN(net_12459), .C1(net_12216), .A(net_2534) );
INV_X4 inst_15805 ( .ZN(net_16030), .A(net_15694) );
NAND2_X2 inst_12093 ( .A2(net_20851), .ZN(net_763), .A1(net_102) );
NAND2_X2 inst_11948 ( .ZN(net_2829), .A2(net_1433), .A1(net_524) );
INV_X4 inst_17587 ( .ZN(net_13530), .A(net_10702) );
NAND2_X2 inst_11447 ( .A1(net_7661), .ZN(net_3272), .A2(net_2359) );
CLKBUF_X2 inst_22080 ( .A(net_21951), .Z(net_21952) );
INV_X2 inst_18884 ( .ZN(net_9719), .A(net_6171) );
INV_X4 inst_12568 ( .ZN(net_18308), .A(net_18202) );
NOR2_X2 inst_4124 ( .A2(net_8483), .ZN(net_7020), .A1(net_4107) );
INV_X4 inst_13078 ( .ZN(net_20140), .A(net_16131) );
INV_X4 inst_15886 ( .A(net_5289), .ZN(net_3710) );
CLKBUF_X2 inst_22386 ( .A(net_22257), .Z(net_22258) );
INV_X4 inst_14740 ( .ZN(net_8486), .A(net_2282) );
INV_X2 inst_19256 ( .A(net_4180), .ZN(net_3200) );
AOI21_X2 inst_20985 ( .ZN(net_18873), .A(net_15300), .B1(net_13686), .B2(net_6502) );
INV_X4 inst_17648 ( .ZN(net_2339), .A(net_508) );
INV_X4 inst_15837 ( .ZN(net_2537), .A(net_1800) );
NAND3_X2 inst_5672 ( .A3(net_19167), .A1(net_19166), .ZN(net_16373), .A2(net_14808) );
INV_X4 inst_17987 ( .A(net_21046), .ZN(net_354) );
NAND2_X2 inst_10273 ( .ZN(net_7969), .A1(net_7968), .A2(net_6216) );
AOI21_X2 inst_20392 ( .ZN(net_15462), .B1(net_14462), .B2(net_14457), .A(net_10082) );
NOR2_X2 inst_3348 ( .ZN(net_18028), .A2(net_18011), .A1(net_17283) );
NAND2_X4 inst_7700 ( .A1(net_20870), .A2(net_814), .ZN(net_802) );
INV_X4 inst_17993 ( .A(net_20950), .ZN(net_199) );
NAND2_X2 inst_7888 ( .ZN(net_18510), .A2(net_18427), .A1(net_17902) );
NOR2_X2 inst_4848 ( .ZN(net_2572), .A2(net_2328), .A1(net_1614) );
NAND2_X4 inst_7044 ( .A2(net_19740), .A1(net_19739), .ZN(net_17815) );
INV_X4 inst_15139 ( .A(net_3307), .ZN(net_3116) );
NAND2_X2 inst_11906 ( .ZN(net_1944), .A2(net_1789), .A1(net_1562) );
NOR2_X2 inst_4820 ( .ZN(net_3361), .A2(net_2991), .A1(net_2557) );
OAI21_X2 inst_1684 ( .ZN(net_15453), .A(net_15452), .B2(net_14382), .B1(net_10177) );
OAI21_X4 inst_1386 ( .A(net_20928), .B2(net_19476), .B1(net_19475), .ZN(net_19012) );
XNOR2_X2 inst_217 ( .A(net_17537), .ZN(net_17535), .B(net_17534) );
NOR2_X2 inst_4852 ( .ZN(net_6942), .A2(net_4037), .A1(net_2532) );
NOR2_X2 inst_4616 ( .ZN(net_6347), .A1(net_3682), .A2(net_3228) );
NAND2_X2 inst_9816 ( .ZN(net_9657), .A1(net_9656), .A2(net_6031) );
INV_X4 inst_15907 ( .ZN(net_11562), .A(net_8785) );
CLKBUF_X2 inst_22730 ( .A(net_21728), .Z(net_22602) );
OAI21_X2 inst_2213 ( .ZN(net_19409), .A(net_11612), .B2(net_5579), .B1(net_3597) );
CLKBUF_X2 inst_21866 ( .A(net_21737), .Z(net_21738) );
XNOR2_X2 inst_672 ( .A(net_21182), .B(net_21118), .ZN(net_147) );
OAI21_X4 inst_1471 ( .ZN(net_14834), .B2(net_13450), .B1(net_8887), .A(net_278) );
INV_X4 inst_15393 ( .A(net_3367), .ZN(net_2545) );
INV_X4 inst_17977 ( .A(net_21017), .ZN(net_576) );
CLKBUF_X2 inst_22263 ( .A(net_21916), .Z(net_22135) );
NAND2_X2 inst_9610 ( .ZN(net_20808), .A1(net_10714), .A2(net_8452) );
NOR2_X2 inst_3826 ( .ZN(net_9753), .A2(net_8906), .A1(net_8199) );
AOI211_X2 inst_21014 ( .ZN(net_15680), .C1(net_15666), .C2(net_14934), .A(net_8320), .B(net_6650) );
NAND2_X4 inst_7523 ( .ZN(net_3970), .A1(net_2314), .A2(net_2058) );
NAND3_X2 inst_6471 ( .ZN(net_11291), .A2(net_11290), .A3(net_9885), .A1(net_5851) );
DFF_X1 inst_19894 ( .D(net_16939), .CK(net_21591), .Q(x636) );
OAI21_X2 inst_1525 ( .A(net_20912), .ZN(net_18046), .B2(net_15934), .B1(net_12575) );
NOR2_X4 inst_3230 ( .ZN(net_3554), .A1(net_3491), .A2(net_1738) );
NAND2_X2 inst_11820 ( .ZN(net_1996), .A1(net_1922), .A2(net_63) );
NAND2_X2 inst_9538 ( .ZN(net_13707), .A1(net_11767), .A2(net_10636) );
CLKBUF_X2 inst_21399 ( .A(net_21270), .Z(net_21271) );
NOR2_X4 inst_3281 ( .ZN(net_3093), .A2(net_1697), .A1(net_1054) );
SDFF_X2 inst_703 ( .Q(net_20959), .SE(net_18862), .SI(net_18836), .D(net_436), .CK(net_22269) );
NAND2_X2 inst_11125 ( .A1(net_9310), .ZN(net_4285), .A2(net_2290) );
AOI21_X2 inst_20654 ( .ZN(net_13038), .B2(net_9752), .B1(net_7703), .A(net_339) );
OAI211_X2 inst_2546 ( .A(net_20483), .ZN(net_10823), .B(net_5342), .C2(net_4635), .C1(net_2710) );
NAND2_X2 inst_9474 ( .A2(net_11560), .ZN(net_11463), .A1(net_8979) );
NAND2_X4 inst_7177 ( .ZN(net_10896), .A1(net_9540), .A2(net_6625) );
NOR2_X2 inst_4693 ( .A1(net_20566), .ZN(net_4159), .A2(net_2054) );
NAND2_X2 inst_9882 ( .ZN(net_9433), .A1(net_7394), .A2(net_6025) );
NAND2_X2 inst_11112 ( .ZN(net_12442), .A2(net_3989), .A1(net_532) );
AOI21_X2 inst_20764 ( .ZN(net_10860), .B2(net_7123), .B1(net_7024), .A(net_607) );
INV_X4 inst_12504 ( .A(net_18615), .ZN(net_18614) );
NAND2_X2 inst_10449 ( .ZN(net_7063), .A1(net_7062), .A2(net_3727) );
INV_X4 inst_15737 ( .ZN(net_4032), .A(net_3446) );
INV_X4 inst_14289 ( .ZN(net_5600), .A(net_5599) );
INV_X4 inst_14786 ( .ZN(net_13968), .A(net_4017) );
NAND3_X2 inst_6539 ( .ZN(net_10576), .A3(net_10575), .A2(net_9035), .A1(net_7416) );
OR2_X4 inst_1067 ( .ZN(net_16501), .A1(net_16237), .A2(net_16163) );
INV_X4 inst_12966 ( .ZN(net_16666), .A(net_16522) );
AOI21_X2 inst_20865 ( .A(net_15300), .ZN(net_8666), .B1(net_8665), .B2(net_4106) );
NAND2_X4 inst_7411 ( .A1(net_19825), .ZN(net_9041), .A2(net_3151) );
NOR2_X2 inst_4787 ( .ZN(net_6053), .A2(net_2829), .A1(net_1376) );
NAND2_X2 inst_11970 ( .ZN(net_5557), .A1(net_1357), .A2(net_117) );
CLKBUF_X2 inst_21382 ( .A(x7698), .Z(net_21254) );
NAND2_X2 inst_9735 ( .ZN(net_13862), .A1(net_9972), .A2(net_9403) );
NAND2_X2 inst_9231 ( .ZN(net_19907), .A2(net_10412), .A1(net_9453) );
OAI21_X2 inst_1824 ( .A(net_14179), .ZN(net_14149), .B2(net_10517), .B1(net_10239) );
INV_X2 inst_19407 ( .ZN(net_1983), .A(net_1982) );
OR2_X2 inst_1214 ( .A1(net_6626), .ZN(net_5360), .A2(net_2978) );
INV_X2 inst_18580 ( .ZN(net_10318), .A(net_10317) );
NAND2_X2 inst_8121 ( .A2(net_18067), .ZN(net_18061), .A1(net_15401) );
INV_X4 inst_15151 ( .ZN(net_3480), .A(net_2318) );
INV_X4 inst_16197 ( .ZN(net_3053), .A(net_1273) );
OAI21_X4 inst_1417 ( .A(net_20944), .ZN(net_20141), .B2(net_19922), .B1(net_19921) );
INV_X2 inst_18510 ( .ZN(net_11621), .A(net_11620) );
NAND2_X2 inst_11103 ( .A1(net_20859), .ZN(net_12041), .A2(net_4341) );
CLKBUF_X2 inst_21534 ( .A(net_21405), .Z(net_21406) );
NAND2_X2 inst_11887 ( .ZN(net_2091), .A2(net_1751), .A1(net_61) );
CLKBUF_X2 inst_22262 ( .A(net_21394), .Z(net_22134) );
INV_X2 inst_19430 ( .A(net_5866), .ZN(net_3640) );
INV_X2 inst_19252 ( .ZN(net_3232), .A(net_3231) );
AOI22_X2 inst_19995 ( .ZN(net_14549), .A1(net_14548), .A2(net_11862), .B1(net_7849), .B2(net_2890) );
CLKBUF_X2 inst_22542 ( .A(net_21431), .Z(net_22414) );
INV_X4 inst_17803 ( .A(net_602), .ZN(net_257) );
INV_X1 inst_19752 ( .A(net_12031), .ZN(net_9796) );
NOR2_X4 inst_3335 ( .A1(net_20005), .ZN(net_836), .A2(net_301) );
NOR2_X4 inst_3073 ( .ZN(net_5919), .A1(net_4749), .A2(net_86) );
OAI21_X2 inst_1980 ( .ZN(net_12115), .A(net_11654), .B1(net_7479), .B2(net_6987) );
NAND2_X2 inst_10488 ( .A2(net_9663), .ZN(net_6933), .A1(net_6399) );
INV_X4 inst_17922 ( .A(net_21238), .ZN(net_56) );
INV_X4 inst_16638 ( .ZN(net_8326), .A(net_7432) );
INV_X4 inst_16792 ( .ZN(net_14793), .A(net_1012) );
NAND3_X2 inst_5868 ( .ZN(net_15315), .A2(net_15314), .A3(net_13039), .A1(net_12103) );
AOI21_X2 inst_20389 ( .ZN(net_15467), .B2(net_14588), .A(net_10979), .B1(net_10683) );
NOR2_X4 inst_2885 ( .ZN(net_9689), .A1(net_9688), .A2(net_6575) );
NAND2_X2 inst_9325 ( .ZN(net_12321), .A1(net_12320), .A2(net_9058) );
NOR2_X2 inst_4795 ( .A1(net_6520), .ZN(net_4722), .A2(net_2020) );
NOR3_X4 inst_2632 ( .ZN(net_13892), .A3(net_11350), .A2(net_10625), .A1(net_8920) );
OAI21_X2 inst_2221 ( .B1(net_13556), .ZN(net_8512), .B2(net_8511), .A(net_7819) );
NAND2_X2 inst_10446 ( .A2(net_8949), .ZN(net_7178), .A1(net_5881) );
OAI21_X2 inst_2082 ( .A(net_14104), .ZN(net_10501), .B1(net_9855), .B2(net_5960) );
INV_X4 inst_12469 ( .ZN(net_18772), .A(net_18771) );
INV_X4 inst_15028 ( .ZN(net_9498), .A(net_3369) );
INV_X4 inst_12907 ( .ZN(net_17046), .A(net_16899) );
INV_X4 inst_15299 ( .ZN(net_5422), .A(net_2693) );
INV_X16 inst_19737 ( .A(net_20868), .ZN(net_504) );
CLKBUF_X2 inst_22048 ( .A(net_21449), .Z(net_21920) );
INV_X4 inst_17197 ( .ZN(net_1028), .A(net_710) );
INV_X2 inst_19630 ( .A(net_20865), .ZN(net_30) );
INV_X4 inst_16204 ( .ZN(net_10405), .A(net_9735) );
INV_X4 inst_13004 ( .A(net_16577), .ZN(net_16543) );
SDFF_X2 inst_692 ( .Q(net_20892), .SI(net_18867), .SE(net_18864), .D(net_654), .CK(net_22048) );
NAND3_X2 inst_6800 ( .ZN(net_5899), .A3(net_3436), .A2(net_2744), .A1(net_2018) );
NAND2_X4 inst_6897 ( .ZN(net_18006), .A2(net_17953), .A1(net_17927) );
INV_X4 inst_14819 ( .A(net_5401), .ZN(net_4932) );
OAI21_X2 inst_1517 ( .ZN(net_18464), .A(net_18421), .B1(net_18420), .B2(net_18419) );
INV_X2 inst_19398 ( .A(net_2913), .ZN(net_2043) );
INV_X4 inst_17245 ( .ZN(net_1584), .A(net_954) );
NAND4_X2 inst_5480 ( .ZN(net_12789), .A1(net_12788), .A4(net_12787), .A2(net_11728), .A3(net_11727) );
XNOR2_X2 inst_70 ( .ZN(net_18757), .A(net_18695), .B(net_17081) );
NAND2_X2 inst_10529 ( .ZN(net_6831), .A1(net_6830), .A2(net_6829) );
CLKBUF_X2 inst_22704 ( .A(net_22575), .Z(net_22576) );
NAND2_X4 inst_6915 ( .A2(net_20236), .A1(net_20235), .ZN(net_17790) );
NAND2_X4 inst_7672 ( .ZN(net_845), .A1(net_174), .A2(net_150) );
NAND2_X4 inst_7587 ( .A1(net_19108), .ZN(net_3131), .A2(net_1533) );
INV_X4 inst_15662 ( .A(net_16011), .ZN(net_2072) );
INV_X4 inst_14161 ( .ZN(net_10139), .A(net_6017) );
INV_X4 inst_15987 ( .ZN(net_2720), .A(net_2232) );
CLKBUF_X2 inst_21840 ( .A(net_21711), .Z(net_21712) );
NAND3_X2 inst_6028 ( .A3(net_19818), .ZN(net_19770), .A1(net_13770), .A2(net_7534) );
NOR2_X2 inst_3768 ( .ZN(net_14289), .A2(net_11792), .A1(net_60) );
INV_X4 inst_16757 ( .ZN(net_19759), .A(net_1038) );
NOR2_X2 inst_4207 ( .ZN(net_7945), .A1(net_6669), .A2(net_3752) );
NAND2_X2 inst_9058 ( .ZN(net_13995), .A1(net_13355), .A2(net_11994) );
NAND2_X2 inst_11308 ( .A1(net_5009), .ZN(net_4441), .A2(net_3312) );
NAND3_X2 inst_6218 ( .ZN(net_13253), .A3(net_10058), .A2(net_9659), .A1(net_9070) );
INV_X2 inst_18550 ( .ZN(net_19996), .A(net_10932) );
CLKBUF_X2 inst_22816 ( .A(net_22687), .Z(net_22688) );
INV_X4 inst_13306 ( .ZN(net_11852), .A(net_10491) );
NOR2_X4 inst_2848 ( .A2(net_20343), .A1(net_20342), .ZN(net_18989) );
INV_X4 inst_12686 ( .ZN(net_17704), .A(net_17703) );
INV_X4 inst_15181 ( .ZN(net_4362), .A(net_2982) );
INV_X2 inst_18922 ( .ZN(net_5923), .A(net_5922) );
CLKBUF_X2 inst_22400 ( .A(net_21353), .Z(net_22272) );
CLKBUF_X2 inst_21742 ( .A(net_21613), .Z(net_21614) );
INV_X4 inst_13866 ( .ZN(net_14209), .A(net_9329) );
INV_X4 inst_16504 ( .ZN(net_19314), .A(net_3505) );
NOR2_X2 inst_3593 ( .ZN(net_12604), .A2(net_12603), .A1(net_10709) );
NAND2_X2 inst_8529 ( .A1(net_20768), .A2(net_17244), .ZN(net_16869) );
NAND2_X4 inst_7509 ( .ZN(net_4091), .A2(net_2168), .A1(net_856) );
NOR2_X4 inst_3176 ( .ZN(net_5613), .A1(net_3138), .A2(net_1848) );
INV_X4 inst_15985 ( .ZN(net_3239), .A(net_1679) );
AOI21_X2 inst_20744 ( .A(net_14628), .ZN(net_11403), .B2(net_9085), .B1(net_5721) );
INV_X4 inst_14830 ( .ZN(net_6872), .A(net_3881) );
INV_X4 inst_12655 ( .ZN(net_17832), .A(net_17831) );
INV_X4 inst_13889 ( .ZN(net_19715), .A(net_7318) );
AOI21_X2 inst_20811 ( .A(net_14628), .ZN(net_10132), .B1(net_10131), .B2(net_6003) );
INV_X4 inst_17358 ( .ZN(net_7917), .A(net_1961) );
INV_X4 inst_13730 ( .A(net_7774), .ZN(net_7771) );
NAND2_X2 inst_10821 ( .ZN(net_11830), .A1(net_7414), .A2(net_5419) );
CLKBUF_X2 inst_22847 ( .A(net_22718), .Z(net_22719) );
OR2_X2 inst_1150 ( .ZN(net_9844), .A1(net_9843), .A2(net_9842) );
INV_X4 inst_17305 ( .ZN(net_6877), .A(net_1020) );
NAND2_X4 inst_7685 ( .ZN(net_1602), .A1(net_1333), .A2(net_148) );
NOR2_X2 inst_4914 ( .ZN(net_4331), .A1(net_1911), .A2(net_1548) );
INV_X4 inst_18086 ( .A(net_20890), .ZN(net_120) );
INV_X4 inst_17789 ( .A(net_4268), .ZN(net_718) );
NAND2_X2 inst_11020 ( .ZN(net_11743), .A1(net_4795), .A2(net_3541) );
NAND2_X2 inst_11355 ( .A2(net_3673), .ZN(net_3619), .A1(net_1935) );
AOI21_X4 inst_20209 ( .ZN(net_19586), .B1(net_19533), .B2(net_13709), .A(net_12728) );
INV_X4 inst_16815 ( .ZN(net_1001), .A(net_1000) );
NAND2_X2 inst_11770 ( .A1(net_14027), .ZN(net_2064), .A2(net_2063) );
NAND2_X2 inst_8715 ( .A1(net_16644), .ZN(net_16207), .A2(net_15997) );
NOR2_X2 inst_4535 ( .A1(net_9396), .ZN(net_5089), .A2(net_2134) );
INV_X4 inst_14810 ( .ZN(net_3965), .A(net_3964) );
NOR2_X2 inst_4499 ( .A2(net_20467), .ZN(net_6573), .A1(net_1808) );
INV_X4 inst_12852 ( .ZN(net_17358), .A(net_17232) );
NAND3_X1 inst_6825 ( .A1(net_12551), .ZN(net_8701), .A2(net_8700), .A3(net_8050) );
NAND2_X2 inst_10979 ( .ZN(net_4965), .A2(net_4801), .A1(net_3096) );
INV_X1 inst_19747 ( .A(net_17353), .ZN(net_17071) );
NAND2_X2 inst_8704 ( .A1(net_16743), .ZN(net_16307), .A2(net_16137) );
INV_X2 inst_19637 ( .A(net_19426), .ZN(net_19425) );
INV_X4 inst_12783 ( .A(net_17493), .ZN(net_17302) );
NAND4_X2 inst_5508 ( .A2(net_11808), .ZN(net_11242), .A3(net_10348), .A4(net_6139), .A1(net_2729) );
INV_X4 inst_12661 ( .ZN(net_17812), .A(net_17811) );
AOI21_X2 inst_20334 ( .ZN(net_19659), .A(net_15880), .B1(net_14816), .B2(net_12143) );
NAND2_X2 inst_8611 ( .ZN(net_19866), .A2(net_16780), .A1(net_9236) );
XNOR2_X2 inst_658 ( .B(net_437), .ZN(net_347), .A(net_346) );
NAND3_X2 inst_6190 ( .ZN(net_13336), .A3(net_13335), .A2(net_11269), .A1(net_2390) );
NAND2_X2 inst_7779 ( .ZN(net_18729), .A1(net_18704), .A2(net_18691) );
INV_X8 inst_12192 ( .ZN(net_16465), .A(net_16341) );
INV_X4 inst_17728 ( .ZN(net_621), .A(net_61) );
NOR2_X2 inst_4520 ( .A2(net_7669), .A1(net_4838), .ZN(net_4134) );
INV_X2 inst_19720 ( .A(net_20785), .ZN(net_20783) );
NAND2_X4 inst_7227 ( .ZN(net_10240), .A2(net_6968), .A1(net_3586) );
INV_X2 inst_19564 ( .ZN(net_1394), .A(net_1261) );
INV_X4 inst_15090 ( .ZN(net_14605), .A(net_3251) );
NAND2_X2 inst_9626 ( .ZN(net_20329), .A1(net_11691), .A2(net_7339) );
INV_X2 inst_19426 ( .A(net_10398), .ZN(net_1811) );
NAND2_X2 inst_11391 ( .ZN(net_8088), .A2(net_2551), .A1(net_2079) );
INV_X4 inst_13581 ( .ZN(net_10767), .A(net_9043) );
OAI21_X2 inst_2128 ( .ZN(net_20687), .A(net_10000), .B1(net_9999), .B2(net_5254) );
AOI21_X2 inst_20965 ( .ZN(net_5306), .A(net_5305), .B1(net_5289), .B2(net_5269) );
CLKBUF_X2 inst_22060 ( .A(net_21297), .Z(net_21932) );
CLKBUF_X2 inst_22378 ( .A(net_22249), .Z(net_22250) );
NAND2_X2 inst_10452 ( .ZN(net_7042), .A2(net_7041), .A1(net_6406) );
NAND2_X4 inst_7384 ( .ZN(net_5339), .A1(net_4242), .A2(net_3426) );
INV_X4 inst_14472 ( .ZN(net_4899), .A(net_4898) );
NAND2_X2 inst_10086 ( .ZN(net_13150), .A1(net_8629), .A2(net_7845) );
NAND2_X2 inst_9887 ( .ZN(net_9420), .A1(net_6736), .A2(net_5882) );
INV_X4 inst_18066 ( .A(net_21171), .ZN(net_595) );
NAND2_X2 inst_11385 ( .ZN(net_8567), .A2(net_3233), .A1(net_573) );
NAND2_X2 inst_8289 ( .A1(net_20206), .ZN(net_17619), .A2(net_17618) );
NAND2_X2 inst_9313 ( .ZN(net_19979), .A1(net_14241), .A2(net_9019) );
NAND2_X2 inst_10833 ( .A1(net_5714), .ZN(net_5484), .A2(net_5483) );
NOR2_X2 inst_4455 ( .ZN(net_4676), .A2(net_4675), .A1(net_2067) );
NAND2_X2 inst_11402 ( .ZN(net_5079), .A2(net_2287), .A1(net_703) );
NAND2_X2 inst_7911 ( .ZN(net_18463), .A1(net_18418), .A2(net_18368) );
INV_X4 inst_17236 ( .ZN(net_1155), .A(net_228) );
NAND2_X2 inst_7907 ( .ZN(net_18471), .A2(net_18394), .A1(net_18329) );
SDFF_X2 inst_929 ( .Q(net_21228), .D(net_16503), .SE(net_263), .CK(net_21633), .SI(x7088) );
OAI21_X4 inst_1397 ( .B2(net_19691), .B1(net_19690), .ZN(net_16261), .A(net_16260) );
AOI21_X4 inst_20143 ( .ZN(net_15853), .B2(net_15307), .B1(net_15107), .A(net_14307) );
AOI21_X2 inst_20678 ( .ZN(net_12452), .B2(net_10958), .B1(net_6736), .A(net_4891) );
INV_X2 inst_19456 ( .ZN(net_2054), .A(net_1078) );
INV_X4 inst_17327 ( .A(net_9131), .ZN(net_571) );
NOR2_X4 inst_3303 ( .ZN(net_1453), .A1(net_1176), .A2(net_1175) );
INV_X4 inst_13115 ( .ZN(net_15609), .A(net_15339) );
NAND3_X2 inst_6181 ( .ZN(net_13499), .A3(net_9437), .A1(net_9187), .A2(net_8841) );
INV_X2 inst_19166 ( .ZN(net_3869), .A(net_3868) );
INV_X4 inst_12938 ( .A(net_17487), .ZN(net_17371) );
NAND3_X2 inst_6478 ( .ZN(net_11275), .A3(net_10570), .A2(net_8394), .A1(net_7784) );
OAI21_X2 inst_1938 ( .ZN(net_12913), .B1(net_10960), .A(net_9301), .B2(net_6622) );
NAND2_X2 inst_11870 ( .A1(net_20868), .ZN(net_1639), .A2(net_1162) );
NAND2_X2 inst_9435 ( .A1(net_19465), .ZN(net_11590), .A2(net_11589) );
NAND2_X4 inst_6888 ( .A2(net_19342), .A1(net_19341), .ZN(net_18170) );
INV_X4 inst_16020 ( .ZN(net_2861), .A(net_1643) );
INV_X2 inst_19224 ( .ZN(net_8958), .A(net_3441) );
OAI21_X2 inst_2095 ( .A(net_14563), .ZN(net_10121), .B2(net_5973), .B1(net_4746) );
INV_X4 inst_15659 ( .ZN(net_2715), .A(net_2561) );
INV_X2 inst_18848 ( .A(net_11794), .ZN(net_6650) );
AOI211_X2 inst_21000 ( .ZN(net_15937), .C1(net_15936), .B(net_15253), .C2(net_15173), .A(net_14416) );
INV_X2 inst_19193 ( .ZN(net_3639), .A(net_3638) );
NAND3_X2 inst_5794 ( .ZN(net_15730), .A3(net_15067), .A2(net_10870), .A1(net_6352) );
INV_X4 inst_14103 ( .ZN(net_9777), .A(net_6175) );
NAND2_X2 inst_8896 ( .ZN(net_15106), .A2(net_13889), .A1(net_750) );
NAND3_X2 inst_5652 ( .ZN(net_16551), .A3(net_16407), .A2(net_16087), .A1(net_11011) );
NAND2_X2 inst_8262 ( .ZN(net_19294), .A2(net_17681), .A1(net_101) );
AOI21_X2 inst_20898 ( .ZN(net_7728), .B2(net_7727), .A(net_4863), .B1(net_4391) );
INV_X2 inst_19642 ( .A(net_19438), .ZN(net_19437) );
NAND3_X4 inst_5631 ( .A1(net_19278), .ZN(net_3767), .A2(net_2712), .A3(net_2050) );
XNOR2_X1 inst_683 ( .B(net_21143), .ZN(net_17528), .A(net_17527) );
NAND2_X2 inst_11813 ( .ZN(net_3038), .A2(net_1042), .A1(net_131) );
INV_X4 inst_17144 ( .ZN(net_15020), .A(net_12916) );
NAND2_X2 inst_9094 ( .ZN(net_13786), .A1(net_13785), .A2(net_11621) );
NAND2_X2 inst_9411 ( .A2(net_14844), .ZN(net_11658), .A1(net_8359) );
NAND2_X2 inst_8720 ( .A1(net_20920), .ZN(net_16171), .A2(net_15922) );
INV_X4 inst_17418 ( .ZN(net_4099), .A(net_2746) );
NAND2_X2 inst_12103 ( .ZN(net_472), .A2(net_189), .A1(net_133) );
NAND3_X2 inst_5893 ( .A2(net_19894), .A1(net_19893), .ZN(net_15201), .A3(net_14037) );
NOR2_X2 inst_3881 ( .ZN(net_19070), .A1(net_14962), .A2(net_9314) );
INV_X2 inst_18730 ( .ZN(net_8046), .A(net_8045) );
NOR2_X2 inst_4778 ( .ZN(net_11255), .A2(net_2899), .A1(net_1937) );
INV_X4 inst_14580 ( .ZN(net_4518), .A(net_4517) );
INV_X4 inst_17884 ( .ZN(net_333), .A(net_76) );
NAND2_X4 inst_7663 ( .A1(net_20868), .ZN(net_2170), .A2(net_938) );
NAND4_X2 inst_5325 ( .ZN(net_15724), .A4(net_14967), .A1(net_14068), .A2(net_13174), .A3(net_8784) );
NOR2_X2 inst_4576 ( .ZN(net_5254), .A1(net_4726), .A2(net_2839) );
SDFF_X2 inst_747 ( .Q(net_20874), .SE(net_18581), .SI(net_18540), .D(net_11892), .CK(net_21913) );
INV_X4 inst_15493 ( .ZN(net_11318), .A(net_9510) );
CLKBUF_X2 inst_21687 ( .A(net_21558), .Z(net_21559) );
NAND3_X2 inst_6685 ( .ZN(net_7713), .A2(net_7712), .A3(net_7711), .A1(net_2949) );
NAND2_X2 inst_9070 ( .ZN(net_13977), .A2(net_12204), .A1(net_5682) );
NOR2_X2 inst_3806 ( .A1(net_10968), .ZN(net_9840), .A2(net_2938) );
INV_X2 inst_18594 ( .ZN(net_10127), .A(net_10126) );
NOR2_X2 inst_4486 ( .ZN(net_4317), .A2(net_3135), .A1(net_810) );
INV_X4 inst_15964 ( .ZN(net_10829), .A(net_9894) );
INV_X4 inst_12893 ( .A(net_17022), .ZN(net_16806) );
INV_X4 inst_17747 ( .ZN(net_367), .A(net_225) );
NAND2_X2 inst_11362 ( .ZN(net_5896), .A2(net_1997), .A1(net_338) );
AOI21_X2 inst_20536 ( .ZN(net_14494), .B2(net_11525), .A(net_11302), .B1(net_10031) );
INV_X4 inst_14946 ( .ZN(net_6133), .A(net_3517) );
CLKBUF_X2 inst_22305 ( .A(net_21559), .Z(net_22177) );
NOR3_X2 inst_2775 ( .A2(net_14612), .A3(net_10945), .ZN(net_7773), .A1(net_7772) );
NAND3_X4 inst_5589 ( .ZN(net_18881), .A2(net_13593), .A1(net_12718), .A3(net_12550) );
INV_X4 inst_15324 ( .ZN(net_4959), .A(net_1971) );
INV_X2 inst_19040 ( .ZN(net_8011), .A(net_6641) );
INV_X8 inst_12334 ( .ZN(net_1990), .A(net_954) );
XNOR2_X2 inst_305 ( .B(net_21131), .ZN(net_17095), .A(net_17092) );
NAND3_X2 inst_6795 ( .ZN(net_19662), .A1(net_3457), .A3(net_3456), .A2(net_2160) );
AOI21_X4 inst_20166 ( .B1(net_19957), .ZN(net_15633), .A(net_12862), .B2(net_1046) );
INV_X4 inst_13516 ( .ZN(net_10899), .A(net_9395) );
OAI21_X2 inst_1595 ( .B1(net_21220), .ZN(net_16213), .B2(net_15903), .A(net_15797) );
NAND2_X2 inst_7881 ( .ZN(net_18522), .A2(net_18491), .A1(net_17872) );
NAND3_X2 inst_5651 ( .ZN(net_16704), .A3(net_16433), .A2(net_16250), .A1(net_9556) );
NAND2_X2 inst_7867 ( .ZN(net_18553), .A2(net_18511), .A1(net_18483) );
INV_X4 inst_15922 ( .ZN(net_13418), .A(net_4113) );
NAND2_X2 inst_10926 ( .ZN(net_7935), .A1(net_5459), .A2(net_3779) );
INV_X4 inst_13578 ( .ZN(net_9108), .A(net_9107) );
INV_X8 inst_12319 ( .ZN(net_967), .A(net_163) );
NAND2_X2 inst_8079 ( .ZN(net_18152), .A2(net_18086), .A1(net_16584) );
NAND3_X2 inst_6585 ( .ZN(net_10430), .A2(net_10429), .A3(net_10428), .A1(net_3835) );
INV_X4 inst_13069 ( .ZN(net_16293), .A(net_16222) );
INV_X4 inst_15595 ( .ZN(net_3017), .A(net_2237) );
NAND2_X2 inst_7774 ( .ZN(net_18736), .A2(net_18701), .A1(net_16992) );
SDFF_X2 inst_963 ( .QN(net_21098), .D(net_719), .SE(net_263), .CK(net_22597), .SI(x1425) );
INV_X4 inst_17986 ( .A(net_21185), .ZN(net_95) );
INV_X4 inst_16787 ( .ZN(net_1015), .A(net_238) );
AOI21_X2 inst_20467 ( .ZN(net_14998), .B1(net_13418), .B2(net_13000), .A(net_8900) );
OAI21_X2 inst_1614 ( .ZN(net_16103), .A(net_15847), .B2(net_12908), .B1(net_8264) );
CLKBUF_X2 inst_22361 ( .A(net_22232), .Z(net_22233) );
OAI21_X4 inst_1502 ( .ZN(net_19624), .B1(net_10608), .A(net_7402), .B2(net_1810) );
CLKBUF_X2 inst_21433 ( .A(net_21304), .Z(net_21305) );
NAND4_X2 inst_5436 ( .ZN(net_20268), .A4(net_13920), .A3(net_12480), .A2(net_10259), .A1(net_7951) );
NAND3_X2 inst_6115 ( .ZN(net_13870), .A3(net_13099), .A1(net_11455), .A2(net_8769) );
CLKBUF_X2 inst_21860 ( .A(net_21563), .Z(net_21732) );
NOR2_X2 inst_4091 ( .ZN(net_7254), .A1(net_7253), .A2(net_7252) );
INV_X4 inst_16732 ( .ZN(net_2285), .A(net_953) );
NAND2_X4 inst_7602 ( .ZN(net_2568), .A1(net_2283), .A2(net_1159) );
NAND2_X4 inst_6989 ( .A2(net_19105), .A1(net_19104), .ZN(net_17894) );
NAND3_X2 inst_6807 ( .A1(net_7439), .ZN(net_3046), .A3(net_3045), .A2(net_703) );
INV_X4 inst_15854 ( .ZN(net_2504), .A(net_1816) );
OAI21_X2 inst_1568 ( .B2(net_19467), .B1(net_19466), .ZN(net_16407), .A(net_16359) );
NAND2_X2 inst_11439 ( .A2(net_10819), .ZN(net_3320), .A1(net_1750) );
CLKBUF_X2 inst_21944 ( .A(net_21815), .Z(net_21816) );
NAND3_X2 inst_6177 ( .ZN(net_13541), .A3(net_12960), .A1(net_8472), .A2(net_3064) );
NAND2_X2 inst_8487 ( .A1(net_17767), .A2(net_17371), .ZN(net_16972) );
NOR2_X2 inst_3366 ( .A1(net_21138), .ZN(net_20104), .A2(net_16864) );
SDFF_X2 inst_873 ( .Q(net_21119), .SI(net_17035), .SE(net_945), .CK(net_21543), .D(x4416) );
NAND2_X2 inst_9258 ( .A1(net_15833), .ZN(net_12642), .A2(net_12641) );
INV_X8 inst_12223 ( .A(net_6418), .ZN(net_6250) );
NAND3_X2 inst_6454 ( .ZN(net_11719), .A3(net_11718), .A1(net_9511), .A2(net_5105) );
INV_X4 inst_13439 ( .ZN(net_12974), .A(net_9814) );
NAND2_X2 inst_10022 ( .A2(net_9055), .ZN(net_8763), .A1(net_8762) );
NAND2_X2 inst_10164 ( .ZN(net_11865), .A1(net_8246), .A2(net_8245) );
INV_X4 inst_16614 ( .A(net_4990), .ZN(net_1657) );
NAND2_X2 inst_8563 ( .A1(net_21116), .ZN(net_20453), .A2(net_16562) );
NOR2_X2 inst_3767 ( .ZN(net_10301), .A1(net_10300), .A2(net_5532) );
NAND2_X2 inst_10282 ( .ZN(net_19156), .A2(net_11315), .A1(net_3828) );
CLKBUF_X2 inst_22440 ( .A(net_22311), .Z(net_22312) );
NAND2_X2 inst_8839 ( .ZN(net_15470), .A2(net_14765), .A1(net_13074) );
DFF_X1 inst_19888 ( .D(net_16966), .CK(net_22354), .Q(x763) );
NOR2_X2 inst_4431 ( .ZN(net_4894), .A1(net_4037), .A2(net_3490) );
NAND2_X2 inst_8679 ( .A2(net_16762), .ZN(net_16454), .A1(net_16447) );
NOR2_X2 inst_3371 ( .ZN(net_16693), .A2(net_16656), .A1(net_9256) );
NOR2_X4 inst_3052 ( .ZN(net_8044), .A1(net_4405), .A2(net_168) );
INV_X4 inst_15920 ( .ZN(net_6736), .A(net_4952) );
NAND2_X4 inst_6982 ( .ZN(net_17578), .A1(net_16913), .A2(net_16723) );
INV_X4 inst_17210 ( .A(net_6207), .ZN(net_3368) );
INV_X2 inst_19611 ( .A(net_21230), .ZN(net_50) );
INV_X4 inst_16942 ( .ZN(net_10082), .A(net_333) );
NOR2_X4 inst_2907 ( .ZN(net_8825), .A2(net_8824), .A1(net_8148) );
INV_X4 inst_13548 ( .ZN(net_9175), .A(net_9174) );
NOR2_X2 inst_4072 ( .ZN(net_18978), .A2(net_5210), .A1(net_4609) );
NAND3_X2 inst_5901 ( .ZN(net_15146), .A3(net_13402), .A2(net_10399), .A1(net_5744) );
NOR2_X4 inst_3000 ( .ZN(net_9361), .A1(net_5909), .A2(net_5877) );
OR2_X2 inst_1163 ( .ZN(net_20242), .A1(net_13076), .A2(net_8975) );
NAND2_X2 inst_9668 ( .ZN(net_19697), .A2(net_12286), .A1(net_12033) );
CLKBUF_X2 inst_22558 ( .A(net_22429), .Z(net_22430) );
NAND2_X2 inst_10641 ( .ZN(net_20406), .A2(net_4050), .A1(net_2556) );
AOI211_X2 inst_21048 ( .ZN(net_12857), .C1(net_9374), .B(net_9372), .C2(net_5327), .A(net_5144) );
NAND2_X2 inst_8282 ( .ZN(net_17626), .A1(net_17625), .A2(net_17611) );
INV_X2 inst_18399 ( .ZN(net_20659), .A(net_16439) );
AOI211_X4 inst_20991 ( .ZN(net_16083), .B(net_15545), .C2(net_14208), .A(net_12594), .C1(net_1693) );
NOR2_X4 inst_3239 ( .ZN(net_4125), .A2(net_2744), .A1(net_1802) );
CLKBUF_X2 inst_22773 ( .A(net_22644), .Z(net_22645) );
CLKBUF_X2 inst_22022 ( .A(net_21893), .Z(net_21894) );
OAI21_X2 inst_2314 ( .ZN(net_5730), .B1(net_3941), .B2(net_3218), .A(net_975) );
INV_X4 inst_12885 ( .A(net_16859), .ZN(net_16814) );
NOR2_X4 inst_2812 ( .A2(net_20104), .A1(net_20103), .ZN(net_17603) );
INV_X2 inst_19500 ( .A(net_6495), .ZN(net_2180) );
NOR2_X2 inst_4743 ( .A2(net_4214), .ZN(net_3042), .A1(net_3041) );
INV_X4 inst_15607 ( .ZN(net_2198), .A(net_2197) );
NOR2_X4 inst_3197 ( .A2(net_19726), .ZN(net_7120), .A1(net_3023) );
NOR2_X2 inst_4651 ( .A2(net_9289), .ZN(net_3345), .A1(net_1893) );
NAND2_X2 inst_10126 ( .A1(net_14038), .ZN(net_8354), .A2(net_5159) );
CLKBUF_X2 inst_22427 ( .A(net_22298), .Z(net_22299) );
DFF_X1 inst_19862 ( .D(net_17106), .CK(net_21340), .Q(x173) );
INV_X4 inst_13640 ( .ZN(net_10354), .A(net_8180) );
CLKBUF_X2 inst_21847 ( .A(net_21718), .Z(net_21719) );
NAND2_X2 inst_8006 ( .ZN(net_18303), .A2(net_18273), .A1(net_17298) );
INV_X4 inst_14988 ( .ZN(net_12216), .A(net_3400) );
CLKBUF_X2 inst_21569 ( .A(net_21412), .Z(net_21441) );
OR2_X4 inst_1083 ( .ZN(net_5597), .A2(net_5596), .A1(net_2343) );
CLKBUF_X2 inst_21867 ( .A(net_21738), .Z(net_21739) );
NOR2_X2 inst_4073 ( .ZN(net_7598), .A1(net_7597), .A2(net_7596) );
NAND3_X2 inst_6123 ( .ZN(net_13841), .A2(net_13840), .A3(net_10092), .A1(net_8636) );
OAI211_X2 inst_2466 ( .C1(net_15058), .ZN(net_14088), .B(net_13319), .C2(net_9051), .A(net_3283) );
AOI211_X4 inst_20994 ( .ZN(net_13463), .C1(net_13462), .B(net_9065), .C2(net_9028), .A(net_4454) );
NAND2_X2 inst_11979 ( .A1(net_1692), .ZN(net_1322), .A2(net_970) );
CLKBUF_X2 inst_22223 ( .A(net_22094), .Z(net_22095) );
NAND2_X2 inst_11877 ( .ZN(net_3172), .A2(net_1194), .A1(net_621) );
NAND2_X2 inst_12070 ( .ZN(net_1844), .A2(net_170), .A1(net_90) );
INV_X4 inst_13615 ( .A(net_8894), .ZN(net_8374) );
CLKBUF_X2 inst_22774 ( .A(net_22354), .Z(net_22646) );
SDFF_X2 inst_696 ( .Q(net_20921), .SI(net_18849), .SE(net_18581), .D(net_698), .CK(net_21302) );
NAND2_X2 inst_9719 ( .A2(net_10428), .ZN(net_10161), .A1(net_10160) );
CLKBUF_X2 inst_22325 ( .A(net_22196), .Z(net_22197) );
NAND2_X2 inst_11890 ( .A1(net_10714), .ZN(net_1597), .A2(net_1596) );
INV_X4 inst_15555 ( .A(net_2993), .ZN(net_2324) );
NAND2_X2 inst_10755 ( .A2(net_11718), .ZN(net_5693), .A1(net_4283) );
NAND2_X2 inst_12059 ( .A1(net_21238), .ZN(net_1300), .A2(net_90) );
NOR2_X2 inst_5055 ( .ZN(net_2231), .A1(net_1327), .A2(net_857) );
AOI21_X4 inst_20178 ( .ZN(net_19303), .B1(net_19079), .B2(net_14476), .A(net_12116) );
NAND3_X2 inst_6128 ( .A3(net_19910), .A1(net_19909), .ZN(net_19620), .A2(net_5212) );
CLKBUF_X2 inst_21812 ( .A(net_21683), .Z(net_21684) );
AOI22_X2 inst_20009 ( .ZN(net_12492), .B1(net_9843), .A2(net_7513), .A1(net_7394), .B2(net_3357) );
NAND2_X2 inst_10778 ( .ZN(net_5612), .A2(net_5611), .A1(net_3915) );
NOR2_X2 inst_3969 ( .ZN(net_8412), .A1(net_8411), .A2(net_8410) );
NAND2_X2 inst_11712 ( .ZN(net_2983), .A2(net_1153), .A1(net_1033) );
OAI21_X1 inst_2363 ( .ZN(net_7247), .A(net_7246), .B2(net_6633), .B1(net_2734) );
NAND2_X2 inst_9909 ( .ZN(net_9331), .A1(net_9330), .A2(net_9329) );
NAND3_X2 inst_6014 ( .ZN(net_14408), .A2(net_14407), .A3(net_14336), .A1(net_12555) );
NAND3_X2 inst_6257 ( .A2(net_20770), .ZN(net_13000), .A3(net_12999), .A1(net_6282) );
NOR2_X2 inst_4029 ( .A1(net_7992), .ZN(net_7991), .A2(net_6581) );
OAI21_X2 inst_1629 ( .ZN(net_20622), .A(net_16242), .B1(net_15432), .B2(net_15153) );
INV_X4 inst_16999 ( .ZN(net_1036), .A(net_303) );
CLKBUF_X2 inst_22012 ( .A(net_21883), .Z(net_21884) );
INV_X4 inst_17061 ( .ZN(net_3174), .A(net_448) );
INV_X4 inst_15583 ( .A(net_15666), .ZN(net_2267) );
INV_X1 inst_19763 ( .ZN(net_20648), .A(net_1587) );
NOR2_X2 inst_3424 ( .ZN(net_20400), .A2(net_15060), .A1(net_14991) );
INV_X4 inst_17840 ( .ZN(net_900), .A(net_790) );
NAND2_X1 inst_12138 ( .ZN(net_17354), .A1(net_17353), .A2(net_17212) );
AOI21_X4 inst_20155 ( .B2(net_20247), .B1(net_20246), .ZN(net_19471), .A(net_15245) );
INV_X4 inst_13923 ( .ZN(net_8219), .A(net_5561) );
AOI21_X2 inst_20565 ( .B2(net_20078), .ZN(net_19049), .A(net_8412), .B1(net_8411) );
INV_X4 inst_15895 ( .ZN(net_9541), .A(net_1773) );
OAI211_X2 inst_2580 ( .ZN(net_7678), .A(net_7677), .B(net_7676), .C1(net_2747), .C2(net_1539) );
CLKBUF_X2 inst_21386 ( .A(net_21257), .Z(net_21258) );
NAND2_X2 inst_11342 ( .A1(net_4512), .ZN(net_3676), .A2(net_3675) );
INV_X4 inst_16799 ( .A(net_5458), .ZN(net_4704) );
INV_X4 inst_14213 ( .ZN(net_5898), .A(net_5897) );
INV_X8 inst_12268 ( .ZN(net_19952), .A(net_1796) );
INV_X4 inst_17103 ( .ZN(net_1485), .A(net_621) );
NAND3_X2 inst_5840 ( .ZN(net_15496), .A1(net_14799), .A3(net_14154), .A2(net_13869) );
INV_X4 inst_15290 ( .ZN(net_4804), .A(net_1885) );
OAI21_X2 inst_2054 ( .ZN(net_10842), .A(net_7417), .B1(net_5664), .B2(net_1705) );
INV_X8 inst_12216 ( .ZN(net_7506), .A(net_6074) );
INV_X4 inst_13448 ( .ZN(net_9757), .A(net_9756) );
OAI22_X2 inst_1259 ( .B1(net_21162), .ZN(net_17532), .A1(net_17426), .B2(net_17143), .A2(net_17003) );
INV_X4 inst_18216 ( .A(net_21049), .ZN(net_697) );
INV_X2 inst_19412 ( .A(net_2860), .ZN(net_1968) );
INV_X4 inst_16148 ( .ZN(net_9940), .A(net_7836) );
NAND2_X2 inst_7821 ( .ZN(net_20032), .A2(net_18616), .A1(net_17052) );
OAI21_X2 inst_1796 ( .ZN(net_14507), .B2(net_11595), .B1(net_10313), .A(net_320) );
NAND2_X2 inst_10702 ( .ZN(net_11161), .A1(net_7489), .A2(net_6088) );
INV_X2 inst_18573 ( .A(net_12315), .ZN(net_10706) );
NAND2_X4 inst_7649 ( .ZN(net_1141), .A1(net_990), .A2(net_329) );
INV_X8 inst_12318 ( .ZN(net_1013), .A(net_722) );
XNOR2_X2 inst_535 ( .ZN(net_1675), .B(net_1674), .A(net_517) );
NAND2_X2 inst_11341 ( .A2(net_4203), .ZN(net_3677), .A1(net_85) );
AOI21_X2 inst_20941 ( .A(net_14186), .ZN(net_6412), .B1(net_4198), .B2(net_2766) );
INV_X4 inst_12970 ( .A(net_16517), .ZN(net_16516) );
NAND2_X2 inst_7853 ( .ZN(net_18586), .A2(net_18578), .A1(net_8283) );
NAND2_X2 inst_10059 ( .ZN(net_13154), .A1(net_8685), .A2(net_8684) );
INV_X4 inst_16589 ( .ZN(net_7198), .A(net_1145) );
OAI211_X2 inst_2427 ( .C2(net_19616), .C1(net_19615), .ZN(net_15169), .A(net_14410), .B(net_10104) );
NAND2_X2 inst_11670 ( .ZN(net_2381), .A2(net_2380), .A1(net_1645) );
NAND2_X2 inst_8603 ( .A1(net_21129), .A2(net_19452), .ZN(net_16671) );
NAND2_X2 inst_10496 ( .ZN(net_16009), .A2(net_6948), .A1(net_6924) );
CLKBUF_X2 inst_22594 ( .A(net_22045), .Z(net_22466) );
NOR2_X4 inst_3317 ( .ZN(net_1309), .A1(net_972), .A2(net_249) );
INV_X4 inst_14616 ( .ZN(net_7995), .A(net_4418) );
INV_X4 inst_17399 ( .ZN(net_4917), .A(net_846) );
NAND3_X2 inst_6079 ( .ZN(net_13971), .A3(net_13970), .A2(net_12836), .A1(net_12467) );
INV_X4 inst_13245 ( .ZN(net_13163), .A(net_12218) );
NAND2_X2 inst_11348 ( .A1(net_4918), .A2(net_4009), .ZN(net_3652) );
NAND2_X4 inst_7206 ( .A2(net_20077), .ZN(net_14361), .A1(net_7890) );
NOR2_X4 inst_3168 ( .ZN(net_5534), .A2(net_2744), .A1(net_2421) );
NOR2_X2 inst_3855 ( .ZN(net_9486), .A1(net_9485), .A2(net_9425) );
NAND2_X2 inst_8589 ( .A2(net_20072), .ZN(net_16711), .A1(net_16490) );
NOR2_X4 inst_3318 ( .ZN(net_1778), .A2(net_970), .A1(net_63) );
NAND2_X2 inst_10594 ( .A2(net_12952), .A1(net_9735), .ZN(net_6638) );
INV_X4 inst_12771 ( .A(net_17515), .ZN(net_17335) );
NAND2_X2 inst_10299 ( .A1(net_11681), .ZN(net_7897), .A2(net_4757) );
AOI21_X2 inst_20959 ( .B1(net_5516), .ZN(net_5332), .B2(net_5230), .A(net_4170) );
AOI21_X2 inst_20928 ( .ZN(net_7088), .B1(net_7087), .A(net_4255), .B2(net_4116) );
AOI21_X2 inst_20540 ( .B2(net_20031), .B1(net_20030), .ZN(net_14473), .A(net_14472) );
CLKBUF_X2 inst_22355 ( .A(net_22226), .Z(net_22227) );
NAND4_X4 inst_5176 ( .ZN(net_16665), .A1(net_16353), .A4(net_16176), .A3(net_15887), .A2(net_10824) );
INV_X4 inst_12672 ( .ZN(net_17745), .A(net_17744) );
INV_X2 inst_19145 ( .ZN(net_6815), .A(net_5573) );
OAI22_X1 inst_1322 ( .A1(net_19422), .B2(net_19421), .ZN(net_17116), .B1(net_17115), .A2(net_16799) );
INV_X4 inst_16483 ( .ZN(net_10917), .A(net_5701) );
NAND2_X2 inst_11862 ( .A1(net_21106), .ZN(net_1656), .A2(net_1351) );
INV_X4 inst_17380 ( .ZN(net_1617), .A(net_955) );
CLKBUF_X2 inst_21505 ( .A(net_21350), .Z(net_21377) );
CLKBUF_X2 inst_21440 ( .A(net_21311), .Z(net_21312) );
NAND2_X2 inst_10954 ( .ZN(net_10654), .A1(net_8639), .A2(net_5091) );
INV_X4 inst_14891 ( .A(net_6801), .ZN(net_3653) );
INV_X4 inst_14004 ( .A(net_9935), .ZN(net_9827) );
NAND2_X2 inst_10712 ( .A1(net_10737), .ZN(net_8802), .A2(net_5964) );
INV_X4 inst_14237 ( .ZN(net_9106), .A(net_5814) );
NAND2_X2 inst_10248 ( .ZN(net_15427), .A2(net_5031), .A1(net_60) );
INV_X4 inst_15471 ( .ZN(net_11747), .A(net_10947) );
INV_X4 inst_17029 ( .ZN(net_14734), .A(net_909) );
AOI21_X2 inst_20299 ( .ZN(net_16122), .B2(net_15724), .A(net_15576), .B1(net_7319) );
NAND2_X4 inst_7668 ( .ZN(net_1370), .A1(net_880), .A2(net_108) );
CLKBUF_X2 inst_21770 ( .A(net_21641), .Z(net_21642) );
NAND2_X2 inst_8379 ( .A2(net_17571), .ZN(net_17347), .A1(net_17346) );
NAND2_X2 inst_10156 ( .ZN(net_8265), .A1(net_8264), .A2(net_5056) );
NOR2_X2 inst_3493 ( .ZN(net_18924), .A1(net_13398), .A2(net_9772) );
NAND2_X2 inst_9776 ( .A1(net_10467), .ZN(net_9789), .A2(net_8554) );
NAND2_X2 inst_10413 ( .A1(net_9638), .ZN(net_7251), .A2(net_7250) );
INV_X4 inst_13151 ( .ZN(net_14890), .A(net_14375) );
NOR2_X2 inst_4622 ( .ZN(net_3610), .A1(net_3609), .A2(net_1996) );
CLKBUF_X2 inst_21481 ( .A(net_21352), .Z(net_21353) );
NOR2_X2 inst_3487 ( .ZN(net_14286), .A2(net_13485), .A1(net_1307) );
NOR2_X2 inst_3597 ( .ZN(net_12583), .A2(net_12582), .A1(net_4134) );
NAND2_X2 inst_11783 ( .ZN(net_2010), .A1(net_2009), .A2(net_2008) );
INV_X4 inst_14421 ( .ZN(net_6185), .A(net_5051) );
INV_X4 inst_14555 ( .ZN(net_5839), .A(net_4588) );
NAND2_X2 inst_8210 ( .ZN(net_17857), .A1(net_17693), .A2(net_17571) );
NAND2_X2 inst_10661 ( .ZN(net_19015), .A1(net_13026), .A2(net_6301) );
CLKBUF_X2 inst_22503 ( .A(net_22374), .Z(net_22375) );
NAND2_X2 inst_11757 ( .ZN(net_11225), .A2(net_2097), .A1(net_170) );
CLKBUF_X2 inst_22711 ( .A(net_22582), .Z(net_22583) );
INV_X4 inst_13422 ( .ZN(net_11503), .A(net_10133) );
NOR3_X4 inst_2607 ( .A3(net_19472), .A1(net_19471), .ZN(net_19366), .A2(net_12170) );
INV_X4 inst_16287 ( .A(net_14678), .ZN(net_1340) );
NAND2_X2 inst_8133 ( .ZN(net_18038), .A2(net_18027), .A1(net_18019) );
INV_X4 inst_13893 ( .ZN(net_11880), .A(net_7293) );
NAND2_X2 inst_11395 ( .ZN(net_3496), .A2(net_2531), .A1(net_1848) );
CLKBUF_X2 inst_22477 ( .A(net_22348), .Z(net_22349) );
NAND2_X2 inst_7791 ( .ZN(net_18714), .A2(net_18713), .A1(net_17440) );
NOR3_X2 inst_2690 ( .ZN(net_14345), .A2(net_13824), .A3(net_13788), .A1(net_10130) );
DFF_X1 inst_19918 ( .D(net_16621), .CK(net_22784), .Q(x1227) );
NAND2_X2 inst_8689 ( .ZN(net_16391), .A2(net_16308), .A1(net_15947) );
AOI21_X4 inst_20227 ( .B1(net_19497), .ZN(net_19040), .B2(net_13699), .A(net_8526) );
CLKBUF_X2 inst_22274 ( .A(net_21647), .Z(net_22146) );
NAND2_X2 inst_10467 ( .ZN(net_8359), .A2(net_7000), .A1(net_732) );
CLKBUF_X2 inst_21632 ( .A(net_21503), .Z(net_21504) );
INV_X4 inst_16167 ( .ZN(net_6626), .A(net_6325) );
OAI21_X2 inst_1544 ( .ZN(net_17874), .B1(net_17683), .B2(net_17660), .A(net_17655) );
CLKBUF_X2 inst_22250 ( .A(net_21783), .Z(net_22122) );
AOI21_X2 inst_20414 ( .ZN(net_15277), .A(net_15276), .B2(net_14184), .B1(net_9031) );
DFF_X1 inst_19853 ( .D(net_17160), .CK(net_21601), .Q(x668) );
NAND3_X2 inst_6261 ( .ZN(net_12993), .A1(net_12992), .A3(net_12991), .A2(net_9795) );
NAND2_X2 inst_9771 ( .ZN(net_20109), .A1(net_10449), .A2(net_9799) );
NOR2_X4 inst_3148 ( .ZN(net_4589), .A1(net_3566), .A2(net_758) );
INV_X4 inst_17721 ( .ZN(net_807), .A(net_287) );
NOR2_X2 inst_4761 ( .ZN(net_4267), .A2(net_2991), .A1(net_165) );
NAND4_X4 inst_5180 ( .A2(net_18939), .A1(net_18938), .ZN(net_16985), .A4(net_16279), .A3(net_16278) );
NOR2_X4 inst_3026 ( .ZN(net_7769), .A1(net_5234), .A2(net_3356) );
NAND2_X4 inst_6952 ( .A2(net_20158), .A1(net_20157), .ZN(net_17507) );
NAND2_X2 inst_8573 ( .ZN(net_16733), .A1(net_16732), .A2(net_16562) );
INV_X4 inst_17017 ( .A(net_15370), .ZN(net_15369) );
NOR2_X2 inst_3639 ( .ZN(net_12103), .A1(net_11546), .A2(net_7342) );
INV_X4 inst_13646 ( .A(net_8931), .ZN(net_8161) );
NAND2_X4 inst_7226 ( .ZN(net_9199), .A1(net_3586), .A2(net_3491) );
NAND2_X2 inst_9194 ( .ZN(net_13108), .A2(net_13107), .A1(net_10340) );
NAND2_X2 inst_10411 ( .ZN(net_13192), .A2(net_7260), .A1(net_6845) );
INV_X4 inst_13130 ( .ZN(net_15269), .A(net_14883) );
INV_X4 inst_14241 ( .A(net_9506), .ZN(net_5784) );
INV_X4 inst_12769 ( .ZN(net_17338), .A(net_17337) );
SDFF_X2 inst_752 ( .Q(net_20908), .SE(net_18584), .SI(net_18534), .D(net_11871), .CK(net_22694) );
NOR2_X4 inst_3245 ( .ZN(net_4287), .A1(net_2934), .A2(net_2275) );
NOR2_X4 inst_3202 ( .A2(net_20495), .ZN(net_5393), .A1(net_3095) );
NOR2_X2 inst_4279 ( .ZN(net_6108), .A2(net_6107), .A1(net_4477) );
INV_X4 inst_18125 ( .A(net_21067), .ZN(net_668) );
OAI21_X4 inst_1384 ( .A(net_20896), .B2(net_19549), .B1(net_19548), .ZN(net_16345) );
INV_X4 inst_16116 ( .ZN(net_6237), .A(net_1290) );
OAI21_X2 inst_2118 ( .ZN(net_10023), .A(net_8286), .B2(net_7952), .B1(net_2989) );
AND2_X2 inst_21273 ( .ZN(net_19072), .A1(net_15463), .A2(net_14200) );
INV_X4 inst_16112 ( .ZN(net_2149), .A(net_1836) );
NAND2_X2 inst_7749 ( .ZN(net_18779), .A2(net_18758), .A1(net_18734) );
INV_X2 inst_19554 ( .ZN(net_19287), .A(net_932) );
AOI21_X4 inst_20220 ( .ZN(net_14103), .A(net_11417), .B2(net_10571), .B1(net_588) );
INV_X4 inst_18347 ( .ZN(net_20845), .A(net_20780) );
NAND2_X2 inst_8817 ( .ZN(net_15579), .A2(net_14846), .A1(net_12638) );
NOR2_X2 inst_5048 ( .ZN(net_3234), .A1(net_1842), .A2(net_946) );
INV_X2 inst_18866 ( .A(net_8344), .ZN(net_6286) );
INV_X2 inst_19485 ( .ZN(net_1623), .A(net_1336) );
NAND2_X2 inst_11470 ( .ZN(net_7023), .A1(net_3148), .A2(net_3147) );
INV_X4 inst_12693 ( .ZN(net_17643), .A(net_17642) );
NOR2_X2 inst_4356 ( .ZN(net_20025), .A2(net_4321), .A1(net_3104) );
INV_X2 inst_18753 ( .ZN(net_20121), .A(net_6472) );
INV_X4 inst_18226 ( .A(net_21102), .ZN(net_599) );
AOI21_X2 inst_20460 ( .B1(net_15666), .ZN(net_15033), .A(net_13913), .B2(net_6453) );
INV_X4 inst_16761 ( .ZN(net_1035), .A(net_1034) );
NAND2_X2 inst_11707 ( .ZN(net_2286), .A1(net_2285), .A2(net_1735) );
NAND2_X2 inst_9975 ( .ZN(net_10315), .A1(net_8877), .A2(net_7828) );
INV_X8 inst_12250 ( .ZN(net_5291), .A(net_1957) );
AND2_X4 inst_21262 ( .A1(net_1376), .ZN(net_1166), .A2(net_227) );
NAND4_X2 inst_5329 ( .ZN(net_15572), .A4(net_14207), .A1(net_11998), .A2(net_10696), .A3(net_9930) );
OAI211_X2 inst_2539 ( .ZN(net_10832), .B(net_10831), .C2(net_9698), .C1(net_3497), .A(net_1892) );
NAND2_X2 inst_10141 ( .ZN(net_19335), .A2(net_6958), .A1(net_4434) );
INV_X4 inst_13496 ( .ZN(net_10936), .A(net_7910) );
NOR3_X2 inst_2797 ( .A2(net_12179), .A3(net_4039), .ZN(net_2677), .A1(net_2676) );
CLKBUF_X2 inst_22868 ( .A(net_21782), .Z(net_22740) );
NOR2_X2 inst_3431 ( .ZN(net_19394), .A2(net_14404), .A1(net_13826) );
INV_X4 inst_13193 ( .ZN(net_14126), .A(net_13465) );
OAI21_X2 inst_2085 ( .ZN(net_10412), .B2(net_9746), .A(net_5694), .B1(net_1199) );
INV_X4 inst_17062 ( .ZN(net_15664), .A(net_11968) );
NAND2_X2 inst_11097 ( .ZN(net_4342), .A2(net_4337), .A1(net_3030) );
INV_X2 inst_19677 ( .A(net_20511), .ZN(net_20510) );
NAND4_X2 inst_5264 ( .A2(net_20264), .A1(net_20263), .A4(net_20200), .ZN(net_19651), .A3(net_14705) );
INV_X2 inst_19518 ( .ZN(net_2104), .A(net_1122) );
INV_X4 inst_12910 ( .ZN(net_17220), .A(net_16909) );
NAND2_X4 inst_7069 ( .A1(net_20358), .ZN(net_16206), .A2(net_16035) );
NAND3_X2 inst_6150 ( .ZN(net_13681), .A3(net_13607), .A2(net_10957), .A1(net_5692) );
INV_X4 inst_14230 ( .ZN(net_10834), .A(net_5829) );
XNOR2_X2 inst_556 ( .B(net_16462), .ZN(net_698), .A(net_697) );
NAND2_X2 inst_11779 ( .ZN(net_2027), .A2(net_253), .A1(x6280) );
NOR2_X2 inst_3632 ( .A1(net_13184), .A2(net_13114), .ZN(net_12197) );
AOI21_X2 inst_20885 ( .ZN(net_7817), .B2(net_7665), .B1(net_2997), .A(net_1124) );
NOR2_X1 inst_5147 ( .ZN(net_11653), .A2(net_11478), .A1(net_10701) );
INV_X4 inst_13758 ( .ZN(net_10995), .A(net_7613) );
INV_X4 inst_12573 ( .ZN(net_18231), .A(net_18198) );
DFF_X1 inst_19856 ( .D(net_18872), .CK(net_21983), .Q(x990) );
INV_X2 inst_19729 ( .A(net_20802), .ZN(net_20801) );
NAND2_X2 inst_9650 ( .ZN(net_10363), .A1(net_10063), .A2(net_7761) );
INV_X4 inst_15641 ( .ZN(net_3098), .A(net_2124) );
INV_X4 inst_16457 ( .ZN(net_1222), .A(net_1221) );
NOR2_X4 inst_3300 ( .ZN(net_1718), .A1(net_1699), .A2(net_988) );
NAND2_X4 inst_7597 ( .ZN(net_2546), .A1(net_1751), .A2(net_1384) );
INV_X4 inst_12728 ( .ZN(net_17479), .A(net_17478) );
NOR2_X2 inst_3822 ( .ZN(net_9778), .A2(net_9777), .A1(net_5065) );
NAND2_X2 inst_8757 ( .A1(net_16404), .ZN(net_15909), .A2(net_15516) );
NAND2_X2 inst_9603 ( .ZN(net_13053), .A1(net_10737), .A2(net_9316) );
NAND2_X4 inst_7522 ( .ZN(net_4132), .A1(net_2960), .A2(net_1059) );
NOR2_X2 inst_4593 ( .A1(net_7962), .ZN(net_4765), .A2(net_2774) );
AOI21_X2 inst_20840 ( .ZN(net_9273), .A(net_7599), .B1(net_7580), .B2(net_5989) );
NAND3_X2 inst_6070 ( .ZN(net_14124), .A1(net_11655), .A3(net_10552), .A2(net_8638) );
INV_X4 inst_17769 ( .ZN(net_1384), .A(net_889) );
NOR2_X4 inst_3307 ( .ZN(net_1590), .A1(net_939), .A2(net_110) );
OAI21_X2 inst_1587 ( .ZN(net_19480), .A(net_16359), .B2(net_15941), .B1(net_10601) );
NAND4_X2 inst_5452 ( .ZN(net_13467), .A4(net_10582), .A2(net_9159), .A1(net_5638), .A3(net_4415) );
OR2_X2 inst_1185 ( .ZN(net_4622), .A1(net_4621), .A2(net_1875) );
INV_X4 inst_16262 ( .ZN(net_2195), .A(net_2171) );
NAND2_X2 inst_8742 ( .ZN(net_19503), .A1(net_15991), .A2(net_15814) );
XNOR2_X2 inst_457 ( .ZN(net_13297), .B(net_13296), .A(net_9713) );
INV_X4 inst_13715 ( .ZN(net_11748), .A(net_7828) );
INV_X4 inst_16213 ( .ZN(net_2034), .A(net_1937) );
OAI21_X2 inst_1738 ( .ZN(net_15065), .A(net_15064), .B1(net_13496), .B2(net_11793) );
NOR2_X4 inst_2802 ( .ZN(net_18602), .A2(net_18599), .A1(net_16195) );
INV_X2 inst_19457 ( .A(net_2240), .ZN(net_1508) );
NOR2_X2 inst_4171 ( .A2(net_9887), .A1(net_9131), .ZN(net_8753) );
INV_X4 inst_15169 ( .ZN(net_12915), .A(net_3016) );
NAND2_X2 inst_11276 ( .ZN(net_13147), .A2(net_3367), .A1(net_1790) );
DFF_X1 inst_19859 ( .D(net_17255), .CK(net_22065), .Q(x424) );
INV_X4 inst_16385 ( .ZN(net_19324), .A(net_107) );
NAND2_X4 inst_7204 ( .ZN(net_10254), .A2(net_8175), .A1(net_874) );
NAND3_X4 inst_5529 ( .A3(net_19405), .A1(net_19404), .ZN(net_17660), .A2(net_16042) );
INV_X4 inst_14984 ( .ZN(net_16037), .A(net_15889) );
NAND2_X2 inst_8953 ( .ZN(net_14721), .A1(net_14720), .A2(net_13316) );
NAND2_X2 inst_10250 ( .A1(net_11391), .ZN(net_8009), .A2(net_5004) );
INV_X4 inst_16259 ( .ZN(net_6876), .A(net_4288) );
NAND3_X2 inst_6103 ( .ZN(net_13905), .A1(net_12049), .A3(net_11387), .A2(net_9679) );
CLKBUF_X2 inst_22333 ( .A(net_21577), .Z(net_22205) );
INV_X4 inst_16953 ( .ZN(net_1193), .A(net_907) );
XNOR2_X2 inst_146 ( .ZN(net_18043), .A(net_18014), .B(net_17667) );
INV_X4 inst_15588 ( .ZN(net_7712), .A(net_2261) );
NOR2_X2 inst_3999 ( .ZN(net_8227), .A1(net_8226), .A2(net_8225) );
INV_X2 inst_18710 ( .ZN(net_11856), .A(net_8231) );
INV_X2 inst_18703 ( .ZN(net_11372), .A(net_10428) );
INV_X4 inst_12501 ( .A(net_18617), .ZN(net_18616) );
XNOR2_X2 inst_326 ( .B(net_21127), .ZN(net_17695), .A(net_17024) );
SDFF_X2 inst_817 ( .Q(net_21225), .SI(net_17769), .SE(net_125), .CK(net_21479), .D(x7198) );
NAND2_X2 inst_10589 ( .ZN(net_6658), .A2(net_4778), .A1(net_4264) );
INV_X4 inst_12550 ( .ZN(net_18335), .A(net_18261) );
OAI21_X2 inst_2194 ( .A(net_14563), .ZN(net_8584), .B2(net_8583), .B1(net_3215) );
NAND2_X2 inst_10789 ( .ZN(net_19337), .A1(net_13091), .A2(net_3123) );
INV_X4 inst_16365 ( .ZN(net_2439), .A(net_1288) );
INV_X2 inst_18419 ( .ZN(net_15624), .A(net_15386) );
INV_X2 inst_18698 ( .A(net_10433), .ZN(net_9784) );
INV_X2 inst_18691 ( .ZN(net_8519), .A(net_8518) );
NOR2_X4 inst_3293 ( .A1(net_19537), .ZN(net_2291), .A2(net_1134) );
INV_X4 inst_15825 ( .ZN(net_1868), .A(net_1052) );
CLKBUF_X2 inst_22238 ( .A(net_22109), .Z(net_22110) );
CLKBUF_X2 inst_21763 ( .A(net_21334), .Z(net_21635) );
INV_X2 inst_18809 ( .ZN(net_7369), .A(net_7368) );
INV_X4 inst_16808 ( .ZN(net_7976), .A(net_1759) );
NOR2_X2 inst_3793 ( .ZN(net_10077), .A2(net_6324), .A1(net_5696) );
AOI21_X2 inst_20324 ( .ZN(net_19780), .B2(net_15309), .B1(net_14476), .A(net_13979) );
INV_X4 inst_18333 ( .A(net_20570), .ZN(net_20569) );
XNOR2_X2 inst_108 ( .ZN(net_18520), .A(net_18404), .B(net_17023) );
NAND2_X2 inst_11143 ( .ZN(net_4227), .A2(net_4226), .A1(net_2136) );
INV_X4 inst_16475 ( .ZN(net_1212), .A(net_1211) );
NOR2_X2 inst_4799 ( .ZN(net_6792), .A1(net_1489), .A2(net_1234) );
NOR2_X2 inst_3778 ( .A1(net_11562), .ZN(net_11522), .A2(net_7943) );
NOR2_X2 inst_3940 ( .ZN(net_20345), .A2(net_8649), .A1(net_4958) );
NAND3_X2 inst_6503 ( .ZN(net_10814), .A2(net_7368), .A3(net_6311), .A1(net_3573) );
INV_X2 inst_19689 ( .ZN(net_20537), .A(net_20536) );
XNOR2_X2 inst_638 ( .B(net_16470), .ZN(net_425), .A(net_424) );
NAND2_X2 inst_11937 ( .ZN(net_1459), .A1(net_1176), .A2(net_1107) );
NAND2_X2 inst_7786 ( .ZN(net_18724), .A2(net_18723), .A1(net_17733) );
NAND2_X2 inst_10311 ( .ZN(net_9381), .A1(net_7849), .A2(net_4867) );
CLKBUF_X2 inst_21621 ( .A(net_21492), .Z(net_21493) );
CLKBUF_X2 inst_21447 ( .A(net_21313), .Z(net_21319) );
INV_X4 inst_18139 ( .A(net_20849), .ZN(net_1469) );
NOR2_X2 inst_5008 ( .A1(net_2274), .ZN(net_1290), .A2(net_878) );
NOR2_X4 inst_3275 ( .ZN(net_1702), .A1(net_1096), .A2(net_110) );
NAND2_X2 inst_9237 ( .ZN(net_12709), .A1(net_12708), .A2(net_12707) );
OAI21_X4 inst_1466 ( .ZN(net_18921), .A(net_14103), .B2(net_13302), .B1(net_588) );
OAI21_X2 inst_1726 ( .ZN(net_15091), .A(net_14791), .B2(net_12904), .B1(net_8711) );
NOR2_X4 inst_2841 ( .ZN(net_14627), .A2(net_13305), .A1(net_9540) );
NAND2_X4 inst_7157 ( .ZN(net_11558), .A2(net_9571), .A1(net_9570) );
INV_X4 inst_15591 ( .ZN(net_16287), .A(net_16011) );
CLKBUF_X2 inst_22324 ( .A(net_22195), .Z(net_22196) );
INV_X4 inst_14251 ( .A(net_13157), .ZN(net_10496) );
NAND2_X4 inst_7118 ( .ZN(net_12388), .A1(net_11020), .A2(net_10000) );
INV_X4 inst_16170 ( .A(net_1666), .ZN(net_1446) );
NAND2_X2 inst_10892 ( .ZN(net_9010), .A1(net_5402), .A2(net_5401) );
INV_X4 inst_14576 ( .ZN(net_5810), .A(net_4535) );
SDFF_X2 inst_905 ( .Q(net_21154), .D(net_16850), .SE(net_263), .CK(net_22212), .SI(x5568) );
INV_X4 inst_16426 ( .ZN(net_1876), .A(net_1250) );
INV_X4 inst_14677 ( .ZN(net_10701), .A(net_4309) );
INV_X4 inst_15991 ( .A(net_2219), .ZN(net_1935) );
NAND2_X2 inst_11571 ( .ZN(net_6434), .A1(net_6316), .A2(net_3246) );
CLKBUF_X2 inst_21931 ( .A(net_21338), .Z(net_21803) );
INV_X2 inst_19628 ( .A(net_21107), .ZN(net_33) );
INV_X4 inst_14860 ( .ZN(net_6898), .A(net_3779) );
NOR2_X2 inst_4214 ( .ZN(net_8690), .A1(net_6637), .A2(net_4926) );
INV_X4 inst_12753 ( .ZN(net_17410), .A(net_17409) );
INV_X4 inst_18242 ( .A(net_21065), .ZN(net_619) );
NOR2_X2 inst_3834 ( .ZN(net_9697), .A2(net_9696), .A1(net_6313) );
INV_X4 inst_16687 ( .A(net_13089), .ZN(net_1774) );
NOR2_X2 inst_3651 ( .ZN(net_11671), .A2(net_11670), .A1(net_11009) );
AOI21_X4 inst_20196 ( .B1(net_19943), .ZN(net_15098), .B2(net_14214), .A(net_13703) );
OAI21_X2 inst_1759 ( .B2(net_20083), .B1(net_20082), .ZN(net_18973), .A(net_11395) );
AOI21_X2 inst_20778 ( .ZN(net_19224), .B1(net_10569), .A(net_7136), .B2(net_6403) );
NOR3_X4 inst_2615 ( .A3(net_19807), .A1(net_19806), .ZN(net_18985), .A2(net_7773) );
NAND2_X2 inst_11792 ( .ZN(net_3275), .A1(net_1962), .A2(net_1961) );
NAND4_X2 inst_5485 ( .A2(net_19888), .A1(net_19887), .ZN(net_12404), .A4(net_5726), .A3(net_5493) );
INV_X4 inst_13859 ( .A(net_9386), .ZN(net_7461) );
NAND2_X4 inst_7017 ( .ZN(net_17243), .A1(net_16601), .A2(net_16466) );
NOR2_X2 inst_3463 ( .A2(net_19945), .A1(net_19944), .ZN(net_19113) );
INV_X4 inst_16055 ( .ZN(net_2206), .A(net_1590) );
INV_X4 inst_17867 ( .A(net_972), .ZN(net_295) );
AOI22_X2 inst_20025 ( .ZN(net_9941), .A1(net_9940), .B1(net_8184), .A2(net_4674), .B2(net_3510) );
NAND2_X4 inst_7617 ( .ZN(net_1793), .A2(net_1333), .A1(net_927) );
NAND3_X2 inst_6375 ( .ZN(net_12042), .A1(net_12041), .A3(net_9818), .A2(net_7606) );
NAND2_X2 inst_11115 ( .A1(net_20563), .ZN(net_5539), .A2(net_4316) );
INV_X4 inst_12492 ( .ZN(net_18669), .A(net_18654) );
NOR2_X2 inst_4055 ( .ZN(net_7841), .A2(net_7840), .A1(net_5166) );
INV_X4 inst_16463 ( .ZN(net_2317), .A(net_1219) );
OAI22_X4 inst_1247 ( .ZN(net_17665), .B2(net_17590), .A2(net_17224), .B1(net_16843), .A1(net_16642) );
NAND4_X2 inst_5284 ( .A4(net_19051), .A1(net_19050), .ZN(net_15953), .A2(net_10704), .A3(net_7117) );
INV_X2 inst_18942 ( .ZN(net_5741), .A(net_5740) );
INV_X4 inst_13275 ( .ZN(net_12463), .A(net_11188) );
INV_X4 inst_14541 ( .ZN(net_4644), .A(net_4643) );
INV_X4 inst_17140 ( .ZN(net_9785), .A(net_5205) );
AOI21_X2 inst_20777 ( .ZN(net_10589), .B1(net_9131), .A(net_8013), .B2(net_6428) );
OAI21_X4 inst_1493 ( .ZN(net_20355), .A(net_9130), .B2(net_5991), .B1(net_2876) );
NOR2_X4 inst_2998 ( .ZN(net_7406), .A1(net_5893), .A2(net_5591) );
NAND2_X2 inst_11734 ( .ZN(net_19676), .A2(net_2449), .A1(net_2195) );
NOR3_X4 inst_2612 ( .ZN(net_19155), .A1(net_15807), .A3(net_15303), .A2(net_11967) );
INV_X4 inst_13348 ( .ZN(net_12710), .A(net_11039) );
INV_X4 inst_14116 ( .ZN(net_6147), .A(net_6146) );
INV_X4 inst_15623 ( .ZN(net_4192), .A(net_2153) );
AOI21_X4 inst_20218 ( .ZN(net_14177), .B2(net_10763), .A(net_10687), .B1(net_1449) );
INV_X2 inst_19206 ( .A(net_5006), .ZN(net_3540) );
OAI21_X4 inst_1362 ( .A(net_20912), .B2(net_19321), .B1(net_19320), .ZN(net_18049) );
NAND2_X2 inst_8881 ( .ZN(net_20588), .A1(net_15183), .A2(net_14597) );
INV_X4 inst_12888 ( .A(net_16870), .ZN(net_16812) );
INV_X4 inst_13798 ( .ZN(net_12467), .A(net_9392) );
INV_X2 inst_19110 ( .A(net_5970), .ZN(net_4465) );
XNOR2_X2 inst_272 ( .ZN(net_17211), .A(net_16835), .B(net_434) );
INV_X4 inst_14311 ( .ZN(net_6795), .A(net_5770) );
NOR2_X2 inst_4718 ( .ZN(net_3130), .A2(net_3082), .A1(net_1376) );
AOI22_X2 inst_20055 ( .ZN(net_3698), .B2(net_3697), .A2(net_2726), .A1(net_1233), .B1(net_933) );
NAND2_X2 inst_9213 ( .ZN(net_13040), .A2(net_11358), .A1(net_4687) );
AOI21_X2 inst_20588 ( .B2(net_20058), .B1(net_20057), .A(net_15616), .ZN(net_14011) );
NOR2_X2 inst_4133 ( .ZN(net_19954), .A2(net_6956), .A1(net_4104) );
SDFF_X2 inst_789 ( .Q(net_20853), .SE(net_18576), .SI(net_18036), .D(net_1512), .CK(net_21801) );
OAI21_X2 inst_1806 ( .ZN(net_14470), .B2(net_12517), .A(net_9620), .B1(net_9472) );
OAI21_X2 inst_1810 ( .B2(net_19926), .B1(net_19925), .ZN(net_14204), .A(net_14203) );
OAI21_X2 inst_1860 ( .ZN(net_13806), .A(net_13805), .B2(net_10604), .B1(net_3266) );
INV_X4 inst_15177 ( .ZN(net_7838), .A(net_2498) );
INV_X4 inst_16636 ( .ZN(net_1999), .A(net_1107) );
INV_X4 inst_15561 ( .ZN(net_10231), .A(net_4931) );
OAI21_X2 inst_1885 ( .A(net_15452), .ZN(net_13520), .B2(net_9025), .B1(net_7045) );
CLKBUF_X2 inst_22294 ( .A(net_22165), .Z(net_22166) );
INV_X4 inst_13232 ( .ZN(net_19088), .A(net_12448) );
NAND2_X2 inst_7926 ( .ZN(net_20720), .A1(net_20018), .A2(net_17876) );
NAND2_X2 inst_11184 ( .ZN(net_6983), .A1(net_4288), .A2(net_1880) );
INV_X2 inst_18505 ( .ZN(net_11932), .A(net_10508) );
INV_X4 inst_14136 ( .A(net_8204), .ZN(net_6090) );
INV_X4 inst_13189 ( .ZN(net_19832), .A(net_13613) );
INV_X2 inst_18981 ( .A(net_8035), .ZN(net_5144) );
NOR2_X2 inst_4885 ( .A2(net_7703), .ZN(net_4334), .A1(net_1435) );
AOI21_X2 inst_20686 ( .B1(net_14743), .ZN(net_12260), .A(net_12259), .B2(net_8516) );
INV_X4 inst_17149 ( .ZN(net_7253), .A(net_5244) );
CLKBUF_X2 inst_22396 ( .A(net_22267), .Z(net_22268) );
INV_X4 inst_18255 ( .A(net_21167), .ZN(net_16879) );
OAI211_X2 inst_2496 ( .ZN(net_12919), .C1(net_12036), .C2(net_11182), .B(net_4534), .A(net_4367) );
NAND2_X2 inst_8393 ( .ZN(net_17409), .A2(net_17018), .A1(net_16872) );
INV_X4 inst_13466 ( .ZN(net_13322), .A(net_9678) );
INV_X4 inst_15158 ( .A(net_11318), .ZN(net_9569) );
NOR2_X2 inst_4381 ( .ZN(net_5326), .A2(net_3974), .A1(net_2336) );
INV_X4 inst_17940 ( .A(net_21038), .ZN(net_716) );
NAND2_X2 inst_11406 ( .ZN(net_6229), .A1(net_2731), .A2(net_2373) );
CLKBUF_X2 inst_21989 ( .A(net_21860), .Z(net_21861) );
NAND2_X2 inst_11280 ( .A2(net_3946), .ZN(net_3858), .A1(net_573) );
NAND2_X2 inst_8229 ( .ZN(net_17969), .A1(net_17605), .A2(net_17601) );
INV_X2 inst_19707 ( .ZN(net_20574), .A(net_20568) );
NOR3_X2 inst_2671 ( .ZN(net_14818), .A2(net_14817), .A1(net_11436), .A3(net_7805) );
INV_X4 inst_17689 ( .ZN(net_2709), .A(net_226) );
INV_X4 inst_16675 ( .ZN(net_5499), .A(net_4526) );
NAND2_X2 inst_9638 ( .A1(net_10875), .ZN(net_10396), .A2(net_10393) );
INV_X4 inst_18118 ( .A(net_21066), .ZN(net_424) );
INV_X4 inst_14713 ( .ZN(net_6039), .A(net_2703) );
INV_X4 inst_13068 ( .ZN(net_19355), .A(net_16224) );
DFF_X1 inst_19831 ( .D(net_17528), .CK(net_21761), .Q(x33) );
OAI21_X4 inst_1355 ( .ZN(net_18351), .B2(net_18299), .A(net_18215), .B1(net_18214) );
NAND3_X2 inst_6612 ( .A3(net_14921), .A2(net_9663), .ZN(net_9078), .A1(net_6927) );
SDFF_X2 inst_877 ( .Q(net_21159), .SI(net_16892), .SE(net_125), .CK(net_22228), .D(x5360) );
NAND2_X2 inst_10267 ( .ZN(net_9523), .A2(net_7881), .A1(net_7659) );
INV_X2 inst_18717 ( .ZN(net_8167), .A(net_8166) );
CLKBUF_X2 inst_22311 ( .A(net_22182), .Z(net_22183) );
NAND3_X2 inst_6563 ( .A2(net_12442), .ZN(net_10483), .A3(net_6789), .A1(net_4790) );
NAND2_X2 inst_10704 ( .ZN(net_8744), .A2(net_6126), .A1(net_3707) );
INV_X4 inst_12698 ( .ZN(net_17630), .A(net_17629) );
NAND2_X4 inst_7372 ( .ZN(net_11822), .A2(net_4305), .A1(net_3077) );
AOI22_X2 inst_20053 ( .ZN(net_3701), .A1(net_3700), .B2(net_3351), .A2(net_1463), .B1(net_1016) );
NAND3_X2 inst_6384 ( .ZN(net_12021), .A2(net_9209), .A1(net_5614), .A3(net_5463) );
INV_X2 inst_19666 ( .A(net_20477), .ZN(net_20476) );
INV_X4 inst_17430 ( .A(net_4770), .ZN(net_4715) );
NAND3_X2 inst_5829 ( .A2(net_20614), .A1(net_20613), .ZN(net_15532), .A3(net_14715) );
INV_X4 inst_14523 ( .A(net_15519), .ZN(net_4772) );
NAND3_X2 inst_5904 ( .ZN(net_15128), .A3(net_13394), .A2(net_11564), .A1(net_9644) );
NAND2_X2 inst_10274 ( .ZN(net_7963), .A1(net_7962), .A2(net_5920) );
NAND2_X2 inst_10734 ( .A2(net_11822), .A1(net_10627), .ZN(net_5772) );
NAND2_X2 inst_11013 ( .ZN(net_20381), .A1(net_4807), .A2(net_2474) );
AND2_X2 inst_21340 ( .A1(net_6696), .ZN(net_3119), .A2(net_3118) );
NAND2_X2 inst_9206 ( .ZN(net_19505), .A2(net_11277), .A1(net_1244) );
AOI21_X2 inst_20838 ( .ZN(net_9283), .B1(net_9282), .A(net_6181), .B2(net_3471) );
OAI21_X2 inst_1894 ( .ZN(net_13365), .B1(net_9851), .B2(net_8513), .A(net_1471) );
INV_X4 inst_13960 ( .ZN(net_6746), .A(net_6745) );
NAND3_X2 inst_6707 ( .ZN(net_7114), .A3(net_7113), .A1(net_4318), .A2(net_3431) );
INV_X4 inst_15401 ( .ZN(net_15926), .A(net_15688) );
NOR2_X2 inst_4643 ( .A1(net_3592), .ZN(net_3392), .A2(net_3391) );
INV_X4 inst_14379 ( .A(net_6807), .ZN(net_6289) );
NAND3_X2 inst_6636 ( .ZN(net_8974), .A3(net_8973), .A2(net_6828), .A1(net_5711) );
CLKBUF_X2 inst_22129 ( .A(net_22000), .Z(net_22001) );
INV_X4 inst_13677 ( .ZN(net_9134), .A(net_8003) );
NOR3_X2 inst_2701 ( .ZN(net_13959), .A1(net_11919), .A2(net_11212), .A3(net_7851) );
NAND2_X2 inst_8321 ( .A1(net_20070), .ZN(net_17562), .A2(net_17561) );
NAND2_X2 inst_9171 ( .ZN(net_13354), .A1(net_13353), .A2(net_10535) );
INV_X4 inst_18078 ( .A(net_21084), .ZN(net_527) );
CLKBUF_X2 inst_21739 ( .A(net_21610), .Z(net_21611) );
NAND2_X2 inst_10385 ( .A2(net_10525), .ZN(net_7329), .A1(net_4001) );
NOR2_X4 inst_3165 ( .ZN(net_3846), .A2(net_2568), .A1(net_993) );
AOI21_X4 inst_20125 ( .ZN(net_19568), .B1(net_19331), .B2(net_15110), .A(net_14012) );
NAND2_X2 inst_11222 ( .ZN(net_6742), .A2(net_3933), .A1(net_1228) );
XNOR2_X2 inst_575 ( .ZN(net_620), .A(net_619), .B(net_618) );
NAND2_X2 inst_11738 ( .ZN(net_2549), .A1(net_2179), .A2(net_2178) );
NAND2_X2 inst_10151 ( .ZN(net_10375), .A1(net_8286), .A2(net_8285) );
INV_X4 inst_16335 ( .ZN(net_2445), .A(net_1301) );
CLKBUF_X2 inst_21873 ( .A(net_21522), .Z(net_21745) );
INV_X4 inst_18130 ( .A(net_21196), .ZN(net_552) );
XNOR2_X2 inst_627 ( .B(net_15957), .ZN(net_457), .A(net_456) );
INV_X4 inst_14606 ( .ZN(net_7815), .A(net_4435) );
NAND2_X4 inst_6831 ( .ZN(net_18827), .A1(net_18775), .A2(net_18751) );
NOR2_X2 inst_4725 ( .ZN(net_3100), .A1(net_2753), .A2(net_763) );
NOR2_X2 inst_3352 ( .ZN(net_17789), .A2(net_17645), .A1(net_17580) );
XNOR2_X2 inst_344 ( .ZN(net_16961), .A(net_16481), .B(net_471) );
AOI21_X4 inst_20139 ( .ZN(net_16042), .B1(net_16041), .A(net_15812), .B2(net_15230) );
NAND2_X4 inst_6928 ( .A2(net_19641), .A1(net_19640), .ZN(net_19428) );
INV_X4 inst_17285 ( .ZN(net_2630), .A(net_703) );
CLKBUF_X2 inst_22232 ( .A(net_22103), .Z(net_22104) );
NOR2_X2 inst_3818 ( .ZN(net_9797), .A2(net_9699), .A1(net_6236) );
NAND3_X2 inst_5975 ( .ZN(net_14748), .A2(net_14747), .A1(net_12391), .A3(net_12331) );
INV_X4 inst_15209 ( .ZN(net_5106), .A(net_2509) );
OAI221_X2 inst_1338 ( .ZN(net_14772), .A(net_14121), .C1(net_13157), .B2(net_11859), .B1(net_4350), .C2(net_3639) );
DFF_X1 inst_19924 ( .QN(net_21115), .D(net_13207), .CK(net_22197) );
INV_X4 inst_17698 ( .ZN(net_1214), .A(net_251) );
OAI211_X2 inst_2430 ( .ZN(net_15141), .B(net_14533), .C1(net_14346), .C2(net_12087), .A(net_6880) );
INV_X4 inst_13093 ( .ZN(net_15879), .A(net_15752) );
CLKBUF_X2 inst_22585 ( .A(net_21327), .Z(net_22457) );
NOR2_X2 inst_4952 ( .ZN(net_3085), .A2(net_1543), .A1(net_222) );
NOR2_X2 inst_3731 ( .ZN(net_12641), .A2(net_11055), .A1(net_10875) );
INV_X4 inst_13932 ( .ZN(net_8782), .A(net_6857) );
NAND2_X4 inst_6899 ( .ZN(net_17995), .A1(net_17896), .A2(net_17847) );
NOR2_X2 inst_4839 ( .ZN(net_2370), .A1(net_1728), .A2(net_706) );
OAI21_X2 inst_2028 ( .ZN(net_11314), .B2(net_9635), .B1(net_6256), .A(net_4032) );
INV_X4 inst_15364 ( .A(net_15522), .ZN(net_3433) );
CLKBUF_X2 inst_21610 ( .A(net_21481), .Z(net_21482) );
INV_X2 inst_19369 ( .ZN(net_2211), .A(net_2210) );
NAND2_X2 inst_8381 ( .ZN(net_17343), .A2(net_17079), .A1(net_16991) );
INV_X4 inst_15038 ( .ZN(net_19299), .A(net_4991) );
AND2_X2 inst_21335 ( .ZN(net_14931), .A1(net_8865), .A2(net_4302) );
INV_X4 inst_16409 ( .ZN(net_1715), .A(net_822) );
INV_X4 inst_16994 ( .A(net_14945), .ZN(net_872) );
INV_X4 inst_14904 ( .ZN(net_7681), .A(net_3600) );
AOI21_X2 inst_20487 ( .ZN(net_14790), .A(net_14557), .B2(net_13251), .B1(net_10044) );
SDFF_X2 inst_722 ( .Q(net_20900), .SE(net_18804), .SI(net_18575), .D(net_594), .CK(net_22262) );
NAND3_X2 inst_6019 ( .ZN(net_20830), .A3(net_12622), .A2(net_12368), .A1(net_8609) );
NAND2_X2 inst_8093 ( .A1(net_20443), .ZN(net_19138), .A2(net_18128) );
NAND2_X2 inst_9502 ( .ZN(net_11342), .A1(net_8270), .A2(net_6764) );
NOR2_X2 inst_4232 ( .ZN(net_6584), .A2(net_6583), .A1(net_3810) );
NOR2_X2 inst_4270 ( .A1(net_7975), .ZN(net_7542), .A2(net_6133) );
NOR2_X4 inst_3010 ( .ZN(net_7952), .A1(net_5652), .A2(net_2273) );
INV_X4 inst_16726 ( .ZN(net_1375), .A(net_876) );
NAND2_X2 inst_8010 ( .ZN(net_18297), .A2(net_18199), .A1(net_17742) );
INV_X4 inst_17151 ( .A(net_2456), .ZN(net_757) );
INV_X8 inst_12282 ( .ZN(net_8222), .A(net_1477) );
NOR2_X4 inst_3133 ( .A1(net_4863), .ZN(net_4822), .A2(net_3829) );
NAND2_X2 inst_8207 ( .ZN(net_17865), .A1(net_17710), .A2(net_17614) );
NAND3_X2 inst_6412 ( .ZN(net_11954), .A2(net_10160), .A1(net_7081), .A3(net_5072) );
OAI211_X2 inst_2588 ( .B(net_6391), .ZN(net_6385), .A(net_6384), .C1(net_2503), .C2(net_1325) );
NAND3_X2 inst_6547 ( .ZN(net_10538), .A3(net_10477), .A2(net_9714), .A1(net_3840) );
INV_X4 inst_15844 ( .ZN(net_7378), .A(net_1840) );
INV_X4 inst_15859 ( .ZN(net_2116), .A(net_1812) );
NAND2_X2 inst_7724 ( .ZN(net_18832), .A2(net_18788), .A1(net_17728) );
INV_X4 inst_17671 ( .A(net_20860), .ZN(net_539) );
NAND2_X4 inst_6994 ( .ZN(net_17348), .A1(net_16738), .A2(net_16592) );
AOI21_X2 inst_20738 ( .B2(net_18979), .B1(net_18978), .ZN(net_11456), .A(net_1266) );
NOR2_X2 inst_4665 ( .ZN(net_4708), .A1(net_2751), .A2(net_2481) );
INV_X4 inst_15379 ( .ZN(net_12339), .A(net_10659) );
INV_X4 inst_18142 ( .A(net_21023), .ZN(net_485) );
INV_X2 inst_19695 ( .A(net_20550), .ZN(net_20549) );
INV_X4 inst_18209 ( .A(net_21073), .ZN(net_479) );
INV_X2 inst_18837 ( .ZN(net_6739), .A(net_6738) );
NAND3_X2 inst_5712 ( .ZN(net_16169), .A3(net_15789), .A2(net_15755), .A1(net_15024) );
NAND3_X4 inst_5562 ( .ZN(net_16000), .A1(net_15698), .A3(net_15627), .A2(net_7142) );
NAND4_X2 inst_5374 ( .ZN(net_15229), .A2(net_14331), .A4(net_14067), .A1(net_12347), .A3(net_10277) );
NOR2_X2 inst_4466 ( .A1(net_5677), .ZN(net_4496), .A2(net_4495) );
CLKBUF_X2 inst_22214 ( .A(net_22085), .Z(net_22086) );
INV_X2 inst_19219 ( .ZN(net_3471), .A(net_3470) );
NAND2_X2 inst_11058 ( .ZN(net_4620), .A2(net_4619), .A1(net_976) );
INV_X4 inst_15543 ( .A(net_16281), .ZN(net_15976) );
NAND2_X2 inst_11035 ( .ZN(net_7731), .A1(net_4264), .A2(net_2805) );
CLKBUF_X2 inst_22350 ( .A(net_22221), .Z(net_22222) );
NOR2_X4 inst_2875 ( .ZN(net_20111), .A2(net_9411), .A1(net_8903) );
NAND2_X2 inst_8447 ( .A1(net_20435), .ZN(net_19397), .A2(net_17103) );
AOI21_X2 inst_20598 ( .ZN(net_13867), .B2(net_10256), .B1(net_7253), .A(net_6557) );
DFF_X1 inst_19922 ( .Q(net_21110), .D(net_14397), .CK(net_22200) );
NAND2_X2 inst_9067 ( .ZN(net_13983), .A1(net_13544), .A2(net_12010) );
NAND2_X2 inst_11084 ( .ZN(net_4414), .A2(net_4413), .A1(net_4200) );
NAND2_X2 inst_10341 ( .ZN(net_7529), .A1(net_7528), .A2(net_4497) );
NAND2_X4 inst_7162 ( .ZN(net_9505), .A1(net_9504), .A2(net_2744) );
NAND2_X2 inst_9396 ( .A2(net_12923), .ZN(net_11703), .A1(net_11702) );
NAND3_X2 inst_6248 ( .ZN(net_13016), .A3(net_9816), .A1(net_8780), .A2(net_3997) );
NOR2_X2 inst_3389 ( .ZN(net_20421), .A2(net_15984), .A1(net_14502) );
SDFF_X2 inst_782 ( .Q(net_20949), .SE(net_18584), .SI(net_18041), .D(net_590), .CK(net_22630) );
CLKBUF_X2 inst_21693 ( .A(net_21442), .Z(net_21565) );
NAND3_X2 inst_5744 ( .A1(net_20418), .ZN(net_20043), .A3(net_11556), .A2(net_6350) );
NOR2_X4 inst_2869 ( .ZN(net_12649), .A1(net_10962), .A2(net_7509) );
NAND2_X2 inst_10546 ( .A1(net_8707), .A2(net_6851), .ZN(net_6764) );
XOR2_X2 inst_6 ( .A(net_21209), .B(net_20507), .Z(net_17593) );
NAND2_X2 inst_10603 ( .ZN(net_10503), .A1(net_6617), .A2(net_6616) );
INV_X4 inst_16181 ( .ZN(net_10142), .A(net_4113) );
OAI211_X2 inst_2486 ( .ZN(net_13256), .C2(net_11091), .B(net_10067), .A(net_9071), .C1(net_1471) );
NAND4_X2 inst_5461 ( .ZN(net_13331), .A1(net_13330), .A2(net_13010), .A4(net_12838), .A3(net_11708) );
OAI211_X2 inst_2410 ( .ZN(net_15525), .C1(net_15524), .B(net_14560), .C2(net_13941), .A(net_10042) );
INV_X2 inst_19406 ( .ZN(net_1985), .A(net_1984) );
NAND2_X2 inst_11832 ( .A2(net_2686), .ZN(net_1845), .A1(net_61) );
CLKBUF_X2 inst_22058 ( .A(net_21929), .Z(net_21930) );
NAND2_X2 inst_8927 ( .ZN(net_14912), .A2(net_13807), .A1(net_11943) );
NAND2_X2 inst_8728 ( .ZN(net_20117), .A2(net_15773), .A1(net_15681) );
INV_X4 inst_16670 ( .ZN(net_9579), .A(net_8097) );
CLKBUF_X2 inst_22486 ( .A(net_22357), .Z(net_22358) );
INV_X4 inst_12760 ( .ZN(net_17392), .A(net_17391) );
INV_X4 inst_17674 ( .ZN(net_9617), .A(net_242) );
INV_X4 inst_14650 ( .A(net_15561), .ZN(net_4370) );
NAND2_X2 inst_11726 ( .ZN(net_4306), .A2(net_2231), .A1(net_2050) );
INV_X4 inst_17601 ( .A(net_337), .ZN(net_323) );
INV_X4 inst_13030 ( .ZN(net_16734), .A(net_16718) );
AND2_X2 inst_21295 ( .ZN(net_19124), .A1(net_12226), .A2(net_10746) );
NAND2_X2 inst_8108 ( .A1(net_20504), .ZN(net_18110), .A2(net_18086) );
NAND2_X2 inst_8211 ( .ZN(net_17850), .A1(net_17694), .A2(net_17599) );
NAND3_X2 inst_6031 ( .ZN(net_14368), .A3(net_14327), .A2(net_12406), .A1(net_11112) );
CLKBUF_X2 inst_21725 ( .A(net_21303), .Z(net_21597) );
AOI21_X2 inst_20502 ( .ZN(net_14648), .B2(net_12098), .B1(net_8836), .A(net_7693) );
NAND2_X2 inst_7729 ( .ZN(net_18821), .A2(net_18790), .A1(net_17842) );
AOI22_X2 inst_20043 ( .A1(net_9378), .ZN(net_7073), .A2(net_7072), .B1(net_7071), .B2(net_4070) );
SDFF_X2 inst_1026 ( .QN(net_21018), .D(net_574), .SE(net_253), .CK(net_21886), .SI(x2713) );
OAI22_X2 inst_1320 ( .A1(net_6947), .B1(net_5308), .ZN(net_4199), .B2(net_4198), .A2(net_3294) );
INV_X4 inst_15638 ( .ZN(net_14496), .A(net_11345) );
CLKBUF_X2 inst_22008 ( .A(net_21595), .Z(net_21880) );
NAND3_X2 inst_6250 ( .ZN(net_13013), .A1(net_13012), .A3(net_12891), .A2(net_4007) );
NAND2_X2 inst_11289 ( .ZN(net_4824), .A2(net_3834), .A1(net_168) );
CLKBUF_X2 inst_22896 ( .A(net_22767), .Z(net_22768) );
NAND3_X4 inst_5576 ( .A2(net_19283), .A1(net_19282), .ZN(net_15739), .A3(net_15106) );
INV_X4 inst_12826 ( .ZN(net_18470), .A(net_17154) );
NAND4_X4 inst_5246 ( .ZN(net_20118), .A2(net_19183), .A1(net_19182), .A4(net_4559), .A3(net_4372) );
XNOR2_X2 inst_95 ( .ZN(net_18549), .A(net_18448), .B(net_17501) );
NOR2_X2 inst_3376 ( .ZN(net_16493), .A2(net_16391), .A1(net_14492) );
CLKBUF_X2 inst_22468 ( .A(net_22339), .Z(net_22340) );
NOR2_X4 inst_2921 ( .ZN(net_9589), .A1(net_8057), .A2(net_761) );
INV_X4 inst_13058 ( .ZN(net_16371), .A(net_16329) );
NAND2_X2 inst_10622 ( .A1(net_11297), .ZN(net_8645), .A2(net_6579) );
NAND2_X2 inst_10499 ( .A1(net_13198), .ZN(net_6923), .A2(net_6922) );
AND2_X4 inst_21195 ( .A1(net_11886), .A2(net_10435), .ZN(net_10234) );
AOI21_X2 inst_20681 ( .ZN(net_20359), .B1(net_20265), .A(net_9977), .B2(net_8836) );
INV_X4 inst_14794 ( .ZN(net_4002), .A(net_4001) );
INV_X2 inst_18358 ( .A(net_18390), .ZN(net_18350) );
NOR2_X2 inst_4009 ( .ZN(net_8078), .A1(net_6064), .A2(net_3001) );
NAND2_X2 inst_9766 ( .ZN(net_9823), .A1(net_9822), .A2(net_5585) );
NAND2_X2 inst_10870 ( .A1(net_9146), .ZN(net_5431), .A2(net_3555) );
NAND2_X2 inst_8071 ( .A2(net_20794), .ZN(net_20324), .A1(net_17103) );
AOI21_X2 inst_20358 ( .ZN(net_15686), .A(net_15184), .B1(net_14600), .B2(net_14581) );
NAND2_X2 inst_8297 ( .ZN(net_17606), .A2(net_17418), .A1(net_13298) );
NOR2_X2 inst_4900 ( .A1(net_14378), .ZN(net_1993), .A2(net_1068) );
INV_X4 inst_13325 ( .ZN(net_11326), .A(net_10013) );
NAND3_X2 inst_5837 ( .ZN(net_15510), .A2(net_14725), .A1(net_14639), .A3(net_14577) );
NAND4_X2 inst_5394 ( .ZN(net_14823), .A4(net_13360), .A1(net_12041), .A2(net_11488), .A3(net_8960) );
NAND2_X4 inst_7194 ( .A2(net_20211), .ZN(net_9818), .A1(net_9478) );
INV_X4 inst_13883 ( .A(net_9536), .ZN(net_9212) );
AOI21_X4 inst_20130 ( .B1(net_20084), .ZN(net_16118), .A(net_15350), .B2(net_2573) );
NAND2_X4 inst_7537 ( .ZN(net_19462), .A1(net_2315), .A2(net_1270) );
INV_X4 inst_17317 ( .ZN(net_14014), .A(net_13530) );
NAND2_X2 inst_10407 ( .A2(net_11766), .ZN(net_7265), .A1(net_7264) );
AOI221_X2 inst_20093 ( .ZN(net_14347), .B1(net_14346), .C1(net_13274), .B2(net_12624), .A(net_9474), .C2(net_9272) );
INV_X2 inst_19126 ( .ZN(net_5147), .A(net_3130) );
AOI21_X2 inst_20375 ( .ZN(net_19937), .B2(net_19409), .B1(net_19408), .A(net_15166) );
INV_X8 inst_12369 ( .ZN(net_4394), .A(net_304) );
INV_X2 inst_19154 ( .ZN(net_6936), .A(net_4044) );
NAND2_X2 inst_8955 ( .A1(net_14731), .ZN(net_14718), .A2(net_13214) );
NOR2_X2 inst_4901 ( .A1(net_4394), .ZN(net_4175), .A2(net_1116) );
INV_X4 inst_14758 ( .ZN(net_6931), .A(net_4063) );
NOR2_X2 inst_3590 ( .A1(net_19996), .ZN(net_12611), .A2(net_7219) );
INV_X2 inst_19319 ( .A(net_3758), .ZN(net_2616) );
INV_X2 inst_18783 ( .A(net_8475), .ZN(net_7505) );
INV_X4 inst_18071 ( .A(net_21025), .ZN(net_650) );
INV_X4 inst_17594 ( .A(net_20876), .ZN(net_2253) );
INV_X2 inst_18830 ( .ZN(net_6780), .A(net_6779) );
NAND2_X2 inst_8145 ( .ZN(net_18020), .A2(net_17963), .A1(net_17592) );
NAND2_X2 inst_9252 ( .A1(net_15664), .ZN(net_12663), .A2(net_12662) );
INV_X2 inst_19305 ( .ZN(net_2738), .A(net_2737) );
NOR2_X2 inst_4974 ( .ZN(net_2453), .A2(net_1561), .A1(net_1376) );
NAND2_X2 inst_8582 ( .A2(net_20072), .ZN(net_16720), .A1(net_16519) );
NAND2_X2 inst_10836 ( .ZN(net_15565), .A1(net_5482), .A2(net_5481) );
INV_X4 inst_18189 ( .A(net_21144), .ZN(net_631) );
CLKBUF_X2 inst_21917 ( .A(net_21788), .Z(net_21789) );
OAI211_X2 inst_2476 ( .ZN(net_13622), .A(net_13621), .C2(net_13620), .C1(net_13565), .B(net_10992) );
INV_X4 inst_16660 ( .ZN(net_19757), .A(net_1084) );
NAND2_X2 inst_12078 ( .A2(net_2712), .ZN(net_787), .A1(net_271) );
NAND2_X2 inst_8116 ( .A2(net_20442), .ZN(net_19207), .A1(net_16662) );
INV_X4 inst_18305 ( .A(net_20495), .ZN(net_20490) );
NOR2_X2 inst_4502 ( .ZN(net_5383), .A1(net_4250), .A2(net_4249) );
AOI21_X2 inst_20696 ( .ZN(net_12156), .B2(net_8040), .A(net_6922), .B1(net_5415) );
INV_X4 inst_14258 ( .ZN(net_8762), .A(net_5746) );
NAND3_X4 inst_5624 ( .A1(net_20753), .ZN(net_11568), .A3(net_8278), .A2(net_8068) );
NAND2_X4 inst_7451 ( .ZN(net_6674), .A2(net_3060), .A1(net_2529) );
INV_X2 inst_19328 ( .ZN(net_4336), .A(net_2552) );
INV_X2 inst_19226 ( .ZN(net_6019), .A(net_3431) );
NAND2_X4 inst_7458 ( .ZN(net_9295), .A2(net_2828), .A1(net_2827) );
INV_X4 inst_14072 ( .A(net_7992), .ZN(net_7576) );
SDFF_X2 inst_1036 ( .QN(net_21003), .D(net_1874), .SE(net_263), .CK(net_21879), .SI(x3001) );
CLKBUF_X2 inst_22560 ( .A(net_22375), .Z(net_22432) );
NAND2_X2 inst_10094 ( .A1(net_10488), .ZN(net_8617), .A2(net_7893) );
NAND2_X2 inst_10334 ( .A1(net_9903), .ZN(net_7582), .A2(net_7581) );
NAND2_X2 inst_8653 ( .A1(net_21109), .ZN(net_16555), .A2(net_16554) );
NAND3_X2 inst_5694 ( .ZN(net_16257), .A3(net_15952), .A2(net_12302), .A1(net_11730) );
INV_X4 inst_14700 ( .ZN(net_18585), .A(net_18025) );
NAND2_X1 inst_12141 ( .A2(net_20434), .ZN(net_19398), .A1(net_17104) );
NOR2_X2 inst_4613 ( .ZN(net_6353), .A1(net_3356), .A2(net_2651) );
NAND3_X2 inst_5852 ( .ZN(net_15422), .A3(net_14394), .A2(net_11168), .A1(net_5885) );
AOI22_X2 inst_19966 ( .ZN(net_15927), .A1(net_15926), .A2(net_15231), .B2(net_13850), .B1(net_3338) );
OAI211_X4 inst_2376 ( .B(net_20608), .A(net_20607), .ZN(net_16222), .C1(net_15880), .C2(net_15479) );
CLKBUF_X2 inst_22649 ( .A(net_22520), .Z(net_22521) );
NAND2_X2 inst_7925 ( .ZN(net_18448), .A1(net_18340), .A2(net_18284) );
NAND2_X4 inst_7496 ( .A1(net_20875), .ZN(net_7109), .A2(net_2325) );
NAND2_X4 inst_7050 ( .ZN(net_16420), .A1(net_16344), .A2(net_16247) );
NOR2_X2 inst_4360 ( .ZN(net_5558), .A1(net_5557), .A2(net_5556) );
INV_X2 inst_19086 ( .ZN(net_4574), .A(net_4573) );
SDFF_X2 inst_860 ( .Q(net_21157), .D(net_17172), .SE(net_263), .CK(net_21476), .SI(x5464) );
XNOR2_X2 inst_563 ( .ZN(net_677), .A(net_676), .B(net_675) );
INV_X4 inst_14074 ( .ZN(net_6228), .A(net_6227) );
NOR2_X2 inst_3962 ( .ZN(net_19892), .A1(net_8590), .A2(net_5296) );
SDFF_X2 inst_943 ( .QN(net_21044), .D(net_467), .SE(net_263), .CK(net_22527), .SI(x2260) );
NAND4_X2 inst_5314 ( .ZN(net_20191), .A4(net_15083), .A2(net_14480), .A1(net_14366), .A3(net_10658) );
INV_X4 inst_15714 ( .A(net_15842), .ZN(net_13138) );
CLKBUF_X2 inst_22341 ( .A(net_21336), .Z(net_22213) );
INV_X2 inst_18979 ( .ZN(net_5156), .A(net_5155) );
NOR2_X2 inst_4711 ( .ZN(net_9834), .A1(net_6812), .A2(net_1585) );
OAI21_X2 inst_1964 ( .A(net_14476), .ZN(net_12357), .B1(net_7641), .B2(net_7358) );
NAND2_X1 inst_12151 ( .A1(net_11878), .A2(net_10620), .ZN(net_10327) );
NAND2_X4 inst_7464 ( .ZN(net_4735), .A2(net_3402), .A1(net_2146) );
OAI21_X2 inst_1765 ( .ZN(net_14703), .B2(net_12039), .A(net_11541), .B1(net_9789) );
CLKBUF_X2 inst_21684 ( .A(net_21497), .Z(net_21556) );
INV_X2 inst_18908 ( .ZN(net_7497), .A(net_6048) );
INV_X2 inst_18657 ( .A(net_11104), .ZN(net_9210) );
CLKBUF_X2 inst_22418 ( .A(net_22289), .Z(net_22290) );
INV_X4 inst_13525 ( .ZN(net_14211), .A(net_9332) );
NAND3_X2 inst_6357 ( .ZN(net_12090), .A3(net_11912), .A1(net_8374), .A2(net_3999) );
NAND2_X2 inst_11944 ( .A2(net_1563), .ZN(net_1440), .A1(net_165) );
INV_X4 inst_17279 ( .ZN(net_7439), .A(net_152) );
INV_X4 inst_16231 ( .ZN(net_15677), .A(net_10252) );
XNOR2_X2 inst_178 ( .ZN(net_17772), .A(net_17771), .B(net_9240) );
INV_X2 inst_18588 ( .ZN(net_11577), .A(net_10232) );
NAND2_X2 inst_9179 ( .ZN(net_13338), .A1(net_10709), .A2(net_10579) );
INV_X2 inst_19323 ( .ZN(net_2599), .A(net_2598) );
AOI21_X2 inst_20790 ( .ZN(net_10543), .B2(net_8712), .B1(net_7018), .A(net_816) );
NAND2_X2 inst_8257 ( .A2(net_17851), .ZN(net_17696), .A1(net_17695) );
NAND3_X2 inst_5941 ( .ZN(net_14903), .A2(net_14902), .A3(net_14873), .A1(net_10021) );
INV_X4 inst_13562 ( .ZN(net_12361), .A(net_9150) );
OR2_X2 inst_1148 ( .A1(net_9925), .ZN(net_9850), .A2(net_9849) );
NOR2_X2 inst_3919 ( .A2(net_10499), .A1(net_10415), .ZN(net_8797) );
INV_X4 inst_17643 ( .ZN(net_606), .A(net_275) );
CLKBUF_X2 inst_22142 ( .A(net_22013), .Z(net_22014) );
NAND2_X2 inst_10292 ( .ZN(net_7916), .A1(net_7915), .A2(net_5902) );
NOR2_X2 inst_4350 ( .ZN(net_19305), .A1(net_3846), .A2(net_2935) );
NAND2_X2 inst_8270 ( .ZN(net_17654), .A1(net_17653), .A2(net_17550) );
AOI21_X2 inst_20446 ( .ZN(net_15102), .A(net_15058), .B1(net_14314), .B2(net_13111) );
INV_X2 inst_18467 ( .A(net_13819), .ZN(net_12729) );
CLKBUF_X2 inst_21644 ( .A(net_21515), .Z(net_21516) );
AOI21_X2 inst_20648 ( .ZN(net_13069), .B2(net_11582), .B1(net_11366), .A(net_8300) );
NAND2_X2 inst_9659 ( .A1(net_11384), .ZN(net_10334), .A2(net_7759) );
NAND3_X2 inst_6004 ( .ZN(net_14427), .A3(net_12452), .A1(net_7856), .A2(net_2749) );
SDFF_X2 inst_842 ( .Q(net_21146), .SI(net_17318), .SE(net_125), .CK(net_22162), .D(x3416) );
CLKBUF_X2 inst_22289 ( .A(net_22160), .Z(net_22161) );
OAI21_X2 inst_2068 ( .ZN(net_10660), .A(net_10659), .B2(net_8655), .B1(net_6341) );
NAND2_X2 inst_9897 ( .ZN(net_13802), .A2(net_12757), .A1(net_2884) );
INV_X2 inst_19652 ( .A(net_20076), .ZN(net_20075) );
XNOR2_X2 inst_551 ( .B(net_11872), .ZN(net_715), .A(net_714) );
NAND2_X2 inst_9697 ( .ZN(net_10223), .A2(net_9576), .A1(net_8460) );
INV_X4 inst_17577 ( .ZN(net_866), .A(net_761) );
OAI21_X2 inst_2101 ( .A(net_12712), .ZN(net_10065), .B1(net_9250), .B2(net_6171) );
XNOR2_X2 inst_353 ( .A(net_16983), .ZN(net_16933), .B(net_16094) );
INV_X2 inst_19132 ( .A(net_4902), .ZN(net_4191) );
NOR2_X2 inst_3808 ( .ZN(net_9836), .A1(net_8397), .A2(net_5931) );
INV_X4 inst_15721 ( .ZN(net_2551), .A(net_1709) );
INV_X2 inst_18819 ( .ZN(net_6974), .A(net_6973) );
OAI21_X2 inst_1940 ( .B1(net_12911), .ZN(net_12850), .A(net_8353), .B2(net_761) );
NAND3_X2 inst_6286 ( .ZN(net_12845), .A3(net_12844), .A2(net_10575), .A1(net_9780) );
INV_X4 inst_16770 ( .ZN(net_15366), .A(net_15077) );
NOR2_X2 inst_4632 ( .A2(net_5288), .ZN(net_4517), .A1(net_3546) );
NAND2_X2 inst_8492 ( .A1(net_19444), .ZN(net_16955), .A2(net_16954) );
NAND2_X2 inst_10400 ( .ZN(net_13815), .A1(net_11645), .A2(net_6858) );
INV_X4 inst_13456 ( .A(net_11941), .ZN(net_11487) );
INV_X4 inst_15025 ( .A(net_14078), .ZN(net_3370) );
NAND3_X2 inst_6212 ( .ZN(net_13270), .A3(net_8857), .A2(net_8078), .A1(net_8058) );
INV_X4 inst_13917 ( .A(net_11943), .ZN(net_8247) );
NOR2_X2 inst_4041 ( .ZN(net_11775), .A1(net_7903), .A2(net_7902) );
INV_X4 inst_13761 ( .ZN(net_10975), .A(net_9640) );
NAND2_X2 inst_9559 ( .ZN(net_13679), .A2(net_10995), .A1(net_10031) );
INV_X4 inst_14184 ( .ZN(net_11218), .A(net_5983) );
INV_X4 inst_13869 ( .A(net_9460), .ZN(net_9115) );
INV_X4 inst_14588 ( .ZN(net_5783), .A(net_4477) );
NAND3_X2 inst_6745 ( .ZN(net_6386), .A2(net_4974), .A3(net_4136), .A1(net_3003) );
NAND2_X2 inst_11321 ( .ZN(net_6552), .A1(net_3758), .A2(net_3757) );
CLKBUF_X2 inst_21954 ( .A(net_21346), .Z(net_21826) );
AOI21_X4 inst_20113 ( .B2(net_20944), .B1(net_19993), .ZN(net_16318), .A(net_12130) );
CLKBUF_X2 inst_21659 ( .A(net_21530), .Z(net_21531) );
INV_X4 inst_14064 ( .ZN(net_9761), .A(net_7781) );
AOI21_X2 inst_20714 ( .ZN(net_12043), .A(net_8325), .B2(net_7737), .B1(net_7230) );
INV_X2 inst_18824 ( .A(net_8965), .ZN(net_6881) );
INV_X4 inst_17626 ( .ZN(net_1289), .A(net_1080) );
INV_X4 inst_13980 ( .ZN(net_7880), .A(net_5394) );
AND3_X2 inst_21130 ( .ZN(net_15428), .A2(net_15427), .A1(net_14988), .A3(net_8218) );
INV_X4 inst_12624 ( .ZN(net_20651), .A(net_17984) );
NAND2_X4 inst_7134 ( .ZN(net_14535), .A1(net_9735), .A2(net_9614) );
NOR2_X2 inst_3370 ( .ZN(net_17616), .A2(net_16498), .A1(net_16430) );
NAND2_X2 inst_10168 ( .ZN(net_9711), .A1(net_8232), .A2(net_6159) );
INV_X4 inst_15301 ( .ZN(net_3428), .A(net_2688) );
NAND2_X2 inst_8993 ( .ZN(net_14459), .A1(net_14458), .A2(net_12946) );
NAND3_X2 inst_6579 ( .ZN(net_10443), .A3(net_10442), .A1(net_6697), .A2(net_5828) );
NAND2_X4 inst_7210 ( .ZN(net_11979), .A1(net_6068), .A2(net_4207) );
SDFF_X2 inst_901 ( .Q(net_21214), .SI(net_16765), .SE(net_125), .CK(net_22281), .D(x7558) );
NAND2_X2 inst_10992 ( .ZN(net_4925), .A2(net_4076), .A1(net_1058) );
NAND2_X4 inst_7261 ( .ZN(net_7861), .A2(net_7597), .A1(net_4879) );
NAND3_X2 inst_6094 ( .ZN(net_13929), .A3(net_13854), .A1(net_12545), .A2(net_9649) );
CLKBUF_X2 inst_22597 ( .A(net_22007), .Z(net_22469) );
INV_X4 inst_13821 ( .ZN(net_10894), .A(net_7510) );
NAND2_X2 inst_9957 ( .ZN(net_19851), .A1(net_8918), .A2(net_5606) );
NAND2_X2 inst_10863 ( .ZN(net_10488), .A1(net_5435), .A2(net_5434) );
INV_X2 inst_19718 ( .ZN(net_20780), .A(net_20779) );
INV_X4 inst_14843 ( .ZN(net_6624), .A(net_3849) );
OAI211_X2 inst_2403 ( .ZN(net_20612), .C1(net_15864), .B(net_15331), .A(net_13672), .C2(net_13245) );
NOR2_X2 inst_4948 ( .ZN(net_2669), .A1(net_2202), .A2(net_1219) );
NAND2_X2 inst_9104 ( .A1(net_14751), .ZN(net_13732), .A2(net_11715) );
INV_X4 inst_14545 ( .A(net_14083), .ZN(net_5758) );
AND3_X2 inst_21139 ( .A2(net_12137), .ZN(net_11262), .A3(net_5198), .A1(net_4245) );
CLKBUF_X2 inst_21825 ( .A(net_21696), .Z(net_21697) );
NOR2_X4 inst_3098 ( .ZN(net_5519), .A1(net_4207), .A2(net_4206) );
INV_X4 inst_13834 ( .ZN(net_9163), .A(net_7493) );
NAND2_X2 inst_10679 ( .A1(net_10114), .ZN(net_6183), .A2(net_6182) );
CLKBUF_X2 inst_22761 ( .A(net_22632), .Z(net_22633) );
NAND3_X2 inst_6144 ( .ZN(net_19147), .A1(net_12360), .A2(net_9111), .A3(net_6664) );
NOR2_X2 inst_5013 ( .A1(net_20548), .ZN(net_6097), .A2(net_1259) );
CLKBUF_X2 inst_21422 ( .A(net_21245), .Z(net_21294) );
CLKBUF_X2 inst_22381 ( .A(net_22252), .Z(net_22253) );
NAND2_X2 inst_12034 ( .ZN(net_974), .A1(net_973), .A2(net_525) );
CLKBUF_X2 inst_21572 ( .A(net_21443), .Z(net_21444) );
NAND3_X2 inst_5910 ( .ZN(net_15023), .A3(net_13040), .A2(net_12596), .A1(net_10666) );
SDFF_X2 inst_928 ( .Q(net_21156), .D(net_16505), .SE(net_263), .CK(net_21517), .SI(x5505) );
INV_X4 inst_15782 ( .ZN(net_3211), .A(net_1631) );
NAND2_X2 inst_10695 ( .A1(net_9401), .ZN(net_6072), .A2(net_6071) );
INV_X4 inst_17828 ( .ZN(net_931), .A(net_106) );
OAI21_X2 inst_1539 ( .ZN(net_17904), .B2(net_17851), .A(net_17700), .B1(net_17699) );
NOR3_X2 inst_2662 ( .ZN(net_19870), .A2(net_19000), .A1(net_18999), .A3(net_12045) );
INV_X4 inst_16309 ( .A(net_7129), .ZN(net_5509) );
INV_X4 inst_18035 ( .A(net_20850), .ZN(net_102) );
OAI21_X2 inst_1718 ( .B2(net_20269), .B1(net_20268), .ZN(net_19264), .A(net_14104) );
INV_X2 inst_18912 ( .ZN(net_6022), .A(net_6021) );
NAND2_X2 inst_9424 ( .ZN(net_11618), .A1(net_11617), .A2(net_9685) );
NAND2_X2 inst_8549 ( .ZN(net_16795), .A1(net_16794), .A2(net_16451) );
INV_X2 inst_18385 ( .ZN(net_17189), .A(net_16911) );
NAND2_X2 inst_11126 ( .A1(net_7129), .ZN(net_5452), .A2(net_4313) );
INV_X4 inst_16779 ( .ZN(net_10590), .A(net_5414) );
NAND2_X4 inst_7654 ( .ZN(net_1348), .A1(net_981), .A2(net_916) );
AND2_X4 inst_21217 ( .ZN(net_11368), .A2(net_6019), .A1(net_5265) );
OAI22_X2 inst_1296 ( .A1(net_13095), .A2(net_12910), .ZN(net_11851), .B1(net_10389), .B2(net_7043) );
INV_X4 inst_14443 ( .A(net_6436), .ZN(net_4988) );
NOR2_X2 inst_3671 ( .ZN(net_20229), .A1(net_11493), .A2(net_11492) );
INV_X4 inst_17781 ( .A(net_6078), .ZN(net_142) );
NAND2_X2 inst_7978 ( .ZN(net_18346), .A2(net_18245), .A1(net_17260) );
AND2_X2 inst_21330 ( .ZN(net_19821), .A1(net_9360), .A2(net_5210) );
INV_X4 inst_13121 ( .ZN(net_15472), .A(net_15210) );
AND4_X2 inst_21097 ( .A4(net_13746), .ZN(net_13649), .A2(net_13648), .A1(net_8384), .A3(net_3749) );
NOR2_X2 inst_4513 ( .A2(net_7700), .A1(net_5435), .ZN(net_4186) );
CLKBUF_X2 inst_22525 ( .A(net_22396), .Z(net_22397) );
AOI21_X2 inst_20403 ( .ZN(net_15350), .B2(net_13773), .B1(net_12362), .A(net_2573) );
CLKBUF_X2 inst_21446 ( .A(net_21317), .Z(net_21318) );
INV_X4 inst_15078 ( .ZN(net_3636), .A(net_3268) );
NAND3_X2 inst_6290 ( .A3(net_20292), .ZN(net_12834), .A1(net_12833), .A2(net_12752) );
NAND2_X2 inst_10855 ( .ZN(net_5881), .A1(net_5458), .A2(net_2858) );
INV_X4 inst_17339 ( .ZN(net_555), .A(net_170) );
NOR2_X2 inst_4452 ( .ZN(net_10068), .A1(net_5157), .A2(net_2824) );
NAND2_X2 inst_10633 ( .A1(net_20124), .ZN(net_19110), .A2(net_4410) );
CLKBUF_X2 inst_22844 ( .A(net_21847), .Z(net_22716) );
NAND2_X2 inst_9954 ( .A1(net_9829), .ZN(net_8932), .A2(net_8931) );
NOR2_X2 inst_4151 ( .A1(net_7260), .ZN(net_6903), .A2(net_6902) );
OAI21_X2 inst_1825 ( .ZN(net_14143), .B2(net_10519), .B1(net_10215), .A(net_1006) );
OAI21_X2 inst_1606 ( .ZN(net_16148), .B2(net_15717), .A(net_15370), .B1(net_12851) );
NOR2_X4 inst_2851 ( .ZN(net_13288), .A2(net_10722), .A1(net_10647) );
AND2_X2 inst_21276 ( .ZN(net_13809), .A1(net_13808), .A2(net_13705) );
NAND3_X4 inst_5619 ( .ZN(net_12622), .A2(net_11465), .A3(net_11464), .A1(net_9745) );
NOR2_X2 inst_5126 ( .ZN(net_267), .A1(net_129), .A2(net_128) );
XNOR2_X2 inst_410 ( .ZN(net_16623), .A(net_16622), .B(net_15960) );
XNOR2_X2 inst_316 ( .A(net_17086), .ZN(net_17072), .B(net_16680) );
OR2_X2 inst_1174 ( .A1(net_11214), .ZN(net_5890), .A2(net_5889) );
INV_X4 inst_12860 ( .ZN(net_17044), .A(net_16893) );
AOI21_X4 inst_20168 ( .B1(net_19343), .ZN(net_15627), .B2(net_14279), .A(net_9736) );
SDFF_X2 inst_1023 ( .QN(net_21014), .D(net_641), .SE(net_263), .CK(net_21832), .SI(x2802) );
INV_X4 inst_16665 ( .ZN(net_4840), .A(net_61) );
CLKBUF_X2 inst_22543 ( .A(net_22414), .Z(net_22415) );
INV_X4 inst_17509 ( .A(net_6669), .ZN(net_2344) );
XNOR2_X1 inst_678 ( .ZN(net_18650), .A(net_18649), .B(net_17019) );
NAND2_X2 inst_8515 ( .ZN(net_16915), .A1(net_16783), .A2(net_16590) );
INV_X4 inst_17429 ( .A(net_3890), .ZN(net_1759) );
INV_X2 inst_19505 ( .ZN(net_2079), .A(net_1236) );
NOR2_X2 inst_4359 ( .ZN(net_5566), .A1(net_5565), .A2(net_5564) );
INV_X4 inst_16936 ( .ZN(net_5570), .A(net_925) );
CLKBUF_X2 inst_22373 ( .A(net_22244), .Z(net_22245) );
NAND2_X4 inst_7310 ( .ZN(net_12245), .A1(net_5481), .A2(net_4194) );
INV_X4 inst_13177 ( .ZN(net_14352), .A(net_13868) );
INV_X4 inst_15765 ( .A(net_3196), .ZN(net_2783) );
CLKBUF_X2 inst_21805 ( .A(net_21676), .Z(net_21677) );
NAND2_X2 inst_8033 ( .ZN(net_18337), .A2(net_18186), .A1(net_18161) );
INV_X8 inst_12191 ( .ZN(net_16574), .A(net_16379) );
AOI21_X2 inst_20457 ( .ZN(net_15040), .A(net_15039), .B2(net_12827), .B1(net_9266) );
OAI21_X2 inst_1946 ( .ZN(net_12591), .B1(net_11204), .B2(net_9189), .A(net_8393) );
NAND2_X2 inst_10472 ( .A2(net_7113), .ZN(net_6987), .A1(net_6986) );
NAND2_X2 inst_8686 ( .ZN(net_16848), .A2(net_16365), .A1(net_13656) );
NAND4_X2 inst_5322 ( .ZN(net_15729), .A4(net_14971), .A1(net_14969), .A2(net_14669), .A3(net_13808) );
NAND2_X2 inst_9226 ( .ZN(net_19354), .A2(net_10163), .A1(net_4522) );
NAND2_X2 inst_9786 ( .A1(net_11681), .ZN(net_11102), .A2(net_9750) );
NAND2_X2 inst_9073 ( .ZN(net_19972), .A1(net_12146), .A2(net_10176) );
NOR2_X2 inst_3457 ( .A2(net_20253), .A1(net_20252), .ZN(net_19649) );
INV_X4 inst_12996 ( .A(net_16802), .ZN(net_16487) );
XNOR2_X1 inst_688 ( .A(net_16979), .ZN(net_16934), .B(net_16098) );
CLKBUF_X2 inst_21579 ( .A(net_21450), .Z(net_21451) );
OAI211_X2 inst_2549 ( .ZN(net_10820), .B(net_10819), .C2(net_10818), .A(net_3227), .C1(net_2745) );
CLKBUF_X2 inst_22514 ( .A(net_22385), .Z(net_22386) );
AND2_X2 inst_21355 ( .A1(net_2345), .ZN(net_2122), .A2(net_2121) );
NOR2_X2 inst_3641 ( .ZN(net_12058), .A2(net_10047), .A1(net_8017) );
NOR2_X2 inst_4894 ( .A2(net_20859), .ZN(net_2055), .A1(net_1969) );
AOI21_X2 inst_20963 ( .ZN(net_5310), .A(net_5309), .B1(net_5308), .B2(net_3811) );
OAI211_X2 inst_2387 ( .C1(net_19076), .ZN(net_16294), .A(net_16111), .C2(net_15708), .B(net_15634) );
INV_X4 inst_15372 ( .ZN(net_13848), .A(net_3758) );
INV_X4 inst_16099 ( .ZN(net_2980), .A(net_1514) );
INV_X4 inst_12980 ( .ZN(net_19677), .A(net_16429) );
INV_X4 inst_13351 ( .ZN(net_12624), .A(net_10988) );
INV_X4 inst_14416 ( .ZN(net_7753), .A(net_5070) );
NOR2_X2 inst_4391 ( .ZN(net_6302), .A1(net_5200), .A2(net_3254) );
INV_X4 inst_12474 ( .ZN(net_18753), .A(net_18752) );
NAND2_X2 inst_10137 ( .ZN(net_8327), .A1(net_8326), .A2(net_8325) );
NAND2_X2 inst_10017 ( .ZN(net_12013), .A1(net_10037), .A2(net_8151) );
NAND2_X2 inst_10163 ( .ZN(net_10213), .A2(net_8249), .A1(net_6930) );
NAND3_X2 inst_6423 ( .ZN(net_11940), .A3(net_10235), .A2(net_9190), .A1(net_6382) );
NOR2_X4 inst_3156 ( .ZN(net_4369), .A2(net_3915), .A1(net_3136) );
NOR3_X2 inst_2747 ( .ZN(net_12559), .A2(net_7147), .A1(net_7106), .A3(net_6213) );
INV_X4 inst_13744 ( .ZN(net_9227), .A(net_7633) );
OR2_X2 inst_1220 ( .A1(net_6207), .ZN(net_5675), .A2(net_2829) );
OAI21_X4 inst_1456 ( .A(net_15366), .ZN(net_15293), .B1(net_14857), .B2(net_5723) );
OAI21_X2 inst_2181 ( .A(net_9909), .ZN(net_8844), .B2(net_4819), .B1(net_2662) );
NAND2_X2 inst_8554 ( .ZN(net_19839), .A2(net_16777), .A1(net_5567) );
NAND2_X2 inst_8909 ( .ZN(net_20658), .A1(net_14966), .A2(net_13668) );
INV_X4 inst_16904 ( .ZN(net_10105), .A(net_1253) );
NAND2_X2 inst_8965 ( .A1(net_15858), .ZN(net_14672), .A2(net_13263) );
CLKBUF_X2 inst_22455 ( .A(net_22326), .Z(net_22327) );
NOR2_X1 inst_5154 ( .A2(net_9537), .A1(net_7472), .ZN(net_7435) );
NOR2_X2 inst_4195 ( .A1(net_6842), .ZN(net_6713), .A2(net_6583) );
NAND2_X2 inst_10593 ( .A2(net_7065), .ZN(net_6640), .A1(net_6639) );
NAND2_X2 inst_8473 ( .ZN(net_17016), .A1(net_17015), .A2(net_17014) );
NAND2_X2 inst_9305 ( .ZN(net_19326), .A1(net_10816), .A2(net_9217) );
INV_X4 inst_13605 ( .ZN(net_10974), .A(net_8520) );
NOR2_X2 inst_4440 ( .ZN(net_4809), .A2(net_3131), .A1(net_1231) );
NAND2_X4 inst_7072 ( .A2(net_20844), .A1(net_20843), .ZN(net_19475) );
NAND3_X2 inst_5959 ( .ZN(net_14843), .A2(net_14642), .A3(net_14197), .A1(net_9097) );
NAND2_X2 inst_11607 ( .ZN(net_2619), .A1(net_2618), .A2(net_2617) );
INV_X4 inst_17292 ( .ZN(net_774), .A(net_227) );
NAND2_X2 inst_9149 ( .A1(net_13703), .ZN(net_13402), .A2(net_10640) );
NOR2_X2 inst_4199 ( .ZN(net_19549), .A1(net_11476), .A2(net_9988) );
INV_X4 inst_18174 ( .A(net_21019), .ZN(net_402) );
INV_X4 inst_13588 ( .A(net_10747), .ZN(net_8909) );
INV_X4 inst_14370 ( .ZN(net_9485), .A(net_6742) );
INV_X4 inst_12718 ( .ZN(net_20705), .A(net_17926) );
NAND2_X2 inst_8902 ( .ZN(net_19877), .A1(net_15664), .A2(net_13960) );
NAND3_X2 inst_5749 ( .ZN(net_19045), .A1(net_15816), .A3(net_15455), .A2(net_6768) );
NAND3_X2 inst_6225 ( .ZN(net_13236), .A3(net_13128), .A2(net_9457), .A1(net_5631) );
INV_X4 inst_12754 ( .ZN(net_17598), .A(net_17408) );
NOR2_X2 inst_4420 ( .A1(net_9387), .ZN(net_6141), .A2(net_4987) );
INV_X4 inst_14209 ( .ZN(net_20239), .A(net_5919) );
INV_X4 inst_13795 ( .ZN(net_13490), .A(net_7560) );
SDFF_X1 inst_1057 ( .QN(net_21067), .D(net_668), .SE(net_263), .CK(net_21749), .SI(x1963) );
INV_X4 inst_14097 ( .ZN(net_11379), .A(net_6184) );
NAND2_X2 inst_10359 ( .ZN(net_11971), .A1(net_7432), .A2(net_4561) );
INV_X4 inst_15225 ( .ZN(net_4284), .A(net_2859) );
NAND2_X2 inst_8843 ( .ZN(net_15438), .A2(net_15022), .A1(net_1946) );
INV_X4 inst_17118 ( .ZN(net_11214), .A(net_8868) );
NAND4_X4 inst_5191 ( .A4(net_18918), .A1(net_18917), .ZN(net_16512), .A3(net_16175), .A2(net_14358) );
INV_X4 inst_14565 ( .ZN(net_6215), .A(net_4559) );
AOI21_X2 inst_20895 ( .B1(net_10037), .ZN(net_7783), .A(net_4171), .B2(net_3660) );
NAND3_X4 inst_5602 ( .A3(net_19662), .ZN(net_19082), .A1(net_14448), .A2(net_9945) );
INV_X4 inst_16497 ( .ZN(net_1734), .A(net_1193) );
NAND2_X2 inst_10743 ( .ZN(net_19309), .A1(net_5719), .A2(net_5471) );
INV_X4 inst_17487 ( .ZN(net_3002), .A(net_938) );
SDFF_X2 inst_748 ( .Q(net_20897), .SE(net_18584), .SI(net_18538), .D(net_651), .CK(net_21495) );
NAND2_X2 inst_10610 ( .ZN(net_6602), .A1(net_6601), .A2(net_6600) );
NOR2_X4 inst_2839 ( .ZN(net_20373), .A2(net_19673), .A1(net_19672) );
NAND2_X2 inst_8609 ( .A2(net_16780), .A1(net_16757), .ZN(net_16626) );
NAND3_X2 inst_6730 ( .ZN(net_6486), .A2(net_6485), .A1(net_4190), .A3(net_1621) );
INV_X2 inst_19448 ( .A(net_2060), .ZN(net_1601) );
INV_X4 inst_17097 ( .ZN(net_1495), .A(net_796) );
NAND2_X2 inst_11373 ( .ZN(net_3569), .A1(net_3334), .A2(net_2415) );
NOR2_X2 inst_4582 ( .ZN(net_4860), .A2(net_2851), .A1(net_601) );
NAND2_X2 inst_9266 ( .A2(net_12614), .ZN(net_12613), .A1(net_12612) );
AOI21_X2 inst_20814 ( .A(net_20921), .ZN(net_10084), .B2(net_6043), .B1(net_5295) );
INV_X4 inst_16973 ( .ZN(net_3696), .A(net_903) );
INV_X4 inst_18152 ( .A(net_21214), .ZN(net_790) );
NAND3_X4 inst_5532 ( .A3(net_20445), .ZN(net_17586), .A2(net_16123), .A1(net_14304) );
NOR2_X2 inst_4526 ( .ZN(net_5549), .A2(net_2868), .A1(net_168) );
INV_X4 inst_15700 ( .ZN(net_3514), .A(net_2013) );
NAND2_X2 inst_11070 ( .ZN(net_5922), .A2(net_4864), .A1(net_242) );
INV_X4 inst_17406 ( .A(net_14308), .ZN(net_1030) );
NOR2_X2 inst_4587 ( .ZN(net_4796), .A2(net_3814), .A1(net_3742) );
OAI21_X2 inst_1986 ( .ZN(net_12051), .B1(net_12050), .A(net_10874), .B2(net_7747) );
CLKBUF_X2 inst_21941 ( .A(net_21812), .Z(net_21813) );
OAI21_X2 inst_1949 ( .ZN(net_12575), .B2(net_12574), .A(net_9612), .B1(net_7119) );
NAND3_X2 inst_6170 ( .ZN(net_13613), .A2(net_13582), .A1(net_12381), .A3(net_9564) );
NAND3_X2 inst_5726 ( .ZN(net_16105), .A1(net_15849), .A2(net_10186), .A3(net_8265) );
NAND2_X2 inst_10644 ( .ZN(net_6364), .A1(net_6363), .A2(net_6362) );
NAND2_X1 inst_12163 ( .ZN(net_848), .A1(net_315), .A2(net_129) );
INV_X4 inst_15899 ( .ZN(net_13462), .A(net_6639) );
NAND3_X2 inst_5867 ( .ZN(net_15325), .A3(net_13638), .A2(net_11421), .A1(net_8893) );
NAND2_X2 inst_8243 ( .ZN(net_17803), .A2(net_17555), .A1(net_17467) );
NOR2_X4 inst_2911 ( .ZN(net_9794), .A1(net_8351), .A2(net_8334) );
INV_X4 inst_13770 ( .ZN(net_9216), .A(net_7599) );
AOI21_X2 inst_20635 ( .B1(net_19479), .ZN(net_13342), .B2(net_10785), .A(net_9666) );
AOI21_X2 inst_20474 ( .ZN(net_19270), .A(net_14945), .B1(net_14295), .B2(net_12668) );
OAI21_X2 inst_1859 ( .ZN(net_13807), .B1(net_11092), .A(net_9023), .B2(net_6675) );
NAND2_X2 inst_7734 ( .ZN(net_18814), .A2(net_18768), .A1(net_17636) );
NAND2_X2 inst_8238 ( .ZN(net_17749), .A2(net_17681), .A1(net_17549) );
NOR2_X4 inst_2815 ( .A1(net_20632), .ZN(net_20103), .A2(net_745) );
INV_X4 inst_15818 ( .A(net_11443), .ZN(net_10659) );
AOI21_X2 inst_20748 ( .ZN(net_11373), .A(net_11372), .B1(net_7196), .B2(net_5669) );
NAND2_X2 inst_8267 ( .A1(net_17681), .A2(net_17660), .ZN(net_17657) );
NAND3_X2 inst_5754 ( .ZN(net_16003), .A1(net_15693), .A3(net_15136), .A2(net_10007) );
NOR2_X2 inst_4208 ( .A1(net_6730), .ZN(net_6666), .A2(net_6665) );
NAND2_X2 inst_8426 ( .A1(net_20071), .ZN(net_17180), .A2(net_16615) );
NOR2_X2 inst_3605 ( .A2(net_20211), .ZN(net_19086), .A1(net_12372) );
XNOR2_X2 inst_651 ( .B(net_16794), .ZN(net_377), .A(net_376) );
NAND2_X2 inst_9617 ( .A1(net_14751), .ZN(net_10693), .A2(net_8474) );
INV_X4 inst_15977 ( .ZN(net_2039), .A(net_1684) );
INV_X2 inst_19212 ( .A(net_4859), .ZN(net_3503) );
NAND2_X2 inst_11392 ( .A1(net_20851), .ZN(net_6137), .A2(net_3516) );
OR2_X2 inst_1157 ( .A1(net_10672), .ZN(net_8289), .A2(net_8288) );
NAND2_X2 inst_11560 ( .A2(net_7397), .A1(net_2827), .ZN(net_2821) );
CLKBUF_X2 inst_21462 ( .A(net_21333), .Z(net_21334) );
NAND2_X2 inst_8065 ( .A2(net_18187), .ZN(net_18186), .A1(net_17679) );
NAND2_X2 inst_9993 ( .ZN(net_19587), .A1(net_10504), .A2(net_6496) );
NAND2_X2 inst_8408 ( .A1(net_20433), .ZN(net_18933), .A2(net_17236) );
INV_X4 inst_13395 ( .ZN(net_10670), .A(net_10669) );
CLKBUF_X2 inst_22195 ( .A(net_22066), .Z(net_22067) );
INV_X4 inst_16414 ( .ZN(net_4108), .A(net_3276) );
NOR2_X2 inst_3528 ( .ZN(net_13590), .A1(net_13589), .A2(net_13588) );
AOI211_X2 inst_21071 ( .A(net_20486), .B(net_10886), .ZN(net_7692), .C2(net_4634), .C1(net_3646) );
OAI21_X2 inst_2061 ( .ZN(net_10696), .B1(net_10695), .B2(net_6890), .A(net_652) );
AND2_X4 inst_21231 ( .ZN(net_19695), .A1(net_7917), .A2(net_4170) );
NOR2_X2 inst_4255 ( .ZN(net_6333), .A2(net_6332), .A1(net_3816) );
INV_X4 inst_13486 ( .ZN(net_9527), .A(net_7986) );
NAND3_X2 inst_6138 ( .ZN(net_13720), .A3(net_12705), .A2(net_10539), .A1(net_6830) );
INV_X4 inst_14981 ( .A(net_15889), .ZN(net_4466) );
NAND4_X2 inst_5272 ( .A2(net_19326), .A1(net_19325), .ZN(net_16117), .A4(net_15038), .A3(net_9621) );
INV_X4 inst_15242 ( .ZN(net_3498), .A(net_2817) );
INV_X4 inst_17980 ( .A(net_20852), .ZN(net_131) );
OAI21_X2 inst_2262 ( .A(net_7237), .ZN(net_7165), .B1(net_4157), .B2(net_3337) );
NOR2_X4 inst_3288 ( .ZN(net_2610), .A1(net_1139), .A2(net_225) );
AOI21_X4 inst_20200 ( .B1(net_19774), .ZN(net_14999), .B2(net_14605), .A(net_10400) );
INV_X2 inst_18898 ( .ZN(net_6096), .A(net_6095) );
OR2_X2 inst_1160 ( .ZN(net_7451), .A1(net_7450), .A2(net_7449) );
OAI21_X4 inst_1394 ( .ZN(net_19068), .A(net_16395), .B1(net_15990), .B2(net_15233) );
NAND2_X2 inst_9131 ( .ZN(net_13526), .A1(net_13525), .A2(net_10835) );
INV_X4 inst_13724 ( .ZN(net_12800), .A(net_7800) );
CLKBUF_X2 inst_21438 ( .A(net_21309), .Z(net_21310) );
INV_X4 inst_17951 ( .A(net_21095), .ZN(net_558) );
NAND2_X2 inst_10767 ( .A1(net_20528), .ZN(net_5634), .A2(net_4141) );
CLKBUF_X2 inst_21654 ( .A(net_21525), .Z(net_21526) );
OAI21_X2 inst_1876 ( .ZN(net_13692), .A(net_13691), .B2(net_12066), .B1(net_4350) );
DFF_X2 inst_19771 ( .QN(net_20876), .D(net_18580), .CK(net_21931) );
INV_X2 inst_18517 ( .A(net_14541), .ZN(net_12651) );
INV_X4 inst_12869 ( .ZN(net_17125), .A(net_16969) );
OAI22_X2 inst_1315 ( .B2(net_11861), .ZN(net_7076), .A1(net_7075), .A2(net_7074), .B1(net_60) );
INV_X4 inst_17179 ( .ZN(net_5658), .A(net_493) );
NOR2_X2 inst_5035 ( .A2(net_3402), .ZN(net_1126), .A1(net_146) );
NOR2_X2 inst_4759 ( .ZN(net_5494), .A2(net_2080), .A1(net_428) );
OAI211_X2 inst_2392 ( .ZN(net_16163), .C1(net_15971), .A(net_15908), .B(net_15820), .C2(net_15474) );
NOR2_X2 inst_4678 ( .A2(net_6524), .ZN(net_6379), .A1(net_1582) );
NAND2_X2 inst_9531 ( .ZN(net_12383), .A1(net_10445), .A2(net_9343) );
NOR2_X2 inst_3667 ( .ZN(net_12653), .A2(net_11547), .A1(net_7394) );
INV_X4 inst_13513 ( .ZN(net_13007), .A(net_9403) );
NAND2_X2 inst_7972 ( .A2(net_19864), .A1(net_19863), .ZN(net_18354) );
NOR2_X2 inst_4434 ( .ZN(net_6026), .A2(net_4870), .A1(net_154) );
INV_X4 inst_14775 ( .A(net_9525), .ZN(net_6799) );
INV_X2 inst_18841 ( .A(net_7192), .ZN(net_6718) );
NAND3_X2 inst_6380 ( .A2(net_12063), .ZN(net_12032), .A3(net_10565), .A1(net_9650) );
NOR2_X2 inst_4967 ( .ZN(net_1591), .A2(net_1276), .A1(net_168) );
NAND2_X4 inst_7217 ( .ZN(net_9351), .A2(net_7915), .A1(net_7837) );
INV_X4 inst_14953 ( .A(net_4855), .ZN(net_3504) );
INV_X2 inst_19331 ( .A(net_4289), .ZN(net_2534) );
CLKBUF_X2 inst_22903 ( .A(net_22693), .Z(net_22775) );
NAND3_X2 inst_6785 ( .ZN(net_4231), .A1(net_4230), .A2(net_3171), .A3(net_2562) );
NAND2_X2 inst_10792 ( .ZN(net_14402), .A1(net_8190), .A2(net_5543) );
XNOR2_X2 inst_656 ( .B(net_16833), .ZN(net_355), .A(net_354) );
NAND2_X2 inst_10866 ( .A2(net_20779), .ZN(net_20238), .A1(net_5432) );
INV_X4 inst_13993 ( .ZN(net_6448), .A(net_5281) );
NAND2_X4 inst_6900 ( .ZN(net_17993), .A1(net_17895), .A2(net_17846) );
NAND2_X2 inst_9690 ( .ZN(net_10241), .A1(net_10240), .A2(net_9721) );
XOR2_X2 inst_45 ( .A(net_21128), .Z(net_528), .B(net_527) );
INV_X4 inst_15351 ( .A(net_4230), .ZN(net_3686) );
NAND2_X2 inst_9551 ( .ZN(net_11024), .A2(net_7634), .A1(net_6889) );
INV_X4 inst_12500 ( .ZN(net_18645), .A(net_18617) );
INV_X4 inst_15125 ( .ZN(net_3948), .A(net_3149) );
XNOR2_X2 inst_458 ( .ZN(net_13295), .B(net_13294), .A(net_9237) );
NOR2_X4 inst_3093 ( .ZN(net_6980), .A2(net_4256), .A1(net_85) );
OAI21_X2 inst_1562 ( .B1(net_20708), .ZN(net_17208), .A(net_16910), .B2(net_16909) );
NAND2_X2 inst_9934 ( .ZN(net_9149), .A2(net_7105), .A1(net_117) );
NOR2_X2 inst_4148 ( .A2(net_12409), .A1(net_8739), .ZN(net_6907) );
NAND2_X2 inst_11814 ( .A1(net_3645), .ZN(net_2521), .A2(net_2497) );
INV_X4 inst_17407 ( .ZN(net_3060), .A(net_225) );
NAND3_X4 inst_5539 ( .ZN(net_20711), .A3(net_19804), .A1(net_19803), .A2(net_16156) );
NAND2_X2 inst_8644 ( .A2(net_16574), .ZN(net_16570), .A1(net_16569) );
SDFF_X2 inst_741 ( .Q(net_20898), .SE(net_18585), .SI(net_18537), .D(net_689), .CK(net_21441) );
INV_X2 inst_18440 ( .ZN(net_19606), .A(net_13258) );
INV_X4 inst_18063 ( .A(net_21083), .ZN(net_729) );
NAND2_X2 inst_9377 ( .ZN(net_11980), .A1(net_11018), .A2(net_8698) );
AOI21_X4 inst_20105 ( .B2(net_20896), .B1(net_19651), .ZN(net_16387), .A(net_13767) );
INV_X4 inst_16976 ( .ZN(net_1451), .A(net_886) );
NAND2_X4 inst_7195 ( .ZN(net_9817), .A1(net_8372), .A2(net_7976) );
NAND2_X2 inst_8700 ( .A2(net_20968), .A1(net_20611), .ZN(net_20273) );
NAND2_X2 inst_9338 ( .ZN(net_12276), .A1(net_12275), .A2(net_9281) );
CLKBUF_X2 inst_22935 ( .A(net_22806), .Z(net_22807) );
NAND2_X2 inst_10178 ( .A1(net_9349), .ZN(net_8196), .A2(net_8195) );
INV_X4 inst_12964 ( .ZN(net_16669), .A(net_16524) );
NAND2_X2 inst_8124 ( .A2(net_18070), .ZN(net_18054), .A1(net_15892) );
INV_X4 inst_17349 ( .ZN(net_9466), .A(net_6863) );
NOR2_X4 inst_2828 ( .A2(net_19783), .A1(net_19782), .ZN(net_15978) );
NAND2_X2 inst_7769 ( .A2(net_18745), .ZN(net_18744), .A1(net_17427) );
INV_X4 inst_13560 ( .ZN(net_10723), .A(net_9156) );
NOR2_X2 inst_4745 ( .A1(net_6112), .A2(net_3083), .ZN(net_3040) );
NOR2_X2 inst_3877 ( .ZN(net_9355), .A2(net_9354), .A1(net_8080) );
NAND2_X2 inst_9859 ( .ZN(net_9499), .A1(net_9498), .A2(net_6555) );
INV_X4 inst_16236 ( .A(net_13619), .ZN(net_11430) );
AND2_X4 inst_21236 ( .ZN(net_6730), .A2(net_3864), .A1(net_90) );
INV_X4 inst_17300 ( .ZN(net_988), .A(net_292) );
NAND2_X4 inst_7320 ( .A2(net_20851), .ZN(net_9900), .A1(net_4462) );
OR2_X4 inst_1131 ( .A2(net_20539), .ZN(net_3816), .A1(net_146) );
INV_X2 inst_19415 ( .ZN(net_1913), .A(net_1912) );
INV_X4 inst_14617 ( .ZN(net_6246), .A(net_4415) );
SDFF_X2 inst_691 ( .Q(net_20891), .SI(net_18868), .SE(net_18859), .D(net_627), .CK(net_22051) );
INV_X4 inst_14538 ( .ZN(net_4653), .A(net_4652) );
CLKBUF_X2 inst_21469 ( .A(net_21276), .Z(net_21341) );
INV_X2 inst_18523 ( .ZN(net_11140), .A(net_9839) );
NAND2_X2 inst_11769 ( .A1(net_2585), .A2(net_2445), .ZN(net_2065) );
NAND3_X2 inst_6402 ( .A3(net_20115), .ZN(net_20061), .A1(net_11979), .A2(net_7182) );
INV_X4 inst_12845 ( .A(net_17498), .ZN(net_17080) );
SDFF_X2 inst_770 ( .Q(net_20965), .SE(net_18862), .SI(net_18477), .D(net_800), .CK(net_21488) );
XNOR2_X2 inst_565 ( .B(net_17522), .ZN(net_666), .A(net_665) );
INV_X4 inst_15912 ( .ZN(net_1750), .A(net_1749) );
XNOR2_X2 inst_622 ( .B(net_9712), .A(net_557), .ZN(net_471) );
OAI21_X2 inst_1971 ( .ZN(net_12204), .A(net_12203), .B2(net_7824), .B1(net_5558) );
DFF_X1 inst_19909 ( .D(net_16776), .CK(net_21579), .Q(x585) );
NAND2_X4 inst_7418 ( .ZN(net_11041), .A2(net_4090), .A1(net_2540) );
INV_X8 inst_12342 ( .ZN(net_1803), .A(net_1730) );
INV_X4 inst_14345 ( .ZN(net_7837), .A(net_5339) );
INV_X4 inst_17772 ( .ZN(net_15362), .A(net_14714) );
INV_X4 inst_17206 ( .A(net_3542), .ZN(net_1357) );
INV_X4 inst_14531 ( .A(net_4724), .ZN(net_4723) );
XNOR2_X2 inst_409 ( .B(net_21147), .ZN(net_16624), .A(net_16378) );
NAND2_X2 inst_11679 ( .ZN(net_10837), .A1(net_4324), .A2(net_2345) );
INV_X8 inst_12323 ( .ZN(net_786), .A(net_106) );
INV_X4 inst_17181 ( .A(net_2431), .ZN(net_2361) );
NAND3_X2 inst_6672 ( .ZN(net_7761), .A2(net_7745), .A3(net_6893), .A1(net_4210) );
NAND3_X2 inst_5813 ( .ZN(net_15644), .A1(net_15032), .A3(net_14302), .A2(net_13231) );
CLKBUF_X2 inst_21904 ( .A(net_21739), .Z(net_21776) );
INV_X4 inst_15611 ( .ZN(net_4123), .A(net_1396) );
NAND2_X2 inst_8013 ( .ZN(net_18293), .A2(net_18242), .A1(net_17385) );
INV_X4 inst_12933 ( .ZN(net_17129), .A(net_16642) );
NOR2_X2 inst_3506 ( .ZN(net_13976), .A2(net_12202), .A1(net_10075) );
INV_X4 inst_17478 ( .ZN(net_439), .A(net_438) );
NAND2_X2 inst_9220 ( .ZN(net_19377), .A1(net_12976), .A2(net_10275) );
INV_X2 inst_18880 ( .ZN(net_6190), .A(net_6189) );
NAND2_X4 inst_7396 ( .A1(net_19491), .ZN(net_5357), .A2(net_4099) );
NAND2_X4 inst_7092 ( .ZN(net_14778), .A2(net_14130), .A1(net_13433) );
NAND2_X2 inst_11947 ( .ZN(net_7044), .A1(net_3929), .A2(net_1328) );
NAND2_X2 inst_11389 ( .ZN(net_6832), .A2(net_3525), .A1(net_2109) );
NAND2_X2 inst_7795 ( .ZN(net_18707), .A2(net_18692), .A1(net_17410) );
INV_X4 inst_15198 ( .ZN(net_3669), .A(net_2916) );
AOI21_X2 inst_20611 ( .ZN(net_13696), .A(net_13695), .B1(net_8981), .B2(net_6414) );
XNOR2_X2 inst_663 ( .A(net_21191), .B(net_21127), .ZN(net_283) );
NOR2_X4 inst_3227 ( .A1(net_20557), .ZN(net_3902), .A2(net_2561) );
NAND2_X2 inst_8949 ( .A1(net_15107), .ZN(net_14726), .A2(net_13233) );
INV_X4 inst_16493 ( .ZN(net_1670), .A(net_1187) );
NOR2_X2 inst_4224 ( .ZN(net_10646), .A2(net_7723), .A1(net_2969) );
AND3_X4 inst_21121 ( .ZN(net_12745), .A3(net_12744), .A2(net_10195), .A1(net_9499) );
CLKBUF_X2 inst_22624 ( .A(net_21876), .Z(net_22496) );
INV_X2 inst_19247 ( .A(net_4236), .ZN(net_3265) );
CLKBUF_X2 inst_22163 ( .A(net_22034), .Z(net_22035) );
NAND2_X4 inst_7279 ( .ZN(net_7565), .A2(net_4591), .A1(net_3134) );
OAI21_X2 inst_2290 ( .ZN(net_6519), .A(net_6518), .B2(net_1980), .B1(net_1016) );
INV_X4 inst_17463 ( .ZN(net_945), .A(net_253) );
INV_X2 inst_19675 ( .A(net_20500), .ZN(net_20499) );
NAND2_X2 inst_11913 ( .A1(net_20493), .ZN(net_2562), .A2(net_1640) );
INV_X2 inst_19476 ( .A(net_15692), .ZN(net_1411) );
NOR2_X2 inst_5070 ( .ZN(net_10381), .A1(net_761), .A2(net_44) );
NAND3_X2 inst_5797 ( .ZN(net_15719), .A1(net_15062), .A3(net_14995), .A2(net_13520) );
CLKBUF_X2 inst_21922 ( .A(net_21793), .Z(net_21794) );
INV_X4 inst_14640 ( .ZN(net_4630), .A(net_4380) );
NOR3_X4 inst_2621 ( .A3(net_19204), .A1(net_19203), .ZN(net_15475), .A2(net_11565) );
INV_X4 inst_15743 ( .ZN(net_2763), .A(net_1944) );
NAND2_X2 inst_9159 ( .ZN(net_13382), .A1(net_12366), .A2(net_10434) );
CLKBUF_X2 inst_22881 ( .A(net_22752), .Z(net_22753) );
NAND2_X2 inst_10815 ( .ZN(net_7275), .A1(net_5516), .A2(net_5515) );
INV_X4 inst_14454 ( .ZN(net_9885), .A(net_4954) );
INV_X2 inst_18559 ( .ZN(net_10863), .A(net_10862) );
INV_X4 inst_16598 ( .ZN(net_1795), .A(net_1008) );
NAND2_X2 inst_11928 ( .ZN(net_2423), .A2(net_1477), .A1(net_238) );
NAND2_X2 inst_9358 ( .A1(net_13544), .ZN(net_12152), .A2(net_12151) );
NAND2_X4 inst_7699 ( .ZN(net_419), .A2(net_325), .A1(net_248) );
OAI21_X2 inst_1647 ( .A(net_16242), .ZN(net_15907), .B2(net_15181), .B1(net_15079) );
NOR2_X4 inst_3263 ( .ZN(net_4321), .A1(net_2909), .A2(net_2328) );
NAND2_X2 inst_12114 ( .ZN(net_231), .A1(net_230), .A2(net_229) );
OAI21_X4 inst_1376 ( .ZN(net_20791), .B1(net_16395), .A(net_16293), .B2(net_16199) );
NOR2_X4 inst_2882 ( .ZN(net_18895), .A1(net_9854), .A2(net_7048) );
NAND2_X2 inst_10507 ( .ZN(net_11799), .A2(net_6922), .A1(net_81) );
INV_X4 inst_12605 ( .A(net_18099), .ZN(net_18094) );
INV_X4 inst_18325 ( .A(net_20923), .ZN(net_20540) );
NAND2_X2 inst_8182 ( .ZN(net_17930), .A2(net_17912), .A1(net_17904) );
NAND2_X2 inst_11483 ( .ZN(net_8507), .A2(net_3120), .A1(net_2127) );
CLKBUF_X2 inst_22450 ( .A(net_22321), .Z(net_22322) );
NAND2_X2 inst_10654 ( .ZN(net_11908), .A2(net_6315), .A1(net_1916) );
DFF_X1 inst_19900 ( .D(net_16852), .CK(net_22351), .Q(x675) );
NAND3_X2 inst_6188 ( .ZN(net_13465), .A3(net_9132), .A2(net_7938), .A1(net_4346) );
NAND2_X2 inst_10742 ( .ZN(net_9151), .A2(net_5539), .A1(net_4754) );
OAI21_X2 inst_1659 ( .A(net_15840), .ZN(net_15786), .B2(net_14780), .B1(net_5151) );
CLKBUF_X2 inst_21775 ( .A(net_21646), .Z(net_21647) );
INV_X4 inst_17331 ( .ZN(net_5506), .A(net_655) );
AOI21_X2 inst_20872 ( .ZN(net_8557), .A(net_8556), .B2(net_8501), .B1(net_1386) );
NAND2_X2 inst_8184 ( .ZN(net_17928), .A1(net_17864), .A2(net_17801) );
NAND3_X2 inst_5702 ( .ZN(net_19834), .A3(net_15907), .A2(net_14285), .A1(net_13831) );
XNOR2_X2 inst_398 ( .A(net_16764), .ZN(net_16754), .B(net_481) );
AOI21_X4 inst_20233 ( .B2(net_20679), .B1(net_20678), .ZN(net_12728), .A(net_308) );
XNOR2_X2 inst_436 ( .ZN(net_16098), .A(net_16097), .B(net_15589) );
NAND2_X2 inst_11766 ( .ZN(net_9959), .A1(net_6092), .A2(net_2075) );
INV_X4 inst_13265 ( .ZN(net_12654), .A(net_12653) );
NAND3_X2 inst_6529 ( .ZN(net_10605), .A3(net_10604), .A2(net_10454), .A1(net_9634) );
NAND2_X2 inst_9852 ( .ZN(net_9519), .A1(net_9518), .A2(net_6979) );
INV_X2 inst_19280 ( .ZN(net_5193), .A(net_2938) );
NOR2_X2 inst_3705 ( .ZN(net_11089), .A1(net_11088), .A2(net_7379) );
INV_X2 inst_19077 ( .ZN(net_4599), .A(net_4598) );
INV_X4 inst_17990 ( .A(net_21179), .ZN(net_488) );
NAND3_X2 inst_6746 ( .A2(net_8334), .ZN(net_5819), .A1(net_5818), .A3(net_5165) );
OAI21_X2 inst_2231 ( .ZN(net_8185), .A(net_8184), .B1(net_7124), .B2(net_3604) );
XNOR2_X2 inst_144 ( .B(net_21199), .A(net_20218), .ZN(net_18179) );
INV_X2 inst_18891 ( .ZN(net_6116), .A(net_6115) );
NAND2_X2 inst_9750 ( .ZN(net_10058), .A1(net_8851), .A2(net_6975) );
NAND2_X2 inst_10565 ( .ZN(net_13883), .A1(net_6712), .A2(net_6597) );
INV_X4 inst_13660 ( .ZN(net_9615), .A(net_8113) );
INV_X4 inst_18230 ( .A(net_20925), .ZN(net_108) );
NAND2_X4 inst_6912 ( .A2(net_19920), .A1(net_19919), .ZN(net_17800) );
INV_X4 inst_17524 ( .A(net_731), .ZN(net_398) );
NOR2_X2 inst_4857 ( .ZN(net_2613), .A1(net_2280), .A2(net_2279) );
CLKBUF_X2 inst_22182 ( .A(net_22053), .Z(net_22054) );
NAND2_X2 inst_9763 ( .A1(net_20511), .ZN(net_19360), .A2(net_4725) );
INV_X4 inst_16892 ( .ZN(net_2996), .A(net_951) );
NAND3_X4 inst_5555 ( .ZN(net_19658), .A3(net_15919), .A2(net_15260), .A1(net_13832) );
NAND2_X2 inst_10026 ( .A2(net_8780), .ZN(net_8755), .A1(net_5831) );
NOR2_X2 inst_4447 ( .A1(net_4783), .ZN(net_4782), .A2(net_2722) );
NAND3_X2 inst_6194 ( .ZN(net_19554), .A3(net_9860), .A1(net_8403), .A2(net_5659) );
NAND2_X2 inst_8493 ( .ZN(net_20157), .A1(net_19444), .A2(net_16564) );
INV_X4 inst_15694 ( .A(net_2674), .ZN(net_2021) );
INV_X4 inst_17818 ( .ZN(net_242), .A(net_152) );
AOI21_X2 inst_20833 ( .ZN(net_9687), .A(net_7357), .B2(net_4483), .B1(net_2893) );
NAND3_X2 inst_6329 ( .ZN(net_12481), .A3(net_12480), .A1(net_9674), .A2(net_6225) );
INV_X4 inst_12470 ( .ZN(net_20296), .A(net_18769) );
INV_X2 inst_19575 ( .ZN(net_796), .A(net_139) );
INV_X4 inst_16065 ( .ZN(net_2510), .A(net_2296) );
INV_X4 inst_15878 ( .ZN(net_1838), .A(net_1788) );
INV_X4 inst_14937 ( .ZN(net_4553), .A(net_3537) );
CLKBUF_X2 inst_21522 ( .A(net_21393), .Z(net_21394) );
AOI21_X2 inst_20803 ( .B2(net_19676), .ZN(net_10347), .A(net_9754), .B1(net_7633) );
OAI21_X4 inst_1360 ( .B2(net_20639), .B1(net_20638), .A(net_18067), .ZN(net_18055) );
INV_X4 inst_15871 ( .ZN(net_2887), .A(net_1027) );
INV_X4 inst_16578 ( .ZN(net_1522), .A(net_1156) );
XNOR2_X2 inst_466 ( .B(net_21191), .ZN(net_12874), .A(net_11178) );
NOR2_X2 inst_3981 ( .ZN(net_8386), .A1(net_7769), .A2(net_4796) );
INV_X4 inst_18237 ( .A(net_20999), .ZN(net_2132) );
NAND4_X4 inst_5205 ( .A3(net_18926), .A1(net_18925), .ZN(net_16762), .A4(net_16248), .A2(net_15830) );
INV_X4 inst_14742 ( .ZN(net_6810), .A(net_5752) );
NAND2_X2 inst_10073 ( .A1(net_14962), .ZN(net_8653), .A2(net_8242) );
NOR2_X4 inst_3038 ( .ZN(net_8066), .A1(net_3643), .A2(net_1076) );
NAND2_X4 inst_7605 ( .ZN(net_4216), .A2(net_1404), .A1(net_1403) );
INV_X4 inst_14154 ( .A(net_7248), .ZN(net_6025) );
INV_X2 inst_19282 ( .ZN(net_2933), .A(net_2932) );
NAND2_X4 inst_7542 ( .A1(net_20181), .ZN(net_4026), .A2(net_1861) );
INV_X4 inst_16863 ( .ZN(net_9360), .A(net_961) );
NOR2_X2 inst_3864 ( .ZN(net_12804), .A1(net_9387), .A2(net_9386) );
CLKBUF_X2 inst_22552 ( .A(net_22423), .Z(net_22424) );
INV_X4 inst_15482 ( .ZN(net_9843), .A(net_9541) );
INV_X4 inst_12735 ( .A(net_17586), .ZN(net_17455) );
INV_X4 inst_15596 ( .A(net_3171), .ZN(net_2228) );
NAND2_X4 inst_7406 ( .ZN(net_6705), .A2(net_2869), .A1(net_222) );
NAND2_X2 inst_9757 ( .ZN(net_19742), .A2(net_10004), .A1(net_1915) );
INV_X2 inst_19606 ( .A(net_21213), .ZN(net_104) );
INV_X2 inst_18566 ( .ZN(net_13713), .A(net_7573) );
CLKBUF_X2 inst_22017 ( .A(net_21888), .Z(net_21889) );
AOI21_X2 inst_20760 ( .ZN(net_11153), .B1(net_10231), .B2(net_7469), .A(net_3166) );
NAND2_X4 inst_7283 ( .A1(net_20671), .ZN(net_5729), .A2(net_1961) );
NAND4_X4 inst_5214 ( .A3(net_20141), .A1(net_20140), .ZN(net_16619), .A4(net_16261), .A2(net_14495) );
CLKBUF_X2 inst_22958 ( .A(net_22154), .Z(net_22830) );
INV_X4 inst_15170 ( .ZN(net_14669), .A(net_3015) );
INV_X4 inst_13331 ( .ZN(net_13014), .A(net_11136) );
NOR2_X2 inst_4794 ( .ZN(net_4717), .A1(net_2964), .A2(net_2674) );
INV_X4 inst_13838 ( .ZN(net_10919), .A(net_7485) );
NAND2_X2 inst_10804 ( .ZN(net_14384), .A1(net_6924), .A2(net_5467) );
INV_X4 inst_13688 ( .A(net_7965), .ZN(net_7964) );
NOR2_X2 inst_3829 ( .A1(net_12179), .ZN(net_11096), .A2(net_6149) );
NAND2_X2 inst_7883 ( .ZN(net_18517), .A1(net_18473), .A2(net_17741) );
INV_X4 inst_14465 ( .ZN(net_7866), .A(net_4923) );
INV_X4 inst_17755 ( .ZN(net_661), .A(net_304) );
NAND2_X2 inst_9012 ( .ZN(net_19691), .A1(net_14303), .A2(net_12650) );
INV_X4 inst_13414 ( .ZN(net_10294), .A(net_10293) );
INV_X4 inst_14621 ( .ZN(net_5840), .A(net_2537) );
CLKBUF_X2 inst_22756 ( .A(net_22627), .Z(net_22628) );
NAND2_X2 inst_10325 ( .ZN(net_9315), .A2(net_6028), .A1(net_6007) );
NAND2_X2 inst_10971 ( .A1(net_9098), .ZN(net_4977), .A2(net_4877) );
INV_X4 inst_13918 ( .A(net_10523), .ZN(net_8242) );
INV_X4 inst_15791 ( .ZN(net_5664), .A(net_1901) );
CLKBUF_X2 inst_22206 ( .A(net_21327), .Z(net_22078) );
INV_X4 inst_17811 ( .ZN(net_263), .A(net_125) );
NAND2_X2 inst_8161 ( .ZN(net_17975), .A2(net_17893), .A1(net_17844) );
OAI21_X2 inst_2168 ( .ZN(net_8930), .B2(net_6148), .B1(net_1305), .A(net_70) );
NAND2_X4 inst_7241 ( .ZN(net_10437), .A2(net_7941), .A1(net_6998) );
INV_X4 inst_15060 ( .ZN(net_3305), .A(net_3304) );
INV_X2 inst_18889 ( .ZN(net_9716), .A(net_6129) );
NOR2_X2 inst_4322 ( .ZN(net_5864), .A1(net_3637), .A2(net_2173) );
OR2_X4 inst_1078 ( .ZN(net_10462), .A1(net_9131), .A2(net_6632) );
NAND3_X2 inst_6497 ( .ZN(net_20654), .A2(net_7367), .A3(net_6432), .A1(net_3957) );
AND2_X4 inst_21162 ( .A1(net_20763), .ZN(net_13773), .A2(net_13772) );
AOI21_X2 inst_20960 ( .ZN(net_5331), .B1(net_5330), .B2(net_4188), .A(net_4164) );
NOR2_X2 inst_3557 ( .ZN(net_13017), .A2(net_10344), .A1(net_8896) );
SDFF_X2 inst_1039 ( .QN(net_20995), .D(net_1866), .SE(net_263), .CK(net_21825), .SI(x3106) );
OAI21_X2 inst_1992 ( .ZN(net_20614), .B2(net_11733), .A(net_11443), .B1(net_10493) );
INV_X4 inst_16679 ( .ZN(net_20181), .A(net_1075) );
NAND4_X2 inst_5449 ( .ZN(net_13527), .A1(net_7553), .A3(net_7520), .A4(net_7460), .A2(net_5680) );
NOR2_X2 inst_4048 ( .ZN(net_9394), .A1(net_6009), .A2(net_4286) );
NAND2_X4 inst_7549 ( .ZN(net_3109), .A2(net_276), .A1(net_123) );
NOR2_X2 inst_4003 ( .ZN(net_8142), .A2(net_8141), .A1(net_2302) );
NAND2_X4 inst_6868 ( .ZN(net_18269), .A2(net_18263), .A1(net_17739) );
AOI21_X2 inst_20546 ( .ZN(net_14396), .B1(net_14395), .B2(net_12468), .A(net_4781) );
NOR2_X2 inst_5033 ( .ZN(net_1804), .A2(net_1138), .A1(net_761) );
NAND2_X2 inst_8306 ( .A2(net_21209), .A1(net_20230), .ZN(net_19188) );
INV_X4 inst_15512 ( .ZN(net_14612), .A(net_2408) );
CLKBUF_X2 inst_21996 ( .A(net_21867), .Z(net_21868) );
INV_X4 inst_13966 ( .ZN(net_8731), .A(net_6709) );
NAND2_X2 inst_8846 ( .ZN(net_19311), .A2(net_15091), .A1(net_14927) );
NAND4_X2 inst_5363 ( .A4(net_19224), .A1(net_19223), .ZN(net_15286), .A3(net_11231), .A2(net_10703) );
INV_X4 inst_17128 ( .ZN(net_8924), .A(net_4890) );
NOR2_X2 inst_3542 ( .ZN(net_14200), .A2(net_13367), .A1(net_10405) );
INV_X4 inst_15529 ( .A(net_3118), .ZN(net_2385) );
INV_X4 inst_16547 ( .ZN(net_15880), .A(net_14046) );
NAND3_X2 inst_6300 ( .ZN(net_12810), .A2(net_12809), .A1(net_10916), .A3(net_7279) );
XNOR2_X2 inst_115 ( .ZN(net_18498), .A(net_18413), .B(net_17116) );
CLKBUF_X2 inst_21991 ( .A(net_21862), .Z(net_21863) );
NOR2_X2 inst_4691 ( .ZN(net_3909), .A2(net_3696), .A1(net_3182) );
NOR2_X2 inst_3726 ( .ZN(net_10895), .A2(net_10894), .A1(net_8025) );
NOR2_X4 inst_3045 ( .ZN(net_8295), .A1(net_5055), .A2(net_955) );
NAND2_X2 inst_9801 ( .ZN(net_11693), .A2(net_9699), .A1(net_8785) );
INV_X4 inst_12741 ( .ZN(net_17438), .A(net_17437) );
CLKBUF_X2 inst_22640 ( .A(net_22157), .Z(net_22512) );
AOI21_X2 inst_20319 ( .ZN(net_15925), .B1(net_15924), .B2(net_15229), .A(net_14951) );
INV_X2 inst_18877 ( .ZN(net_6203), .A(net_6202) );
NAND3_X2 inst_6113 ( .ZN(net_19713), .A3(net_11303), .A1(net_8290), .A2(net_6914) );
OAI22_X2 inst_1263 ( .B1(net_21140), .ZN(net_17391), .A1(net_17113), .B2(net_16954), .A2(net_16946) );
INV_X2 inst_19299 ( .ZN(net_2784), .A(net_2783) );
INV_X2 inst_19657 ( .A(net_20434), .ZN(net_20433) );
CLKBUF_X2 inst_21374 ( .A(net_21245), .Z(net_21246) );
INV_X4 inst_16699 ( .ZN(net_7244), .A(net_1147) );
NAND2_X2 inst_8047 ( .ZN(net_18229), .A2(net_18179), .A1(net_17607) );
NOR2_X4 inst_3330 ( .A2(net_386), .ZN(net_247), .A1(net_246) );
NAND2_X2 inst_10225 ( .ZN(net_10365), .A1(net_8067), .A2(net_8066) );
NAND2_X4 inst_7374 ( .ZN(net_5770), .A1(net_4301), .A2(net_3076) );
OAI21_X4 inst_1445 ( .B2(net_19697), .B1(net_19696), .ZN(net_15746), .A(net_15699) );
NAND2_X2 inst_11907 ( .ZN(net_1558), .A2(net_1418), .A1(net_222) );
INV_X4 inst_16728 ( .ZN(net_6301), .A(net_1053) );
NOR2_X2 inst_3990 ( .A2(net_20779), .ZN(net_19860), .A1(net_8287) );
INV_X4 inst_17500 ( .A(net_10683), .ZN(net_421) );
NAND2_X2 inst_8976 ( .ZN(net_14513), .A1(net_14367), .A2(net_12846) );
INV_X4 inst_18318 ( .ZN(net_20527), .A(net_16469) );
INV_X4 inst_13156 ( .ZN(net_14871), .A(net_14328) );
NAND3_X2 inst_5982 ( .ZN(net_19872), .A2(net_14547), .A3(net_13980), .A1(net_13380) );
NAND2_X2 inst_12115 ( .ZN(net_1043), .A2(net_856), .A1(net_225) );
NAND2_X2 inst_7931 ( .ZN(net_18440), .A1(net_18439), .A2(net_18438) );
INV_X4 inst_15945 ( .ZN(net_1714), .A(net_1233) );
INV_X4 inst_16744 ( .ZN(net_3314), .A(net_1349) );
NAND2_X2 inst_7932 ( .ZN(net_18437), .A1(net_18411), .A2(net_17568) );
OAI21_X2 inst_1512 ( .B2(net_19626), .B1(net_19625), .ZN(net_18583), .A(net_18582) );
NAND2_X2 inst_10366 ( .ZN(net_10865), .A1(net_6636), .A2(net_5829) );
NAND4_X4 inst_5160 ( .ZN(net_18604), .A2(net_18596), .A1(net_18591), .A4(net_16064), .A3(net_16032) );
NAND2_X2 inst_8733 ( .ZN(net_16056), .A2(net_15782), .A1(net_15486) );
INV_X4 inst_13209 ( .ZN(net_13725), .A(net_12983) );
INV_X4 inst_14395 ( .ZN(net_10174), .A(net_6781) );
INV_X2 inst_19523 ( .A(net_5256), .ZN(net_2008) );
INV_X2 inst_19260 ( .ZN(net_20656), .A(net_15976) );
INV_X2 inst_18791 ( .A(net_9573), .ZN(net_7480) );
NAND2_X2 inst_10727 ( .A2(net_20575), .ZN(net_7368), .A1(net_3436) );
AOI21_X2 inst_20510 ( .ZN(net_14629), .B1(net_14628), .A(net_12073), .B2(net_11953) );
NAND2_X4 inst_7692 ( .ZN(net_20582), .A2(net_646), .A1(net_105) );
INV_X4 inst_16017 ( .ZN(net_9510), .A(net_1650) );
INV_X4 inst_14822 ( .ZN(net_4921), .A(net_3912) );
OAI21_X2 inst_2299 ( .ZN(net_6417), .B2(net_5859), .A(net_5118), .B1(net_2016) );
NAND2_X2 inst_11691 ( .ZN(net_4854), .A1(net_2585), .A2(net_2326) );
INV_X8 inst_12441 ( .ZN(net_20494), .A(net_20493) );
INV_X2 inst_19184 ( .ZN(net_3741), .A(net_3740) );
NAND2_X4 inst_7504 ( .ZN(net_2268), .A1(net_2139), .A2(net_1022) );
NAND4_X2 inst_5292 ( .ZN(net_15931), .A4(net_15188), .A1(net_14018), .A3(net_13044), .A2(net_11601) );
CLKBUF_X2 inst_22055 ( .A(net_21489), .Z(net_21927) );
INV_X4 inst_16829 ( .ZN(net_1124), .A(net_112) );
NAND2_X4 inst_7578 ( .ZN(net_3110), .A2(net_834), .A1(net_216) );
NAND2_X2 inst_8166 ( .ZN(net_17965), .A1(net_17886), .A2(net_17840) );
INV_X8 inst_12366 ( .A(net_20868), .ZN(net_3026) );
INV_X4 inst_14963 ( .A(net_5035), .ZN(net_3442) );
CLKBUF_X2 inst_22126 ( .A(net_21997), .Z(net_21998) );
OAI21_X2 inst_1642 ( .ZN(net_20096), .A(net_16187), .B2(net_15238), .B1(net_14252) );
CLKBUF_X2 inst_22189 ( .A(net_22053), .Z(net_22061) );
INV_X4 inst_12703 ( .ZN(net_17797), .A(net_17708) );
CLKBUF_X2 inst_22138 ( .A(net_22009), .Z(net_22010) );
INV_X4 inst_13434 ( .ZN(net_19831), .A(net_8427) );
XNOR2_X2 inst_199 ( .A(net_17673), .ZN(net_17670), .B(net_7651) );
INV_X4 inst_12540 ( .ZN(net_20018), .A(net_18353) );
INV_X4 inst_13259 ( .ZN(net_12702), .A(net_12701) );
NAND3_X2 inst_6764 ( .ZN(net_5359), .A3(net_5358), .A2(net_1916), .A1(net_804) );
NAND2_X4 inst_6976 ( .A2(net_20405), .A1(net_20404), .ZN(net_17328) );
INV_X4 inst_13313 ( .ZN(net_14449), .A(net_10324) );
NOR2_X2 inst_4875 ( .ZN(net_2205), .A2(net_2204), .A1(net_1643) );
INV_X4 inst_14274 ( .ZN(net_5661), .A(net_5660) );
INV_X2 inst_19341 ( .A(net_8559), .ZN(net_2451) );
INV_X4 inst_16956 ( .ZN(net_9966), .A(net_5308) );
INV_X4 inst_18163 ( .A(net_21069), .ZN(net_793) );
INV_X4 inst_14252 ( .ZN(net_5759), .A(net_5758) );
INV_X4 inst_15412 ( .A(net_14038), .ZN(net_10279) );
CLKBUF_X2 inst_22688 ( .A(net_21824), .Z(net_22560) );
CLKBUF_X2 inst_22533 ( .A(net_21289), .Z(net_22405) );
NOR2_X2 inst_4114 ( .A2(net_12935), .ZN(net_7060), .A1(net_7059) );
XNOR2_X2 inst_540 ( .B(net_942), .ZN(net_854), .A(net_853) );
OAI21_X2 inst_2356 ( .A(net_9031), .ZN(net_2959), .B1(net_2523), .B2(net_1837) );
SDFF_X2 inst_998 ( .QN(net_21085), .D(net_591), .SE(net_263), .CK(net_22584), .SI(x1651) );
NAND2_X2 inst_7989 ( .ZN(net_19948), .A1(net_18326), .A2(net_18325) );
NAND3_X2 inst_6044 ( .ZN(net_14261), .A3(net_12278), .A2(net_11115), .A1(net_3770) );
NAND3_X2 inst_5952 ( .ZN(net_14879), .A3(net_14878), .A1(net_8691), .A2(net_5998) );
NOR2_X4 inst_3209 ( .A2(net_20494), .ZN(net_5443), .A1(net_3023) );
INV_X4 inst_13989 ( .A(net_13655), .ZN(net_6544) );
AOI21_X2 inst_20943 ( .ZN(net_6398), .B1(net_2644), .B2(net_2328), .A(net_2322) );
NAND2_X2 inst_9730 ( .ZN(net_13049), .A1(net_10114), .A2(net_9332) );
INV_X8 inst_12298 ( .ZN(net_1456), .A(net_705) );
INV_X4 inst_14042 ( .ZN(net_7619), .A(net_6261) );
DFF_X1 inst_19795 ( .D(net_18249), .CK(net_22405), .Q(x771) );
CLKBUF_X2 inst_21553 ( .A(net_21285), .Z(net_21425) );
NAND2_X2 inst_9792 ( .ZN(net_9718), .A1(net_9717), .A2(net_9716) );
CLKBUF_X2 inst_21558 ( .A(net_21429), .Z(net_21430) );
NAND2_X2 inst_9242 ( .ZN(net_12690), .A2(net_12689), .A1(net_12373) );
NAND2_X2 inst_10205 ( .ZN(net_8118), .A1(net_8117), .A2(net_4665) );
NAND2_X2 inst_11442 ( .ZN(net_12830), .A1(net_3293), .A2(net_3292) );
NOR2_X2 inst_5090 ( .A2(net_897), .ZN(net_835), .A1(net_834) );
NAND3_X2 inst_6720 ( .A2(net_14572), .A3(net_10690), .ZN(net_6531), .A1(net_6530) );
XNOR2_X2 inst_192 ( .ZN(net_17680), .A(net_17679), .B(net_942) );
INV_X4 inst_14400 ( .A(net_6732), .ZN(net_5115) );
NOR3_X2 inst_2715 ( .ZN(net_13507), .A3(net_9971), .A2(net_9175), .A1(net_2793) );
NOR2_X2 inst_4242 ( .ZN(net_7793), .A2(net_6646), .A1(net_60) );
INV_X4 inst_13059 ( .ZN(net_16364), .A(net_16321) );
NOR2_X2 inst_4126 ( .ZN(net_6994), .A1(net_6993), .A2(net_6992) );
NAND2_X4 inst_7434 ( .ZN(net_6725), .A2(net_3384), .A1(net_3108) );
AND2_X2 inst_21269 ( .ZN(net_18149), .A2(net_18147), .A1(net_18086) );
NOR2_X2 inst_4178 ( .A2(net_10937), .ZN(net_8126), .A1(net_6720) );
NOR2_X2 inst_3547 ( .ZN(net_13106), .A1(net_13105), .A2(net_10885) );
NAND2_X2 inst_8741 ( .A1(net_16259), .ZN(net_15993), .A2(net_15823) );
INV_X4 inst_12720 ( .ZN(net_17711), .A(net_17618) );
NAND3_X2 inst_6558 ( .A2(net_11598), .A3(net_10553), .ZN(net_10508), .A1(net_3689) );
INV_X2 inst_18901 ( .ZN(net_9601), .A(net_8087) );
NAND2_X2 inst_9739 ( .ZN(net_10103), .A2(net_9383), .A1(net_9037) );
NAND2_X4 inst_7234 ( .A1(net_20440), .ZN(net_8697), .A2(net_4945) );
XNOR2_X2 inst_486 ( .B(net_21200), .ZN(net_10495), .A(net_7323) );
INV_X4 inst_12977 ( .A(net_16701), .ZN(net_16694) );
INV_X4 inst_15117 ( .ZN(net_5989), .A(net_2105) );
INV_X4 inst_13365 ( .ZN(net_12328), .A(net_10911) );
OR2_X2 inst_1240 ( .A2(net_20875), .ZN(net_961), .A1(net_34) );
NAND4_X2 inst_5445 ( .ZN(net_13877), .A1(net_13876), .A3(net_13479), .A2(net_12383), .A4(net_6452) );
CLKBUF_X2 inst_22608 ( .A(net_22479), .Z(net_22480) );
NAND3_X2 inst_6597 ( .ZN(net_9902), .A2(net_7488), .A3(net_5140), .A1(net_3927) );
AOI22_X2 inst_19971 ( .ZN(net_15691), .A2(net_15051), .B1(net_14554), .B2(net_11394), .A1(net_1850) );
INV_X2 inst_18740 ( .ZN(net_10385), .A(net_7909) );
INV_X4 inst_15941 ( .ZN(net_2052), .A(net_1716) );
CLKBUF_X2 inst_21418 ( .A(net_21249), .Z(net_21290) );
CLKBUF_X2 inst_22746 ( .A(net_22617), .Z(net_22618) );
NAND2_X2 inst_9186 ( .A1(net_14303), .ZN(net_13131), .A2(net_10332) );
OAI21_X2 inst_1521 ( .B2(net_20220), .ZN(net_18198), .A(net_18111), .B1(net_18085) );
INV_X2 inst_19472 ( .A(net_2606), .ZN(net_1437) );
NAND3_X2 inst_6620 ( .A3(net_10306), .ZN(net_9058), .A2(net_9033), .A1(net_6784) );
INV_X4 inst_13692 ( .ZN(net_10140), .A(net_7932) );
NAND2_X2 inst_9679 ( .A1(net_14361), .ZN(net_10268), .A2(net_10267) );
INV_X4 inst_12976 ( .A(net_16510), .ZN(net_16509) );
NOR2_X2 inst_4845 ( .A1(net_2636), .A2(net_2485), .ZN(net_2352) );
OAI22_X2 inst_1306 ( .ZN(net_9920), .B1(net_8190), .A1(net_7156), .B2(net_5133), .A2(net_4662) );
OAI211_X2 inst_2563 ( .ZN(net_9879), .A(net_9878), .C1(net_7844), .C2(net_7755), .B(net_6111) );
NAND2_X2 inst_10766 ( .ZN(net_5636), .A1(net_5635), .A2(net_4143) );
NAND2_X2 inst_11208 ( .ZN(net_4031), .A1(net_4030), .A2(net_4029) );
INV_X4 inst_18007 ( .A(net_21238), .ZN(net_81) );
NAND2_X2 inst_9931 ( .ZN(net_20624), .A2(net_7112), .A1(net_1959) );
INV_X4 inst_15640 ( .ZN(net_4315), .A(net_3162) );
OAI21_X4 inst_1407 ( .A(net_20872), .B2(net_19707), .B1(net_19706), .ZN(net_16182) );
INV_X4 inst_12916 ( .A(net_16669), .ZN(net_16668) );
NAND2_X2 inst_8096 ( .A1(net_20506), .ZN(net_18125), .A2(net_18124) );
INV_X4 inst_13128 ( .ZN(net_15275), .A(net_14905) );
INV_X4 inst_13803 ( .A(net_9709), .ZN(net_7550) );
NAND2_X4 inst_7018 ( .ZN(net_17633), .A1(net_16583), .A2(net_16456) );
CLKBUF_X2 inst_22650 ( .A(net_22521), .Z(net_22522) );
INV_X4 inst_16176 ( .ZN(net_10898), .A(net_4056) );
NAND2_X2 inst_9132 ( .ZN(net_13523), .A1(net_12133), .A2(net_10806) );
NAND3_X2 inst_6052 ( .ZN(net_14236), .A2(net_14235), .A1(net_12600), .A3(net_11459) );
NAND2_X2 inst_11526 ( .ZN(net_2972), .A2(net_2971), .A1(net_1019) );
INV_X4 inst_17862 ( .ZN(net_315), .A(net_131) );
NAND2_X4 inst_6965 ( .ZN(net_17419), .A1(net_17013), .A2(net_16869) );
NAND2_X2 inst_11051 ( .A2(net_20466), .ZN(net_8665), .A1(net_4707) );
NAND2_X2 inst_9687 ( .ZN(net_19754), .A2(net_10246), .A1(net_9395) );
NAND2_X2 inst_10217 ( .ZN(net_12093), .A2(net_9485), .A1(net_573) );
NOR2_X2 inst_5099 ( .ZN(net_10063), .A2(net_788), .A1(net_70) );
CLKBUF_X2 inst_21662 ( .A(net_21316), .Z(net_21534) );
NAND2_X2 inst_11116 ( .ZN(net_6829), .A1(net_2996), .A2(net_1966) );
NAND3_X2 inst_6134 ( .ZN(net_13737), .A3(net_12603), .A2(net_11085), .A1(net_8413) );
XNOR2_X2 inst_584 ( .B(net_1896), .ZN(net_587), .A(net_586) );
NAND2_X2 inst_9561 ( .A2(net_19644), .ZN(net_12646), .A1(net_10974) );
CLKBUF_X2 inst_21856 ( .A(net_21495), .Z(net_21728) );
XNOR2_X2 inst_470 ( .ZN(net_12265), .B(net_12264), .A(net_7741) );
NAND2_X2 inst_8668 ( .A2(net_16619), .ZN(net_16472), .A1(net_618) );
INV_X4 inst_15566 ( .A(net_3007), .ZN(net_2290) );
INV_X4 inst_12917 ( .ZN(net_16667), .A(net_16666) );
CLKBUF_X2 inst_21515 ( .A(net_21376), .Z(net_21387) );
NAND2_X2 inst_8138 ( .A1(net_20166), .ZN(net_18030), .A2(net_17879) );
NOR2_X2 inst_4490 ( .ZN(net_8075), .A2(net_4306), .A1(net_3275) );
OAI21_X2 inst_1752 ( .A(net_15087), .ZN(net_14796), .B1(net_13441), .B2(net_13257) );
INV_X4 inst_18221 ( .A(net_20902), .ZN(net_164) );
INV_X4 inst_16394 ( .ZN(net_8199), .A(net_5516) );
NAND3_X2 inst_6816 ( .ZN(net_4420), .A3(net_1454), .A2(net_375), .A1(x7654) );
NOR2_X2 inst_4333 ( .A1(net_13940), .A2(net_13885), .ZN(net_13119) );
OR3_X2 inst_1063 ( .ZN(net_2680), .A1(net_2486), .A3(net_1922), .A2(net_75) );
CLKBUF_X2 inst_22721 ( .A(net_22592), .Z(net_22593) );
NOR3_X2 inst_2700 ( .ZN(net_19824), .A3(net_11342), .A1(net_8880), .A2(net_8781) );
CLKBUF_X2 inst_21404 ( .A(net_21275), .Z(net_21276) );
NOR2_X4 inst_3252 ( .ZN(net_3012), .A2(net_1743), .A1(net_190) );
AOI22_X2 inst_19973 ( .ZN(net_15668), .A2(net_15017), .B2(net_11289), .B1(net_6587), .A1(net_852) );
INV_X4 inst_13542 ( .ZN(net_10769), .A(net_9199) );
NOR2_X2 inst_4565 ( .A1(net_7487), .ZN(net_3899), .A2(net_3898) );
NOR2_X2 inst_4755 ( .ZN(net_11221), .A2(net_7091), .A1(net_1732) );
CLKBUF_X2 inst_22617 ( .A(net_22488), .Z(net_22489) );
CLKBUF_X2 inst_22733 ( .A(net_22604), .Z(net_22605) );
INV_X2 inst_19100 ( .ZN(net_19961), .A(net_7727) );
NAND4_X2 inst_5276 ( .A2(net_20224), .A1(net_20223), .A4(net_20130), .ZN(net_19087), .A3(net_13939) );
INV_X4 inst_18203 ( .A(net_20896), .ZN(net_16368) );
INV_X4 inst_17375 ( .ZN(net_14945), .A(net_13362) );
OR2_X2 inst_1167 ( .ZN(net_7051), .A2(net_7050), .A1(net_6589) );
NAND2_X2 inst_9452 ( .A1(net_14554), .ZN(net_12629), .A2(net_11515) );
CLKBUF_X2 inst_22811 ( .A(net_22682), .Z(net_22683) );
NAND2_X4 inst_6879 ( .ZN(net_18232), .A1(net_18122), .A2(net_18109) );
INV_X4 inst_17931 ( .A(net_21024), .ZN(net_426) );
NAND2_X2 inst_8767 ( .ZN(net_15877), .A1(net_15810), .A2(net_15423) );
INV_X4 inst_14595 ( .ZN(net_14070), .A(net_11786) );
OAI22_X2 inst_1303 ( .B1(net_13709), .ZN(net_10505), .A1(net_10504), .A2(net_10503), .B2(net_10502) );
OAI21_X2 inst_1623 ( .A(net_21228), .ZN(net_16068), .B2(net_15478), .B1(net_6649) );
NOR2_X2 inst_4088 ( .ZN(net_8806), .A1(net_5962), .A2(net_5562) );
INV_X4 inst_12788 ( .ZN(net_18291), .A(net_17293) );
AOI21_X2 inst_20773 ( .A(net_14227), .B2(net_13883), .ZN(net_10632), .B1(net_10631) );
NAND3_X2 inst_6163 ( .A2(net_20763), .ZN(net_13635), .A3(net_12689), .A1(net_10925) );
NOR2_X2 inst_4922 ( .ZN(net_11208), .A1(net_6538), .A2(net_1844) );
NAND2_X2 inst_8369 ( .ZN(net_19018), .A1(net_17371), .A2(net_17209) );
CLKBUF_X2 inst_22301 ( .A(net_21836), .Z(net_22173) );
NOR2_X2 inst_3452 ( .ZN(net_14877), .A2(net_13763), .A1(net_10138) );
NAND2_X2 inst_10183 ( .ZN(net_8182), .A1(net_8181), .A2(net_6302) );
INV_X4 inst_17708 ( .A(net_826), .ZN(net_208) );
OAI21_X2 inst_1516 ( .ZN(net_18503), .B1(net_18470), .A(net_18391), .B2(net_18390) );
INV_X2 inst_19047 ( .ZN(net_4746), .A(net_4745) );
INV_X4 inst_14695 ( .ZN(net_18581), .A(net_18025) );
XNOR2_X2 inst_386 ( .ZN(net_16782), .A(net_16780), .B(net_12875) );
NAND2_X2 inst_8497 ( .ZN(net_17083), .A1(net_16617), .A2(net_16477) );
INV_X8 inst_12372 ( .ZN(net_1270), .A(net_931) );
INV_X4 inst_15110 ( .ZN(net_4251), .A(net_3199) );
NAND2_X4 inst_7255 ( .ZN(net_8736), .A2(net_6177), .A1(net_4939) );
NAND2_X2 inst_10543 ( .ZN(net_10484), .A1(net_6788), .A2(net_5667) );
INV_X4 inst_16914 ( .ZN(net_1625), .A(net_762) );
NAND2_X2 inst_9863 ( .ZN(net_9492), .A1(net_6601), .A2(net_6196) );
CLKBUF_X2 inst_21478 ( .A(net_21349), .Z(net_21350) );
INV_X2 inst_18780 ( .ZN(net_7518), .A(net_7517) );
NAND2_X2 inst_8089 ( .ZN(net_18133), .A2(net_18106), .A1(net_17022) );
NAND2_X2 inst_7826 ( .ZN(net_18643), .A1(net_18642), .A2(net_18632) );
NAND2_X2 inst_11040 ( .ZN(net_11263), .A1(net_4737), .A2(net_4736) );
INV_X4 inst_16220 ( .ZN(net_2416), .A(net_1605) );
NAND4_X4 inst_5225 ( .ZN(net_16556), .A4(net_16184), .A2(net_16021), .A1(net_15987), .A3(net_15874) );
INV_X4 inst_16620 ( .A(net_1451), .ZN(net_1116) );
NAND4_X2 inst_5320 ( .A2(net_19917), .A1(net_19916), .ZN(net_15768), .A4(net_14101), .A3(net_8843) );
NOR3_X2 inst_2778 ( .ZN(net_7734), .A2(net_5309), .A1(net_4505), .A3(net_2131) );
NAND2_X2 inst_9826 ( .ZN(net_9627), .A1(net_9626), .A2(net_9625) );
NAND2_X2 inst_10173 ( .A1(net_8798), .ZN(net_8208), .A2(net_8207) );
NAND2_X2 inst_11883 ( .ZN(net_5300), .A1(net_3844), .A2(net_836) );
NAND4_X4 inst_5223 ( .A4(net_18878), .A1(net_18877), .ZN(net_16340), .A2(net_16022), .A3(net_15735) );
NAND4_X2 inst_5468 ( .ZN(net_13221), .A2(net_13220), .A1(net_11705), .A4(net_10036), .A3(net_9875) );
INV_X2 inst_19072 ( .ZN(net_4627), .A(net_4626) );
INV_X4 inst_17265 ( .ZN(net_3844), .A(net_193) );
NAND2_X2 inst_9599 ( .ZN(net_10760), .A1(net_10759), .A2(net_7371) );
NAND2_X2 inst_8716 ( .ZN(net_20095), .A2(net_15998), .A1(net_13083) );
NAND2_X2 inst_10060 ( .ZN(net_8683), .A1(net_8682), .A2(net_8681) );
NAND2_X2 inst_11064 ( .A2(net_5649), .ZN(net_4525), .A1(net_3463) );
SDFF_X2 inst_811 ( .Q(net_21121), .SI(net_17830), .SE(net_125), .CK(net_21567), .D(x4345) );
INV_X8 inst_12375 ( .ZN(net_287), .A(net_128) );
CLKBUF_X2 inst_21393 ( .A(net_21253), .Z(net_21265) );
INV_X2 inst_19578 ( .ZN(net_907), .A(net_204) );
NAND2_X2 inst_9591 ( .ZN(net_12626), .A1(net_10864), .A2(net_9134) );
INV_X4 inst_16447 ( .ZN(net_15110), .A(net_10683) );
AND2_X4 inst_21252 ( .A1(net_20897), .ZN(net_8117), .A2(net_308) );
NOR2_X2 inst_3909 ( .ZN(net_8859), .A2(net_6498), .A1(net_4078) );
INV_X4 inst_18296 ( .A(net_20469), .ZN(net_20467) );
OAI21_X2 inst_1869 ( .ZN(net_13730), .B2(net_12666), .B1(net_10799), .A(net_1399) );
SDFF_X2 inst_897 ( .Q(net_21118), .D(net_16755), .SE(net_263), .CK(net_21533), .SI(x4444) );
AOI21_X2 inst_20527 ( .ZN(net_14550), .B1(net_13032), .B2(net_11926), .A(net_6263) );
NOR2_X2 inst_3945 ( .A1(net_12050), .ZN(net_8628), .A2(net_6389) );
INV_X4 inst_15592 ( .ZN(net_12478), .A(net_2243) );
OR2_X2 inst_1201 ( .A2(net_6429), .ZN(net_3778), .A1(net_3777) );
NAND2_X2 inst_11656 ( .ZN(net_3336), .A1(net_2431), .A2(net_2291) );
CLKBUF_X2 inst_22329 ( .A(net_21774), .Z(net_22201) );
NAND2_X2 inst_8760 ( .ZN(net_19139), .A2(net_15539), .A1(net_15275) );
DFF_X1 inst_19890 ( .D(net_16883), .CK(net_21975), .Q(x923) );
NAND3_X2 inst_5899 ( .ZN(net_15161), .A3(net_13936), .A2(net_11175), .A1(net_9091) );
NAND2_X2 inst_9294 ( .ZN(net_12407), .A1(net_12406), .A2(net_12405) );
INV_X4 inst_18331 ( .A(net_20563), .ZN(net_20562) );
OAI21_X2 inst_1927 ( .A(net_14720), .ZN(net_12955), .B1(net_12954), .B2(net_9720) );
AOI22_X2 inst_19991 ( .ZN(net_14752), .B1(net_14751), .A1(net_14085), .A2(net_12281), .B2(net_5663) );
XNOR2_X2 inst_184 ( .A(net_17777), .ZN(net_17764), .B(net_17763) );
OAI21_X2 inst_1847 ( .ZN(net_20723), .A(net_14014), .B2(net_10318), .B1(net_4713) );
NAND2_X2 inst_8878 ( .ZN(net_15210), .A1(net_14283), .A2(net_14196) );
INV_X8 inst_12270 ( .ZN(net_11526), .A(net_10323) );
INV_X4 inst_16312 ( .ZN(net_9861), .A(net_112) );
NAND2_X4 inst_6921 ( .A2(net_20462), .ZN(net_19604), .A1(net_17100) );
NAND2_X2 inst_8775 ( .ZN(net_15824), .A2(net_15327), .A1(net_14942) );
AOI21_X4 inst_20240 ( .ZN(net_11155), .B1(net_7464), .A(net_2370), .B2(net_1173) );
NAND2_X2 inst_7742 ( .ZN(net_18798), .A2(net_18767), .A1(net_17637) );
NAND2_X2 inst_9409 ( .ZN(net_11662), .A1(net_11661), .A2(net_11099) );
NAND2_X2 inst_9125 ( .ZN(net_13533), .A2(net_13532), .A1(net_10955) );
NAND2_X2 inst_10919 ( .ZN(net_5992), .A1(net_4865), .A2(net_2638) );
INV_X4 inst_15950 ( .ZN(net_2366), .A(net_1710) );
INV_X4 inst_17270 ( .ZN(net_1397), .A(net_280) );
INV_X4 inst_17654 ( .A(net_602), .ZN(net_532) );
CLKBUF_X2 inst_21753 ( .A(net_21624), .Z(net_21625) );
INV_X2 inst_19372 ( .ZN(net_19286), .A(net_1834) );
OAI21_X2 inst_2114 ( .A(net_10714), .ZN(net_10035), .B2(net_10034), .B1(net_6191) );
NOR3_X2 inst_2784 ( .ZN(net_6447), .A1(net_6446), .A2(net_6445), .A3(net_6444) );
NAND3_X2 inst_6330 ( .ZN(net_12470), .A2(net_7815), .A3(net_7569), .A1(net_4986) );
INV_X4 inst_13817 ( .ZN(net_12520), .A(net_7521) );
INV_X4 inst_13001 ( .A(net_16780), .ZN(net_16777) );
INV_X4 inst_16105 ( .ZN(net_2124), .A(net_1502) );
NAND2_X2 inst_9036 ( .A1(net_14636), .ZN(net_14062), .A2(net_11831) );
NAND2_X2 inst_10538 ( .ZN(net_8768), .A1(net_7325), .A2(net_6841) );
NAND2_X4 inst_7149 ( .ZN(net_9639), .A2(net_9638), .A1(net_9274) );
INV_X4 inst_16627 ( .ZN(net_19660), .A(net_1301) );
INV_X4 inst_13458 ( .A(net_10221), .ZN(net_9722) );
INV_X4 inst_13697 ( .A(net_7927), .ZN(net_7922) );
NOR2_X2 inst_4377 ( .ZN(net_5379), .A2(net_5378), .A1(net_4074) );
NOR2_X2 inst_4301 ( .A1(net_9571), .ZN(net_5941), .A2(net_5940) );
INV_X4 inst_16046 ( .ZN(net_15684), .A(net_13525) );
INV_X4 inst_13432 ( .ZN(net_20678), .A(net_9869) );
NAND2_X2 inst_8537 ( .A2(net_20216), .A1(net_17359), .ZN(net_16855) );
INV_X4 inst_16188 ( .ZN(net_12551), .A(net_11016) );
INV_X4 inst_15018 ( .ZN(net_20401), .A(net_15926) );
NOR2_X2 inst_5106 ( .A1(net_761), .ZN(net_759), .A2(net_758) );
OAI21_X4 inst_1410 ( .A(net_20896), .B2(net_19191), .B1(net_19190), .ZN(net_16176) );
INV_X4 inst_14943 ( .ZN(net_8542), .A(net_3524) );
INV_X4 inst_16510 ( .ZN(net_2489), .A(net_1081) );
NAND2_X2 inst_10675 ( .ZN(net_9056), .A1(net_6081), .A2(net_5806) );
NOR2_X2 inst_4424 ( .ZN(net_7948), .A2(net_2765), .A1(net_1163) );
AND2_X2 inst_21356 ( .ZN(net_3941), .A2(net_1481), .A1(net_955) );
NAND2_X4 inst_7028 ( .ZN(net_17571), .A1(net_16566), .A2(net_16563) );
NAND3_X2 inst_5994 ( .ZN(net_14528), .A1(net_13392), .A3(net_7331), .A2(net_4680) );
INV_X2 inst_19067 ( .ZN(net_4636), .A(net_3308) );
NAND2_X2 inst_10210 ( .A1(net_10113), .ZN(net_9608), .A2(net_8101) );
INV_X2 inst_18952 ( .A(net_11656), .ZN(net_5604) );
NAND3_X2 inst_6653 ( .A3(net_13472), .ZN(net_8545), .A1(net_3377), .A2(net_2738) );
INV_X4 inst_18284 ( .A(net_20079), .ZN(net_20078) );
OAI21_X2 inst_2074 ( .ZN(net_10591), .B1(net_10590), .A(net_9759), .B2(net_6442) );
NAND2_X2 inst_11330 ( .A1(net_7396), .ZN(net_3735), .A2(net_3734) );
NAND2_X4 inst_7296 ( .ZN(net_9099), .A1(net_6854), .A2(net_2404) );
NOR2_X2 inst_4823 ( .A2(net_6041), .ZN(net_4313), .A1(net_2532) );
OR2_X2 inst_1236 ( .A1(net_2329), .ZN(net_1580), .A2(net_1261) );
XNOR2_X2 inst_221 ( .ZN(net_17510), .A(net_17500), .B(net_7740) );
AOI21_X2 inst_20395 ( .ZN(net_15459), .B2(net_14451), .B1(net_13983), .A(net_828) );
NOR2_X2 inst_5112 ( .ZN(net_6563), .A1(net_602), .A2(net_304) );
NAND3_X2 inst_5929 ( .ZN(net_14934), .A2(net_14933), .A1(net_13637), .A3(net_11254) );
NOR2_X4 inst_3313 ( .ZN(net_1593), .A2(net_990), .A1(net_241) );
INV_X4 inst_12640 ( .ZN(net_17908), .A(net_17907) );
NOR2_X2 inst_3562 ( .ZN(net_18991), .A2(net_12616), .A1(net_12147) );
NAND2_X2 inst_9545 ( .ZN(net_11046), .A1(net_11045), .A2(net_9869) );
INV_X4 inst_13502 ( .ZN(net_12866), .A(net_9431) );
INV_X2 inst_18635 ( .A(net_11839), .ZN(net_9399) );
OAI21_X2 inst_2334 ( .ZN(net_4686), .A(net_4685), .B1(net_3590), .B2(net_2255) );
NAND2_X2 inst_11967 ( .ZN(net_1835), .A2(net_831), .A1(net_279) );
AND4_X2 inst_21099 ( .A3(net_12907), .ZN(net_12799), .A4(net_12798), .A1(net_12096), .A2(net_8096) );
INV_X4 inst_17261 ( .A(net_10676), .ZN(net_8868) );
OAI21_X2 inst_2210 ( .A(net_13538), .ZN(net_8531), .B1(net_5563), .B2(net_4531) );
NAND3_X2 inst_6040 ( .ZN(net_14323), .A3(net_13780), .A2(net_13306), .A1(net_12367) );
NOR2_X2 inst_5028 ( .ZN(net_4085), .A2(net_860), .A1(net_222) );
OAI211_X2 inst_2590 ( .ZN(net_5512), .B(net_5511), .C2(net_5510), .A(net_2304), .C1(net_25) );
NAND2_X2 inst_11577 ( .A1(net_6604), .ZN(net_6491), .A2(net_2739) );
NAND2_X2 inst_10949 ( .ZN(net_7279), .A2(net_5114), .A1(net_112) );
NAND2_X2 inst_10435 ( .A2(net_13456), .ZN(net_7201), .A1(net_6705) );
NOR2_X2 inst_5025 ( .A2(net_20799), .A1(net_6606), .ZN(net_1575) );
INV_X4 inst_16947 ( .ZN(net_4990), .A(net_4815) );
INV_X2 inst_18739 ( .A(net_11948), .ZN(net_7911) );
INV_X4 inst_13341 ( .ZN(net_12413), .A(net_11084) );
INV_X4 inst_18340 ( .A(net_20711), .ZN(net_20709) );
INV_X4 inst_17900 ( .ZN(net_2246), .A(net_1848) );
CLKBUF_X2 inst_22135 ( .A(net_22006), .Z(net_22007) );
INV_X8 inst_12451 ( .A(net_20923), .ZN(net_20548) );
NOR2_X2 inst_4459 ( .ZN(net_6365), .A1(net_6081), .A2(net_4645) );
INV_X4 inst_15261 ( .ZN(net_11382), .A(net_2772) );
INV_X4 inst_14028 ( .ZN(net_6288), .A(net_6287) );
OR2_X4 inst_1117 ( .ZN(net_7679), .A1(net_790), .A2(net_134) );
NAND2_X4 inst_7343 ( .A2(net_20491), .ZN(net_7887), .A1(net_3562) );
NOR2_X2 inst_4015 ( .ZN(net_11322), .A1(net_8037), .A2(net_6871) );
NAND2_X2 inst_11374 ( .ZN(net_3564), .A1(net_1914), .A2(net_1201) );
INV_X4 inst_13909 ( .ZN(net_8894), .A(net_7014) );
INV_X2 inst_19597 ( .A(net_321), .ZN(net_198) );
NAND2_X4 inst_6887 ( .ZN(net_18204), .A2(net_18103), .A1(net_18088) );
NOR3_X2 inst_2725 ( .ZN(net_13249), .A1(net_10591), .A2(net_10459), .A3(net_9949) );
NAND3_X2 inst_6681 ( .ZN(net_7736), .A1(net_6137), .A3(net_5970), .A2(net_3882) );
NOR2_X2 inst_5141 ( .A2(net_1733), .A1(net_874), .ZN(net_149) );
INV_X4 inst_14476 ( .A(net_8448), .ZN(net_6037) );
NAND2_X2 inst_8204 ( .ZN(net_17917), .A2(net_17719), .A1(net_17626) );
OAI21_X2 inst_1610 ( .ZN(net_16120), .B1(net_16046), .B2(net_15726), .A(net_14488) );
XNOR2_X2 inst_334 ( .B(net_17522), .A(net_17000), .ZN(net_16989) );
INV_X4 inst_13337 ( .A(net_12746), .ZN(net_12422) );
SDFF_X2 inst_1042 ( .QN(net_21047), .D(net_435), .SE(net_263), .CK(net_22494), .SI(x2230) );
INV_X4 inst_14190 ( .A(net_8002), .ZN(net_5978) );
INV_X2 inst_19238 ( .ZN(net_3317), .A(net_2006) );
NAND3_X2 inst_5961 ( .ZN(net_19619), .A3(net_13447), .A2(net_12533), .A1(net_9682) );
INV_X4 inst_15850 ( .ZN(net_2797), .A(net_1825) );
NAND3_X4 inst_5595 ( .ZN(net_19025), .A3(net_12290), .A1(net_11666), .A2(net_4036) );
NAND2_X2 inst_8153 ( .ZN(net_18007), .A1(net_17954), .A2(net_17929) );
INV_X2 inst_19420 ( .ZN(net_2945), .A(net_1845) );
INV_X4 inst_17068 ( .ZN(net_10022), .A(net_6570) );
INV_X2 inst_18497 ( .ZN(net_12309), .A(net_12308) );
NAND2_X2 inst_8058 ( .ZN(net_18203), .A1(net_18145), .A2(net_18120) );
XNOR2_X2 inst_595 ( .A(net_16402), .ZN(net_553), .B(net_552) );
INV_X4 inst_13255 ( .ZN(net_20727), .A(net_11700) );
NOR2_X2 inst_5002 ( .ZN(net_2735), .A2(net_1356), .A1(net_154) );
NAND2_X2 inst_8222 ( .A2(net_17875), .ZN(net_17816), .A1(net_17815) );
NAND3_X2 inst_6343 ( .A3(net_15694), .A2(net_14706), .ZN(net_12251), .A1(net_9057) );
INV_X4 inst_13554 ( .ZN(net_12378), .A(net_9163) );
NAND2_X2 inst_9014 ( .ZN(net_14257), .A2(net_12671), .A1(net_10198) );
INV_X2 inst_19035 ( .ZN(net_4858), .A(net_4857) );
AOI21_X4 inst_20191 ( .ZN(net_20375), .B1(net_15205), .B2(net_14109), .A(net_12256) );
NOR2_X2 inst_4688 ( .A1(net_3334), .ZN(net_3189), .A2(net_1739) );
INV_X4 inst_12658 ( .ZN(net_17819), .A(net_17818) );
INV_X4 inst_15451 ( .ZN(net_2598), .A(net_2491) );
INV_X4 inst_17833 ( .ZN(net_3297), .A(net_102) );
INV_X4 inst_17219 ( .ZN(net_6719), .A(net_703) );
NOR2_X2 inst_4798 ( .A2(net_5256), .ZN(net_3521), .A1(net_1482) );
AOI21_X4 inst_20110 ( .ZN(net_19145), .B1(net_16242), .B2(net_16085), .A(net_16071) );
NOR2_X2 inst_3849 ( .A2(net_12287), .ZN(net_11548), .A1(net_9542) );
INV_X8 inst_12205 ( .ZN(net_11015), .A(net_5763) );
INV_X4 inst_15575 ( .A(net_9903), .ZN(net_7688) );
INV_X4 inst_15840 ( .A(net_14622), .ZN(net_14617) );
INV_X2 inst_19188 ( .A(net_5200), .ZN(net_3685) );
SDFF_X2 inst_1029 ( .QN(net_21065), .D(net_619), .SE(net_253), .CK(net_21705), .SI(x1987) );
NAND4_X2 inst_5413 ( .ZN(net_14586), .A2(net_12451), .A4(net_8522), .A3(net_8023), .A1(net_7032) );
NAND3_X2 inst_6666 ( .ZN(net_8439), .A3(net_8438), .A2(net_4829), .A1(net_3887) );
NAND2_X2 inst_9246 ( .ZN(net_20393), .A2(net_12673), .A1(net_11432) );
NAND2_X4 inst_6841 ( .A2(net_19164), .A1(net_19163), .ZN(net_18692) );
CLKBUF_X2 inst_22226 ( .A(net_22097), .Z(net_22098) );
CLKBUF_X2 inst_22110 ( .A(net_21981), .Z(net_21982) );
NAND2_X4 inst_7032 ( .A2(net_19412), .A1(net_19411), .ZN(net_17166) );
NAND3_X2 inst_6245 ( .A2(net_13481), .ZN(net_13172), .A3(net_13171), .A1(net_7222) );
NAND3_X2 inst_6551 ( .ZN(net_10531), .A3(net_10530), .A2(net_7527), .A1(net_5238) );
NAND3_X2 inst_5767 ( .ZN(net_15902), .A3(net_15383), .A2(net_13993), .A1(net_10234) );
INV_X4 inst_13048 ( .A(net_17290), .ZN(net_17177) );
NAND2_X2 inst_10067 ( .A2(net_13776), .ZN(net_10128), .A1(net_8664) );
NAND3_X2 inst_6443 ( .ZN(net_11803), .A2(net_9315), .A3(net_7919), .A1(net_5518) );
INV_X2 inst_19546 ( .ZN(net_923), .A(net_922) );
INV_X4 inst_14404 ( .A(net_6799), .ZN(net_5103) );
OAI21_X2 inst_1534 ( .ZN(net_17991), .A(net_17891), .B1(net_17890), .B2(net_17889) );
NAND2_X2 inst_9985 ( .A1(net_10054), .ZN(net_8850), .A2(net_6505) );
CLKBUF_X2 inst_22792 ( .A(net_22663), .Z(net_22664) );
XNOR2_X2 inst_319 ( .ZN(net_17042), .A(net_16647), .B(net_713) );
NAND2_X2 inst_9108 ( .ZN(net_13706), .A1(net_13705), .A2(net_10230) );
OAI211_X2 inst_2422 ( .ZN(net_15271), .C1(net_15270), .C2(net_14847), .B(net_13800), .A(net_10265) );
INV_X4 inst_12745 ( .ZN(net_17429), .A(net_17428) );
NAND2_X2 inst_10688 ( .ZN(net_7514), .A2(net_6153), .A1(net_6092) );
XNOR2_X2 inst_649 ( .B(net_16404), .ZN(net_383), .A(net_382) );
INV_X2 inst_18724 ( .ZN(net_20274), .A(net_8104) );
NAND3_X2 inst_5790 ( .ZN(net_15740), .A1(net_15125), .A3(net_15003), .A2(net_8853) );
INV_X2 inst_18676 ( .ZN(net_9105), .A(net_9104) );
INV_X4 inst_15166 ( .A(net_10386), .ZN(net_3828) );
CLKBUF_X2 inst_21806 ( .A(net_21677), .Z(net_21678) );
OAI211_X2 inst_2597 ( .C2(net_6537), .B(net_5367), .ZN(net_5251), .C1(net_5250), .A(net_2056) );
NAND2_X2 inst_8504 ( .A2(net_20498), .ZN(net_16927), .A1(net_15294) );
INV_X4 inst_16379 ( .A(net_9396), .ZN(net_6625) );
INV_X4 inst_14269 ( .ZN(net_9274), .A(net_5691) );
NAND3_X4 inst_5569 ( .A3(net_20376), .A1(net_20375), .ZN(net_15921), .A2(net_14180) );
NAND4_X4 inst_5185 ( .A4(net_19136), .A1(net_19135), .ZN(net_16732), .A3(net_15761), .A2(net_10828) );
INV_X8 inst_12227 ( .ZN(net_4590), .A(net_2818) );
NAND3_X2 inst_6059 ( .ZN(net_14199), .A1(net_13968), .A3(net_12261), .A2(net_11215) );
OAI21_X2 inst_1575 ( .A(net_20952), .ZN(net_19969), .B2(net_16048), .B1(net_12585) );
INV_X4 inst_17453 ( .ZN(net_7455), .A(net_86) );
CLKBUF_X2 inst_22027 ( .A(net_21395), .Z(net_21899) );
NAND2_X2 inst_9644 ( .A1(net_20205), .ZN(net_19723), .A2(net_749) );
INV_X2 inst_19653 ( .ZN(net_20100), .A(net_20077) );
INV_X4 inst_16300 ( .ZN(net_5900), .A(net_2199) );
NAND3_X4 inst_5522 ( .ZN(net_18633), .A2(net_18593), .A3(net_18592), .A1(net_15875) );
OAI22_X2 inst_1258 ( .B1(net_21136), .A2(net_20713), .B2(net_20710), .ZN(net_17591), .A1(net_16836) );
NOR2_X4 inst_3141 ( .ZN(net_5226), .A1(net_3717), .A2(net_2585) );
NAND2_X2 inst_10148 ( .ZN(net_8294), .A1(net_8293), .A2(net_6189) );
NOR2_X2 inst_3921 ( .ZN(net_8787), .A2(net_8136), .A1(net_8008) );
INV_X4 inst_16820 ( .A(net_8220), .ZN(net_7298) );
OAI21_X2 inst_1957 ( .ZN(net_12534), .A(net_11260), .B1(net_9903), .B2(net_7468) );
NOR2_X1 inst_5151 ( .A1(net_15108), .A2(net_13620), .ZN(net_8017) );
NAND2_X2 inst_9524 ( .ZN(net_11125), .A1(net_11124), .A2(net_11065) );
INV_X4 inst_13860 ( .ZN(net_12273), .A(net_11209) );
NAND2_X4 inst_7446 ( .ZN(net_4060), .A1(net_3121), .A2(net_955) );
NAND2_X2 inst_10456 ( .ZN(net_7029), .A2(net_7028), .A1(net_4260) );
AOI211_X2 inst_21055 ( .C1(net_13700), .ZN(net_11755), .A(net_11754), .B(net_11753), .C2(net_11001) );
INV_X4 inst_13813 ( .ZN(net_7535), .A(net_7534) );
NOR2_X2 inst_4624 ( .ZN(net_3605), .A1(net_2117), .A2(net_1129) );
NAND2_X2 inst_7811 ( .ZN(net_18738), .A1(net_18654), .A2(net_17774) );
INV_X8 inst_12458 ( .ZN(net_20787), .A(net_17045) );
NAND2_X2 inst_11257 ( .A2(net_20868), .ZN(net_3913), .A1(net_2814) );
CLKBUF_X2 inst_21703 ( .A(net_21574), .Z(net_21575) );
AND3_X2 inst_21143 ( .ZN(net_8549), .A3(net_8444), .A1(net_6284), .A2(net_4249) );
INV_X2 inst_18597 ( .ZN(net_9980), .A(net_9979) );
NAND3_X2 inst_6062 ( .ZN(net_14182), .A3(net_13716), .A1(net_12474), .A2(net_6192) );
NAND2_X2 inst_9254 ( .ZN(net_14295), .A1(net_12885), .A2(net_12649) );
NAND2_X4 inst_7428 ( .ZN(net_5937), .A1(net_3491), .A2(net_2552) );
NAND2_X2 inst_7778 ( .A1(net_19719), .ZN(net_18777), .A2(net_18730) );
NAND3_X2 inst_6608 ( .ZN(net_9292), .A2(net_9291), .A3(net_3320), .A1(net_2393) );
NOR2_X4 inst_2983 ( .ZN(net_11388), .A2(net_6150), .A1(net_4549) );
INV_X1 inst_19759 ( .A(net_5393), .ZN(net_3417) );
NAND2_X4 inst_7421 ( .ZN(net_7702), .A1(net_3542), .A2(net_2087) );
INV_X4 inst_13233 ( .ZN(net_13476), .A(net_12445) );
INV_X4 inst_13584 ( .A(net_10746), .ZN(net_8914) );
NAND2_X2 inst_8862 ( .A1(net_15864), .ZN(net_15342), .A2(net_14385) );
NAND2_X2 inst_9969 ( .A1(net_11984), .ZN(net_8892), .A2(net_8368) );
INV_X4 inst_12881 ( .A(net_16919), .ZN(net_16823) );
INV_X2 inst_19353 ( .ZN(net_2378), .A(net_2377) );
OR2_X4 inst_1120 ( .ZN(net_6520), .A2(net_222), .A1(net_98) );
AOI21_X2 inst_20367 ( .ZN(net_15634), .B2(net_14429), .A(net_11867), .B1(net_238) );
NAND3_X2 inst_6238 ( .ZN(net_13208), .A3(net_9978), .A2(net_5781), .A1(net_5762) );
INV_X4 inst_12986 ( .A(net_16996), .ZN(net_16641) );
INV_X4 inst_16035 ( .A(net_10309), .ZN(net_1986) );
AOI21_X2 inst_20263 ( .B2(net_20880), .ZN(net_18069), .A(net_18051), .B1(net_16117) );
NAND2_X2 inst_8545 ( .A1(net_17487), .ZN(net_16816), .A2(net_16815) );
INV_X4 inst_15029 ( .ZN(net_4583), .A(net_3565) );
NOR2_X4 inst_3184 ( .ZN(net_5485), .A1(net_3115), .A2(net_1592) );
NAND3_X2 inst_6398 ( .ZN(net_11992), .A2(net_10520), .A3(net_8144), .A1(net_7985) );
NAND2_X2 inst_9715 ( .ZN(net_10171), .A1(net_10170), .A2(net_7709) );
SDFF_X2 inst_947 ( .QN(net_21017), .D(net_576), .SE(net_263), .CK(net_21900), .SI(x2745) );
SDFF_X2 inst_731 ( .Q(net_20937), .SE(net_18585), .SI(net_18564), .D(net_11883), .CK(net_22762) );
INV_X4 inst_15381 ( .ZN(net_3567), .A(net_3380) );
NAND2_X2 inst_10909 ( .A2(net_6692), .ZN(net_5912), .A1(net_5370) );
INV_X4 inst_13788 ( .ZN(net_9201), .A(net_7567) );
INV_X4 inst_15005 ( .A(net_4438), .ZN(net_3387) );
OAI211_X2 inst_2459 ( .ZN(net_14212), .A(net_14211), .B(net_14210), .C2(net_14209), .C1(net_6363) );
DFF_X1 inst_19812 ( .QN(net_21193), .D(net_18004), .CK(net_21446) );
NAND2_X4 inst_7165 ( .ZN(net_12816), .A1(net_9512), .A2(net_8868) );
XNOR2_X2 inst_301 ( .A(net_20707), .ZN(net_17114), .B(net_17113) );
XNOR2_X2 inst_363 ( .B(net_21178), .ZN(net_16877), .A(net_16876) );
OAI21_X2 inst_2141 ( .ZN(net_9970), .A(net_9969), .B1(net_9968), .B2(net_9967) );
CLKBUF_X2 inst_22033 ( .A(net_21904), .Z(net_21905) );
NAND2_X2 inst_12041 ( .ZN(net_953), .A2(net_386), .A1(net_290) );
CLKBUF_X2 inst_22179 ( .A(net_22050), .Z(net_22051) );
NAND3_X2 inst_6609 ( .ZN(net_9288), .A2(net_5848), .A1(net_4202), .A3(net_1579) );
NAND2_X4 inst_7079 ( .A2(net_20746), .A1(net_20745), .ZN(net_15806) );
INV_X4 inst_13213 ( .ZN(net_19052), .A(net_12820) );
NAND2_X2 inst_7870 ( .ZN(net_18546), .A1(net_18503), .A2(net_18221) );
INV_X4 inst_14021 ( .ZN(net_10348), .A(net_8249) );
INV_X2 inst_19000 ( .A(net_8444), .ZN(net_5056) );
NOR2_X2 inst_4706 ( .ZN(net_5618), .A1(net_3929), .A2(net_1879) );
NOR2_X2 inst_4348 ( .ZN(net_19056), .A2(net_6299), .A1(net_4224) );
AOI21_X2 inst_20608 ( .ZN(net_20328), .B1(net_14966), .A(net_12679), .B2(net_10842) );
NOR2_X2 inst_3729 ( .ZN(net_10887), .A1(net_9932), .A2(net_7505) );
INV_X4 inst_14312 ( .ZN(net_5497), .A(net_5496) );
NAND2_X2 inst_8521 ( .ZN(net_16907), .A2(net_16734), .A1(net_16632) );
NAND2_X4 inst_7548 ( .ZN(net_2014), .A1(net_1798), .A2(net_1797) );
NAND2_X2 inst_10430 ( .A1(net_11572), .ZN(net_7212), .A2(net_7192) );
NAND2_X2 inst_8345 ( .ZN(net_19096), .A1(net_17483), .A2(net_17213) );
NAND2_X2 inst_9282 ( .ZN(net_12557), .A2(net_9718), .A1(net_7394) );
CLKBUF_X2 inst_21470 ( .A(net_21341), .Z(net_21342) );
NOR3_X2 inst_2650 ( .ZN(net_15492), .A3(net_14576), .A2(net_14253), .A1(net_13489) );
NAND2_X2 inst_11687 ( .A2(net_19418), .ZN(net_2335), .A1(net_1719) );
INV_X4 inst_14559 ( .A(net_4569), .ZN(net_4568) );
INV_X4 inst_16102 ( .ZN(net_2913), .A(net_1507) );
NOR2_X2 inst_4508 ( .A1(net_6945), .A2(net_6391), .ZN(net_5182) );
INV_X4 inst_16791 ( .ZN(net_3929), .A(net_1747) );
NAND2_X2 inst_7943 ( .ZN(net_18421), .A1(net_18420), .A2(net_18419) );
INV_X4 inst_16134 ( .ZN(net_10875), .A(net_1478) );
NAND2_X2 inst_11626 ( .ZN(net_4047), .A2(net_2295), .A1(net_2274) );
NAND2_X2 inst_9490 ( .ZN(net_14333), .A1(net_11442), .A2(net_10912) );
CLKBUF_X2 inst_22473 ( .A(net_22344), .Z(net_22345) );
NAND2_X2 inst_11666 ( .ZN(net_10844), .A1(net_4052), .A2(net_1488) );
INV_X4 inst_18315 ( .ZN(net_20517), .A(net_20516) );
NOR2_X4 inst_3189 ( .ZN(net_5709), .A1(net_3108), .A2(net_2462) );
AOI21_X2 inst_20938 ( .ZN(net_6467), .B2(net_6466), .B1(net_1589), .A(net_99) );
NAND2_X2 inst_8918 ( .ZN(net_14959), .A2(net_13715), .A1(net_9909) );
INV_X4 inst_12818 ( .ZN(net_17195), .A(net_17194) );
NAND2_X4 inst_6855 ( .A2(net_19949), .A1(net_19948), .ZN(net_18467) );
NAND3_X2 inst_5985 ( .ZN(net_19678), .A2(net_14541), .A3(net_14449), .A1(net_13382) );
NAND3_X4 inst_5548 ( .ZN(net_17517), .A3(net_16286), .A2(net_16212), .A1(net_11911) );
INV_X4 inst_14188 ( .ZN(net_5980), .A(net_5979) );
NAND2_X2 inst_10902 ( .ZN(net_6595), .A2(net_5384), .A1(net_4715) );
XNOR2_X1 inst_684 ( .ZN(net_17331), .B(net_17330), .A(net_17275) );
INV_X2 inst_19362 ( .A(net_3173), .ZN(net_2251) );
NAND3_X2 inst_6263 ( .A1(net_20751), .ZN(net_12975), .A2(net_12612), .A3(net_10433) );
NOR2_X2 inst_4400 ( .ZN(net_6277), .A2(net_4332), .A1(net_154) );
INV_X2 inst_19682 ( .A(net_20523), .ZN(net_20522) );
NOR2_X4 inst_3177 ( .A2(net_20565), .ZN(net_5593), .A1(net_1230) );
INV_X8 inst_12187 ( .ZN(net_17126), .A(net_16428) );
CLKBUF_X2 inst_22799 ( .A(net_22670), .Z(net_22671) );
NOR2_X2 inst_4930 ( .ZN(net_10164), .A1(net_989), .A2(net_120) );
NAND2_X2 inst_10437 ( .ZN(net_7197), .A1(net_7196), .A2(net_5249) );
NAND2_X2 inst_7965 ( .ZN(net_18368), .A1(net_18326), .A2(net_18287) );
AOI21_X2 inst_20624 ( .ZN(net_20321), .B1(net_14038), .B2(net_8950), .A(net_5555) );
INV_X2 inst_18585 ( .ZN(net_10283), .A(net_10282) );
NAND2_X2 inst_11857 ( .ZN(net_19574), .A2(net_1668), .A1(net_749) );
OR2_X2 inst_1138 ( .ZN(net_11514), .A2(net_11513), .A1(net_449) );
AOI21_X2 inst_20335 ( .ZN(net_20102), .B2(net_14818), .A(net_12275), .B1(net_8032) );
CLKBUF_X2 inst_22718 ( .A(net_22111), .Z(net_22590) );
NAND3_X2 inst_6568 ( .ZN(net_10473), .A3(net_10472), .A2(net_4768), .A1(net_3222) );
AND2_X4 inst_21244 ( .A1(net_6525), .A2(net_3462), .ZN(net_2792) );
SDFF_X2 inst_1004 ( .QN(net_20984), .D(net_382), .SE(net_263), .CK(net_22664), .SI(x3268) );
XNOR2_X2 inst_189 ( .ZN(net_17799), .A(net_17442), .B(net_17112) );
NAND2_X2 inst_9316 ( .ZN(net_12347), .A1(net_10930), .A2(net_8996) );
OAI211_X2 inst_2450 ( .ZN(net_14576), .B(net_12537), .C2(net_11191), .A(net_8849), .C1(net_3383) );
INV_X4 inst_13248 ( .ZN(net_12840), .A(net_11827) );
DFF_X1 inst_19821 ( .D(net_17680), .CK(net_21622), .Q(x719) );
NAND2_X4 inst_7437 ( .ZN(net_4410), .A1(net_3719), .A2(net_1970) );
NAND2_X2 inst_8597 ( .A1(net_20215), .A2(net_17233), .ZN(net_16686) );
INV_X4 inst_16190 ( .ZN(net_7988), .A(net_5077) );
NAND2_X4 inst_7430 ( .ZN(net_6612), .A1(net_3418), .A2(net_2154) );
XNOR2_X2 inst_62 ( .ZN(net_18815), .A(net_18755), .B(net_17764) );
NAND2_X2 inst_9529 ( .A2(net_19419), .ZN(net_11111), .A1(net_9138) );
NAND2_X2 inst_11006 ( .A2(net_9897), .A1(net_7975), .ZN(net_4884) );
NOR2_X2 inst_4696 ( .ZN(net_7058), .A2(net_2585), .A1(net_2250) );
NOR2_X2 inst_3743 ( .ZN(net_10617), .A2(net_8569), .A1(net_6737) );
INV_X4 inst_16247 ( .ZN(net_9735), .A(net_5918) );
NOR2_X4 inst_2860 ( .A2(net_13383), .ZN(net_12660), .A1(net_10972) );
NAND4_X4 inst_5194 ( .ZN(net_17763), .A1(net_16318), .A4(net_16043), .A2(net_15685), .A3(net_14859) );
INV_X4 inst_17713 ( .ZN(net_3356), .A(net_992) );
NAND2_X2 inst_8387 ( .A1(net_21139), .A2(net_19457), .ZN(net_17291) );
INV_X4 inst_14496 ( .ZN(net_7803), .A(net_6629) );
CLKBUF_X2 inst_21885 ( .A(net_21756), .Z(net_21757) );
NAND3_X2 inst_5888 ( .ZN(net_15227), .A3(net_14125), .A2(net_7794), .A1(net_2064) );
NAND2_X2 inst_11266 ( .A2(net_4669), .ZN(net_3896), .A1(net_2139) );
INV_X4 inst_17344 ( .A(net_9131), .ZN(net_6743) );
NAND2_X2 inst_11162 ( .ZN(net_7028), .A2(net_5230), .A1(net_4179) );
INV_X4 inst_13956 ( .A(net_6755), .ZN(net_6754) );
NAND2_X4 inst_7344 ( .ZN(net_7885), .A2(net_5333), .A1(net_4862) );
NAND2_X2 inst_8252 ( .ZN(net_17710), .A1(net_17530), .A2(net_17202) );
INV_X8 inst_12416 ( .A(net_20900), .ZN(net_1645) );
NOR2_X2 inst_4482 ( .A1(net_8748), .ZN(net_4338), .A2(net_4337) );
INV_X4 inst_15462 ( .ZN(net_15183), .A(net_2528) );
AOI21_X2 inst_20957 ( .B1(net_9146), .ZN(net_5335), .A(net_4169), .B2(net_3656) );
INV_X2 inst_19532 ( .ZN(net_19648), .A(net_1056) );
DFF_X1 inst_19788 ( .D(net_18659), .CK(net_22126), .Q(x563) );
INV_X4 inst_16713 ( .ZN(net_10233), .A(net_7325) );
DFF_X1 inst_19907 ( .D(net_16756), .CK(net_21582), .Q(x615) );
NAND2_X2 inst_7903 ( .ZN(net_18479), .A1(net_18478), .A2(net_18374) );
INV_X4 inst_18051 ( .A(net_21233), .ZN(net_227) );
SDFF_X2 inst_791 ( .Q(net_20885), .SE(net_18804), .SI(net_18031), .D(net_453), .CK(net_21800) );
INV_X4 inst_18016 ( .A(net_20990), .ZN(net_2472) );
NAND2_X2 inst_10427 ( .A2(net_9028), .ZN(net_7220), .A1(net_7219) );
INV_X4 inst_13371 ( .ZN(net_19909), .A(net_10899) );
OAI21_X2 inst_2021 ( .B1(net_13999), .B2(net_11927), .ZN(net_11334), .A(net_8971) );
NAND2_X2 inst_9631 ( .ZN(net_13879), .A1(net_10490), .A2(net_9344) );
INV_X2 inst_18424 ( .ZN(net_15264), .A(net_14864) );
NOR2_X2 inst_4379 ( .A1(net_10550), .ZN(net_5356), .A2(net_5355) );
NAND3_X2 inst_5668 ( .A3(net_20750), .A1(net_20749), .ZN(net_16381), .A2(net_16023) );
INV_X4 inst_13326 ( .ZN(net_11303), .A(net_11302) );
NOR2_X2 inst_5086 ( .A2(net_928), .ZN(net_851), .A1(net_83) );
INV_X4 inst_15107 ( .ZN(net_4934), .A(net_3211) );
INV_X4 inst_12811 ( .ZN(net_17207), .A(net_17206) );
INV_X4 inst_17983 ( .A(net_21187), .ZN(net_17097) );
INV_X4 inst_14670 ( .ZN(net_6421), .A(net_5465) );
NAND2_X2 inst_8576 ( .ZN(net_16728), .A2(net_16612), .A1(net_16486) );
INV_X4 inst_14399 ( .ZN(net_11315), .A(net_5116) );
NAND2_X2 inst_11924 ( .ZN(net_2049), .A1(net_1501), .A2(net_1316) );
INV_X4 inst_13020 ( .ZN(net_16488), .A(net_16422) );
NAND2_X2 inst_11888 ( .A1(net_2712), .ZN(net_1600), .A2(net_1599) );
CLKBUF_X2 inst_21863 ( .A(net_21311), .Z(net_21735) );
AOI21_X2 inst_20554 ( .ZN(net_14297), .A(net_13703), .B2(net_12424), .B1(net_5085) );
AOI21_X2 inst_20727 ( .ZN(net_11922), .B1(net_10672), .A(net_9920), .B2(net_5741) );
NAND2_X2 inst_7848 ( .A2(net_18601), .ZN(net_18595), .A1(net_15509) );
NAND2_X2 inst_8142 ( .ZN(net_18023), .A2(net_17991), .A1(net_17880) );
NAND3_X2 inst_6143 ( .A1(net_13840), .ZN(net_13690), .A3(net_11028), .A2(net_7410) );
INV_X2 inst_19231 ( .ZN(net_3366), .A(net_3365) );
NAND2_X4 inst_7304 ( .ZN(net_10567), .A2(net_5521), .A1(net_5472) );
INV_X4 inst_12864 ( .ZN(net_16993), .A(net_16992) );
CLKBUF_X2 inst_21732 ( .A(net_21603), .Z(net_21604) );
NOR2_X2 inst_4404 ( .A1(net_7903), .A2(net_7703), .ZN(net_5128) );
NAND2_X2 inst_8937 ( .ZN(net_14842), .A1(net_14511), .A2(net_13579) );
INV_X4 inst_18119 ( .A(net_21140), .ZN(net_17113) );
CLKBUF_X2 inst_21591 ( .A(net_21400), .Z(net_21463) );
NAND2_X2 inst_9054 ( .A1(net_15372), .ZN(net_14004), .A2(net_12008) );
NAND2_X2 inst_8154 ( .ZN(net_18002), .A2(net_17945), .A1(net_7386) );
NAND3_X2 inst_6581 ( .A3(net_12041), .ZN(net_10439), .A2(net_8087), .A1(net_7504) );
CLKBUF_X2 inst_22284 ( .A(net_21316), .Z(net_22156) );
INV_X4 inst_17651 ( .A(net_926), .ZN(net_338) );
NAND2_X2 inst_11261 ( .ZN(net_11801), .A1(net_3906), .A2(net_2057) );
INV_X4 inst_16130 ( .ZN(net_3331), .A(net_1208) );
INV_X2 inst_18395 ( .A(net_17010), .ZN(net_16876) );
NAND3_X2 inst_6716 ( .ZN(net_8916), .A1(net_7812), .A2(net_6876), .A3(net_5060) );
INV_X4 inst_15046 ( .ZN(net_13444), .A(net_9636) );
INV_X2 inst_19390 ( .ZN(net_2083), .A(net_2082) );
NAND3_X4 inst_5541 ( .ZN(net_17170), .A1(net_16493), .A3(net_15890), .A2(net_15272) );
AOI21_X2 inst_20709 ( .ZN(net_12101), .A(net_12100), .B1(net_12099), .B2(net_12088) );
AOI21_X2 inst_20844 ( .A(net_10142), .ZN(net_9262), .B1(net_5240), .B2(net_4585) );
INV_X4 inst_16430 ( .ZN(net_8842), .A(net_8293) );
NOR2_X2 inst_4018 ( .A1(net_14600), .A2(net_11743), .ZN(net_8030) );
NAND3_X2 inst_5636 ( .ZN(net_20392), .A1(net_18210), .A3(net_17478), .A2(net_17360) );
OAI21_X2 inst_2219 ( .B1(net_9861), .B2(net_9738), .ZN(net_8514), .A(net_5364) );
INV_X4 inst_17854 ( .ZN(net_4478), .A(net_824) );
NAND2_X2 inst_8331 ( .A1(net_21186), .A2(net_20508), .ZN(net_17519) );
NAND2_X2 inst_8884 ( .ZN(net_15152), .A2(net_14695), .A1(net_13774) );
CLKBUF_X2 inst_22569 ( .A(net_22297), .Z(net_22441) );
CLKBUF_X2 inst_21891 ( .A(net_21762), .Z(net_21763) );
OAI22_X2 inst_1284 ( .ZN(net_15117), .B1(net_14653), .A2(net_13252), .B2(net_12799), .A1(net_8978) );
XNOR2_X2 inst_546 ( .ZN(net_728), .A(net_727), .B(net_726) );
INV_X2 inst_18970 ( .ZN(net_9942), .A(net_5228) );
OAI211_X2 inst_2465 ( .ZN(net_14111), .C2(net_13880), .B(net_10461), .A(net_6791), .C1(net_60) );
SDFF_X2 inst_704 ( .Q(net_20858), .SE(net_18837), .SI(net_18825), .D(net_425), .CK(net_22033) );
NAND2_X2 inst_9301 ( .ZN(net_12379), .A1(net_12378), .A2(net_7517) );
INV_X4 inst_16128 ( .ZN(net_2731), .A(net_1372) );
NOR2_X2 inst_4542 ( .ZN(net_6922), .A1(net_3988), .A2(net_3940) );
AOI211_X2 inst_21082 ( .ZN(net_5263), .B(net_4838), .C1(net_2471), .C2(net_1905), .A(net_1827) );
NAND2_X4 inst_7084 ( .A2(net_20683), .A1(net_20682), .ZN(net_15646) );
NAND3_X4 inst_5558 ( .A3(net_19337), .A1(net_19336), .ZN(net_19212), .A2(net_15500) );
NAND2_X2 inst_8285 ( .A2(net_20464), .ZN(net_19772), .A1(net_17527) );
CLKBUF_X2 inst_22795 ( .A(net_22666), .Z(net_22667) );
OAI21_X2 inst_2226 ( .B2(net_10429), .ZN(net_8466), .A(net_4971), .B1(net_571) );
INV_X4 inst_15538 ( .A(net_3073), .ZN(net_2367) );
NAND4_X2 inst_5467 ( .A1(net_20099), .ZN(net_13222), .A4(net_12431), .A3(net_10246), .A2(net_8881) );
INV_X4 inst_17113 ( .ZN(net_14731), .A(net_13058) );
INV_X2 inst_18915 ( .ZN(net_5997), .A(net_5996) );
INV_X4 inst_17299 ( .ZN(net_14657), .A(net_609) );
INV_X4 inst_16652 ( .A(net_5591), .ZN(net_4207) );
INV_X4 inst_17926 ( .A(net_21036), .ZN(net_356) );
NAND2_X4 inst_6986 ( .ZN(net_17852), .A1(net_16856), .A2(net_16687) );
NAND2_X2 inst_11476 ( .ZN(net_3126), .A2(net_3061), .A1(net_110) );
AND2_X2 inst_21282 ( .ZN(net_18928), .A1(net_14547), .A2(net_7322) );
NAND2_X2 inst_8983 ( .ZN(net_14497), .A1(net_14496), .A2(net_12969) );
NAND2_X2 inst_11523 ( .A1(net_6879), .A2(net_3224), .ZN(net_2977) );
INV_X4 inst_17054 ( .ZN(net_5169), .A(net_825) );
INV_X4 inst_13885 ( .ZN(net_7331), .A(net_7330) );
NAND4_X4 inst_5211 ( .ZN(net_20076), .A2(net_16211), .A1(net_16150), .A3(net_16031), .A4(net_15946) );
NAND2_X2 inst_11467 ( .A2(net_3253), .A1(net_3168), .ZN(net_3161) );
OAI221_X2 inst_1342 ( .ZN(net_13927), .C1(net_13926), .B1(net_13926), .B2(net_13226), .A(net_10187), .C2(net_9283) );
NOR2_X4 inst_2971 ( .ZN(net_7624), .A2(net_4490), .A1(net_624) );
NOR2_X2 inst_4549 ( .A1(net_4264), .ZN(net_3967), .A2(net_3966) );
CLKBUF_X2 inst_21958 ( .A(net_21829), .Z(net_21830) );
CLKBUF_X2 inst_21639 ( .A(net_21510), .Z(net_21511) );
NAND2_X4 inst_7483 ( .ZN(net_4022), .A2(net_2439), .A1(net_1881) );
NAND3_X2 inst_6012 ( .ZN(net_14411), .A2(net_14410), .A3(net_13761), .A1(net_12552) );
NAND2_X2 inst_10551 ( .ZN(net_19107), .A2(net_4973), .A1(net_3297) );
NOR2_X2 inst_3933 ( .ZN(net_19746), .A2(net_6949), .A1(net_6717) );
OAI21_X2 inst_1656 ( .A(net_16743), .ZN(net_15796), .B1(net_14835), .B2(net_14821) );
NAND3_X2 inst_5881 ( .A2(net_16037), .ZN(net_15272), .A1(net_14261), .A3(net_13655) );
CLKBUF_X2 inst_22660 ( .A(net_22527), .Z(net_22532) );
OAI21_X2 inst_1881 ( .ZN(net_13546), .B1(net_13509), .A(net_10920), .B2(net_9813) );
INV_X2 inst_18894 ( .A(net_7952), .ZN(net_6102) );
INV_X2 inst_18729 ( .ZN(net_8056), .A(net_8055) );
AOI221_X2 inst_20089 ( .ZN(net_15650), .C1(net_15649), .B1(net_15012), .C2(net_13682), .A(net_10448), .B2(net_8642) );
NAND3_X4 inst_5590 ( .A1(net_19371), .ZN(net_18900), .A2(net_12640), .A3(net_12157) );
NOR2_X4 inst_3034 ( .A1(net_20257), .ZN(net_8325), .A2(net_809) );
XNOR2_X2 inst_295 ( .B(net_21144), .A(net_17485), .ZN(net_17128) );
INV_X4 inst_15507 ( .ZN(net_12070), .A(net_10672) );
INV_X2 inst_18812 ( .A(net_10004), .ZN(net_7322) );
INV_X4 inst_17700 ( .ZN(net_3780), .A(net_309) );
INV_X4 inst_17665 ( .A(net_20875), .ZN(net_4945) );
NAND2_X2 inst_8971 ( .ZN(net_14519), .A2(net_12867), .A1(net_8031) );
INV_X4 inst_13018 ( .ZN(net_16489), .A(net_16424) );
XNOR2_X2 inst_607 ( .A(net_16404), .ZN(net_517), .B(net_516) );
NAND3_X2 inst_6484 ( .ZN(net_11201), .A3(net_9586), .A2(net_6612), .A1(net_4193) );
OAI211_X2 inst_2432 ( .ZN(net_15025), .B(net_15024), .A(net_13036), .C2(net_11355), .C1(net_3484) );
AOI21_X2 inst_20575 ( .B1(net_20339), .ZN(net_14106), .B2(net_11505), .A(net_4186) );
NOR2_X2 inst_4263 ( .ZN(net_6230), .A2(net_6229), .A1(net_5217) );
INV_X4 inst_14698 ( .ZN(net_18804), .A(net_18025) );
NAND3_X2 inst_6693 ( .ZN(net_7701), .A2(net_7700), .A3(net_4566), .A1(net_3706) );
NOR2_X2 inst_5061 ( .A2(net_2636), .ZN(net_994), .A1(net_993) );
NAND2_X2 inst_8273 ( .ZN(net_17736), .A1(net_17476), .A2(net_17354) );
NAND2_X4 inst_7614 ( .ZN(net_2293), .A2(net_1025), .A1(net_343) );
NAND2_X2 inst_10130 ( .ZN(net_12033), .A2(net_8344), .A1(net_6610) );
NOR2_X2 inst_4343 ( .ZN(net_5662), .A1(net_5129), .A2(net_2941) );
NAND2_X2 inst_8560 ( .A1(net_21131), .ZN(net_20619), .A2(net_16562) );
INV_X4 inst_16352 ( .ZN(net_1605), .A(net_858) );
AOI21_X2 inst_20679 ( .B1(net_20569), .ZN(net_12449), .B2(net_6213), .A(net_3042) );
INV_X4 inst_15399 ( .ZN(net_15974), .A(net_15183) );
NAND3_X2 inst_5684 ( .A3(net_20354), .A1(net_20353), .ZN(net_16321), .A2(net_14288) );
NAND2_X2 inst_11537 ( .ZN(net_2924), .A2(net_1912), .A1(net_761) );
NAND3_X2 inst_6627 ( .A3(net_9075), .ZN(net_9040), .A2(net_9039), .A1(net_4504) );
NAND2_X2 inst_11841 ( .ZN(net_2098), .A2(net_1563), .A1(net_168) );
CLKBUF_X2 inst_22495 ( .A(net_22366), .Z(net_22367) );
XNOR2_X2 inst_235 ( .B(net_21128), .A(net_20711), .ZN(net_17520) );
NAND2_X2 inst_11493 ( .ZN(net_7093), .A2(net_3088), .A1(net_1790) );
NAND2_X2 inst_8610 ( .ZN(net_19840), .A2(net_16780), .A1(net_5568) );
INV_X1 inst_19756 ( .ZN(net_6060), .A(net_6059) );
INV_X8 inst_12257 ( .ZN(net_4272), .A(net_2433) );
NAND3_X2 inst_5643 ( .ZN(net_17340), .A3(net_16894), .A2(net_16039), .A1(net_13818) );
NAND3_X2 inst_6750 ( .A1(net_5852), .ZN(net_5795), .A3(net_3319), .A2(net_81) );
INV_X4 inst_12555 ( .ZN(net_18288), .A(net_18247) );
NAND2_X2 inst_8217 ( .ZN(net_17961), .A1(net_17811), .A2(net_17642) );
NAND2_X2 inst_8370 ( .ZN(net_19097), .A1(net_17370), .A2(net_17214) );
NAND2_X2 inst_12051 ( .ZN(net_1251), .A2(net_323), .A1(net_192) );
NOR2_X2 inst_4338 ( .ZN(net_5692), .A2(net_5421), .A1(net_5397) );
NAND2_X2 inst_8806 ( .ZN(net_15648), .A2(net_14998), .A1(net_7301) );
INV_X4 inst_16784 ( .ZN(net_3792), .A(net_3047) );
NAND2_X2 inst_8194 ( .ZN(net_17893), .A2(net_17829), .A1(net_6374) );
NOR2_X4 inst_2835 ( .ZN(net_15487), .A2(net_14797), .A1(net_12214) );
INV_X4 inst_12846 ( .A(net_17245), .ZN(net_17079) );
INV_X4 inst_16907 ( .ZN(net_4773), .A(net_3915) );
NOR3_X2 inst_2731 ( .ZN(net_12849), .A3(net_11906), .A1(net_11128), .A2(net_8145) );
NAND2_X2 inst_10399 ( .ZN(net_7281), .A1(net_7280), .A2(net_7279) );
NAND2_X2 inst_11136 ( .ZN(net_4262), .A2(net_4261), .A1(net_1992) );
NAND2_X2 inst_8663 ( .A2(net_20766), .ZN(net_19639), .A1(net_5294) );
CLKBUF_X2 inst_21426 ( .A(net_21297), .Z(net_21298) );
INV_X4 inst_17971 ( .A(net_20865), .ZN(net_78) );
CLKBUF_X2 inst_22861 ( .A(net_22732), .Z(net_22733) );
AND2_X4 inst_21174 ( .A1(net_12497), .ZN(net_12318), .A2(net_12317) );
NOR2_X2 inst_4813 ( .ZN(net_9929), .A1(net_2559), .A2(net_1436) );
AOI22_X2 inst_20037 ( .ZN(net_7660), .A1(net_7659), .A2(net_6000), .B1(net_5516), .B2(net_2184) );
INV_X4 inst_16960 ( .ZN(net_2007), .A(net_903) );
NAND2_X2 inst_9725 ( .ZN(net_13117), .A1(net_12675), .A2(net_10140) );
AOI211_X2 inst_21080 ( .B(net_6321), .ZN(net_5266), .A(net_5265), .C1(net_2992), .C2(net_2006) );
INV_X2 inst_18488 ( .ZN(net_13422), .A(net_12360) );
INV_X4 inst_15348 ( .A(net_3766), .ZN(net_2593) );
INV_X4 inst_18178 ( .A(net_21206), .ZN(net_16599) );
XNOR2_X2 inst_477 ( .ZN(net_11877), .A(net_11876), .B(net_2473) );
NOR2_X2 inst_3398 ( .ZN(net_15856), .A2(net_15620), .A1(net_12292) );
NOR2_X2 inst_3576 ( .ZN(net_13598), .A1(net_13538), .A2(net_12705) );
XNOR2_X2 inst_423 ( .ZN(net_16505), .A(net_16501), .B(net_1674) );
NAND2_X2 inst_10006 ( .A2(net_11763), .ZN(net_8810), .A1(net_5040) );
INV_X4 inst_17367 ( .ZN(net_12393), .A(net_178) );
SDFF_X2 inst_835 ( .Q(net_21195), .SI(net_17505), .SE(net_125), .CK(net_22316), .D(x6224) );
NOR2_X4 inst_3082 ( .ZN(net_5902), .A1(net_5556), .A2(net_4737) );
NOR2_X2 inst_4137 ( .ZN(net_20407), .A2(net_6939), .A1(net_5062) );
NAND2_X4 inst_6852 ( .A2(net_20154), .A1(net_20153), .ZN(net_18496) );
OR2_X4 inst_1112 ( .ZN(net_6321), .A2(net_143), .A1(net_112) );
NOR2_X2 inst_4081 ( .ZN(net_14441), .A2(net_7221), .A1(net_2589) );
NAND2_X2 inst_9678 ( .ZN(net_12950), .A2(net_10269), .A1(net_10031) );
INV_X4 inst_14571 ( .ZN(net_5820), .A(net_4544) );
NAND2_X2 inst_8869 ( .ZN(net_19838), .A1(net_15297), .A2(net_14244) );
INV_X2 inst_18924 ( .ZN(net_5916), .A(net_5915) );
OAI21_X2 inst_1817 ( .ZN(net_14163), .A(net_11783), .B2(net_10621), .B1(net_7019) );
NAND2_X2 inst_10375 ( .A1(net_18025), .ZN(net_7391), .A2(net_383) );
INV_X4 inst_17997 ( .A(net_21093), .ZN(net_452) );
NAND2_X2 inst_11056 ( .ZN(net_4649), .A2(net_4619), .A1(net_2925) );
INV_X2 inst_19045 ( .ZN(net_4755), .A(net_4754) );
NAND2_X2 inst_10081 ( .A1(net_11451), .ZN(net_8638), .A2(net_8637) );
INV_X4 inst_14715 ( .ZN(net_4455), .A(net_4200) );
NOR2_X4 inst_2871 ( .A1(net_19281), .ZN(net_12336), .A2(net_874) );
NAND2_X4 inst_7475 ( .ZN(net_3553), .A2(net_1752), .A1(net_1064) );
INV_X4 inst_17669 ( .ZN(net_5250), .A(net_2123) );
NOR2_X2 inst_3629 ( .ZN(net_12270), .A2(net_9110), .A1(net_3072) );
AOI21_X2 inst_20756 ( .ZN(net_11215), .B1(net_11214), .B2(net_9807), .A(net_3386) );
DFF_X1 inst_19844 ( .D(net_17405), .CK(net_21606), .Q(x603) );
INV_X4 inst_16297 ( .ZN(net_15506), .A(net_15156) );
INV_X4 inst_12593 ( .ZN(net_20297), .A(net_18116) );
INV_X2 inst_19385 ( .ZN(net_2128), .A(net_2127) );
INV_X4 inst_13370 ( .A(net_11554), .ZN(net_10904) );
INV_X2 inst_19567 ( .ZN(net_19644), .A(net_8868) );
NAND2_X2 inst_9946 ( .A1(net_15692), .ZN(net_9027), .A2(net_5703) );
INV_X4 inst_15427 ( .A(net_5714), .ZN(net_3678) );
AND2_X2 inst_21364 ( .ZN(net_2190), .A2(net_2094), .A1(net_896) );
NAND2_X4 inst_7129 ( .ZN(net_14536), .A2(net_10233), .A1(net_9678) );
NOR2_X2 inst_4414 ( .A1(net_5776), .ZN(net_5038), .A2(net_5037) );
INV_X2 inst_18845 ( .A(net_7305), .ZN(net_6667) );
NAND2_X2 inst_10052 ( .A1(net_11472), .ZN(net_8692), .A2(net_8147) );
CLKBUF_X2 inst_21795 ( .A(net_21666), .Z(net_21667) );
NOR2_X4 inst_3085 ( .ZN(net_5667), .A2(net_4256), .A1(net_809) );
NAND2_X2 inst_8648 ( .A2(net_16614), .ZN(net_16565), .A1(net_16564) );
INV_X4 inst_15337 ( .ZN(net_15224), .A(net_5486) );
NAND2_X4 inst_7620 ( .ZN(net_1703), .A2(net_1327), .A1(net_374) );
INV_X4 inst_16345 ( .ZN(net_14675), .A(net_14600) );
CLKBUF_X2 inst_21466 ( .A(net_21244), .Z(net_21338) );
INV_X2 inst_19005 ( .A(net_6878), .ZN(net_5026) );
INV_X4 inst_16438 ( .ZN(net_2683), .A(net_1240) );
INV_X4 inst_13768 ( .ZN(net_10928), .A(net_7604) );
NAND3_X2 inst_5661 ( .ZN(net_16426), .A3(net_16307), .A2(net_16276), .A1(net_14953) );
NAND2_X2 inst_9918 ( .A2(net_12471), .ZN(net_9298), .A1(net_3335) );
NAND2_X2 inst_11541 ( .A1(net_10521), .ZN(net_2918), .A2(net_2917) );
AND2_X2 inst_21308 ( .ZN(net_13319), .A1(net_10631), .A2(net_8670) );
INV_X4 inst_14120 ( .A(net_6168), .ZN(net_6139) );
NOR2_X2 inst_4292 ( .ZN(net_5990), .A2(net_5989), .A1(net_5958) );
OAI211_X2 inst_2449 ( .ZN(net_14623), .C1(net_14622), .B(net_11977), .A(net_8634), .C2(net_5314) );
NAND2_X2 inst_12083 ( .ZN(net_2773), .A1(net_303), .A2(net_279) );
NAND3_X2 inst_6570 ( .A2(net_20087), .ZN(net_19796), .A1(net_10619), .A3(net_8811) );
INV_X4 inst_14709 ( .ZN(net_4647), .A(net_4241) );
AOI21_X2 inst_20450 ( .ZN(net_15074), .B1(net_14509), .A(net_14293), .B2(net_13015) );
INV_X4 inst_13096 ( .ZN(net_15874), .A(net_15738) );
CLKBUF_X2 inst_21746 ( .A(net_21324), .Z(net_21618) );
OAI21_X4 inst_1431 ( .A(net_16368), .ZN(net_16021), .B1(net_15465), .B2(net_15417) );
NOR2_X2 inst_3760 ( .ZN(net_13105), .A1(net_13070), .A2(net_12033) );
AOI221_X2 inst_20080 ( .B1(net_20688), .ZN(net_16055), .C1(net_16054), .B2(net_15840), .C2(net_15376), .A(net_15276) );
OAI21_X4 inst_1398 ( .A(net_20960), .ZN(net_20623), .B2(net_19345), .B1(net_19344) );
INV_X4 inst_12841 ( .ZN(net_18493), .A(net_17243) );
CLKBUF_X2 inst_21964 ( .A(net_21835), .Z(net_21836) );
NAND2_X4 inst_7639 ( .ZN(net_1143), .A2(net_1142), .A1(net_208) );
INV_X2 inst_18514 ( .ZN(net_12679), .A(net_11577) );
NAND2_X4 inst_7122 ( .A1(net_20597), .A2(net_11018), .ZN(net_10963) );
NAND2_X2 inst_8477 ( .ZN(net_20064), .A1(net_17011), .A2(net_17010) );
NOR2_X4 inst_2849 ( .A1(net_19065), .ZN(net_14857), .A2(net_13576) );
OAI211_X2 inst_2440 ( .ZN(net_14864), .B(net_14863), .C1(net_12504), .A(net_6978), .C2(net_6757) );
INV_X4 inst_13808 ( .ZN(net_9185), .A(net_7656) );
AOI21_X2 inst_20876 ( .ZN(net_8458), .B1(net_8457), .B2(net_7258), .A(net_4894) );
NAND2_X2 inst_9261 ( .ZN(net_20183), .A1(net_15107), .A2(net_12635) );
INV_X4 inst_15533 ( .ZN(net_14086), .A(net_9516) );
NOR2_X4 inst_3327 ( .ZN(net_332), .A1(net_153), .A2(net_37) );
NAND2_X2 inst_10241 ( .ZN(net_10260), .A1(net_7427), .A2(net_6109) );
OAI21_X2 inst_2134 ( .ZN(net_9987), .A(net_9581), .B1(net_8191), .B2(net_5966) );
OAI21_X2 inst_1744 ( .ZN(net_14967), .A(net_14966), .B2(net_12711), .B1(net_8895) );
CLKBUF_X2 inst_22042 ( .A(net_21407), .Z(net_21914) );
INV_X2 inst_19214 ( .ZN(net_3487), .A(net_3486) );
NOR2_X2 inst_4805 ( .ZN(net_3353), .A2(net_2720), .A1(net_90) );
NAND3_X4 inst_5628 ( .A3(net_8644), .ZN(net_5930), .A2(net_4701), .A1(net_2439) );
NAND2_X2 inst_11958 ( .ZN(net_1390), .A2(net_1389), .A1(net_63) );
NOR2_X2 inst_4117 ( .ZN(net_7049), .A1(net_7048), .A2(net_6553) );
NAND2_X2 inst_11311 ( .ZN(net_6727), .A1(net_3867), .A2(net_2378) );
NAND2_X2 inst_9329 ( .ZN(net_13574), .A2(net_9127), .A1(net_8981) );
NAND2_X2 inst_10047 ( .ZN(net_14740), .A1(net_12320), .A2(net_8703) );
NAND2_X2 inst_11198 ( .ZN(net_6992), .A1(net_4863), .A2(net_2825) );
INV_X4 inst_16480 ( .ZN(net_7844), .A(net_5984) );
NAND2_X2 inst_11639 ( .ZN(net_2786), .A2(net_2089), .A1(net_2074) );
NAND2_X4 inst_6940 ( .A2(net_19154), .A1(net_19153), .ZN(net_17588) );
NAND2_X2 inst_11954 ( .A1(net_3780), .ZN(net_3113), .A2(net_200) );
INV_X4 inst_17354 ( .ZN(net_3675), .A(net_352) );
SDFF_X2 inst_712 ( .Q(net_20925), .SE(net_18865), .SI(net_18811), .D(net_617), .CK(net_22022) );
INV_X4 inst_14271 ( .ZN(net_5731), .A(net_5670) );
INV_X8 inst_12436 ( .ZN(net_20445), .A(net_16709) );
NOR2_X4 inst_3111 ( .ZN(net_6579), .A1(net_2855), .A2(net_1544) );
INV_X2 inst_18455 ( .ZN(net_13407), .A(net_13406) );
OAI21_X2 inst_2035 ( .ZN(net_11306), .B2(net_9779), .B1(net_5130), .A(net_4455) );
INV_X4 inst_17121 ( .ZN(net_9917), .A(net_5454) );
AOI21_X2 inst_20786 ( .ZN(net_10551), .B1(net_10550), .A(net_9529), .B2(net_6420) );
INV_X4 inst_16500 ( .ZN(net_6706), .A(net_573) );
CLKBUF_X2 inst_22589 ( .A(net_22460), .Z(net_22461) );
INV_X4 inst_13530 ( .ZN(net_9224), .A(net_9223) );
NAND2_X2 inst_10442 ( .ZN(net_7187), .A2(net_5257), .A1(net_1864) );
NAND2_X2 inst_11569 ( .ZN(net_4974), .A1(net_2887), .A2(net_2769) );
NAND2_X2 inst_11121 ( .ZN(net_14439), .A2(net_4304), .A1(net_2484) );
INV_X4 inst_14686 ( .A(net_11860), .ZN(net_4292) );
INV_X4 inst_16252 ( .ZN(net_6647), .A(net_5438) );
INV_X4 inst_17037 ( .A(net_20859), .ZN(net_4783) );
INV_X4 inst_17023 ( .ZN(net_10759), .A(net_1215) );
INV_X4 inst_12564 ( .ZN(net_18283), .A(net_18196) );
INV_X4 inst_16782 ( .ZN(net_5918), .A(net_5241) );
INV_X4 inst_16529 ( .ZN(net_8273), .A(net_6712) );
NAND3_X2 inst_6483 ( .ZN(net_11227), .A3(net_8348), .A1(net_7512), .A2(net_6039) );
INV_X4 inst_12482 ( .ZN(net_18745), .A(net_18723) );
NAND2_X4 inst_7381 ( .ZN(net_11718), .A2(net_6752), .A1(net_3890) );
XNOR2_X2 inst_525 ( .ZN(net_3582), .B(net_3581), .A(net_2095) );
INV_X2 inst_18735 ( .ZN(net_7943), .A(net_7942) );
CLKBUF_X2 inst_22066 ( .A(net_21937), .Z(net_21938) );
INV_X4 inst_17241 ( .ZN(net_15174), .A(net_14600) );
INV_X4 inst_15360 ( .ZN(net_5550), .A(net_2582) );
NAND2_X2 inst_11774 ( .ZN(net_3749), .A2(net_2053), .A1(net_170) );
INV_X8 inst_12196 ( .ZN(net_16774), .A(net_16338) );
INV_X2 inst_19365 ( .A(net_3175), .ZN(net_2239) );
SDFF_X2 inst_1032 ( .QN(net_21025), .SE(net_17277), .D(net_650), .CK(net_22719), .SI(x2571) );
INV_X8 inst_12424 ( .A(net_20884), .ZN(net_2744) );
NAND2_X2 inst_8985 ( .A1(net_16046), .ZN(net_14488), .A2(net_12743) );
NAND3_X2 inst_6711 ( .ZN(net_7103), .A2(net_7096), .A3(net_4062), .A1(net_3889) );
INV_X4 inst_12638 ( .ZN(net_17913), .A(net_17912) );
AOI21_X2 inst_20901 ( .ZN(net_7718), .B2(net_6172), .B1(net_5243), .A(net_2903) );
INV_X4 inst_16580 ( .ZN(net_6325), .A(net_2996) );
INV_X2 inst_18646 ( .ZN(net_19567), .A(net_9315) );
NAND3_X2 inst_5932 ( .ZN(net_14926), .A1(net_13623), .A3(net_11213), .A2(net_6723) );
NAND2_X4 inst_7585 ( .ZN(net_1559), .A2(net_1193), .A1(net_785) );
NAND2_X2 inst_11682 ( .ZN(net_3142), .A2(net_2343), .A1(net_748) );
NAND2_X2 inst_11148 ( .ZN(net_9964), .A1(net_4212), .A2(net_4083) );
AOI21_X2 inst_20769 ( .ZN(net_10680), .B1(net_9353), .A(net_9148), .B2(net_6957) );
INV_X8 inst_12339 ( .A(net_1645), .ZN(net_825) );
NAND2_X2 inst_11106 ( .ZN(net_11816), .A2(net_2575), .A1(net_86) );
AOI211_X2 inst_21018 ( .ZN(net_15256), .C1(net_14174), .C2(net_14112), .B(net_12108), .A(net_8466) );
INV_X4 inst_17413 ( .ZN(net_2273), .A(net_896) );
OAI21_X2 inst_2269 ( .A(net_9131), .ZN(net_7143), .B2(net_5590), .B1(net_3946) );
OAI21_X2 inst_1780 ( .ZN(net_14666), .B2(net_11936), .B1(net_8761), .A(net_1012) );
INV_X2 inst_18459 ( .ZN(net_13182), .A(net_12222) );
NAND2_X2 inst_11839 ( .ZN(net_1736), .A2(net_1735), .A1(net_247) );
OAI21_X4 inst_1436 ( .B2(net_19358), .B1(net_19357), .A(net_16357), .ZN(net_15920) );
AOI211_X2 inst_21042 ( .ZN(net_13449), .C1(net_13448), .B(net_10285), .C2(net_9879), .A(net_4769) );
SDFF_X2 inst_852 ( .Q(net_21198), .SI(net_17257), .SE(net_125), .CK(net_21545), .D(x6145) );
INV_X4 inst_12792 ( .ZN(net_17958), .A(net_17158) );
AOI21_X2 inst_20321 ( .B1(net_19836), .ZN(net_15863), .B2(net_15831), .A(net_13547) );
NAND3_X2 inst_6663 ( .ZN(net_8449), .A2(net_8448), .A3(net_4528), .A1(net_3956) );
INV_X2 inst_19345 ( .A(net_9514), .ZN(net_2435) );
NOR2_X2 inst_4306 ( .ZN(net_7430), .A2(net_5926), .A1(net_1007) );
OAI21_X4 inst_1474 ( .ZN(net_19820), .B2(net_19236), .B1(net_19235), .A(net_278) );
INV_X4 inst_12528 ( .ZN(net_18427), .A(net_18426) );
INV_X4 inst_17821 ( .A(net_790), .ZN(net_111) );
NAND2_X2 inst_11974 ( .ZN(net_1686), .A2(net_1339), .A1(net_933) );
INV_X4 inst_17563 ( .ZN(net_2618), .A(net_1304) );
OAI21_X2 inst_1920 ( .ZN(net_13027), .A(net_13026), .B1(net_13025), .B2(net_11499) );
NAND2_X2 inst_9022 ( .ZN(net_19788), .A1(net_14160), .A2(net_12247) );
INV_X2 inst_19142 ( .ZN(net_4105), .A(net_4104) );
INV_X4 inst_13269 ( .ZN(net_12568), .A(net_11364) );
INV_X4 inst_18047 ( .A(net_20938), .ZN(net_115) );
INV_X4 inst_12787 ( .A(net_17651), .ZN(net_17580) );
NOR2_X2 inst_4143 ( .ZN(net_8281), .A1(net_7244), .A2(net_3965) );
NOR2_X4 inst_3234 ( .ZN(net_6752), .A1(net_2422), .A2(net_956) );
NAND2_X2 inst_11194 ( .ZN(net_5168), .A1(net_3418), .A2(net_2810) );
NOR3_X2 inst_2639 ( .ZN(net_16001), .A1(net_15703), .A3(net_13718), .A2(net_12859) );
INV_X2 inst_18554 ( .ZN(net_10900), .A(net_10899) );
NAND2_X2 inst_11122 ( .ZN(net_14927), .A1(net_12401), .A2(net_4303) );
INV_X4 inst_15666 ( .ZN(net_5230), .A(net_1600) );
NAND3_X2 inst_5897 ( .ZN(net_20655), .A1(net_14566), .A2(net_12957), .A3(net_12825) );
NAND3_X2 inst_6632 ( .ZN(net_19005), .A2(net_6895), .A3(net_6820), .A1(net_2249) );
OAI211_X2 inst_2542 ( .ZN(net_10827), .B(net_5884), .C2(net_4627), .A(net_3451), .C1(net_1658) );
INV_X4 inst_15864 ( .ZN(net_15071), .A(net_14738) );
CLKBUF_X2 inst_22908 ( .A(net_22578), .Z(net_22780) );
NAND2_X2 inst_11791 ( .ZN(net_6441), .A2(net_1106), .A1(net_573) );
NAND2_X4 inst_6829 ( .A1(net_19955), .ZN(net_18833), .A2(net_17572) );
NAND2_X2 inst_9506 ( .ZN(net_11332), .A1(net_8836), .A2(net_8165) );
NAND2_X4 inst_7567 ( .ZN(net_3225), .A2(net_1662), .A1(net_1661) );
NAND3_X2 inst_6590 ( .ZN(net_9965), .A2(net_9964), .A3(net_9963), .A1(net_5328) );
XNOR2_X2 inst_417 ( .A(net_19446), .ZN(net_16534), .B(net_16470) );
CLKBUF_X2 inst_21844 ( .A(net_21715), .Z(net_21716) );
XNOR2_X2 inst_671 ( .B(net_21159), .A(net_21127), .ZN(net_14910) );
INV_X2 inst_18356 ( .ZN(net_18502), .A(net_18501) );
INV_X4 inst_12733 ( .ZN(net_17679), .A(net_17456) );
INV_X4 inst_13473 ( .ZN(net_11534), .A(net_9630) );
INV_X4 inst_15812 ( .A(net_9940), .ZN(net_8732) );
INV_X4 inst_18083 ( .A(net_21103), .ZN(net_346) );
XOR2_X2 inst_21 ( .B(net_21134), .A(net_16766), .Z(net_16761) );
NAND2_X2 inst_9462 ( .A1(net_14465), .ZN(net_11490), .A2(net_11489) );
INV_X4 inst_14782 ( .A(net_15561), .ZN(net_15537) );
CLKBUF_X2 inst_22089 ( .A(net_21960), .Z(net_21961) );
INV_X2 inst_18364 ( .ZN(net_17990), .A(net_17989) );
INV_X4 inst_17724 ( .ZN(net_1385), .A(net_508) );
INV_X2 inst_18741 ( .ZN(net_9448), .A(net_7908) );
INV_X4 inst_16381 ( .A(net_3505), .ZN(net_1650) );
NAND2_X2 inst_11024 ( .A1(net_20548), .ZN(net_6340), .A2(net_4675) );
NAND2_X2 inst_10286 ( .ZN(net_11724), .A1(net_11296), .A2(net_7947) );
INV_X2 inst_19163 ( .ZN(net_3923), .A(net_3922) );
OAI21_X2 inst_2311 ( .A(net_14700), .ZN(net_5744), .B2(net_5743), .B1(net_2856) );
NOR2_X2 inst_3885 ( .ZN(net_19968), .A2(net_9274), .A1(net_6108) );
NAND2_X4 inst_7703 ( .ZN(net_364), .A2(net_199), .A1(net_82) );
AOI211_X2 inst_21027 ( .C1(net_15524), .ZN(net_14566), .C2(net_12016), .B(net_9086), .A(net_8217) );
INV_X4 inst_17309 ( .ZN(net_8220), .A(net_3201) );
NOR2_X2 inst_3683 ( .A1(net_12428), .ZN(net_11421), .A2(net_6427) );
NOR2_X4 inst_2941 ( .ZN(net_6959), .A2(net_6958), .A1(net_4102) );
INV_X4 inst_13655 ( .ZN(net_11924), .A(net_8147) );
INV_X4 inst_13528 ( .ZN(net_9305), .A(net_7782) );
AOI21_X4 inst_20163 ( .B1(net_19228), .ZN(net_15669), .A(net_12255), .B2(net_750) );
NAND2_X2 inst_9861 ( .A1(net_15012), .ZN(net_9495), .A2(net_5999) );
INV_X8 inst_12351 ( .A(net_20901), .ZN(net_1134) );
NAND2_X2 inst_9203 ( .A1(net_15375), .ZN(net_13075), .A2(net_10289) );
CLKBUF_X2 inst_22423 ( .A(net_22294), .Z(net_22295) );
NAND2_X2 inst_8442 ( .ZN(net_17260), .A2(net_16793), .A1(net_16645) );
INV_X4 inst_17742 ( .A(net_788), .ZN(net_652) );
NAND2_X2 inst_10920 ( .ZN(net_5994), .A1(net_5594), .A2(net_4930) );
NAND2_X2 inst_11930 ( .A2(net_9571), .A1(net_4862), .ZN(net_3326) );
CLKBUF_X2 inst_22786 ( .A(net_22657), .Z(net_22658) );
INV_X2 inst_19635 ( .A(net_19422), .ZN(net_19421) );
INV_X2 inst_18618 ( .ZN(net_9600), .A(net_9599) );
NOR3_X2 inst_2637 ( .A2(net_20222), .A1(net_20221), .ZN(net_16059), .A3(net_15285) );
NAND2_X2 inst_9604 ( .ZN(net_20271), .A1(net_10736), .A2(net_8913) );
INV_X4 inst_16319 ( .ZN(net_1317), .A(net_1316) );
CLKBUF_X2 inst_22812 ( .A(net_22208), .Z(net_22684) );
XNOR2_X2 inst_236 ( .B(net_21122), .ZN(net_17403), .A(net_17402) );
NOR2_X2 inst_4539 ( .ZN(net_5070), .A2(net_4010), .A1(net_165) );
AOI21_X2 inst_20362 ( .ZN(net_15660), .A(net_15659), .B2(net_14937), .B1(net_13751) );
NOR2_X2 inst_3878 ( .ZN(net_11538), .A2(net_11195), .A1(net_9345) );
AOI21_X2 inst_20272 ( .B2(net_20920), .B1(net_19217), .ZN(net_16363), .A(net_13769) );
INV_X4 inst_13295 ( .ZN(net_20127), .A(net_10946) );
DFF_X1 inst_19911 ( .D(net_16845), .CK(net_21578), .Q(x726) );
NAND2_X2 inst_9806 ( .ZN(net_9691), .A2(net_9601), .A1(net_1663) );
SDFF_X2 inst_986 ( .QN(net_21039), .D(net_461), .SE(net_263), .CK(net_22511), .SI(x2344) );
NOR2_X4 inst_3172 ( .ZN(net_7033), .A2(net_3159), .A1(net_874) );
NOR2_X2 inst_4983 ( .ZN(net_12638), .A2(net_1477), .A1(net_1469) );
OAI21_X4 inst_1422 ( .A(net_16385), .ZN(net_16108), .B1(net_15655), .B2(net_15414) );
NAND2_X2 inst_10263 ( .ZN(net_7987), .A2(net_6110), .A1(net_4874) );
NAND2_X2 inst_8337 ( .ZN(net_17509), .A2(net_17230), .A1(net_17111) );
NAND2_X2 inst_9702 ( .ZN(net_19701), .A1(net_10211), .A2(net_10210) );
NAND2_X4 inst_6893 ( .A2(net_18070), .ZN(net_18058), .A1(net_15718) );
NAND2_X2 inst_10522 ( .A1(net_12363), .ZN(net_6852), .A2(net_6851) );
OR2_X2 inst_1221 ( .ZN(net_13648), .A1(net_9014), .A2(net_2987) );
CLKBUF_X2 inst_22266 ( .A(net_21563), .Z(net_22138) );
NAND2_X2 inst_8675 ( .A1(net_19432), .A2(net_16594), .ZN(net_16459) );
INV_X2 inst_19149 ( .ZN(net_4069), .A(net_4068) );
NAND2_X2 inst_7750 ( .ZN(net_18778), .A1(net_18777), .A2(net_18776) );
NAND2_X1 inst_12158 ( .ZN(net_9661), .A1(net_5439), .A2(net_3761) );
INV_X4 inst_15000 ( .A(net_11678), .ZN(net_10945) );
NAND2_X2 inst_7951 ( .ZN(net_20721), .A2(net_18353), .A1(net_17875) );
INV_X4 inst_16005 ( .ZN(net_15842), .A(net_15411) );
INV_X4 inst_15121 ( .A(net_15976), .ZN(net_4189) );
NOR2_X2 inst_5139 ( .A1(net_1271), .A2(net_246), .ZN(net_173) );
INV_X4 inst_16240 ( .ZN(net_19964), .A(net_1372) );
INV_X2 inst_19724 ( .A(net_20793), .ZN(net_20792) );
NOR3_X2 inst_2664 ( .ZN(net_14989), .A3(net_12814), .A1(net_11634), .A2(net_11208) );
NAND2_X2 inst_10793 ( .ZN(net_7270), .A2(net_4265), .A1(net_656) );
INV_X2 inst_19528 ( .A(net_1354), .ZN(net_1032) );
NAND2_X2 inst_8761 ( .ZN(net_19724), .A2(net_15540), .A1(net_14393) );
NAND2_X2 inst_11615 ( .ZN(net_2591), .A2(net_2590), .A1(net_308) );
INV_X4 inst_15463 ( .ZN(net_2471), .A(net_2470) );
NAND3_X2 inst_6757 ( .A2(net_11297), .ZN(net_5678), .A3(net_5677), .A1(net_2550) );
DFF_X1 inst_19841 ( .D(net_17288), .CK(net_21354), .Q(x161) );
INV_X2 inst_19197 ( .A(net_5034), .ZN(net_3626) );
NAND2_X2 inst_8170 ( .ZN(net_17955), .A2(net_17913), .A1(net_17905) );
NAND2_X2 inst_7915 ( .ZN(net_18458), .A2(net_18345), .A1(net_18289) );
NAND3_X2 inst_5862 ( .ZN(net_19867), .A1(net_14178), .A3(net_13733), .A2(net_10375) );
INV_X4 inst_14007 ( .ZN(net_7370), .A(net_3586) );
INV_X2 inst_19138 ( .ZN(net_4140), .A(net_4139) );
NAND2_X2 inst_10966 ( .ZN(net_8225), .A2(net_5057), .A1(net_2585) );
NAND2_X4 inst_7658 ( .ZN(net_1054), .A2(net_935), .A1(net_181) );
INV_X4 inst_18080 ( .A(net_20898), .ZN(net_308) );
NAND2_X2 inst_11381 ( .ZN(net_5889), .A2(net_2285), .A1(net_1606) );
INV_X4 inst_15253 ( .ZN(net_4916), .A(net_2791) );
NAND2_X2 inst_10570 ( .ZN(net_6701), .A2(net_6700), .A1(net_1560) );
AND2_X4 inst_21202 ( .ZN(net_8343), .A1(net_8342), .A2(net_5061) );
NAND2_X2 inst_8051 ( .ZN(net_18217), .A2(net_18144), .A1(net_1701) );
NAND2_X2 inst_8413 ( .A1(net_21109), .ZN(net_17230), .A2(net_16930) );
INV_X4 inst_16090 ( .ZN(net_1527), .A(net_1526) );
NOR2_X2 inst_3932 ( .ZN(net_19285), .A1(net_8651), .A2(net_5478) );
INV_X4 inst_15811 ( .ZN(net_3328), .A(net_1829) );
INV_X4 inst_16162 ( .ZN(net_7528), .A(net_5900) );
CLKBUF_X2 inst_22678 ( .A(net_22549), .Z(net_22550) );
AOI21_X2 inst_20477 ( .A(net_15119), .ZN(net_14947), .B2(net_12723), .B1(net_12586) );
INV_X4 inst_16520 ( .ZN(net_15753), .A(net_14643) );
CLKBUF_X2 inst_21785 ( .A(net_21656), .Z(net_21657) );
INV_X4 inst_13634 ( .ZN(net_11807), .A(net_8219) );
NAND3_X2 inst_6295 ( .ZN(net_12819), .A2(net_10880), .A1(net_8123), .A3(net_7909) );
AOI21_X4 inst_20148 ( .B1(net_19141), .ZN(net_18934), .B2(net_14046), .A(net_12052) );
INV_X4 inst_16736 ( .ZN(net_8748), .A(net_3805) );
INV_X4 inst_17323 ( .ZN(net_1012), .A(net_816) );
AOI211_X2 inst_21063 ( .C1(net_11751), .ZN(net_9891), .B(net_9890), .A(net_7348), .C2(net_6205) );
NAND2_X2 inst_11433 ( .ZN(net_6835), .A2(net_3339), .A1(net_1910) );
NAND2_X2 inst_11429 ( .A1(net_10514), .ZN(net_10131), .A2(net_3751) );
INV_X4 inst_18136 ( .A(net_21131), .ZN(net_500) );
INV_X2 inst_18590 ( .ZN(net_10167), .A(net_10166) );
INV_X4 inst_15980 ( .ZN(net_13070), .A(net_8202) );
CLKBUF_X2 inst_22778 ( .A(net_22649), .Z(net_22650) );
NAND4_X2 inst_5512 ( .ZN(net_10775), .A2(net_10774), .A3(net_10773), .A4(net_7143), .A1(net_7082) );
INV_X4 inst_13112 ( .ZN(net_15632), .A(net_15396) );
NAND2_X2 inst_11973 ( .A1(net_4324), .ZN(net_3393), .A2(net_154) );
INV_X8 inst_12265 ( .ZN(net_4242), .A(net_1571) );
NOR2_X2 inst_3781 ( .A1(net_13785), .A2(net_13458), .ZN(net_10130) );
NAND2_X2 inst_9081 ( .ZN(net_13828), .A1(net_13827), .A2(net_13819) );
NOR2_X2 inst_3552 ( .A1(net_13565), .ZN(net_13067), .A2(net_11226) );
OAI21_X2 inst_1702 ( .ZN(net_15298), .A(net_15297), .B2(net_13601), .B1(net_12582) );
OAI22_X2 inst_1277 ( .ZN(net_16282), .B1(net_16281), .A2(net_16001), .B2(net_14987), .A1(net_4135) );
INV_X4 inst_17802 ( .ZN(net_8596), .A(net_862) );
NOR2_X2 inst_4076 ( .ZN(net_7490), .A1(net_7489), .A2(net_7488) );
OAI21_X2 inst_2092 ( .ZN(net_10201), .B2(net_9465), .A(net_7230), .B1(net_2843) );
NAND3_X4 inst_5586 ( .ZN(net_15380), .A3(net_14052), .A2(net_11567), .A1(net_9639) );
INV_X4 inst_13784 ( .ZN(net_20597), .A(net_7571) );
OAI21_X4 inst_1440 ( .A(net_20889), .ZN(net_15836), .B1(net_15296), .B2(net_13143) );
NAND2_X2 inst_9415 ( .ZN(net_11649), .A2(net_9298), .A1(net_1889) );
INV_X4 inst_13611 ( .ZN(net_20809), .A(net_7063) );
INV_X4 inst_15522 ( .ZN(net_3656), .A(net_1444) );
NAND2_X2 inst_9854 ( .ZN(net_12911), .A2(net_9514), .A1(net_7549) );
INV_X4 inst_13734 ( .ZN(net_7691), .A(net_7690) );
NOR2_X2 inst_3355 ( .ZN(net_20317), .A2(net_17554), .A1(net_17542) );
NAND2_X1 inst_12148 ( .A1(net_17290), .A2(net_16721), .ZN(net_16456) );
NAND2_X2 inst_8179 ( .A1(net_17958), .ZN(net_17934), .A2(net_17933) );
NAND3_X2 inst_6213 ( .ZN(net_13267), .A2(net_13266), .A3(net_13179), .A1(net_10023) );
INV_X4 inst_17214 ( .ZN(net_948), .A(net_242) );
NAND2_X2 inst_8354 ( .ZN(net_17464), .A2(net_17463), .A1(net_17058) );
OAI21_X2 inst_1591 ( .A(net_20848), .B2(net_20147), .B1(net_20146), .ZN(net_16249) );
NOR2_X2 inst_3697 ( .ZN(net_11152), .A1(net_11151), .A2(net_11150) );
CLKBUF_X2 inst_22447 ( .A(net_22318), .Z(net_22319) );
NAND4_X2 inst_5470 ( .ZN(net_13217), .A3(net_11710), .A2(net_11688), .A1(net_8440), .A4(net_7150) );
NAND2_X2 inst_7827 ( .A2(net_20523), .ZN(net_18641), .A1(net_16919) );
NAND2_X2 inst_8312 ( .A1(net_21113), .ZN(net_17583), .A2(net_17338) );
OAI211_X2 inst_2570 ( .B(net_10575), .A(net_9693), .ZN(net_9019), .C1(net_9018), .C2(net_1497) );
INV_X4 inst_12856 ( .ZN(net_17059), .A(net_17058) );
INV_X2 inst_18375 ( .A(net_17607), .ZN(net_17281) );
NOR2_X2 inst_4960 ( .ZN(net_3129), .A2(net_2110), .A1(net_252) );
INV_X4 inst_16811 ( .ZN(net_5716), .A(net_253) );
INV_X4 inst_14205 ( .ZN(net_9573), .A(net_7887) );
NAND2_X2 inst_9098 ( .ZN(net_13775), .A1(net_13774), .A2(net_12499) );
NOR2_X2 inst_3719 ( .ZN(net_20716), .A1(net_11020), .A2(net_9354) );
INV_X2 inst_19560 ( .A(net_2179), .ZN(net_837) );
INV_X2 inst_19553 ( .A(net_2942), .ZN(net_887) );
NOR2_X2 inst_4095 ( .ZN(net_13082), .A2(net_10534), .A1(net_10142) );
XNOR2_X2 inst_74 ( .ZN(net_18735), .B(net_18734), .A(net_17897) );
INV_X4 inst_15926 ( .ZN(net_9926), .A(net_9861) );
CLKBUF_X2 inst_21645 ( .A(net_21516), .Z(net_21517) );
AOI22_X2 inst_20010 ( .ZN(net_12477), .A1(net_11318), .B1(net_9458), .A2(net_9178), .B2(net_6801) );
OAI21_X2 inst_2244 ( .ZN(net_7363), .B2(net_5700), .B1(net_5437), .A(net_320) );
INV_X4 inst_13357 ( .ZN(net_13650), .A(net_10960) );
INV_X2 inst_18760 ( .A(net_12248), .ZN(net_7630) );
INV_X4 inst_14739 ( .ZN(net_12488), .A(net_5575) );
NOR2_X4 inst_3284 ( .ZN(net_2282), .A1(net_1230), .A2(net_61) );
NAND2_X2 inst_11435 ( .ZN(net_5491), .A2(net_3084), .A1(net_388) );
CLKBUF_X2 inst_22041 ( .A(net_21912), .Z(net_21913) );
AOI21_X4 inst_20184 ( .B1(net_19147), .ZN(net_15302), .B2(net_15301), .A(net_8600) );
INV_X2 inst_18652 ( .ZN(net_9221), .A(net_9220) );
NAND3_X2 inst_5719 ( .ZN(net_16137), .A3(net_15686), .A2(net_14318), .A1(net_13696) );
NAND3_X2 inst_5648 ( .ZN(net_16893), .A3(net_16525), .A2(net_16361), .A1(net_15425) );
NOR2_X2 inst_4512 ( .ZN(net_6665), .A2(net_3838), .A1(net_1102) );
INV_X4 inst_14265 ( .A(net_8997), .ZN(net_5724) );
CLKBUF_X2 inst_22443 ( .A(net_22314), .Z(net_22315) );
AOI21_X2 inst_20533 ( .ZN(net_14503), .B1(net_12629), .B2(net_10226), .A(net_652) );
AOI21_X2 inst_20483 ( .B1(net_14949), .ZN(net_14850), .B2(net_13228), .A(net_8694) );
INV_X4 inst_16946 ( .ZN(net_1298), .A(net_809) );
AOI211_X2 inst_20995 ( .C2(net_21236), .C1(net_19762), .ZN(net_16319), .A(net_15280), .B(net_12384) );
NAND2_X2 inst_8483 ( .A2(net_17371), .ZN(net_16976), .A1(net_4661) );
INV_X2 inst_18936 ( .ZN(net_9810), .A(net_7401) );
NAND3_X2 inst_5991 ( .ZN(net_14530), .A3(net_13965), .A1(net_13397), .A2(net_4688) );
NAND2_X2 inst_11234 ( .ZN(net_8256), .A1(net_4502), .A2(net_3085) );
INV_X4 inst_13619 ( .ZN(net_9814), .A(net_8368) );
NAND2_X4 inst_6949 ( .ZN(net_17611), .A1(net_17180), .A2(net_17054) );
INV_X4 inst_17919 ( .A(net_21032), .ZN(net_505) );
INV_X4 inst_16506 ( .ZN(net_9937), .A(net_3929) );
NAND3_X2 inst_5709 ( .ZN(net_16197), .A2(net_15861), .A3(net_15673), .A1(net_5361) );
NAND2_X2 inst_11401 ( .A2(net_3906), .ZN(net_3461), .A1(net_1978) );
CLKBUF_X2 inst_22482 ( .A(net_22353), .Z(net_22354) );
INV_X4 inst_16573 ( .ZN(net_15334), .A(net_14949) );
NAND4_X2 inst_5335 ( .ZN(net_15528), .A4(net_14484), .A3(net_11738), .A2(net_8658), .A1(net_4445) );
OAI211_X2 inst_2397 ( .ZN(net_16081), .B(net_15552), .C1(net_15369), .C2(net_12966), .A(net_11370) );
AOI222_X1 inst_20068 ( .ZN(net_11921), .A1(net_10590), .A2(net_8675), .C1(net_7858), .B2(net_7383), .B1(net_7155), .C2(net_2464) );
INV_X4 inst_12802 ( .A(net_17590), .ZN(net_17224) );
INV_X4 inst_13539 ( .ZN(net_13326), .A(net_9203) );
OR2_X4 inst_1090 ( .ZN(net_8413), .A1(net_4151), .A2(net_4150) );
NAND2_X2 inst_9709 ( .A1(net_12809), .ZN(net_10193), .A2(net_10192) );
NAND2_X2 inst_9088 ( .ZN(net_13796), .A2(net_12484), .A1(net_10386) );
OAI211_X4 inst_2372 ( .C2(net_20904), .A(net_20390), .C1(net_18919), .ZN(net_16553), .B(net_10376) );
CLKBUF_X2 inst_22422 ( .A(net_22293), .Z(net_22294) );
OAI211_X2 inst_2575 ( .C1(net_11654), .ZN(net_8491), .C2(net_8490), .A(net_6862), .B(net_4698) );
INV_X4 inst_17437 ( .A(net_1662), .ZN(net_946) );
NOR2_X2 inst_5007 ( .ZN(net_3203), .A2(net_1588), .A1(net_358) );
AOI211_X2 inst_21049 ( .ZN(net_12456), .C1(net_12238), .C2(net_9185), .B(net_8324), .A(net_5436) );
NAND2_X2 inst_10923 ( .A2(net_7725), .ZN(net_5235), .A1(net_60) );
INV_X4 inst_12496 ( .A(net_18645), .ZN(net_18629) );
INV_X4 inst_13521 ( .ZN(net_9347), .A(net_9346) );
NAND3_X2 inst_5655 ( .A3(net_18880), .A1(net_18879), .ZN(net_16541), .A2(net_16112) );
INV_X4 inst_17071 ( .ZN(net_15553), .A(net_1000) );
INV_X4 inst_16534 ( .A(net_9254), .ZN(net_8739) );
NAND2_X2 inst_11874 ( .ZN(net_2165), .A2(net_1293), .A1(net_63) );
NAND3_X2 inst_5874 ( .A3(net_20835), .A1(net_20834), .ZN(net_15305), .A2(net_12536) );
INV_X2 inst_19490 ( .A(net_10063), .ZN(net_1307) );
NOR2_X4 inst_3126 ( .A1(net_19805), .ZN(net_5687), .A2(net_225) );
INV_X4 inst_12547 ( .ZN(net_18344), .A(net_18287) );
NAND2_X2 inst_8028 ( .ZN(net_18267), .A2(net_18231), .A1(net_17894) );
XNOR2_X2 inst_503 ( .A(net_17097), .ZN(net_8994), .B(net_5668) );
NAND2_X2 inst_8770 ( .ZN(net_15862), .A2(net_15453), .A1(net_13062) );
NAND2_X2 inst_12107 ( .A2(net_21219), .ZN(net_982), .A1(net_215) );
INV_X2 inst_19220 ( .ZN(net_5734), .A(net_4406) );
NAND4_X2 inst_5340 ( .ZN(net_15495), .A4(net_14507), .A2(net_13934), .A1(net_13096), .A3(net_10109) );
NAND2_X2 inst_8724 ( .A1(net_16644), .ZN(net_16106), .A2(net_15867) );
OAI21_X2 inst_1936 ( .ZN(net_12926), .B1(net_12925), .B2(net_9251), .A(net_4532) );
NOR2_X4 inst_3193 ( .ZN(net_5386), .A1(net_3136), .A2(net_3086) );
NAND3_X2 inst_6458 ( .ZN(net_11527), .A1(net_11526), .A3(net_10966), .A2(net_9098) );
OAI21_X2 inst_2099 ( .A(net_11997), .ZN(net_10070), .B2(net_4728), .B1(net_3685) );
NOR2_X2 inst_4069 ( .ZN(net_7658), .A1(net_4996), .A2(net_4759) );
NAND4_X2 inst_5433 ( .A3(net_19811), .ZN(net_19786), .A1(net_13616), .A4(net_13307), .A2(net_9655) );
OR2_X4 inst_1097 ( .ZN(net_3335), .A1(net_3334), .A2(net_2940) );
NAND2_X2 inst_11079 ( .ZN(net_6235), .A2(net_4462), .A1(net_1182) );
INV_X4 inst_15268 ( .A(net_3933), .ZN(net_2766) );
DFF_X1 inst_19866 ( .D(net_17108), .CK(net_21339), .Q(x266) );
INV_X4 inst_16710 ( .ZN(net_14663), .A(net_1292) );
NOR2_X4 inst_2888 ( .A1(net_19157), .ZN(net_10652), .A2(net_3297) );
NAND3_X2 inst_6804 ( .ZN(net_12249), .A3(net_3045), .A1(net_1086), .A2(net_703) );
NAND2_X2 inst_9382 ( .ZN(net_19500), .A2(net_8927), .A1(net_7928) );
INV_X4 inst_12633 ( .A(net_17921), .ZN(net_17920) );
INV_X4 inst_12683 ( .ZN(net_17725), .A(net_17724) );
INV_X8 inst_12330 ( .ZN(net_956), .A(net_110) );
SDFF_X2 inst_967 ( .QN(net_21092), .D(net_491), .SE(net_263), .CK(net_21775), .SI(x1510) );
NAND2_X2 inst_9235 ( .ZN(net_12727), .A1(net_12726), .A2(net_11794) );
INV_X4 inst_13117 ( .A(net_21111), .ZN(net_16857) );
AOI21_X4 inst_20140 ( .B1(net_19234), .ZN(net_16031), .B2(net_16030), .A(net_13667) );
INV_X2 inst_18619 ( .ZN(net_9590), .A(net_9589) );
INV_X4 inst_12665 ( .ZN(net_17804), .A(net_17803) );
AOI21_X2 inst_20354 ( .ZN(net_15700), .B1(net_15699), .B2(net_15009), .A(net_14310) );
INV_X4 inst_16553 ( .A(net_10447), .ZN(net_10309) );
NAND2_X2 inst_7863 ( .ZN(net_18558), .A2(net_18515), .A1(net_18489) );
NAND2_X2 inst_11495 ( .ZN(net_7090), .A2(net_3085), .A1(net_2183) );
INV_X8 inst_12200 ( .ZN(net_20004), .A(net_15583) );
NAND2_X2 inst_12029 ( .A1(net_1339), .ZN(net_1226), .A2(net_103) );
INV_X4 inst_16522 ( .ZN(net_2118), .A(net_1535) );
INV_X4 inst_16469 ( .A(net_11045), .ZN(net_7210) );
OR2_X2 inst_1227 ( .ZN(net_11257), .A2(net_2883), .A1(net_2244) );
OAI21_X2 inst_2324 ( .ZN(net_5650), .B1(net_1918), .A(net_1726), .B2(net_1317) );
NAND3_X2 inst_5856 ( .ZN(net_15401), .A1(net_14602), .A2(net_10792), .A3(net_10749) );
NAND2_X2 inst_9443 ( .ZN(net_15385), .A1(net_11549), .A2(net_11548) );
NAND3_X2 inst_5732 ( .A2(net_20367), .ZN(net_19066), .A1(net_14074), .A3(net_5998) );
AOI21_X2 inst_20429 ( .B2(net_19607), .B1(net_19606), .ZN(net_15189), .A(net_10216) );
INV_X2 inst_19613 ( .A(net_20956), .ZN(net_46) );
NOR2_X4 inst_2897 ( .ZN(net_10882), .A2(net_9353), .A1(net_4704) );
INV_X4 inst_15086 ( .ZN(net_5498), .A(net_2446) );
OAI211_X2 inst_2529 ( .C1(net_13274), .ZN(net_11750), .C2(net_10426), .A(net_9604), .B(net_8713) );
INV_X4 inst_15687 ( .ZN(net_2035), .A(net_2034) );
NAND2_X2 inst_11807 ( .ZN(net_4010), .A2(net_2093), .A1(net_221) );
OAI21_X2 inst_1787 ( .A(net_15699), .ZN(net_14649), .B2(net_11809), .B1(net_9922) );
INV_X2 inst_19087 ( .ZN(net_4572), .A(net_4571) );
NAND2_X4 inst_7274 ( .ZN(net_7476), .A1(net_4590), .A2(net_4030) );
INV_X4 inst_12581 ( .ZN(net_18213), .A(net_18183) );
NAND2_X2 inst_9741 ( .ZN(net_13854), .A2(net_7875), .A1(net_761) );
INV_X4 inst_14290 ( .ZN(net_7401), .A(net_5598) );
NAND3_X2 inst_5943 ( .ZN(net_14898), .A2(net_14897), .A3(net_14878), .A1(net_12556) );
INV_X4 inst_17844 ( .ZN(net_300), .A(net_100) );
NAND2_X2 inst_9891 ( .A2(net_10619), .ZN(net_9412), .A1(net_3495) );
CLKBUF_X2 inst_22681 ( .A(net_22552), .Z(net_22553) );
NAND3_X2 inst_6310 ( .ZN(net_12773), .A1(net_11063), .A3(net_8915), .A2(net_6817) );
OAI21_X2 inst_1540 ( .ZN(net_17902), .B2(net_17852), .A(net_17698), .B1(net_17697) );
NAND2_X2 inst_9493 ( .ZN(net_11433), .A2(net_9419), .A1(net_3870) );
NOR3_X2 inst_2742 ( .ZN(net_19631), .A3(net_11042), .A1(net_10193), .A2(net_5353) );
NOR2_X2 inst_3536 ( .A2(net_13716), .ZN(net_13436), .A1(net_9575) );
NAND2_X4 inst_7515 ( .A1(net_19259), .ZN(net_4081), .A2(net_938) );
NAND4_X4 inst_5243 ( .ZN(net_19228), .A2(net_19089), .A1(net_19088), .A3(net_10975), .A4(net_9995) );
INV_X8 inst_12355 ( .A(net_20870), .ZN(net_776) );
OAI21_X2 inst_2346 ( .ZN(net_4344), .A(net_4343), .B1(net_2926), .B2(net_2350) );
INV_X4 inst_12486 ( .ZN(net_18673), .A(net_18672) );
NAND2_X2 inst_12123 ( .ZN(net_380), .A2(net_164), .A1(net_163) );
INV_X4 inst_13653 ( .A(net_8150), .ZN(net_8149) );
INV_X4 inst_15629 ( .ZN(net_10191), .A(net_9023) );
CLKBUF_X2 inst_21608 ( .A(net_21297), .Z(net_21480) );
NAND2_X4 inst_7250 ( .ZN(net_12838), .A2(net_6981), .A1(net_6672) );
INV_X8 inst_12291 ( .ZN(net_1526), .A(net_1074) );
INV_X4 inst_15680 ( .ZN(net_2651), .A(net_2042) );
NAND2_X4 inst_7363 ( .ZN(net_10573), .A1(net_5498), .A2(net_2199) );
NAND2_X2 inst_9746 ( .ZN(net_19416), .A1(net_10122), .A2(net_8381) );
INV_X4 inst_15279 ( .ZN(net_4076), .A(net_2354) );
CLKBUF_X2 inst_21794 ( .A(net_21369), .Z(net_21666) );
INV_X4 inst_17492 ( .A(net_9131), .ZN(net_8676) );
INV_X4 inst_15135 ( .A(net_7109), .ZN(net_3123) );
INV_X4 inst_16801 ( .ZN(net_8674), .A(net_5449) );
AOI221_X2 inst_20082 ( .ZN(net_19201), .B1(net_16011), .C1(net_15897), .C2(net_15324), .B2(net_14839), .A(net_5287) );
NAND2_X4 inst_7171 ( .ZN(net_11554), .A1(net_9843), .A2(net_7559) );
SDFF_X2 inst_1005 ( .QN(net_21099), .D(net_431), .SE(net_263), .CK(net_21765), .SI(x1413) );
INV_X2 inst_18767 ( .A(net_14642), .ZN(net_7600) );
NAND2_X4 inst_6979 ( .ZN(net_20207), .A2(net_19681), .A1(net_19680) );
INV_X4 inst_14895 ( .ZN(net_3635), .A(net_3634) );
OAI21_X2 inst_1580 ( .B2(net_19046), .B1(net_19045), .ZN(net_18913), .A(net_16395) );
OAI21_X2 inst_1842 ( .ZN(net_14021), .B2(net_11304), .B1(net_11143), .A(net_10082) );
INV_X4 inst_17456 ( .A(net_8596), .ZN(net_828) );
INV_X4 inst_17929 ( .A(net_20992), .ZN(net_361) );
NAND2_X4 inst_7534 ( .ZN(net_2601), .A2(net_1991), .A1(net_1679) );
AND2_X2 inst_21314 ( .A2(net_10477), .ZN(net_8804), .A1(net_7282) );
NAND3_X2 inst_6737 ( .ZN(net_6472), .A3(net_6471), .A1(net_4749), .A2(net_2272) );
NOR2_X2 inst_3703 ( .ZN(net_11098), .A1(net_8865), .A2(net_7382) );
OAI221_X2 inst_1333 ( .B1(net_15506), .ZN(net_15478), .A(net_15036), .B2(net_13959), .C2(net_11292), .C1(net_7292) );
AOI21_X4 inst_20257 ( .ZN(net_5304), .B1(net_4150), .B2(net_2723), .A(net_405) );
INV_X4 inst_12613 ( .ZN(net_18099), .A(net_18089) );
NOR2_X2 inst_3953 ( .ZN(net_8603), .A2(net_8602), .A1(net_7072) );
DFF_X1 inst_19808 ( .D(net_18105), .CK(net_22817), .Q(x1103) );
NAND2_X4 inst_7315 ( .ZN(net_8830), .A2(net_6849), .A1(net_5136) );
AOI21_X2 inst_20670 ( .B1(net_13157), .ZN(net_12858), .A(net_10209), .B2(net_6541) );
OAI21_X2 inst_1551 ( .ZN(net_17724), .A(net_17495), .B1(net_17494), .B2(net_17493) );
INV_X4 inst_14505 ( .ZN(net_7832), .A(net_3839) );
AND2_X4 inst_21156 ( .ZN(net_20669), .A1(net_14303), .A2(net_14302) );
NAND2_X2 inst_9579 ( .ZN(net_12607), .A2(net_10928), .A1(net_4468) );
OR2_X4 inst_1088 ( .ZN(net_5801), .A1(net_4520), .A2(net_4495) );
INV_X4 inst_13200 ( .ZN(net_13869), .A(net_13193) );
INV_X4 inst_15238 ( .ZN(net_2833), .A(net_1578) );
NAND2_X2 inst_8692 ( .A1(net_20944), .ZN(net_16362), .A2(net_16202) );
INV_X4 inst_15498 ( .A(net_15058), .ZN(net_10011) );
NAND2_X2 inst_11672 ( .ZN(net_10631), .A2(net_3203), .A1(net_1233) );
INV_X4 inst_13165 ( .ZN(net_14807), .A(net_14217) );
NAND3_X2 inst_5844 ( .A3(net_19118), .A1(net_19117), .ZN(net_15465), .A2(net_10849) );
NAND2_X2 inst_8781 ( .ZN(net_19495), .A2(net_15290), .A1(net_14248) );
INV_X4 inst_13142 ( .ZN(net_15079), .A(net_14677) );
NAND3_X2 inst_6433 ( .A2(net_11924), .ZN(net_11840), .A3(net_11839), .A1(net_8343) );
AOI21_X2 inst_20508 ( .ZN(net_14632), .B1(net_13462), .B2(net_12077), .A(net_6398) );
NAND2_X2 inst_9922 ( .ZN(net_19923), .A2(net_8520), .A1(net_3117) );
INV_X4 inst_12941 ( .A(net_16965), .ZN(net_16959) );
NOR2_X4 inst_2931 ( .A1(net_18903), .ZN(net_11067), .A2(net_4374) );
INV_X2 inst_18795 ( .ZN(net_12337), .A(net_7441) );
NOR2_X2 inst_4768 ( .ZN(net_5270), .A1(net_4711), .A2(net_2975) );
INV_X4 inst_14483 ( .A(net_6550), .ZN(net_6024) );
OAI211_X2 inst_2530 ( .ZN(net_11749), .A(net_11748), .C1(net_11747), .C2(net_11746), .B(net_8046) );
CLKBUF_X2 inst_22244 ( .A(net_22052), .Z(net_22116) );
OAI21_X4 inst_1503 ( .ZN(net_10411), .A(net_9997), .B2(net_9743), .B1(net_1760) );
INV_X8 inst_12234 ( .ZN(net_5698), .A(net_3438) );
NAND3_X2 inst_5656 ( .ZN(net_16983), .A1(net_16392), .A3(net_16162), .A2(net_15841) );
NAND2_X2 inst_7874 ( .A2(net_19693), .A1(net_19692), .ZN(net_18538) );
NOR2_X2 inst_3802 ( .ZN(net_9856), .A2(net_9855), .A1(net_8431) );
NAND2_X2 inst_8317 ( .ZN(net_17640), .A2(net_17377), .A1(net_17249) );
INV_X4 inst_12926 ( .ZN(net_17359), .A(net_17233) );
CLKBUF_X2 inst_22823 ( .A(net_22691), .Z(net_22695) );
NAND2_X2 inst_10718 ( .ZN(net_20824), .A1(net_5259), .A2(net_3412) );
NAND2_X2 inst_11094 ( .ZN(net_10426), .A2(net_2716), .A1(net_662) );
CLKBUF_X2 inst_22916 ( .A(net_22787), .Z(net_22788) );
SDFF_X2 inst_933 ( .QN(net_21001), .D(net_2511), .SE(net_263), .CK(net_21857), .SI(x3014) );
CLKBUF_X2 inst_21982 ( .A(net_21853), .Z(net_21854) );
CLKBUF_X2 inst_22085 ( .A(net_21956), .Z(net_21957) );
INV_X4 inst_13902 ( .ZN(net_9673), .A(net_8057) );
INV_X4 inst_17566 ( .A(net_4205), .ZN(net_359) );
SDFF_X2 inst_1013 ( .QN(net_21035), .D(net_469), .SE(net_263), .CK(net_21954), .SI(x2401) );
INV_X4 inst_14362 ( .ZN(net_11713), .A(net_5226) );
NOR2_X2 inst_3613 ( .ZN(net_12392), .A1(net_12361), .A2(net_11034) );
NAND2_X2 inst_9439 ( .ZN(net_11557), .A1(net_11556), .A2(net_9444) );
NAND2_X2 inst_7790 ( .A2(net_20471), .ZN(net_18716), .A1(net_18715) );
INV_X4 inst_12870 ( .A(net_17658), .ZN(net_17402) );
INV_X4 inst_14054 ( .A(net_8014), .ZN(net_6249) );
NAND2_X2 inst_8481 ( .A1(net_21111), .ZN(net_17004), .A2(net_16812) );
XNOR2_X2 inst_124 ( .ZN(net_18385), .A(net_18310), .B(net_15585) );
NOR2_X2 inst_3515 ( .ZN(net_13818), .A1(net_13695), .A2(net_13132) );
NAND2_X2 inst_10982 ( .A2(net_4961), .ZN(net_4960), .A1(net_4959) );
INV_X2 inst_19112 ( .A(net_5909), .ZN(net_4459) );
INV_X4 inst_13849 ( .ZN(net_11764), .A(net_7469) );
NAND3_X2 inst_6332 ( .ZN(net_12468), .A3(net_12467), .A2(net_8187), .A1(net_4977) );
OAI22_X2 inst_1270 ( .A2(net_18214), .ZN(net_16883), .B2(net_16882), .A1(net_5706), .B1(net_4376) );
NAND2_X2 inst_11593 ( .ZN(net_2684), .A1(net_2683), .A2(net_2682) );
INV_X4 inst_12531 ( .ZN(net_18409), .A(net_18408) );
CLKBUF_X2 inst_22629 ( .A(net_22500), .Z(net_22501) );
NAND2_X2 inst_8001 ( .ZN(net_18309), .A2(net_18308), .A1(net_17633) );
NOR2_X2 inst_3448 ( .ZN(net_14937), .A1(net_14936), .A2(net_13756) );
NAND3_X2 inst_6088 ( .ZN(net_13948), .A1(net_13156), .A3(net_13072), .A2(net_7753) );
NAND2_X2 inst_10123 ( .A1(net_9926), .ZN(net_8367), .A2(net_8366) );
INV_X4 inst_16856 ( .A(net_7173), .ZN(net_968) );
INV_X4 inst_13032 ( .A(net_16721), .ZN(net_16596) );
AND2_X2 inst_21305 ( .ZN(net_20385), .A1(net_14395), .A2(net_9854) );
INV_X4 inst_14561 ( .ZN(net_8404), .A(net_4566) );
INV_X2 inst_19253 ( .A(net_10976), .ZN(net_3227) );
NAND4_X2 inst_5361 ( .ZN(net_20270), .A2(net_13726), .A3(net_11036), .A4(net_10059), .A1(net_9192) );
INV_X4 inst_15602 ( .A(net_3057), .ZN(net_2894) );
INV_X4 inst_12489 ( .ZN(net_18668), .A(net_18667) );
INV_X4 inst_13049 ( .A(net_16602), .ZN(net_16467) );
INV_X4 inst_15620 ( .A(net_2975), .ZN(net_2155) );
OAI21_X2 inst_2156 ( .A(net_10598), .ZN(net_9272), .B2(net_6392), .B1(net_2778) );
INV_X2 inst_18958 ( .A(net_10261), .ZN(net_5501) );
INV_X4 inst_13389 ( .ZN(net_13399), .A(net_10735) );
NAND2_X1 inst_12142 ( .ZN(net_19042), .A2(net_17100), .A1(net_16921) );
INV_X2 inst_18411 ( .ZN(net_19538), .A(net_16080) );
INV_X2 inst_19009 ( .A(net_6848), .ZN(net_5017) );
NAND4_X2 inst_5417 ( .ZN(net_18966), .A2(net_12433), .A1(net_11137), .A4(net_7131), .A3(net_4045) );
NAND2_X4 inst_7009 ( .A2(net_19143), .A1(net_19142), .ZN(net_17141) );
OAI211_X2 inst_2515 ( .ZN(net_12218), .B(net_12217), .C1(net_12216), .C2(net_12215), .A(net_10179) );
INV_X4 inst_17108 ( .ZN(net_4052), .A(net_399) );
AOI221_X2 inst_20076 ( .C1(net_16404), .ZN(net_16158), .B1(net_15818), .C2(net_15507), .A(net_13688), .B2(net_13114) );
INV_X4 inst_15798 ( .A(net_6861), .ZN(net_3758) );
AND2_X4 inst_21177 ( .ZN(net_11639), .A2(net_11638), .A1(net_10606) );
NAND2_X2 inst_8703 ( .A1(net_16404), .ZN(net_16308), .A2(net_16138) );
INV_X4 inst_12900 ( .A(net_16954), .ZN(net_16946) );
XNOR2_X2 inst_117 ( .ZN(net_18487), .A(net_18322), .B(net_17074) );
NAND4_X4 inst_5172 ( .ZN(net_17019), .A1(net_16387), .A4(net_16160), .A2(net_15966), .A3(net_12206) );
DFF_X1 inst_19883 ( .D(net_17132), .CK(net_22793), .Q(x1291) );
INV_X4 inst_13104 ( .ZN(net_15807), .A(net_15611) );
INV_X4 inst_15195 ( .ZN(net_4670), .A(net_2923) );
NOR2_X2 inst_4106 ( .ZN(net_19793), .A2(net_9010), .A1(net_8232) );
XNOR2_X2 inst_465 ( .B(net_21182), .ZN(net_12876), .A(net_12875) );
OAI21_X2 inst_2304 ( .ZN(net_5858), .A(net_3179), .B2(net_2135), .B1(net_844) );
NAND2_X2 inst_11367 ( .ZN(net_4598), .A1(net_2112), .A2(net_1093) );
NAND2_X2 inst_11701 ( .ZN(net_2304), .A2(net_2303), .A1(net_25) );
OAI21_X2 inst_2173 ( .B2(net_20394), .ZN(net_8923), .A(net_8521), .B1(net_8285) );
AND2_X2 inst_21324 ( .A1(net_9968), .ZN(net_6557), .A2(net_6556) );
NAND2_X4 inst_7048 ( .ZN(net_16799), .A1(net_16358), .A2(net_16351) );
CLKBUF_X2 inst_21450 ( .A(net_21295), .Z(net_21322) );
NOR2_X4 inst_3214 ( .ZN(net_3779), .A1(net_2992), .A2(net_252) );
INV_X4 inst_15039 ( .ZN(net_6153), .A(net_3327) );
INV_X4 inst_16722 ( .A(net_1687), .ZN(net_1499) );
OAI21_X2 inst_1905 ( .ZN(net_13135), .B2(net_9319), .B1(net_6894), .A(net_652) );
INV_X4 inst_12940 ( .ZN(net_16974), .A(net_16636) );
AOI21_X2 inst_20632 ( .ZN(net_13386), .A(net_10074), .B2(net_8699), .B1(net_7052) );
NAND2_X2 inst_11917 ( .ZN(net_3073), .A2(net_1456), .A1(net_284) );
INV_X4 inst_16201 ( .ZN(net_14743), .A(net_1688) );
OAI21_X2 inst_2264 ( .A(net_10066), .ZN(net_7160), .B2(net_7159), .B1(net_2358) );
INV_X4 inst_14925 ( .A(net_4833), .ZN(net_3558) );
INV_X2 inst_18999 ( .ZN(net_5063), .A(net_5062) );
INV_X4 inst_17163 ( .A(net_5250), .ZN(net_1004) );
NOR3_X2 inst_2697 ( .ZN(net_14095), .A2(net_12142), .A3(net_10481), .A1(net_8856) );
XOR2_X2 inst_15 ( .B(net_21135), .Z(net_17026), .A(net_17024) );
NAND2_X2 inst_10196 ( .A2(net_8250), .ZN(net_8139), .A1(net_8138) );
NOR2_X2 inst_3747 ( .ZN(net_10527), .A2(net_8510), .A1(net_7027) );
NAND2_X2 inst_11902 ( .ZN(net_6489), .A1(net_3107), .A2(net_1552) );
AOI21_X2 inst_20910 ( .ZN(net_7362), .A(net_6730), .B2(net_4213), .B1(net_81) );
NOR2_X2 inst_3496 ( .ZN(net_14190), .A1(net_13422), .A2(net_9229) );
INV_X4 inst_16025 ( .A(net_10470), .ZN(net_10292) );
INV_X4 inst_13082 ( .ZN(net_16101), .A(net_15988) );
CLKBUF_X2 inst_22652 ( .A(net_22523), .Z(net_22524) );
NAND2_X2 inst_9830 ( .ZN(net_11602), .A1(net_9617), .A2(net_9536) );
CLKBUF_X2 inst_22030 ( .A(net_21901), .Z(net_21902) );
INV_X4 inst_13642 ( .A(net_8811), .ZN(net_8173) );
OAI21_X2 inst_2123 ( .A(net_13091), .ZN(net_10018), .B2(net_5461), .B1(net_4322) );
NAND2_X2 inst_12020 ( .A1(net_20481), .ZN(net_1039), .A2(net_955) );
AOI21_X2 inst_20919 ( .ZN(net_7299), .A(net_7298), .B2(net_3859), .B1(net_3611) );
NOR2_X2 inst_4918 ( .ZN(net_1885), .A2(net_1479), .A1(net_233) );
NAND2_X2 inst_8615 ( .ZN(net_16613), .A2(net_16612), .A1(net_636) );
INV_X4 inst_17879 ( .A(net_153), .ZN(net_80) );
INV_X4 inst_17736 ( .ZN(net_7268), .A(net_1438) );
INV_X4 inst_14668 ( .ZN(net_11897), .A(net_4325) );
INV_X4 inst_17110 ( .ZN(net_5220), .A(net_2361) );
XNOR2_X2 inst_349 ( .B(net_21211), .ZN(net_16939), .A(net_16750) );
NAND2_X2 inst_10690 ( .ZN(net_11249), .A1(net_6089), .A2(net_6088) );
INV_X4 inst_14145 ( .ZN(net_9532), .A(net_6056) );
INV_X4 inst_14381 ( .A(net_9707), .ZN(net_6151) );
NOR2_X2 inst_4249 ( .ZN(net_6411), .A2(net_6410), .A1(net_2379) );
NOR2_X2 inst_4235 ( .ZN(net_13183), .A2(net_11729), .A1(net_8563) );
INV_X4 inst_13940 ( .A(net_10567), .ZN(net_6819) );
INV_X2 inst_18967 ( .ZN(net_5313), .A(net_5312) );
INV_X4 inst_17190 ( .ZN(net_2230), .A(net_225) );
NAND2_X2 inst_11507 ( .A1(net_7917), .ZN(net_3048), .A2(net_1594) );
INV_X4 inst_13629 ( .ZN(net_13279), .A(net_8308) );
NAND2_X2 inst_9570 ( .ZN(net_10961), .A2(net_7603), .A1(net_3628) );
NAND3_X2 inst_6024 ( .ZN(net_14375), .A3(net_13154), .A2(net_12356), .A1(net_7177) );
INV_X4 inst_17030 ( .ZN(net_13452), .A(net_652) );
INV_X4 inst_14876 ( .ZN(net_4652), .A(net_3683) );
INV_X4 inst_17965 ( .A(net_21202), .ZN(net_1896) );
INV_X4 inst_17584 ( .ZN(net_2539), .A(net_1376) );
INV_X4 inst_15725 ( .ZN(net_1964), .A(net_1963) );
OAI21_X2 inst_2252 ( .ZN(net_7296), .A(net_7295), .B2(net_5498), .B1(net_3602) );
INV_X8 inst_12289 ( .A(net_1783), .ZN(net_1765) );
INV_X4 inst_12514 ( .ZN(net_20062), .A(net_18604) );
INV_X4 inst_16095 ( .ZN(net_2694), .A(net_1522) );
INV_X4 inst_17170 ( .ZN(net_6631), .A(net_120) );
NOR2_X2 inst_4229 ( .A2(net_9692), .ZN(net_8737), .A1(net_7116) );
INV_X4 inst_18253 ( .A(net_20883), .ZN(net_107) );
NAND2_X2 inst_12065 ( .A2(net_20495), .ZN(net_5256), .A1(net_1404) );
NOR3_X2 inst_2763 ( .ZN(net_10460), .A3(net_10459), .A2(net_9890), .A1(net_7286) );
NAND2_X2 inst_10301 ( .ZN(net_11832), .A1(net_7892), .A2(net_7881) );
INV_X4 inst_14334 ( .A(net_14972), .ZN(net_5755) );
NAND3_X2 inst_6798 ( .A3(net_20475), .A2(net_10417), .ZN(net_3448), .A1(net_1492) );
NAND2_X2 inst_10554 ( .ZN(net_6729), .A1(net_6728), .A2(net_6727) );
CLKBUF_X2 inst_21389 ( .A(net_21260), .Z(net_21261) );
AOI211_X2 inst_21044 ( .ZN(net_13188), .A(net_13187), .B(net_13186), .C2(net_11470), .C1(net_6544) );
AOI211_X2 inst_21022 ( .ZN(net_14987), .C1(net_14986), .A(net_13776), .B(net_12768), .C2(net_9038) );
AND2_X4 inst_21248 ( .ZN(net_12353), .A2(net_2424), .A1(net_1778) );
SDFF_X2 inst_761 ( .Q(net_20902), .SE(net_18863), .SI(net_18519), .D(net_587), .CK(net_21489) );
NOR2_X2 inst_4867 ( .ZN(net_4166), .A1(net_2274), .A2(net_2241) );
INV_X4 inst_13342 ( .A(net_11489), .ZN(net_11083) );
NOR2_X4 inst_2803 ( .A2(net_19768), .A1(net_19767), .ZN(net_19625) );
AND2_X2 inst_21363 ( .A1(net_1645), .ZN(net_1316), .A2(net_1134) );
NOR2_X2 inst_4120 ( .ZN(net_7040), .A1(net_4835), .A2(net_2906) );
NAND3_X4 inst_5525 ( .ZN(net_18162), .A3(net_18077), .A2(net_16190), .A1(net_10750) );
NAND2_X2 inst_9211 ( .ZN(net_13045), .A1(net_12307), .A2(net_11286) );
NOR2_X2 inst_5097 ( .ZN(net_10056), .A1(net_117), .A2(net_100) );
NAND2_X2 inst_10003 ( .ZN(net_13808), .A1(net_11441), .A2(net_6881) );
INV_X4 inst_16967 ( .ZN(net_5358), .A(net_901) );
CLKBUF_X2 inst_22878 ( .A(net_22749), .Z(net_22750) );
AND2_X4 inst_21228 ( .ZN(net_9905), .A1(net_6598), .A2(net_4928) );
NOR3_X2 inst_2641 ( .ZN(net_19112), .A1(net_15662), .A3(net_13393), .A2(net_7776) );
AOI21_X2 inst_20507 ( .A(net_15174), .ZN(net_14633), .B2(net_11782), .B1(net_11199) );
AOI21_X2 inst_20384 ( .ZN(net_15502), .B1(net_15501), .A(net_14817), .B2(net_14530) );
AOI21_X4 inst_20205 ( .B1(net_19330), .ZN(net_14760), .B2(net_14759), .A(net_8055) );
OAI21_X2 inst_1638 ( .ZN(net_15952), .B2(net_15228), .A(net_14630), .B1(net_9483) );
NAND3_X2 inst_5771 ( .ZN(net_15895), .A2(net_15405), .A3(net_14739), .A1(net_12642) );
NAND2_X2 inst_11450 ( .A2(net_20529), .ZN(net_4309), .A1(net_2282) );
INV_X4 inst_17518 ( .ZN(net_19026), .A(net_2744) );
INV_X2 inst_19062 ( .ZN(net_4689), .A(net_4344) );
NOR2_X4 inst_3220 ( .ZN(net_5400), .A1(net_3311), .A2(net_2650) );
NAND2_X2 inst_9812 ( .ZN(net_9674), .A2(net_9673), .A1(net_761) );
INV_X2 inst_18885 ( .ZN(net_6164), .A(net_6163) );
NAND2_X2 inst_8177 ( .ZN(net_17937), .A2(net_17921), .A1(net_17273) );
CLKBUF_X2 inst_21780 ( .A(net_21581), .Z(net_21652) );
NAND4_X2 inst_5354 ( .ZN(net_19684), .A3(net_14782), .A1(net_14658), .A4(net_12163), .A2(net_7220) );
NAND2_X2 inst_11983 ( .A2(net_20495), .ZN(net_1788), .A1(net_941) );
CLKBUF_X2 inst_21908 ( .A(net_21779), .Z(net_21780) );
NAND2_X4 inst_7560 ( .ZN(net_3034), .A1(net_1708), .A2(net_216) );
NAND4_X2 inst_5373 ( .ZN(net_15230), .A3(net_14858), .A4(net_14076), .A1(net_14073), .A2(net_13483) );
NOR2_X2 inst_4783 ( .ZN(net_11211), .A1(net_2872), .A2(net_2362) );
CLKBUF_X2 inst_21457 ( .A(net_21279), .Z(net_21329) );
NAND2_X2 inst_9047 ( .ZN(net_14042), .A2(net_12084), .A1(net_7237) );
NAND3_X2 inst_6556 ( .A3(net_10562), .ZN(net_10510), .A2(net_10251), .A1(net_3679) );
NOR2_X2 inst_3862 ( .ZN(net_11479), .A1(net_9438), .A2(net_9437) );
CLKBUF_X2 inst_22736 ( .A(net_21877), .Z(net_22608) );
INV_X4 inst_17531 ( .A(net_3491), .ZN(net_3009) );
NAND3_X2 inst_6532 ( .ZN(net_10596), .A3(net_10595), .A1(net_10428), .A2(net_9373) );
NAND4_X2 inst_5304 ( .ZN(net_15868), .A1(net_15299), .A2(net_14874), .A4(net_14523), .A3(net_13811) );
NAND2_X2 inst_10847 ( .ZN(net_6745), .A1(net_4464), .A2(net_4017) );
NAND2_X2 inst_10482 ( .ZN(net_10440), .A2(net_7006), .A1(net_6840) );
INV_X4 inst_14326 ( .ZN(net_7957), .A(net_3938) );
XNOR2_X2 inst_633 ( .ZN(net_16095), .B(net_488), .A(net_437) );
INV_X4 inst_18263 ( .A(net_19437), .ZN(net_19434) );
INV_X4 inst_12837 ( .ZN(net_17480), .A(net_17275) );
CLKBUF_X2 inst_22946 ( .A(net_21368), .Z(net_22818) );
NOR2_X2 inst_4060 ( .ZN(net_9343), .A2(net_7832), .A1(net_4707) );
OAI21_X2 inst_2285 ( .B2(net_7663), .A(net_6962), .ZN(net_6543), .B1(net_2035) );
NAND2_X2 inst_10500 ( .A1(net_14185), .A2(net_11113), .ZN(net_6921) );
NOR2_X2 inst_4478 ( .ZN(net_6952), .A2(net_5292), .A1(net_3697) );
NOR2_X2 inst_3344 ( .ZN(net_18102), .A2(net_18101), .A1(net_13469) );
NOR2_X2 inst_3447 ( .ZN(net_14939), .A2(net_13627), .A1(net_13065) );
NAND2_X2 inst_11878 ( .A1(net_3350), .ZN(net_2940), .A2(net_107) );
INV_X4 inst_15968 ( .ZN(net_7968), .A(net_7427) );
INV_X4 inst_17517 ( .ZN(net_3115), .A(net_1848) );
NAND2_X4 inst_7199 ( .ZN(net_11941), .A1(net_9801), .A2(net_7865) );
NOR2_X2 inst_4862 ( .A1(net_3780), .ZN(net_2257), .A2(net_1398) );
INV_X2 inst_19096 ( .ZN(net_10030), .A(net_4543) );
NOR2_X2 inst_4663 ( .ZN(net_5278), .A1(net_3284), .A2(net_3182) );
INV_X4 inst_15220 ( .ZN(net_5034), .A(net_2869) );
NAND2_X2 inst_10360 ( .ZN(net_10248), .A1(net_6346), .A2(net_5810) );
SDFF_X2 inst_882 ( .Q(net_21203), .SI(net_16961), .SE(net_125), .CK(net_21391), .D(x6012) );
INV_X4 inst_13935 ( .ZN(net_8941), .A(net_6843) );
NAND2_X2 inst_9848 ( .A1(net_11472), .ZN(net_9534), .A2(net_7500) );
INV_X4 inst_13700 ( .ZN(net_9422), .A(net_7883) );
CLKBUF_X2 inst_21527 ( .A(net_21287), .Z(net_21399) );
NOR2_X4 inst_2938 ( .A2(net_12877), .ZN(net_8613), .A1(net_6608) );
NAND2_X2 inst_9116 ( .ZN(net_13570), .A1(net_13569), .A2(net_13568) );
NAND2_X4 inst_6931 ( .A2(net_18995), .A1(net_18994), .ZN(net_17648) );
NOR2_X2 inst_5083 ( .ZN(net_8851), .A1(net_1961), .A2(net_816) );
INV_X4 inst_15627 ( .ZN(net_2813), .A(net_2146) );
INV_X4 inst_15802 ( .ZN(net_9666), .A(net_761) );
NOR2_X2 inst_4855 ( .A1(net_2712), .ZN(net_2298), .A2(net_2045) );
OAI21_X4 inst_1374 ( .B2(net_20004), .B1(net_20003), .ZN(net_16406), .A(net_16395) );
CLKBUF_X2 inst_21493 ( .A(net_21342), .Z(net_21365) );
INV_X4 inst_17893 ( .ZN(net_65), .A(net_64) );
OAI211_X2 inst_2510 ( .ZN(net_12485), .C2(net_10728), .C1(net_8798), .B(net_6063), .A(net_5037) );
NAND2_X2 inst_9046 ( .ZN(net_14043), .A2(net_12075), .A1(net_10168) );
NAND3_X2 inst_6316 ( .ZN(net_12573), .A2(net_11293), .A3(net_7615), .A1(net_4825) );
INV_X4 inst_15882 ( .ZN(net_4511), .A(net_1780) );
AND2_X2 inst_21339 ( .A2(net_12353), .A1(net_11776), .ZN(net_3158) );
INV_X4 inst_16532 ( .ZN(net_10015), .A(net_120) );
INV_X2 inst_19177 ( .ZN(net_19991), .A(net_3801) );
NAND2_X2 inst_11548 ( .ZN(net_2877), .A1(net_2876), .A2(net_2875) );
INV_X4 inst_14199 ( .ZN(net_8324), .A(net_5967) );
CLKBUF_X2 inst_22808 ( .A(net_21918), .Z(net_22680) );
INV_X4 inst_15184 ( .ZN(net_13785), .A(net_11446) );
INV_X2 inst_19274 ( .ZN(net_2990), .A(net_2989) );
INV_X4 inst_16322 ( .ZN(net_2066), .A(net_1314) );
NAND3_X2 inst_6780 ( .ZN(net_4469), .A2(net_4468), .A1(net_3288), .A3(net_905) );
INV_X2 inst_18577 ( .ZN(net_10404), .A(net_10403) );
NOR2_X2 inst_4398 ( .ZN(net_8366), .A2(net_7748), .A1(net_3792) );
NOR2_X2 inst_4165 ( .ZN(net_20748), .A2(net_12409), .A1(net_9254) );
OAI21_X2 inst_2272 ( .B1(net_20579), .A(net_14055), .ZN(net_7139), .B2(net_7138) );
OAI21_X2 inst_1608 ( .A(net_16259), .ZN(net_16145), .B1(net_15750), .B2(net_15237) );
NAND2_X2 inst_11631 ( .A1(net_3458), .ZN(net_2527), .A2(net_1160) );
OAI21_X4 inst_1484 ( .ZN(net_20840), .B2(net_19966), .B1(net_19965), .A(net_14159) );
SDFF_X2 inst_856 ( .Q(net_21133), .D(net_17152), .SE(net_263), .CK(net_21402), .SI(x3863) );
NAND3_X2 inst_5677 ( .A3(net_19890), .A1(net_19889), .ZN(net_16338), .A2(net_16110) );
INV_X2 inst_18537 ( .A(net_13322), .ZN(net_11044) );

endmodule
